module tt_um_risc_v_wg_swc1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire clknet_leaf_0_clk;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire \fpga_top.bus_gather.d_write_data[0] ;
 wire \fpga_top.bus_gather.d_write_data[10] ;
 wire \fpga_top.bus_gather.d_write_data[11] ;
 wire \fpga_top.bus_gather.d_write_data[12] ;
 wire \fpga_top.bus_gather.d_write_data[13] ;
 wire \fpga_top.bus_gather.d_write_data[14] ;
 wire \fpga_top.bus_gather.d_write_data[15] ;
 wire \fpga_top.bus_gather.d_write_data[16] ;
 wire \fpga_top.bus_gather.d_write_data[17] ;
 wire \fpga_top.bus_gather.d_write_data[18] ;
 wire \fpga_top.bus_gather.d_write_data[19] ;
 wire \fpga_top.bus_gather.d_write_data[1] ;
 wire \fpga_top.bus_gather.d_write_data[20] ;
 wire \fpga_top.bus_gather.d_write_data[21] ;
 wire \fpga_top.bus_gather.d_write_data[22] ;
 wire \fpga_top.bus_gather.d_write_data[23] ;
 wire \fpga_top.bus_gather.d_write_data[24] ;
 wire \fpga_top.bus_gather.d_write_data[25] ;
 wire \fpga_top.bus_gather.d_write_data[26] ;
 wire \fpga_top.bus_gather.d_write_data[27] ;
 wire \fpga_top.bus_gather.d_write_data[28] ;
 wire \fpga_top.bus_gather.d_write_data[29] ;
 wire \fpga_top.bus_gather.d_write_data[2] ;
 wire \fpga_top.bus_gather.d_write_data[30] ;
 wire \fpga_top.bus_gather.d_write_data[31] ;
 wire \fpga_top.bus_gather.d_write_data[3] ;
 wire \fpga_top.bus_gather.d_write_data[4] ;
 wire \fpga_top.bus_gather.d_write_data[5] ;
 wire \fpga_top.bus_gather.d_write_data[6] ;
 wire \fpga_top.bus_gather.d_write_data[7] ;
 wire \fpga_top.bus_gather.d_write_data[8] ;
 wire \fpga_top.bus_gather.d_write_data[9] ;
 wire \fpga_top.bus_gather.i_read_adr[10] ;
 wire \fpga_top.bus_gather.i_read_adr[11] ;
 wire \fpga_top.bus_gather.i_read_adr[12] ;
 wire \fpga_top.bus_gather.i_read_adr[13] ;
 wire \fpga_top.bus_gather.i_read_adr[14] ;
 wire \fpga_top.bus_gather.i_read_adr[15] ;
 wire \fpga_top.bus_gather.i_read_adr[16] ;
 wire \fpga_top.bus_gather.i_read_adr[17] ;
 wire \fpga_top.bus_gather.i_read_adr[18] ;
 wire \fpga_top.bus_gather.i_read_adr[19] ;
 wire \fpga_top.bus_gather.i_read_adr[20] ;
 wire \fpga_top.bus_gather.i_read_adr[21] ;
 wire \fpga_top.bus_gather.i_read_adr[22] ;
 wire \fpga_top.bus_gather.i_read_adr[23] ;
 wire \fpga_top.bus_gather.i_read_adr[24] ;
 wire \fpga_top.bus_gather.i_read_adr[25] ;
 wire \fpga_top.bus_gather.i_read_adr[26] ;
 wire \fpga_top.bus_gather.i_read_adr[27] ;
 wire \fpga_top.bus_gather.i_read_adr[28] ;
 wire \fpga_top.bus_gather.i_read_adr[29] ;
 wire \fpga_top.bus_gather.i_read_adr[2] ;
 wire \fpga_top.bus_gather.i_read_adr[30] ;
 wire \fpga_top.bus_gather.i_read_adr[31] ;
 wire \fpga_top.bus_gather.i_read_adr[3] ;
 wire \fpga_top.bus_gather.i_read_adr[4] ;
 wire \fpga_top.bus_gather.i_read_adr[5] ;
 wire \fpga_top.bus_gather.i_read_adr[6] ;
 wire \fpga_top.bus_gather.i_read_adr[7] ;
 wire \fpga_top.bus_gather.i_read_adr[8] ;
 wire \fpga_top.bus_gather.i_read_adr[9] ;
 wire \fpga_top.bus_gather.u_read_adr[10] ;
 wire \fpga_top.bus_gather.u_read_adr[11] ;
 wire \fpga_top.bus_gather.u_read_adr[12] ;
 wire \fpga_top.bus_gather.u_read_adr[13] ;
 wire \fpga_top.bus_gather.u_read_adr[14] ;
 wire \fpga_top.bus_gather.u_read_adr[15] ;
 wire \fpga_top.bus_gather.u_read_adr[16] ;
 wire \fpga_top.bus_gather.u_read_adr[17] ;
 wire \fpga_top.bus_gather.u_read_adr[18] ;
 wire \fpga_top.bus_gather.u_read_adr[19] ;
 wire \fpga_top.bus_gather.u_read_adr[20] ;
 wire \fpga_top.bus_gather.u_read_adr[21] ;
 wire \fpga_top.bus_gather.u_read_adr[22] ;
 wire \fpga_top.bus_gather.u_read_adr[23] ;
 wire \fpga_top.bus_gather.u_read_adr[24] ;
 wire \fpga_top.bus_gather.u_read_adr[25] ;
 wire \fpga_top.bus_gather.u_read_adr[26] ;
 wire \fpga_top.bus_gather.u_read_adr[27] ;
 wire \fpga_top.bus_gather.u_read_adr[28] ;
 wire \fpga_top.bus_gather.u_read_adr[29] ;
 wire \fpga_top.bus_gather.u_read_adr[2] ;
 wire \fpga_top.bus_gather.u_read_adr[30] ;
 wire \fpga_top.bus_gather.u_read_adr[31] ;
 wire \fpga_top.bus_gather.u_read_adr[3] ;
 wire \fpga_top.bus_gather.u_read_adr[4] ;
 wire \fpga_top.bus_gather.u_read_adr[5] ;
 wire \fpga_top.bus_gather.u_read_adr[6] ;
 wire \fpga_top.bus_gather.u_read_adr[7] ;
 wire \fpga_top.bus_gather.u_read_adr[8] ;
 wire \fpga_top.bus_gather.u_read_adr[9] ;
 wire \fpga_top.cmd_ld_ma ;
 wire \fpga_top.cmd_st_ma ;
 wire \fpga_top.cpu_run_state ;
 wire \fpga_top.cpu_start ;
 wire \fpga_top.cpu_start_adr[10] ;
 wire \fpga_top.cpu_start_adr[11] ;
 wire \fpga_top.cpu_start_adr[12] ;
 wire \fpga_top.cpu_start_adr[13] ;
 wire \fpga_top.cpu_start_adr[14] ;
 wire \fpga_top.cpu_start_adr[15] ;
 wire \fpga_top.cpu_start_adr[16] ;
 wire \fpga_top.cpu_start_adr[17] ;
 wire \fpga_top.cpu_start_adr[18] ;
 wire \fpga_top.cpu_start_adr[19] ;
 wire \fpga_top.cpu_start_adr[20] ;
 wire \fpga_top.cpu_start_adr[21] ;
 wire \fpga_top.cpu_start_adr[22] ;
 wire \fpga_top.cpu_start_adr[23] ;
 wire \fpga_top.cpu_start_adr[24] ;
 wire \fpga_top.cpu_start_adr[25] ;
 wire \fpga_top.cpu_start_adr[26] ;
 wire \fpga_top.cpu_start_adr[27] ;
 wire \fpga_top.cpu_start_adr[28] ;
 wire \fpga_top.cpu_start_adr[29] ;
 wire \fpga_top.cpu_start_adr[2] ;
 wire \fpga_top.cpu_start_adr[30] ;
 wire \fpga_top.cpu_start_adr[31] ;
 wire \fpga_top.cpu_start_adr[3] ;
 wire \fpga_top.cpu_start_adr[4] ;
 wire \fpga_top.cpu_start_adr[5] ;
 wire \fpga_top.cpu_start_adr[6] ;
 wire \fpga_top.cpu_start_adr[7] ;
 wire \fpga_top.cpu_start_adr[8] ;
 wire \fpga_top.cpu_start_adr[9] ;
 wire \fpga_top.cpu_top.alu_code[0] ;
 wire \fpga_top.cpu_top.alu_code[1] ;
 wire \fpga_top.cpu_top.alu_code[2] ;
 wire \fpga_top.cpu_top.alui_shamt[0] ;
 wire \fpga_top.cpu_top.alui_shamt[1] ;
 wire \fpga_top.cpu_top.alui_shamt[2] ;
 wire \fpga_top.cpu_top.alui_shamt[3] ;
 wire \fpga_top.cpu_top.alui_shamt[4] ;
 wire \fpga_top.cpu_top.br_ofs[10] ;
 wire \fpga_top.cpu_top.br_ofs[11] ;
 wire \fpga_top.cpu_top.br_ofs[12] ;
 wire \fpga_top.cpu_top.br_ofs[1] ;
 wire \fpga_top.cpu_top.br_ofs[2] ;
 wire \fpga_top.cpu_top.br_ofs[3] ;
 wire \fpga_top.cpu_top.br_ofs[4] ;
 wire \fpga_top.cpu_top.br_ofs[5] ;
 wire \fpga_top.cpu_top.br_ofs[6] ;
 wire \fpga_top.cpu_top.br_ofs[7] ;
 wire \fpga_top.cpu_top.br_ofs[8] ;
 wire \fpga_top.cpu_top.br_ofs[9] ;
 wire \fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[0] ;
 wire \fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[1] ;
 wire \fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[2] ;
 wire \fpga_top.cpu_top.cpu_state_machine.cpu_state[0] ;
 wire \fpga_top.cpu_top.cpu_state_machine.cpu_state[1] ;
 wire \fpga_top.cpu_top.cpu_state_machine.cpu_state[2] ;
 wire \fpga_top.cpu_top.csr_meie ;
 wire \fpga_top.cpu_top.csr_mepc_ex[10] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[11] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[12] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[13] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[14] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[15] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[16] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[17] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[18] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[19] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[20] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[21] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[22] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[23] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[24] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[25] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[26] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[27] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[28] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[29] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[2] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[30] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[31] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[3] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[4] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[5] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[6] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[7] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[8] ;
 wire \fpga_top.cpu_top.csr_mepc_ex[9] ;
 wire \fpga_top.cpu_top.csr_msie ;
 wire \fpga_top.cpu_top.csr_mtie ;
 wire \fpga_top.cpu_top.csr_rmie ;
 wire \fpga_top.cpu_top.csr_uimm[0] ;
 wire \fpga_top.cpu_top.csr_uimm[1] ;
 wire \fpga_top.cpu_top.csr_uimm[2] ;
 wire \fpga_top.cpu_top.csr_uimm[3] ;
 wire \fpga_top.cpu_top.csr_uimm[4] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[0] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[10] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[11] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[1] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[2] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[3] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[4] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[5] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[6] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[7] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[8] ;
 wire \fpga_top.cpu_top.csr_wadr_mon[9] ;
 wire \fpga_top.cpu_top.csr_wdata_mon[0] ;
 wire \fpga_top.cpu_top.csr_wdata_mon[1] ;
 wire \fpga_top.cpu_top.data_rw_mem.data_state[0] ;
 wire \fpga_top.cpu_top.data_rw_mem.data_state[1] ;
 wire \fpga_top.cpu_top.data_rw_mem.data_state[2] ;
 wire \fpga_top.cpu_top.data_rw_mem.dma_io_radr_en ;
 wire \fpga_top.cpu_top.data_rw_mem.dma_io_ren_wb ;
 wire \fpga_top.cpu_top.data_rw_mem.next_data_state[0] ;
 wire \fpga_top.cpu_top.data_rw_mem.next_data_state[1] ;
 wire \fpga_top.cpu_top.data_rw_mem.next_data_state[2] ;
 wire \fpga_top.cpu_top.data_rw_mem.req_hw_dly ;
 wire \fpga_top.cpu_top.data_rw_mem.req_w_dly ;
 wire \fpga_top.cpu_top.data_rw_mem.unsigned_bit_dly ;
 wire \fpga_top.cpu_top.data_rw_mem.wbk_rd_reg_ma ;
 wire \fpga_top.cpu_top.decoder.illegal_ops_inst[0] ;
 wire \fpga_top.cpu_top.decoder.illegal_ops_inst[1] ;
 wire \fpga_top.cpu_top.decoder.illegal_ops_inst[2] ;
 wire \fpga_top.cpu_top.decoder.illegal_ops_inst[3] ;
 wire \fpga_top.cpu_top.decoder.illegal_ops_inst[4] ;
 wire \fpga_top.cpu_top.decoder.illegal_ops_inst[5] ;
 wire \fpga_top.cpu_top.decoder.illegal_ops_inst[6] ;
 wire \fpga_top.cpu_top.execution.alu_sra[31] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mcause[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mcause[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mcause[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mcause[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mcause[4] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mcause[5] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mcause[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mpie ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mpp[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mpp[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[10] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[11] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[12] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[13] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[14] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[15] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[16] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[17] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[18] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[19] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[20] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[21] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[22] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[23] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[24] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[25] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[26] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[27] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[28] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[29] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[30] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[31] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[4] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[5] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[7] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[8] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mscrach[9] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[10] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[11] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[12] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[13] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[14] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[15] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[16] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[17] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[18] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[19] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[20] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[21] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[22] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[23] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[24] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[25] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[26] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[27] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[28] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[29] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[30] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[31] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[7] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[8] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mstatush[9] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[10] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[11] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[12] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[13] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[14] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[15] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[16] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[17] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[18] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[19] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[20] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[21] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[22] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[23] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[24] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[25] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[26] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[27] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[28] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[29] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[30] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[31] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[4] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[5] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[7] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[8] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtval[9] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[10] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[11] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[12] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[13] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[14] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[15] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[16] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[17] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[18] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[19] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[20] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[22] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[23] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[24] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[25] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[26] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[27] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[28] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[29] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[30] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[31] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[4] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[5] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[7] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[8] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_mtvec[9] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[10] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[11] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[12] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[13] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[14] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[15] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[16] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[17] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[18] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[19] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[20] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[21] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[22] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[23] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[24] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[25] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[26] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[27] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[28] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[29] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[30] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[31] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[4] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[5] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[7] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[8] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_rd_data[9] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sie ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_spie ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_spp ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[10] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[11] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[12] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[13] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[14] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[15] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[16] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[17] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[18] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[19] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[20] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[21] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[22] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[23] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[24] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[25] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[26] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[27] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[28] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[29] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[30] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[31] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[4] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[5] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[7] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[8] ;
 wire \fpga_top.cpu_top.execution.csr_array.csr_sscrach[9] ;
 wire \fpga_top.cpu_top.execution.csr_array.frc_cntr_val_leq ;
 wire \fpga_top.cpu_top.execution.csr_array.g_interrupt ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[10] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[11] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[12] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[13] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[14] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[15] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[16] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[17] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[18] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[19] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[20] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[21] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[22] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[23] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[24] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[25] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[26] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[27] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[28] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[29] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[30] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[31] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[4] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[5] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[7] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[8] ;
 wire \fpga_top.cpu_top.execution.csr_array.pc_excep2[9] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[0] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[10] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[11] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[12] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[13] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[14] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[15] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[16] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[17] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[18] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[19] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[1] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[20] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[21] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[22] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[23] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[24] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[25] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[26] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[27] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[28] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[29] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[2] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[30] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[3] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[4] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[5] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[6] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[7] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[8] ;
 wire \fpga_top.cpu_top.execution.csr_array.rs1_sel[9] ;
 wire \fpga_top.cpu_top.inst_mem_read.imr_stat ;
 wire \fpga_top.cpu_top.inst_mem_read.imr_stat_dly ;
 wire \fpga_top.cpu_top.pc_stage.cmd_ebreak_pc_pre ;
 wire \fpga_top.cpu_top.pc_stage.cmd_ecall_pc_pre ;
 wire \fpga_top.cpu_top.pc_stage.cpu_adr_ld ;
 wire \fpga_top.cpu_top.pc_stage.frc_cntr_val_leq_lat ;
 wire \fpga_top.cpu_top.pc_stage.frc_cntr_val_leq_latch ;
 wire \fpga_top.cpu_top.pc_stage.g_interrupt_latch ;
 wire \fpga_top.cpu_top.pc_stage.pc_int_ecall_syn_state ;
 wire \fpga_top.cpu_top.register_file.inst_rs[4] ;
 wire \fpga_top.cpu_top.register_file.inst_rs[5] ;
 wire \fpga_top.cpu_top.register_file.inst_rs[6] ;
 wire \fpga_top.cpu_top.register_file.inst_rs[7] ;
 wire \fpga_top.cpu_top.register_file.inst_rs[8] ;
 wire \fpga_top.cpu_top.register_file.next_rfr_state[0] ;
 wire \fpga_top.cpu_top.register_file.next_rfr_state[1] ;
 wire \fpga_top.cpu_top.register_file.next_rfr_state[2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[0][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[10][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[11][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[12][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[13][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[14][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[15][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[16][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[17][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[18][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[19][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[1][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[20][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[21][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[22][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[23][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[24][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[25][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[26][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[27][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[28][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[29][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[2][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[30][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[31][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[3][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[4][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[5][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[6][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[7][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[8][9] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][0] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][10] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][11] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][12] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][13] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][14] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][15] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][16] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][17] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][18] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][19] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][1] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][20] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][21] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][22] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][23] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][24] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][25] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][26] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][27] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][28] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][29] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][2] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][30] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][31] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][3] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][4] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][5] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][6] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][7] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][8] ;
 wire \fpga_top.cpu_top.register_file.rf_1r1w.ram[9][9] ;
 wire \fpga_top.cpu_top.register_file.rfr_state[0] ;
 wire \fpga_top.cpu_top.register_file.rfr_state[1] ;
 wire \fpga_top.cpu_top.register_file.rfr_state[2] ;
 wire \fpga_top.dbg_bpoint_en[0] ;
 wire \fpga_top.dbg_bpoint_en[1] ;
 wire \fpga_top.dbg_bpoint_en[2] ;
 wire \fpga_top.dma_io_wadr_u[14] ;
 wire \fpga_top.dma_io_wadr_u[15] ;
 wire \fpga_top.interrupter.g_interrupt_dly ;
 wire \fpga_top.interrupter.int0_1lat ;
 wire \fpga_top.interrupter.int0_2lat ;
 wire \fpga_top.interrupter.int0_3lat ;
 wire \fpga_top.interrupter.int_enable_int0 ;
 wire \fpga_top.interrupter.int_enable_rx ;
 wire \fpga_top.interrupter.int_status_int0 ;
 wire \fpga_top.interrupter.int_status_rx ;
 wire \fpga_top.interrupter.re_int_dly[0] ;
 wire \fpga_top.interrupter.re_int_dly[1] ;
 wire \fpga_top.interrupter.re_int_enable ;
 wire \fpga_top.interrupter.re_int_status ;
 wire \fpga_top.io_frc.frc_cmp_val[0] ;
 wire \fpga_top.io_frc.frc_cmp_val[10] ;
 wire \fpga_top.io_frc.frc_cmp_val[11] ;
 wire \fpga_top.io_frc.frc_cmp_val[12] ;
 wire \fpga_top.io_frc.frc_cmp_val[13] ;
 wire \fpga_top.io_frc.frc_cmp_val[14] ;
 wire \fpga_top.io_frc.frc_cmp_val[15] ;
 wire \fpga_top.io_frc.frc_cmp_val[16] ;
 wire \fpga_top.io_frc.frc_cmp_val[17] ;
 wire \fpga_top.io_frc.frc_cmp_val[18] ;
 wire \fpga_top.io_frc.frc_cmp_val[19] ;
 wire \fpga_top.io_frc.frc_cmp_val[1] ;
 wire \fpga_top.io_frc.frc_cmp_val[20] ;
 wire \fpga_top.io_frc.frc_cmp_val[21] ;
 wire \fpga_top.io_frc.frc_cmp_val[22] ;
 wire \fpga_top.io_frc.frc_cmp_val[23] ;
 wire \fpga_top.io_frc.frc_cmp_val[24] ;
 wire \fpga_top.io_frc.frc_cmp_val[25] ;
 wire \fpga_top.io_frc.frc_cmp_val[26] ;
 wire \fpga_top.io_frc.frc_cmp_val[27] ;
 wire \fpga_top.io_frc.frc_cmp_val[28] ;
 wire \fpga_top.io_frc.frc_cmp_val[29] ;
 wire \fpga_top.io_frc.frc_cmp_val[2] ;
 wire \fpga_top.io_frc.frc_cmp_val[30] ;
 wire \fpga_top.io_frc.frc_cmp_val[31] ;
 wire \fpga_top.io_frc.frc_cmp_val[32] ;
 wire \fpga_top.io_frc.frc_cmp_val[33] ;
 wire \fpga_top.io_frc.frc_cmp_val[34] ;
 wire \fpga_top.io_frc.frc_cmp_val[35] ;
 wire \fpga_top.io_frc.frc_cmp_val[36] ;
 wire \fpga_top.io_frc.frc_cmp_val[37] ;
 wire \fpga_top.io_frc.frc_cmp_val[38] ;
 wire \fpga_top.io_frc.frc_cmp_val[39] ;
 wire \fpga_top.io_frc.frc_cmp_val[3] ;
 wire \fpga_top.io_frc.frc_cmp_val[40] ;
 wire \fpga_top.io_frc.frc_cmp_val[41] ;
 wire \fpga_top.io_frc.frc_cmp_val[42] ;
 wire \fpga_top.io_frc.frc_cmp_val[43] ;
 wire \fpga_top.io_frc.frc_cmp_val[44] ;
 wire \fpga_top.io_frc.frc_cmp_val[45] ;
 wire \fpga_top.io_frc.frc_cmp_val[46] ;
 wire \fpga_top.io_frc.frc_cmp_val[47] ;
 wire \fpga_top.io_frc.frc_cmp_val[48] ;
 wire \fpga_top.io_frc.frc_cmp_val[49] ;
 wire \fpga_top.io_frc.frc_cmp_val[4] ;
 wire \fpga_top.io_frc.frc_cmp_val[50] ;
 wire \fpga_top.io_frc.frc_cmp_val[51] ;
 wire \fpga_top.io_frc.frc_cmp_val[52] ;
 wire \fpga_top.io_frc.frc_cmp_val[53] ;
 wire \fpga_top.io_frc.frc_cmp_val[54] ;
 wire \fpga_top.io_frc.frc_cmp_val[55] ;
 wire \fpga_top.io_frc.frc_cmp_val[56] ;
 wire \fpga_top.io_frc.frc_cmp_val[57] ;
 wire \fpga_top.io_frc.frc_cmp_val[58] ;
 wire \fpga_top.io_frc.frc_cmp_val[59] ;
 wire \fpga_top.io_frc.frc_cmp_val[5] ;
 wire \fpga_top.io_frc.frc_cmp_val[60] ;
 wire \fpga_top.io_frc.frc_cmp_val[61] ;
 wire \fpga_top.io_frc.frc_cmp_val[62] ;
 wire \fpga_top.io_frc.frc_cmp_val[63] ;
 wire \fpga_top.io_frc.frc_cmp_val[6] ;
 wire \fpga_top.io_frc.frc_cmp_val[7] ;
 wire \fpga_top.io_frc.frc_cmp_val[8] ;
 wire \fpga_top.io_frc.frc_cmp_val[9] ;
 wire \fpga_top.io_frc.frc_cntr_val[0] ;
 wire \fpga_top.io_frc.frc_cntr_val[10] ;
 wire \fpga_top.io_frc.frc_cntr_val[11] ;
 wire \fpga_top.io_frc.frc_cntr_val[12] ;
 wire \fpga_top.io_frc.frc_cntr_val[13] ;
 wire \fpga_top.io_frc.frc_cntr_val[14] ;
 wire \fpga_top.io_frc.frc_cntr_val[15] ;
 wire \fpga_top.io_frc.frc_cntr_val[16] ;
 wire \fpga_top.io_frc.frc_cntr_val[17] ;
 wire \fpga_top.io_frc.frc_cntr_val[18] ;
 wire \fpga_top.io_frc.frc_cntr_val[19] ;
 wire \fpga_top.io_frc.frc_cntr_val[1] ;
 wire \fpga_top.io_frc.frc_cntr_val[20] ;
 wire \fpga_top.io_frc.frc_cntr_val[21] ;
 wire \fpga_top.io_frc.frc_cntr_val[22] ;
 wire \fpga_top.io_frc.frc_cntr_val[23] ;
 wire \fpga_top.io_frc.frc_cntr_val[24] ;
 wire \fpga_top.io_frc.frc_cntr_val[25] ;
 wire \fpga_top.io_frc.frc_cntr_val[26] ;
 wire \fpga_top.io_frc.frc_cntr_val[27] ;
 wire \fpga_top.io_frc.frc_cntr_val[28] ;
 wire \fpga_top.io_frc.frc_cntr_val[29] ;
 wire \fpga_top.io_frc.frc_cntr_val[2] ;
 wire \fpga_top.io_frc.frc_cntr_val[30] ;
 wire \fpga_top.io_frc.frc_cntr_val[31] ;
 wire \fpga_top.io_frc.frc_cntr_val[32] ;
 wire \fpga_top.io_frc.frc_cntr_val[33] ;
 wire \fpga_top.io_frc.frc_cntr_val[34] ;
 wire \fpga_top.io_frc.frc_cntr_val[35] ;
 wire \fpga_top.io_frc.frc_cntr_val[36] ;
 wire \fpga_top.io_frc.frc_cntr_val[37] ;
 wire \fpga_top.io_frc.frc_cntr_val[38] ;
 wire \fpga_top.io_frc.frc_cntr_val[39] ;
 wire \fpga_top.io_frc.frc_cntr_val[3] ;
 wire \fpga_top.io_frc.frc_cntr_val[40] ;
 wire \fpga_top.io_frc.frc_cntr_val[41] ;
 wire \fpga_top.io_frc.frc_cntr_val[42] ;
 wire \fpga_top.io_frc.frc_cntr_val[43] ;
 wire \fpga_top.io_frc.frc_cntr_val[44] ;
 wire \fpga_top.io_frc.frc_cntr_val[45] ;
 wire \fpga_top.io_frc.frc_cntr_val[46] ;
 wire \fpga_top.io_frc.frc_cntr_val[47] ;
 wire \fpga_top.io_frc.frc_cntr_val[48] ;
 wire \fpga_top.io_frc.frc_cntr_val[49] ;
 wire \fpga_top.io_frc.frc_cntr_val[4] ;
 wire \fpga_top.io_frc.frc_cntr_val[50] ;
 wire \fpga_top.io_frc.frc_cntr_val[51] ;
 wire \fpga_top.io_frc.frc_cntr_val[52] ;
 wire \fpga_top.io_frc.frc_cntr_val[53] ;
 wire \fpga_top.io_frc.frc_cntr_val[54] ;
 wire \fpga_top.io_frc.frc_cntr_val[55] ;
 wire \fpga_top.io_frc.frc_cntr_val[56] ;
 wire \fpga_top.io_frc.frc_cntr_val[57] ;
 wire \fpga_top.io_frc.frc_cntr_val[58] ;
 wire \fpga_top.io_frc.frc_cntr_val[59] ;
 wire \fpga_top.io_frc.frc_cntr_val[5] ;
 wire \fpga_top.io_frc.frc_cntr_val[60] ;
 wire \fpga_top.io_frc.frc_cntr_val[61] ;
 wire \fpga_top.io_frc.frc_cntr_val[62] ;
 wire \fpga_top.io_frc.frc_cntr_val[63] ;
 wire \fpga_top.io_frc.frc_cntr_val[6] ;
 wire \fpga_top.io_frc.frc_cntr_val[7] ;
 wire \fpga_top.io_frc.frc_cntr_val[8] ;
 wire \fpga_top.io_frc.frc_cntr_val[9] ;
 wire \fpga_top.io_frc.frc_cntr_val_rst_lat ;
 wire \fpga_top.io_frc.frc_cntr_val_rst_pre ;
 wire \fpga_top.io_frc.frc_cntrl_val ;
 wire \fpga_top.io_frc.re_frc_cmphi ;
 wire \fpga_top.io_frc.re_frc_cmplo ;
 wire \fpga_top.io_frc.re_frc_cntrl ;
 wire \fpga_top.io_frc.re_frc_dly[0] ;
 wire \fpga_top.io_frc.re_frc_dly[1] ;
 wire \fpga_top.io_frc.re_frc_dly[2] ;
 wire \fpga_top.io_frc.re_frc_dly[3] ;
 wire \fpga_top.io_frc.re_frc_dly[4] ;
 wire \fpga_top.io_frc.re_frc_valhi ;
 wire \fpga_top.io_frc.re_frc_vallo ;
 wire \fpga_top.io_led.dbg_smpl_trgsig ;
 wire \fpga_top.io_led.gpi_init_lat1[0] ;
 wire \fpga_top.io_led.gpi_init_lat1[1] ;
 wire \fpga_top.io_led.gpi_init_lat1[2] ;
 wire \fpga_top.io_led.gpi_init_lat1[3] ;
 wire \fpga_top.io_led.gpi_init_lat1[4] ;
 wire \fpga_top.io_led.gpi_init_lat1[5] ;
 wire \fpga_top.io_led.gpi_init_lat2[0] ;
 wire \fpga_top.io_led.gpi_init_lat2[1] ;
 wire \fpga_top.io_led.gpi_init_lat2[2] ;
 wire \fpga_top.io_led.gpi_init_lat2[3] ;
 wire \fpga_top.io_led.gpi_init_lat2[4] ;
 wire \fpga_top.io_led.gpi_init_lat2[5] ;
 wire \fpga_top.io_led.gpio_in_lat1[0] ;
 wire \fpga_top.io_led.gpio_in_lat1[1] ;
 wire \fpga_top.io_led.gpio_in_lat1[2] ;
 wire \fpga_top.io_led.gpio_in_lat1[3] ;
 wire \fpga_top.io_led.gpio_in_lat2[0] ;
 wire \fpga_top.io_led.gpio_in_lat2[1] ;
 wire \fpga_top.io_led.gpio_in_lat2[2] ;
 wire \fpga_top.io_led.gpio_in_lat2[3] ;
 wire \fpga_top.io_led.led_value[0] ;
 wire \fpga_top.io_led.led_value[1] ;
 wire \fpga_top.io_led.led_value[2] ;
 wire \fpga_top.io_led.re_gpi_value ;
 wire \fpga_top.io_led.re_gpio_en_value ;
 wire \fpga_top.io_led.re_gpio_in_value ;
 wire \fpga_top.io_led.re_gpio_out_value ;
 wire \fpga_top.io_led.re_gpio_value_dly[0] ;
 wire \fpga_top.io_led.re_gpio_value_dly[1] ;
 wire \fpga_top.io_led.re_gpio_value_dly[2] ;
 wire \fpga_top.io_led.re_gpio_value_dly[3] ;
 wire \fpga_top.io_led.re_led_value ;
 wire \fpga_top.io_led.re_led_value_dly ;
 wire \fpga_top.io_spi_lite.bit_sel_org[0] ;
 wire \fpga_top.io_spi_lite.bit_sel_org[1] ;
 wire \fpga_top.io_spi_lite.bit_sel_org[2] ;
 wire \fpga_top.io_spi_lite.cs_all_status ;
 wire \fpga_top.io_spi_lite.miso_bit_cntr[0] ;
 wire \fpga_top.io_spi_lite.miso_bit_cntr[1] ;
 wire \fpga_top.io_spi_lite.miso_bit_cntr[2] ;
 wire \fpga_top.io_spi_lite.miso_byte_org[0] ;
 wire \fpga_top.io_spi_lite.miso_byte_org[1] ;
 wire \fpga_top.io_spi_lite.miso_byte_org[2] ;
 wire \fpga_top.io_spi_lite.miso_byte_org[3] ;
 wire \fpga_top.io_spi_lite.miso_byte_org[4] ;
 wire \fpga_top.io_spi_lite.miso_byte_org[5] ;
 wire \fpga_top.io_spi_lite.miso_byte_org[6] ;
 wire \fpga_top.io_spi_lite.miso_byte_org[7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.radr[0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.radr[1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.radr[2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.radr_early[0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.radr_early[1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.radr_early[2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.rnext ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][3] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][4] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][5] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][6] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][3] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][4] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][5] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][6] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][3] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][4] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][5] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][6] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][3] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][4] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][5] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][6] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][3] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][4] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][5] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][6] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][3] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][4] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][5] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][6] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][3] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][4] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][5] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][6] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][3] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][4] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][5] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][6] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][7] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[0] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[2] ;
 wire \fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wen ;
 wire \fpga_top.io_spi_lite.miso_lat[2] ;
 wire \fpga_top.io_spi_lite.miso_lat[3] ;
 wire \fpga_top.io_spi_lite.miso_lat[4] ;
 wire \fpga_top.io_spi_lite.miso_lat[5] ;
 wire \fpga_top.io_spi_lite.miso_lat[6] ;
 wire \fpga_top.io_spi_lite.miso_lat[7] ;
 wire \fpga_top.io_spi_lite.miso_read_next_byte ;
 wire \fpga_top.io_spi_lite.mosi_fifo.radr[0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.radr[1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.radr[2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.radr_early[0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.radr_early[1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.radr_early[2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][3] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][4] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][5] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][6] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][7] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][3] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][4] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][5] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][6] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][7] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][3] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][4] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][5] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][6] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][7] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][3] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][4] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][5] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][6] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][7] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][3] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][4] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][5] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][6] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][7] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][3] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][4] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][5] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][6] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][7] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][3] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][4] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][5] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][6] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][7] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][2] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][3] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][4] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][5] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][6] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][7] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[0] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[1] ;
 wire \fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[2] ;
 wire \fpga_top.io_spi_lite.mosi_pp_cntr[0] ;
 wire \fpga_top.io_spi_lite.mosi_pp_cntr[1] ;
 wire \fpga_top.io_spi_lite.mosi_pp_cntr[2] ;
 wire \fpga_top.io_spi_lite.mosi_pp_cntr[3] ;
 wire \fpga_top.io_spi_lite.org_mosi ;
 wire \fpga_top.io_spi_lite.org_sck ;
 wire \fpga_top.io_spi_lite.org_sck_dly ;
 wire \fpga_top.io_spi_lite.org_spi_sck ;
 wire \fpga_top.io_spi_lite.re_spi_miso ;
 wire \fpga_top.io_spi_lite.re_spi_mode ;
 wire \fpga_top.io_spi_lite.re_spi_mosi ;
 wire \fpga_top.io_spi_lite.re_spi_sdiv ;
 wire \fpga_top.io_spi_lite.re_spi_value_dly[0] ;
 wire \fpga_top.io_spi_lite.re_spi_value_dly[1] ;
 wire \fpga_top.io_spi_lite.re_spi_value_dly[2] ;
 wire \fpga_top.io_spi_lite.sck_div[0] ;
 wire \fpga_top.io_spi_lite.sck_div[1] ;
 wire \fpga_top.io_spi_lite.sck_div[2] ;
 wire \fpga_top.io_spi_lite.sck_div[3] ;
 wire \fpga_top.io_spi_lite.sck_div[4] ;
 wire \fpga_top.io_spi_lite.sck_div[5] ;
 wire \fpga_top.io_spi_lite.sck_div[6] ;
 wire \fpga_top.io_spi_lite.sck_div[7] ;
 wire \fpga_top.io_spi_lite.sck_div[8] ;
 wire \fpga_top.io_spi_lite.sck_div[9] ;
 wire \fpga_top.io_spi_lite.sel_cs[1] ;
 wire \fpga_top.io_spi_lite.sel_cs[2] ;
 wire \fpga_top.io_spi_lite.sel_cs[3] ;
 wire \fpga_top.io_spi_lite.sel_cs[4] ;
 wire \fpga_top.io_spi_lite.sel_cs[5] ;
 wire \fpga_top.io_spi_lite.sel_cs[6] ;
 wire \fpga_top.io_spi_lite.sel_cs[7] ;
 wire \fpga_top.io_spi_lite.sel_mosi[1] ;
 wire \fpga_top.io_spi_lite.sel_mosi[2] ;
 wire \fpga_top.io_spi_lite.sel_mosi[3] ;
 wire \fpga_top.io_spi_lite.sel_mosi[4] ;
 wire \fpga_top.io_spi_lite.sel_mosi[5] ;
 wire \fpga_top.io_spi_lite.sel_mosi[6] ;
 wire \fpga_top.io_spi_lite.sel_mosi[7] ;
 wire \fpga_top.io_spi_lite.sel_sck[1] ;
 wire \fpga_top.io_spi_lite.sel_sck[2] ;
 wire \fpga_top.io_spi_lite.sel_sck[3] ;
 wire \fpga_top.io_spi_lite.sel_sck[4] ;
 wire \fpga_top.io_spi_lite.sel_sck[5] ;
 wire \fpga_top.io_spi_lite.sel_sck[6] ;
 wire \fpga_top.io_spi_lite.sel_sck[7] ;
 wire \fpga_top.io_spi_lite.spi_mode[0] ;
 wire \fpga_top.io_spi_lite.spi_mode[10] ;
 wire \fpga_top.io_spi_lite.spi_mode[11] ;
 wire \fpga_top.io_spi_lite.spi_mode[12] ;
 wire \fpga_top.io_spi_lite.spi_mode[1] ;
 wire \fpga_top.io_spi_lite.spi_mode[2] ;
 wire \fpga_top.io_spi_lite.spi_mode[4] ;
 wire \fpga_top.io_spi_lite.spi_mode[5] ;
 wire \fpga_top.io_spi_lite.spi_mode[6] ;
 wire \fpga_top.io_spi_lite.spi_mode[7] ;
 wire \fpga_top.io_spi_lite.spi_mode[8] ;
 wire \fpga_top.io_spi_lite.spi_mode[9] ;
 wire \fpga_top.io_spi_lite.spi_mosi ;
 wire \fpga_top.io_spi_lite.spi_mosi_pre ;
 wire \fpga_top.io_spi_lite.spi_sck_div[0] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[1] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[2] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[3] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[4] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[5] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[6] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[7] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[8] ;
 wire \fpga_top.io_spi_lite.spi_sck_div[9] ;
 wire \fpga_top.io_spi_lite.spi_state[0] ;
 wire \fpga_top.io_spi_lite.spi_state[1] ;
 wire \fpga_top.io_uart_out.re_uart_char ;
 wire \fpga_top.io_uart_out.re_uart_full ;
 wire \fpga_top.io_uart_out.re_uart_rdflg_dly[0] ;
 wire \fpga_top.io_uart_out.re_uart_rdflg_dly[1] ;
 wire \fpga_top.io_uart_out.re_uart_rdflg_dly[2] ;
 wire \fpga_top.io_uart_out.re_uart_rdflg_dly[3] ;
 wire \fpga_top.io_uart_out.re_uart_rdflg_dly[4] ;
 wire \fpga_top.io_uart_out.re_uart_rxch ;
 wire \fpga_top.io_uart_out.re_uart_rxec ;
 wire \fpga_top.io_uart_out.re_uart_term ;
 wire \fpga_top.io_uart_out.rout[0] ;
 wire \fpga_top.io_uart_out.rout[1] ;
 wire \fpga_top.io_uart_out.rout[2] ;
 wire \fpga_top.io_uart_out.rout[3] ;
 wire \fpga_top.io_uart_out.rout[4] ;
 wire \fpga_top.io_uart_out.rout[5] ;
 wire \fpga_top.io_uart_out.rout[6] ;
 wire \fpga_top.io_uart_out.rout[7] ;
 wire \fpga_top.io_uart_out.rout_en ;
 wire \fpga_top.io_uart_out.rx_data_latch[0] ;
 wire \fpga_top.io_uart_out.rx_data_latch[1] ;
 wire \fpga_top.io_uart_out.rx_data_latch[2] ;
 wire \fpga_top.io_uart_out.rx_data_latch[3] ;
 wire \fpga_top.io_uart_out.rx_data_latch[4] ;
 wire \fpga_top.io_uart_out.rx_data_latch[5] ;
 wire \fpga_top.io_uart_out.rx_data_latch[6] ;
 wire \fpga_top.io_uart_out.rx_data_latch[7] ;
 wire \fpga_top.io_uart_out.rx_disable_echoback_value ;
 wire \fpga_top.io_uart_out.rx_first_read ;
 wire \fpga_top.io_uart_out.rx_write_error ;
 wire \fpga_top.io_uart_out.uart_io_char[0] ;
 wire \fpga_top.io_uart_out.uart_io_char[1] ;
 wire \fpga_top.io_uart_out.uart_io_char[2] ;
 wire \fpga_top.io_uart_out.uart_io_char[3] ;
 wire \fpga_top.io_uart_out.uart_io_char[4] ;
 wire \fpga_top.io_uart_out.uart_io_char[5] ;
 wire \fpga_top.io_uart_out.uart_io_char[6] ;
 wire \fpga_top.io_uart_out.uart_io_char[7] ;
 wire \fpga_top.io_uart_out.uart_io_we ;
 wire \fpga_top.io_uart_out.uart_term[0] ;
 wire \fpga_top.io_uart_out.uart_term[10] ;
 wire \fpga_top.io_uart_out.uart_term[11] ;
 wire \fpga_top.io_uart_out.uart_term[12] ;
 wire \fpga_top.io_uart_out.uart_term[13] ;
 wire \fpga_top.io_uart_out.uart_term[14] ;
 wire \fpga_top.io_uart_out.uart_term[15] ;
 wire \fpga_top.io_uart_out.uart_term[1] ;
 wire \fpga_top.io_uart_out.uart_term[2] ;
 wire \fpga_top.io_uart_out.uart_term[3] ;
 wire \fpga_top.io_uart_out.uart_term[4] ;
 wire \fpga_top.io_uart_out.uart_term[5] ;
 wire \fpga_top.io_uart_out.uart_term[6] ;
 wire \fpga_top.io_uart_out.uart_term[7] ;
 wire \fpga_top.io_uart_out.uart_term[8] ;
 wire \fpga_top.io_uart_out.uart_term[9] ;
 wire \fpga_top.qspi_if.adr_ofs[0] ;
 wire \fpga_top.qspi_if.adr_ofs[1] ;
 wire \fpga_top.qspi_if.adr_ofs[2] ;
 wire \fpga_top.qspi_if.adr_rw[0] ;
 wire \fpga_top.qspi_if.adr_rw[10] ;
 wire \fpga_top.qspi_if.adr_rw[11] ;
 wire \fpga_top.qspi_if.adr_rw[12] ;
 wire \fpga_top.qspi_if.adr_rw[13] ;
 wire \fpga_top.qspi_if.adr_rw[14] ;
 wire \fpga_top.qspi_if.adr_rw[15] ;
 wire \fpga_top.qspi_if.adr_rw[16] ;
 wire \fpga_top.qspi_if.adr_rw[17] ;
 wire \fpga_top.qspi_if.adr_rw[18] ;
 wire \fpga_top.qspi_if.adr_rw[19] ;
 wire \fpga_top.qspi_if.adr_rw[1] ;
 wire \fpga_top.qspi_if.adr_rw[20] ;
 wire \fpga_top.qspi_if.adr_rw[21] ;
 wire \fpga_top.qspi_if.adr_rw[22] ;
 wire \fpga_top.qspi_if.adr_rw[23] ;
 wire \fpga_top.qspi_if.adr_rw[2] ;
 wire \fpga_top.qspi_if.adr_rw[3] ;
 wire \fpga_top.qspi_if.adr_rw[4] ;
 wire \fpga_top.qspi_if.adr_rw[5] ;
 wire \fpga_top.qspi_if.adr_rw[6] ;
 wire \fpga_top.qspi_if.adr_rw[7] ;
 wire \fpga_top.qspi_if.adr_rw[8] ;
 wire \fpga_top.qspi_if.adr_rw[9] ;
 wire \fpga_top.qspi_if.cmd_ofs[0] ;
 wire \fpga_top.qspi_if.cmd_ofs[1] ;
 wire \fpga_top.qspi_if.cmd_ofs[2] ;
 wire \fpga_top.qspi_if.dbg_2div_cec_lat ;
 wire \fpga_top.qspi_if.dbg_2div_cec_pre ;
 wire \fpga_top.qspi_if.dbg_2div_cew_lat ;
 wire \fpga_top.qspi_if.dbg_2div_cew_pre ;
 wire \fpga_top.qspi_if.dbg_2div_read_half_end ;
 wire \fpga_top.qspi_if.dbg_2div_trt ;
 wire \fpga_top.qspi_if.dbg_2div_wirte_half_end ;
 wire \fpga_top.qspi_if.dbg_reg_2div_cec_read ;
 wire \fpga_top.qspi_if.dbg_reg_2div_cec_write ;
 wire \fpga_top.qspi_if.inner_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/qspi_if.v:768$329.$result[0] ;
 wire \fpga_top.qspi_if.inner_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/qspi_if.v:768$329.$result[1] ;
 wire \fpga_top.qspi_if.inner_state[0] ;
 wire \fpga_top.qspi_if.inner_state[1] ;
 wire \fpga_top.qspi_if.qspi_state[10] ;
 wire \fpga_top.qspi_if.qspi_state[11] ;
 wire \fpga_top.qspi_if.qspi_state[1] ;
 wire \fpga_top.qspi_if.qspi_state[2] ;
 wire \fpga_top.qspi_if.qspi_state[3] ;
 wire \fpga_top.qspi_if.qspi_state[4] ;
 wire \fpga_top.qspi_if.qspi_state[6] ;
 wire \fpga_top.qspi_if.qspi_state[7] ;
 wire \fpga_top.qspi_if.qspi_state[8] ;
 wire \fpga_top.qspi_if.qspi_state[9] ;
 wire \fpga_top.qspi_if.rdcmd0[2] ;
 wire \fpga_top.qspi_if.rdcmd0[4] ;
 wire \fpga_top.qspi_if.rdcmd1[2] ;
 wire \fpga_top.qspi_if.rdcmd1[4] ;
 wire \fpga_top.qspi_if.rdcmd1[7] ;
 wire \fpga_top.qspi_if.rdedge[0] ;
 wire \fpga_top.qspi_if.rdedge[2] ;
 wire \fpga_top.qspi_if.rdwrch[0] ;
 wire \fpga_top.qspi_if.rdwrch[1] ;
 wire \fpga_top.qspi_if.rdwrch[2] ;
 wire \fpga_top.qspi_if.rdwrch[3] ;
 wire \fpga_top.qspi_if.rdwrch[4] ;
 wire \fpga_top.qspi_if.rdwrch[5] ;
 wire \fpga_top.qspi_if.re_qspi_latency0 ;
 wire \fpga_top.qspi_if.re_qspi_latency1 ;
 wire \fpga_top.qspi_if.re_qspi_latency2 ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[0] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[1] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[2] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[3] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[4] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[5] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[6] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[7] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[8] ;
 wire \fpga_top.qspi_if.re_qspi_latency_dly[9] ;
 wire \fpga_top.qspi_if.re_qspi_rdcmd0 ;
 wire \fpga_top.qspi_if.re_qspi_rdcmd1 ;
 wire \fpga_top.qspi_if.re_qspi_rdedge ;
 wire \fpga_top.qspi_if.re_qspi_rdwrch ;
 wire \fpga_top.qspi_if.re_qspi_sckdiv ;
 wire \fpga_top.qspi_if.re_qspi_wrcmd0 ;
 wire \fpga_top.qspi_if.re_qspi_wrcmd1 ;
 wire \fpga_top.qspi_if.read_cntr[0] ;
 wire \fpga_top.qspi_if.read_cntr[1] ;
 wire \fpga_top.qspi_if.read_cntr[2] ;
 wire \fpga_top.qspi_if.read_cntr[3] ;
 wire \fpga_top.qspi_if.read_latency_0[0] ;
 wire \fpga_top.qspi_if.read_latency_0[1] ;
 wire \fpga_top.qspi_if.read_latency_0[2] ;
 wire \fpga_top.qspi_if.read_latency_0[3] ;
 wire \fpga_top.qspi_if.read_latency_1[0] ;
 wire \fpga_top.qspi_if.read_latency_1[1] ;
 wire \fpga_top.qspi_if.read_latency_1[2] ;
 wire \fpga_top.qspi_if.read_latency_1[3] ;
 wire \fpga_top.qspi_if.read_latency_2[0] ;
 wire \fpga_top.qspi_if.read_latency_2[1] ;
 wire \fpga_top.qspi_if.read_latency_2[2] ;
 wire \fpga_top.qspi_if.read_latency_2[3] ;
 wire \fpga_top.qspi_if.rst_cntr[0] ;
 wire \fpga_top.qspi_if.rst_cntr[1] ;
 wire \fpga_top.qspi_if.rst_cntr[2] ;
 wire \fpga_top.qspi_if.rst_cntr[3] ;
 wire \fpga_top.qspi_if.rwait_cntr[0] ;
 wire \fpga_top.qspi_if.rwait_cntr[1] ;
 wire \fpga_top.qspi_if.rwait_cntr[2] ;
 wire \fpga_top.qspi_if.rwait_cntr[3] ;
 wire \fpga_top.qspi_if.sck ;
 wire \fpga_top.qspi_if.sck_cntr[0] ;
 wire \fpga_top.qspi_if.sck_cntr[1] ;
 wire \fpga_top.qspi_if.sck_cntr[2] ;
 wire \fpga_top.qspi_if.sck_cntr[3] ;
 wire \fpga_top.qspi_if.sck_cntr[4] ;
 wire \fpga_top.qspi_if.sck_cntr[5] ;
 wire \fpga_top.qspi_if.sck_cntr[6] ;
 wire \fpga_top.qspi_if.sck_cntr[7] ;
 wire \fpga_top.qspi_if.sck_cntr[8] ;
 wire \fpga_top.qspi_if.sck_cntr[9] ;
 wire \fpga_top.qspi_if.sck_div[1] ;
 wire \fpga_top.qspi_if.sck_div[2] ;
 wire \fpga_top.qspi_if.sck_div[3] ;
 wire \fpga_top.qspi_if.sck_div[4] ;
 wire \fpga_top.qspi_if.sck_div[5] ;
 wire \fpga_top.qspi_if.sck_div[6] ;
 wire \fpga_top.qspi_if.sck_div[7] ;
 wire \fpga_top.qspi_if.sck_div[8] ;
 wire \fpga_top.qspi_if.sck_div[9] ;
 wire \fpga_top.qspi_if.sio_en ;
 wire \fpga_top.qspi_if.sio_in_mt0[0] ;
 wire \fpga_top.qspi_if.sio_in_mt0[1] ;
 wire \fpga_top.qspi_if.sio_in_mt0[2] ;
 wire \fpga_top.qspi_if.sio_in_mt0[3] ;
 wire \fpga_top.qspi_if.sio_in_mt1[0] ;
 wire \fpga_top.qspi_if.sio_in_mt1[1] ;
 wire \fpga_top.qspi_if.sio_in_mt1[2] ;
 wire \fpga_top.qspi_if.sio_in_mt1[3] ;
 wire \fpga_top.qspi_if.sio_in_sync[0] ;
 wire \fpga_top.qspi_if.sio_in_sync[1] ;
 wire \fpga_top.qspi_if.sio_in_sync[2] ;
 wire \fpga_top.qspi_if.sio_in_sync[3] ;
 wire \fpga_top.qspi_if.sio_out_dly[0] ;
 wire \fpga_top.qspi_if.sio_out_dly[1] ;
 wire \fpga_top.qspi_if.sio_out_dly[2] ;
 wire \fpga_top.qspi_if.sio_out_dly[3] ;
 wire \fpga_top.qspi_if.sio_out_enbl_dly ;
 wire \fpga_top.qspi_if.sio_out_enbl_pre ;
 wire \fpga_top.qspi_if.sio_out_pre[0] ;
 wire \fpga_top.qspi_if.sio_out_pre[1] ;
 wire \fpga_top.qspi_if.sio_out_pre[2] ;
 wire \fpga_top.qspi_if.sio_out_pre[3] ;
 wire \fpga_top.qspi_if.wdata[0] ;
 wire \fpga_top.qspi_if.wdata[10] ;
 wire \fpga_top.qspi_if.wdata[11] ;
 wire \fpga_top.qspi_if.wdata[12] ;
 wire \fpga_top.qspi_if.wdata[13] ;
 wire \fpga_top.qspi_if.wdata[14] ;
 wire \fpga_top.qspi_if.wdata[15] ;
 wire \fpga_top.qspi_if.wdata[16] ;
 wire \fpga_top.qspi_if.wdata[17] ;
 wire \fpga_top.qspi_if.wdata[18] ;
 wire \fpga_top.qspi_if.wdata[19] ;
 wire \fpga_top.qspi_if.wdata[1] ;
 wire \fpga_top.qspi_if.wdata[20] ;
 wire \fpga_top.qspi_if.wdata[21] ;
 wire \fpga_top.qspi_if.wdata[22] ;
 wire \fpga_top.qspi_if.wdata[23] ;
 wire \fpga_top.qspi_if.wdata[24] ;
 wire \fpga_top.qspi_if.wdata[25] ;
 wire \fpga_top.qspi_if.wdata[26] ;
 wire \fpga_top.qspi_if.wdata[27] ;
 wire \fpga_top.qspi_if.wdata[28] ;
 wire \fpga_top.qspi_if.wdata[29] ;
 wire \fpga_top.qspi_if.wdata[2] ;
 wire \fpga_top.qspi_if.wdata[30] ;
 wire \fpga_top.qspi_if.wdata[31] ;
 wire \fpga_top.qspi_if.wdata[3] ;
 wire \fpga_top.qspi_if.wdata[4] ;
 wire \fpga_top.qspi_if.wdata[5] ;
 wire \fpga_top.qspi_if.wdata[6] ;
 wire \fpga_top.qspi_if.wdata[7] ;
 wire \fpga_top.qspi_if.wdata[8] ;
 wire \fpga_top.qspi_if.wdata[9] ;
 wire \fpga_top.qspi_if.wdata_ofs[0] ;
 wire \fpga_top.qspi_if.wdata_ofs[1] ;
 wire \fpga_top.qspi_if.wdata_ofs[2] ;
 wire \fpga_top.qspi_if.word_adr[24] ;
 wire \fpga_top.qspi_if.word_adr[25] ;
 wire \fpga_top.qspi_if.word_data[0] ;
 wire \fpga_top.qspi_if.word_data[10] ;
 wire \fpga_top.qspi_if.word_data[11] ;
 wire \fpga_top.qspi_if.word_data[12] ;
 wire \fpga_top.qspi_if.word_data[13] ;
 wire \fpga_top.qspi_if.word_data[14] ;
 wire \fpga_top.qspi_if.word_data[15] ;
 wire \fpga_top.qspi_if.word_data[16] ;
 wire \fpga_top.qspi_if.word_data[17] ;
 wire \fpga_top.qspi_if.word_data[18] ;
 wire \fpga_top.qspi_if.word_data[19] ;
 wire \fpga_top.qspi_if.word_data[1] ;
 wire \fpga_top.qspi_if.word_data[20] ;
 wire \fpga_top.qspi_if.word_data[21] ;
 wire \fpga_top.qspi_if.word_data[22] ;
 wire \fpga_top.qspi_if.word_data[23] ;
 wire \fpga_top.qspi_if.word_data[24] ;
 wire \fpga_top.qspi_if.word_data[25] ;
 wire \fpga_top.qspi_if.word_data[26] ;
 wire \fpga_top.qspi_if.word_data[27] ;
 wire \fpga_top.qspi_if.word_data[28] ;
 wire \fpga_top.qspi_if.word_data[29] ;
 wire \fpga_top.qspi_if.word_data[2] ;
 wire \fpga_top.qspi_if.word_data[30] ;
 wire \fpga_top.qspi_if.word_data[31] ;
 wire \fpga_top.qspi_if.word_data[3] ;
 wire \fpga_top.qspi_if.word_data[4] ;
 wire \fpga_top.qspi_if.word_data[5] ;
 wire \fpga_top.qspi_if.word_data[6] ;
 wire \fpga_top.qspi_if.word_data[7] ;
 wire \fpga_top.qspi_if.word_data[8] ;
 wire \fpga_top.qspi_if.word_data[9] ;
 wire \fpga_top.qspi_if.word_hw ;
 wire \fpga_top.qspi_if.word_w ;
 wire \fpga_top.qspi_if.wrcmd0[0] ;
 wire \fpga_top.qspi_if.wrcmd0[1] ;
 wire \fpga_top.qspi_if.wrcmd0[2] ;
 wire \fpga_top.qspi_if.wrcmd0[6] ;
 wire \fpga_top.qspi_if.wrcmd0[7] ;
 wire \fpga_top.qspi_if.wrcmd1[0] ;
 wire \fpga_top.qspi_if.wrcmd1[1] ;
 wire \fpga_top.qspi_if.wrcmd1[2] ;
 wire \fpga_top.qspi_if.wrcmd1[6] ;
 wire \fpga_top.qspi_if.wrcmd1[7] ;
 wire \fpga_top.qspi_if.wredge[0] ;
 wire \fpga_top.qspi_if.wredge[2] ;
 wire \fpga_top.tx ;
 wire \fpga_top.uart_top.rx_fifo_dvalid ;
 wire \fpga_top.uart_top.rx_fifo_rcntr[0] ;
 wire \fpga_top.uart_top.rx_fifo_rcntr[1] ;
 wire \fpga_top.uart_top.rx_fifo_rcntr[2] ;
 wire \fpga_top.uart_top.trush_running ;
 wire \fpga_top.uart_top.uart_if.byte_data[0] ;
 wire \fpga_top.uart_top.uart_if.byte_data[1] ;
 wire \fpga_top.uart_top.uart_if.byte_data[2] ;
 wire \fpga_top.uart_top.uart_if.byte_data[3] ;
 wire \fpga_top.uart_top.uart_if.byte_data[4] ;
 wire \fpga_top.uart_top.uart_if.byte_data[5] ;
 wire \fpga_top.uart_top.uart_if.byte_data[6] ;
 wire \fpga_top.uart_top.uart_if.byte_data[7] ;
 wire \fpga_top.uart_top.uart_if.next_rx_state[0] ;
 wire \fpga_top.uart_top.uart_if.next_rx_state[1] ;
 wire \fpga_top.uart_top.uart_if.next_rx_state[2] ;
 wire \fpga_top.uart_top.uart_if.next_rx_state[3] ;
 wire \fpga_top.uart_top.uart_if.next_tx_state[0] ;
 wire \fpga_top.uart_top.uart_if.next_tx_state[1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.radr[0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.radr[1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.radr[2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[0][0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[0][1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[0][2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[0][3] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[0][4] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[0][5] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[0][6] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[0][7] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[1][0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[1][1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[1][2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[1][3] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[1][4] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[1][5] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[1][6] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[1][7] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[2][0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[2][1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[2][2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[2][3] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[2][4] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[2][5] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[2][6] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[2][7] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[3][0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[3][1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[3][2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[3][3] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[3][4] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[3][5] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[3][6] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[3][7] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[4][0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[4][1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[4][2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[4][3] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[4][4] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[4][5] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[4][6] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[4][7] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[5][0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[5][1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[5][2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[5][3] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[5][4] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[5][5] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[5][6] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[5][7] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[6][0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[6][1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[6][2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[6][3] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[6][4] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[6][5] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[6][6] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[6][7] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[7][0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[7][1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[7][2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[7][3] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[7][4] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[7][5] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[7][6] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram[7][7] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo_dcntr[0] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo_dcntr[1] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo_dcntr[2] ;
 wire \fpga_top.uart_top.uart_if.rx_fifo_dcntr[3] ;
 wire \fpga_top.uart_top.uart_if.rx_state[0] ;
 wire \fpga_top.uart_top.uart_if.rx_state[1] ;
 wire \fpga_top.uart_top.uart_if.rx_state[2] ;
 wire \fpga_top.uart_top.uart_if.rx_state[3] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[0] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[10] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[11] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[12] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[13] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[14] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[15] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[1] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[2] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[3] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[4] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[5] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[6] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[7] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[8] ;
 wire \fpga_top.uart_top.uart_if.sample_cntr[9] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[0] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[10] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[11] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[12] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[13] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[14] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[15] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[1] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[2] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[3] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[4] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[5] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[6] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[7] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[8] ;
 wire \fpga_top.uart_top.uart_if.tx_cycle_cntr[9] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[0][0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[0][1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[0][2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[0][3] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[0][4] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[0][5] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[0][6] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[0][7] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[1][0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[1][1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[1][2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[1][3] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[1][4] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[1][5] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[1][6] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[1][7] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[2][0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[2][1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[2][2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[2][3] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[2][4] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[2][5] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[2][6] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[2][7] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[3][0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[3][1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[3][2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[3][3] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[3][4] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[3][5] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[3][6] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[3][7] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[4][0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[4][1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[4][2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[4][3] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[4][4] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[4][5] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[4][6] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[4][7] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[5][0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[5][1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[5][2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[5][3] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[5][4] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[5][5] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[5][6] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[5][7] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[6][0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[6][1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[6][2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[6][3] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[6][4] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[6][5] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[6][6] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[6][7] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[7][0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[7][1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[7][2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[7][3] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[7][4] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[7][5] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[7][6] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram[7][7] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram_radr[0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram_radr[1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram_radr[2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo_dcntr[0] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo_dcntr[1] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo_dcntr[2] ;
 wire \fpga_top.uart_top.uart_if.tx_fifo_dcntr[3] ;
 wire \fpga_top.uart_top.uart_if.tx_out_cntr[0] ;
 wire \fpga_top.uart_top.uart_if.tx_out_cntr[1] ;
 wire \fpga_top.uart_top.uart_if.tx_out_cntr[2] ;
 wire \fpga_top.uart_top.uart_if.tx_out_cntr[3] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[1] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[2] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[3] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[4] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[5] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[6] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[7] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[8] ;
 wire \fpga_top.uart_top.uart_if.tx_out_data[9] ;
 wire \fpga_top.uart_top.uart_if.tx_state[0] ;
 wire \fpga_top.uart_top.uart_if.tx_state[1] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_adr[32] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[10] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[11] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[12] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[13] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[14] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[15] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[16] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[17] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[18] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[19] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[20] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[21] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[22] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[23] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[24] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[25] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[26] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[27] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[28] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[29] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[2] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[30] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[31] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[3] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[4] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[5] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[6] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[7] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[8] ;
 wire \fpga_top.uart_top.uart_logics.cmd_read_end[9] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[16] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[17] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[18] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[19] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[20] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[21] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[22] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[23] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[24] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[25] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[26] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[27] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[28] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[29] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[30] ;
 wire \fpga_top.uart_top.uart_logics.cmd_wadr_cntr[31] ;
 wire \fpga_top.uart_top.uart_logics.data_0[0] ;
 wire \fpga_top.uart_top.uart_logics.data_0[10] ;
 wire \fpga_top.uart_top.uart_logics.data_0[11] ;
 wire \fpga_top.uart_top.uart_logics.data_0[12] ;
 wire \fpga_top.uart_top.uart_logics.data_0[13] ;
 wire \fpga_top.uart_top.uart_logics.data_0[14] ;
 wire \fpga_top.uart_top.uart_logics.data_0[15] ;
 wire \fpga_top.uart_top.uart_logics.data_0[16] ;
 wire \fpga_top.uart_top.uart_logics.data_0[17] ;
 wire \fpga_top.uart_top.uart_logics.data_0[18] ;
 wire \fpga_top.uart_top.uart_logics.data_0[19] ;
 wire \fpga_top.uart_top.uart_logics.data_0[1] ;
 wire \fpga_top.uart_top.uart_logics.data_0[20] ;
 wire \fpga_top.uart_top.uart_logics.data_0[21] ;
 wire \fpga_top.uart_top.uart_logics.data_0[22] ;
 wire \fpga_top.uart_top.uart_logics.data_0[23] ;
 wire \fpga_top.uart_top.uart_logics.data_0[24] ;
 wire \fpga_top.uart_top.uart_logics.data_0[25] ;
 wire \fpga_top.uart_top.uart_logics.data_0[26] ;
 wire \fpga_top.uart_top.uart_logics.data_0[27] ;
 wire \fpga_top.uart_top.uart_logics.data_0[28] ;
 wire \fpga_top.uart_top.uart_logics.data_0[29] ;
 wire \fpga_top.uart_top.uart_logics.data_0[2] ;
 wire \fpga_top.uart_top.uart_logics.data_0[30] ;
 wire \fpga_top.uart_top.uart_logics.data_0[31] ;
 wire \fpga_top.uart_top.uart_logics.data_0[3] ;
 wire \fpga_top.uart_top.uart_logics.data_0[4] ;
 wire \fpga_top.uart_top.uart_logics.data_0[5] ;
 wire \fpga_top.uart_top.uart_logics.data_0[6] ;
 wire \fpga_top.uart_top.uart_logics.data_0[7] ;
 wire \fpga_top.uart_top.uart_logics.data_0[8] ;
 wire \fpga_top.uart_top.uart_logics.data_0[9] ;
 wire \fpga_top.uart_top.uart_logics.dma_io_data_en ;
 wire \fpga_top.uart_top.uart_logics.next_status_dump[0] ;
 wire \fpga_top.uart_top.uart_logics.next_status_dump[1] ;
 wire \fpga_top.uart_top.uart_logics.next_status_dump[2] ;
 wire \fpga_top.uart_top.uart_logics.radr_enable ;
 wire \fpga_top.uart_top.uart_logics.rdata_snd_wait ;
 wire \fpga_top.uart_top.uart_logics.rdata_snd_wait_dly ;
 wire \fpga_top.uart_top.uart_logics.status_dump[0] ;
 wire \fpga_top.uart_top.uart_logics.status_dump[1] ;
 wire \fpga_top.uart_top.uart_logics.status_dump[2] ;
 wire \fpga_top.uart_top.uart_logics.trash_cond_dly ;
 wire \fpga_top.uart_top.uart_logics.write_stat ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[10] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[11] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[12] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[13] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[14] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[15] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[16] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[17] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[18] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[19] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[20] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[21] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[22] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[23] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[24] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[25] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[26] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[27] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[28] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[29] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[2] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[30] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[31] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[3] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[4] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[5] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[6] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[7] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[8] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint[9] ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint_en ;
 wire \fpga_top.uart_top.uart_rec_char.bpoint_ld ;
 wire \fpga_top.uart_top.uart_rec_char.cmd_status[0] ;
 wire \fpga_top.uart_top.uart_rec_char.cmd_status[1] ;
 wire \fpga_top.uart_top.uart_rec_char.cmd_status[2] ;
 wire \fpga_top.uart_top.uart_rec_char.cmd_status[3] ;
 wire \fpga_top.uart_top.uart_rec_char.cmd_status[4] ;
 wire \fpga_top.uart_top.uart_rec_char.data_cntr[0] ;
 wire \fpga_top.uart_top.uart_rec_char.data_cntr[1] ;
 wire \fpga_top.uart_top.uart_rec_char.data_cntr[2] ;
 wire \fpga_top.uart_top.uart_rec_char.data_cntr[3] ;
 wire \fpga_top.uart_top.uart_rec_char.data_en ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[0] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[10] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[11] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[12] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[13] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[14] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[15] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[16] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[17] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[18] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[19] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[1] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[20] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[21] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[22] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[23] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[24] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[25] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[26] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[27] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[2] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[3] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[4] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[5] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[6] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[7] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[8] ;
 wire \fpga_top.uart_top.uart_rec_char.data_word[9] ;
 wire \fpga_top.uart_top.uart_rec_char.g_crlf ;
 wire \fpga_top.uart_top.uart_rec_char.g_crlf_dly ;
 wire \fpga_top.uart_top.uart_rec_char.g_crlf_dly2 ;
 wire \fpga_top.uart_top.uart_rec_char.next_cmd_status[0] ;
 wire \fpga_top.uart_top.uart_rec_char.next_cmd_status[1] ;
 wire \fpga_top.uart_top.uart_rec_char.next_cmd_status[2] ;
 wire \fpga_top.uart_top.uart_rec_char.next_cmd_status[3] ;
 wire \fpga_top.uart_top.uart_rec_char.next_cmd_status[4] ;
 wire \fpga_top.uart_top.uart_rec_char.pdata[0] ;
 wire \fpga_top.uart_top.uart_rec_char.pdata[1] ;
 wire \fpga_top.uart_top.uart_rec_char.pdata[2] ;
 wire \fpga_top.uart_top.uart_rec_char.pdata[3] ;
 wire \fpga_top.uart_top.uart_rec_char.pdata[4] ;
 wire \fpga_top.uart_top.uart_rec_char.pdata[5] ;
 wire \fpga_top.uart_top.uart_rec_char.pdata[6] ;
 wire \fpga_top.uart_top.uart_rec_char.pdata[7] ;
 wire \fpga_top.uart_top.uart_rec_char.word_valid ;
 wire \fpga_top.uart_top.uart_rec_char.word_valid_pre ;
 wire \fpga_top.uart_top.uart_send_char.send_cntr[0] ;
 wire \fpga_top.uart_top.uart_send_char.send_cntr[1] ;
 wire \fpga_top.uart_top.uart_send_char.send_cntr[2] ;
 wire \fpga_top.uart_top.uart_send_char.send_cntr[3] ;
 wire \fpga_top.uart_top.uart_send_char.send_cntr[4] ;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_leaf_327_clk;
 wire clknet_leaf_328_clk;
 wire clknet_leaf_329_clk;
 wire clknet_leaf_330_clk;
 wire clknet_leaf_331_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0_0_clk;
 wire clknet_5_1_0_clk;
 wire clknet_5_2_0_clk;
 wire clknet_5_3_0_clk;
 wire clknet_5_4_0_clk;
 wire clknet_5_5_0_clk;
 wire clknet_5_6_0_clk;
 wire clknet_5_7_0_clk;
 wire clknet_5_8_0_clk;
 wire clknet_5_9_0_clk;
 wire clknet_5_10_0_clk;
 wire clknet_5_11_0_clk;
 wire clknet_5_12_0_clk;
 wire clknet_5_13_0_clk;
 wire clknet_5_14_0_clk;
 wire clknet_5_15_0_clk;
 wire clknet_5_16_0_clk;
 wire clknet_5_17_0_clk;
 wire clknet_5_18_0_clk;
 wire clknet_5_19_0_clk;
 wire clknet_5_20_0_clk;
 wire clknet_5_21_0_clk;
 wire clknet_5_22_0_clk;
 wire clknet_5_23_0_clk;
 wire clknet_5_24_0_clk;
 wire clknet_5_25_0_clk;
 wire clknet_5_26_0_clk;
 wire clknet_5_27_0_clk;
 wire clknet_5_28_0_clk;
 wire clknet_5_29_0_clk;
 wire clknet_5_30_0_clk;
 wire clknet_5_31_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6203;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net6319;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6325;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;

 sg13g2_inv_1 _12296_ (.Y(_00141_),
    .A(net1));
 sg13g2_inv_1 _12297_ (.Y(_06497_),
    .A(_00114_));
 sg13g2_inv_2 _12298_ (.Y(_06498_),
    .A(_00111_));
 sg13g2_inv_1 _12299_ (.Y(_06499_),
    .A(_00108_));
 sg13g2_inv_2 _12300_ (.Y(_06500_),
    .A(_00090_));
 sg13g2_inv_2 _12301_ (.Y(_06501_),
    .A(net5424));
 sg13g2_inv_1 _12302_ (.Y(_06502_),
    .A(net3855));
 sg13g2_inv_1 _12303_ (.Y(_06503_),
    .A(net3386));
 sg13g2_inv_2 _12304_ (.Y(_06504_),
    .A(net5616));
 sg13g2_inv_4 _12305_ (.A(net5615),
    .Y(_06505_));
 sg13g2_inv_1 _12306_ (.Y(_06506_),
    .A(net3138));
 sg13g2_inv_4 _12307_ (.A(net6303),
    .Y(_06507_));
 sg13g2_inv_4 _12308_ (.A(net6449),
    .Y(_06508_));
 sg13g2_inv_2 _12309_ (.Y(_06509_),
    .A(\fpga_top.bus_gather.u_read_adr[9] ));
 sg13g2_inv_2 _12310_ (.Y(_06510_),
    .A(net1954));
 sg13g2_inv_2 _12311_ (.Y(_06511_),
    .A(net6364));
 sg13g2_inv_1 _12312_ (.Y(_06512_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[7] ));
 sg13g2_inv_2 _12313_ (.Y(_06513_),
    .A(net6149));
 sg13g2_inv_8 _12314_ (.Y(_06514_),
    .A(net6315));
 sg13g2_inv_2 _12315_ (.Y(_06515_),
    .A(net6255));
 sg13g2_inv_1 _12316_ (.Y(_06516_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[16] ));
 sg13g2_inv_1 _12317_ (.Y(_06517_),
    .A(net6231));
 sg13g2_inv_2 _12318_ (.Y(_06518_),
    .A(net6257));
 sg13g2_inv_1 _12319_ (.Y(_06519_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[13] ));
 sg13g2_inv_1 _12320_ (.Y(_06520_),
    .A(\fpga_top.bus_gather.u_read_adr[13] ));
 sg13g2_inv_1 _12321_ (.Y(_06521_),
    .A(net6301));
 sg13g2_inv_2 _12322_ (.Y(_06522_),
    .A(\fpga_top.bus_gather.u_read_adr[11] ));
 sg13g2_inv_2 _12323_ (.Y(_06523_),
    .A(net6341));
 sg13g2_inv_1 _12324_ (.Y(_06524_),
    .A(net3688));
 sg13g2_inv_1 _12325_ (.Y(_06525_),
    .A(net5614));
 sg13g2_inv_1 _12326_ (.Y(_06526_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[19] ));
 sg13g2_inv_2 _12327_ (.Y(_06527_),
    .A(net6264));
 sg13g2_inv_1 _12328_ (.Y(_06528_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[18] ));
 sg13g2_inv_2 _12329_ (.Y(_06529_),
    .A(net6289));
 sg13g2_inv_2 _12330_ (.Y(_06530_),
    .A(net6239));
 sg13g2_inv_2 _12331_ (.Y(_06531_),
    .A(net6319));
 sg13g2_inv_2 _12332_ (.Y(_06532_),
    .A(net3901));
 sg13g2_inv_1 _12333_ (.Y(_06533_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[22] ));
 sg13g2_inv_1 _12334_ (.Y(_06534_),
    .A(net6317));
 sg13g2_inv_1 _12335_ (.Y(_06535_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[29] ));
 sg13g2_inv_1 _12336_ (.Y(_06536_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[28] ));
 sg13g2_inv_1 _12337_ (.Y(_06537_),
    .A(net3833));
 sg13g2_inv_1 _12338_ (.Y(_06538_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[26] ));
 sg13g2_inv_1 _12339_ (.Y(_06539_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[31] ));
 sg13g2_inv_1 _12340_ (.Y(_06540_),
    .A(net6524));
 sg13g2_inv_1 _12341_ (.Y(_06541_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[30] ));
 sg13g2_inv_2 _12342_ (.Y(_06542_),
    .A(\fpga_top.uart_top.uart_rec_char.pdata[0] ));
 sg13g2_inv_1 _12343_ (.Y(_06543_),
    .A(net5627));
 sg13g2_inv_2 _12344_ (.Y(_06544_),
    .A(\fpga_top.uart_top.uart_rec_char.pdata[4] ));
 sg13g2_inv_1 _12345_ (.Y(_06545_),
    .A(net3944));
 sg13g2_inv_4 _12346_ (.A(net5634),
    .Y(_06546_));
 sg13g2_inv_2 _12347_ (.Y(_06547_),
    .A(\fpga_top.bus_gather.i_read_adr[2] ));
 sg13g2_inv_4 _12348_ (.A(\fpga_top.cpu_top.alui_shamt[2] ),
    .Y(_06548_));
 sg13g2_inv_8 _12349_ (.Y(_06549_),
    .A(net5571));
 sg13g2_inv_4 _12350_ (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[5] ),
    .Y(_06550_));
 sg13g2_inv_1 _12351_ (.Y(_06551_),
    .A(net5582));
 sg13g2_inv_4 _12352_ (.A(net5583),
    .Y(_06552_));
 sg13g2_inv_2 _12353_ (.Y(_06553_),
    .A(net5579));
 sg13g2_inv_4 _12354_ (.A(\fpga_top.cpu_top.br_ofs[7] ),
    .Y(_06554_));
 sg13g2_inv_4 _12355_ (.A(net6615),
    .Y(_06555_));
 sg13g2_inv_4 _12356_ (.A(net5570),
    .Y(_06556_));
 sg13g2_inv_4 _12357_ (.A(\fpga_top.cpu_top.br_ofs[10] ),
    .Y(_06557_));
 sg13g2_inv_4 _12358_ (.A(\fpga_top.cpu_top.br_ofs[5] ),
    .Y(_06558_));
 sg13g2_inv_8 _12359_ (.Y(_06559_),
    .A(net6520));
 sg13g2_inv_4 _12360_ (.A(\fpga_top.cpu_top.br_ofs[1] ),
    .Y(_06560_));
 sg13g2_inv_4 _12361_ (.A(net3303),
    .Y(_06561_));
 sg13g2_inv_8 _12362_ (.Y(_06562_),
    .A(net3695));
 sg13g2_inv_4 _12363_ (.A(net5572),
    .Y(_06563_));
 sg13g2_inv_4 _12364_ (.A(\fpga_top.cpu_top.br_ofs[11] ),
    .Y(_06564_));
 sg13g2_inv_2 _12365_ (.Y(_06565_),
    .A(net5810));
 sg13g2_inv_4 _12366_ (.A(net5803),
    .Y(_06566_));
 sg13g2_inv_2 _12367_ (.Y(_06567_),
    .A(net5800));
 sg13g2_inv_4 _12368_ (.A(\fpga_top.cpu_top.alui_shamt[3] ),
    .Y(_06568_));
 sg13g2_inv_2 _12369_ (.Y(_06569_),
    .A(\fpga_top.cpu_top.br_ofs[3] ));
 sg13g2_inv_4 _12370_ (.A(net3571),
    .Y(_06570_));
 sg13g2_inv_2 _12371_ (.Y(_06571_),
    .A(net5798));
 sg13g2_inv_4 _12372_ (.A(net5797),
    .Y(_06572_));
 sg13g2_inv_4 _12373_ (.A(net5790),
    .Y(_06573_));
 sg13g2_inv_4 _12374_ (.A(net5786),
    .Y(_06574_));
 sg13g2_inv_4 _12375_ (.A(\fpga_top.cpu_top.alui_shamt[4] ),
    .Y(_06575_));
 sg13g2_inv_2 _12376_ (.Y(_06576_),
    .A(\fpga_top.cpu_top.br_ofs[4] ));
 sg13g2_inv_4 _12377_ (.A(net3633),
    .Y(_06577_));
 sg13g2_inv_4 _12378_ (.A(net5777),
    .Y(_06578_));
 sg13g2_inv_4 _12379_ (.A(net5774),
    .Y(_06579_));
 sg13g2_inv_4 _12380_ (.A(net5760),
    .Y(_06580_));
 sg13g2_inv_2 _12381_ (.Y(_06581_),
    .A(net5756));
 sg13g2_inv_8 _12382_ (.Y(_06582_),
    .A(net5754));
 sg13g2_inv_1 _12383_ (.Y(_06583_),
    .A(net1568));
 sg13g2_inv_4 _12384_ (.A(net6538),
    .Y(_06584_));
 sg13g2_inv_1 _12385_ (.Y(_06585_),
    .A(net1528));
 sg13g2_inv_4 _12386_ (.A(net2160),
    .Y(_06586_));
 sg13g2_inv_4 _12387_ (.A(net6483),
    .Y(_06587_));
 sg13g2_inv_4 _12388_ (.A(net5596),
    .Y(_06588_));
 sg13g2_inv_1 _12389_ (.Y(_06589_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[6] ));
 sg13g2_inv_4 _12390_ (.A(net6493),
    .Y(_06590_));
 sg13g2_inv_2 _12391_ (.Y(_06591_),
    .A(net2768));
 sg13g2_inv_4 _12392_ (.A(net6506),
    .Y(_06592_));
 sg13g2_inv_4 _12393_ (.A(net2938),
    .Y(_06593_));
 sg13g2_inv_8 _12394_ (.Y(_06594_),
    .A(net6535));
 sg13g2_inv_2 _12395_ (.Y(_06595_),
    .A(net3657));
 sg13g2_inv_1 _12396_ (.Y(_06596_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[11] ));
 sg13g2_inv_8 _12397_ (.Y(_06597_),
    .A(\fpga_top.bus_gather.i_read_adr[11] ));
 sg13g2_inv_1 _12398_ (.Y(_06598_),
    .A(\fpga_top.bus_gather.d_write_data[12] ));
 sg13g2_inv_8 _12399_ (.Y(_06599_),
    .A(\fpga_top.bus_gather.i_read_adr[12] ));
 sg13g2_inv_1 _12400_ (.Y(_06600_),
    .A(\fpga_top.bus_gather.d_write_data[13] ));
 sg13g2_inv_4 _12401_ (.A(net6564),
    .Y(_06601_));
 sg13g2_inv_1 _12402_ (.Y(_06602_),
    .A(\fpga_top.bus_gather.d_write_data[14] ));
 sg13g2_inv_8 _12403_ (.Y(_06603_),
    .A(net6504));
 sg13g2_inv_4 _12404_ (.A(net3505),
    .Y(_06604_));
 sg13g2_inv_8 _12405_ (.Y(_06605_),
    .A(net6519));
 sg13g2_inv_1 _12406_ (.Y(_06606_),
    .A(net6125));
 sg13g2_inv_1 _12407_ (.Y(_06607_),
    .A(net1563));
 sg13g2_inv_2 _12408_ (.Y(_06608_),
    .A(\fpga_top.cpu_top.csr_uimm[1] ));
 sg13g2_inv_2 _12409_ (.Y(_06609_),
    .A(net3351));
 sg13g2_inv_1 _12410_ (.Y(_06610_),
    .A(\fpga_top.bus_gather.d_write_data[17] ));
 sg13g2_inv_8 _12411_ (.Y(_06611_),
    .A(net6557));
 sg13g2_inv_1 _12412_ (.Y(_06612_),
    .A(\fpga_top.bus_gather.d_write_data[18] ));
 sg13g2_inv_1 _12413_ (.Y(_06613_),
    .A(net1707));
 sg13g2_inv_8 _12414_ (.Y(_06614_),
    .A(\fpga_top.bus_gather.i_read_adr[18] ));
 sg13g2_inv_2 _12415_ (.Y(_06615_),
    .A(net2720));
 sg13g2_inv_8 _12416_ (.Y(_06616_),
    .A(\fpga_top.bus_gather.d_write_data[19] ));
 sg13g2_inv_8 _12417_ (.Y(_06617_),
    .A(net6579));
 sg13g2_inv_4 _12418_ (.A(\fpga_top.cpu_top.csr_uimm[4] ),
    .Y(_06618_));
 sg13g2_inv_8 _12419_ (.Y(_06619_),
    .A(net4038));
 sg13g2_inv_8 _12420_ (.Y(_06620_),
    .A(net6558));
 sg13g2_inv_1 _12421_ (.Y(_06621_),
    .A(net3794));
 sg13g2_inv_1 _12422_ (.Y(_06622_),
    .A(\fpga_top.bus_gather.d_write_data[21] ));
 sg13g2_inv_4 _12423_ (.A(net6562),
    .Y(_06623_));
 sg13g2_inv_8 _12424_ (.Y(_06624_),
    .A(\fpga_top.bus_gather.d_write_data[22] ));
 sg13g2_inv_1 _12425_ (.Y(_06625_),
    .A(\fpga_top.bus_gather.d_write_data[23] ));
 sg13g2_inv_8 _12426_ (.Y(_06626_),
    .A(\fpga_top.bus_gather.i_read_adr[23] ));
 sg13g2_inv_2 _12427_ (.Y(_06627_),
    .A(net2993));
 sg13g2_inv_1 _12428_ (.Y(_06628_),
    .A(\fpga_top.bus_gather.d_write_data[24] ));
 sg13g2_inv_8 _12429_ (.Y(_06629_),
    .A(net6549));
 sg13g2_inv_1 _12430_ (.Y(_06630_),
    .A(\fpga_top.bus_gather.d_write_data[25] ));
 sg13g2_inv_8 _12431_ (.Y(_06631_),
    .A(net6413));
 sg13g2_inv_1 _12432_ (.Y(_06632_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[26] ));
 sg13g2_inv_1 _12433_ (.Y(_06633_),
    .A(\fpga_top.bus_gather.d_write_data[26] ));
 sg13g2_inv_8 _12434_ (.Y(_06634_),
    .A(net6530));
 sg13g2_inv_1 _12435_ (.Y(_06635_),
    .A(\fpga_top.bus_gather.d_write_data[27] ));
 sg13g2_inv_8 _12436_ (.Y(_06636_),
    .A(\fpga_top.bus_gather.i_read_adr[27] ));
 sg13g2_inv_1 _12437_ (.Y(_06637_),
    .A(net3967));
 sg13g2_inv_1 _12438_ (.Y(_06638_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[28] ));
 sg13g2_inv_8 _12439_ (.Y(_06639_),
    .A(\fpga_top.bus_gather.d_write_data[28] ));
 sg13g2_inv_1 _12440_ (.Y(_06640_),
    .A(\fpga_top.bus_gather.d_write_data[29] ));
 sg13g2_inv_8 _12441_ (.Y(_06641_),
    .A(\fpga_top.bus_gather.i_read_adr[29] ));
 sg13g2_inv_1 _12442_ (.Y(_06642_),
    .A(\fpga_top.bus_gather.d_write_data[30] ));
 sg13g2_inv_8 _12443_ (.Y(_06643_),
    .A(\fpga_top.bus_gather.i_read_adr[30] ));
 sg13g2_inv_2 _12444_ (.Y(_06644_),
    .A(net2630));
 sg13g2_inv_1 _12445_ (.Y(_06645_),
    .A(\fpga_top.bus_gather.d_write_data[31] ));
 sg13g2_inv_8 _12446_ (.Y(_06646_),
    .A(net6490));
 sg13g2_inv_1 _12447_ (.Y(_06647_),
    .A(\fpga_top.cmd_st_ma ));
 sg13g2_inv_1 _12448_ (.Y(_06648_),
    .A(net3181));
 sg13g2_inv_1 _12449_ (.Y(_06649_),
    .A(\fpga_top.io_spi_lite.spi_mode[1] ));
 sg13g2_inv_1 _12450_ (.Y(_06650_),
    .A(\fpga_top.qspi_if.sck_div[1] ));
 sg13g2_inv_1 _12451_ (.Y(_06651_),
    .A(\fpga_top.qspi_if.sck_cntr[2] ));
 sg13g2_inv_1 _12452_ (.Y(_06652_),
    .A(net6394));
 sg13g2_inv_2 _12453_ (.Y(_06653_),
    .A(net3857));
 sg13g2_inv_1 _12454_ (.Y(_06654_),
    .A(\fpga_top.qspi_if.sck_cntr[4] ));
 sg13g2_inv_2 _12455_ (.Y(_06655_),
    .A(\fpga_top.qspi_if.sck_div[5] ));
 sg13g2_inv_1 _12456_ (.Y(_06656_),
    .A(\fpga_top.qspi_if.sck_cntr[6] ));
 sg13g2_inv_1 _12457_ (.Y(_06657_),
    .A(\fpga_top.qspi_if.sck_div[6] ));
 sg13g2_inv_1 _12458_ (.Y(_06658_),
    .A(\fpga_top.qspi_if.sck_div[7] ));
 sg13g2_inv_1 _12459_ (.Y(_06659_),
    .A(\fpga_top.qspi_if.sck_cntr[8] ));
 sg13g2_inv_1 _12460_ (.Y(_06660_),
    .A(net3079));
 sg13g2_inv_1 _12461_ (.Y(_06661_),
    .A(net5629));
 sg13g2_inv_1 _12462_ (.Y(_06662_),
    .A(net6481));
 sg13g2_inv_1 _12463_ (.Y(_06663_),
    .A(net1378));
 sg13g2_inv_1 _12464_ (.Y(_06664_),
    .A(net3981));
 sg13g2_inv_2 _12465_ (.Y(_06665_),
    .A(net5665));
 sg13g2_inv_2 _12466_ (.Y(_06666_),
    .A(net6402));
 sg13g2_inv_2 _12467_ (.Y(_06667_),
    .A(net6370));
 sg13g2_inv_2 _12468_ (.Y(_06668_),
    .A(net3937));
 sg13g2_inv_4 _12469_ (.A(net6238),
    .Y(_06669_));
 sg13g2_inv_2 _12470_ (.Y(_06670_),
    .A(net4035));
 sg13g2_inv_1 _12471_ (.Y(_06671_),
    .A(net6194));
 sg13g2_inv_1 _12472_ (.Y(_06672_),
    .A(net6350));
 sg13g2_inv_1 _12473_ (.Y(_06673_),
    .A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[1] ));
 sg13g2_inv_1 _12474_ (.Y(_06674_),
    .A(net6283));
 sg13g2_inv_4 _12475_ (.A(net6516),
    .Y(_06675_));
 sg13g2_inv_2 _12476_ (.Y(_06676_),
    .A(\fpga_top.qspi_if.rdedge[2] ));
 sg13g2_inv_1 _12477_ (.Y(_06677_),
    .A(\fpga_top.qspi_if.rdedge[0] ));
 sg13g2_inv_1 _12478_ (.Y(_06678_),
    .A(\fpga_top.io_uart_out.rx_first_read ));
 sg13g2_inv_4 _12479_ (.A(net5652),
    .Y(_06679_));
 sg13g2_inv_1 _12480_ (.Y(_06680_),
    .A(net6489));
 sg13g2_inv_4 _12481_ (.A(\fpga_top.cpu_top.csr_wdata_mon[1] ),
    .Y(_06681_));
 sg13g2_inv_1 _12482_ (.Y(_06682_),
    .A(net3968));
 sg13g2_inv_4 _12483_ (.A(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .Y(_06683_));
 sg13g2_inv_4 _12484_ (.A(net5664),
    .Y(_06684_));
 sg13g2_inv_2 _12485_ (.Y(_06685_),
    .A(net6143));
 sg13g2_inv_1 _12486_ (.Y(_06686_),
    .A(net6335));
 sg13g2_inv_1 _12487_ (.Y(_06687_),
    .A(net6179));
 sg13g2_inv_2 _12488_ (.Y(_06688_),
    .A(net3848));
 sg13g2_inv_2 _12489_ (.Y(_06689_),
    .A(net3930));
 sg13g2_inv_1 _12490_ (.Y(_06690_),
    .A(net6197));
 sg13g2_inv_1 _12491_ (.Y(_06691_),
    .A(\fpga_top.io_frc.frc_cmp_val[7] ));
 sg13g2_inv_1 _12492_ (.Y(_06692_),
    .A(\fpga_top.io_frc.frc_cmp_val[6] ));
 sg13g2_inv_1 _12493_ (.Y(_06693_),
    .A(net6330));
 sg13g2_inv_1 _12494_ (.Y(_06694_),
    .A(\fpga_top.io_frc.frc_cmp_val[5] ));
 sg13g2_inv_1 _12495_ (.Y(_06695_),
    .A(net6321));
 sg13g2_inv_1 _12496_ (.Y(_06696_),
    .A(net3980));
 sg13g2_inv_2 _12497_ (.Y(_06697_),
    .A(net3902));
 sg13g2_inv_2 _12498_ (.Y(_06698_),
    .A(\fpga_top.io_frc.frc_cmp_val[15] ));
 sg13g2_inv_2 _12499_ (.Y(_06699_),
    .A(net4051));
 sg13g2_inv_1 _12500_ (.Y(_06700_),
    .A(\fpga_top.io_frc.frc_cmp_val[14] ));
 sg13g2_inv_4 _12501_ (.A(net3745),
    .Y(_06701_));
 sg13g2_inv_1 _12502_ (.Y(_06702_),
    .A(\fpga_top.io_frc.frc_cmp_val[13] ));
 sg13g2_inv_1 _12503_ (.Y(_06703_),
    .A(net6250));
 sg13g2_inv_1 _12504_ (.Y(_06704_),
    .A(\fpga_top.io_frc.frc_cmp_val[12] ));
 sg13g2_inv_2 _12505_ (.Y(_06705_),
    .A(\fpga_top.io_frc.frc_cmp_val[11] ));
 sg13g2_inv_1 _12506_ (.Y(_06706_),
    .A(net4016));
 sg13g2_inv_2 _12507_ (.Y(_06707_),
    .A(net3858));
 sg13g2_inv_1 _12508_ (.Y(_06708_),
    .A(net4028));
 sg13g2_inv_1 _12509_ (.Y(_06709_),
    .A(\fpga_top.io_frc.frc_cmp_val[9] ));
 sg13g2_inv_2 _12510_ (.Y(_06710_),
    .A(net6129));
 sg13g2_inv_1 _12511_ (.Y(_06711_),
    .A(\fpga_top.io_frc.frc_cmp_val[8] ));
 sg13g2_inv_4 _12512_ (.A(net6086),
    .Y(_06712_));
 sg13g2_inv_1 _12513_ (.Y(_06713_),
    .A(net4055));
 sg13g2_inv_2 _12514_ (.Y(_06714_),
    .A(net6136));
 sg13g2_inv_1 _12515_ (.Y(_06715_),
    .A(net6347));
 sg13g2_inv_1 _12516_ (.Y(_06716_),
    .A(\fpga_top.io_frc.frc_cmp_val[28] ));
 sg13g2_inv_2 _12517_ (.Y(_06717_),
    .A(net3862));
 sg13g2_inv_2 _12518_ (.Y(_06718_),
    .A(net4040));
 sg13g2_inv_2 _12519_ (.Y(_06719_),
    .A(net6181));
 sg13g2_inv_1 _12520_ (.Y(_06720_),
    .A(\fpga_top.io_frc.frc_cmp_val[25] ));
 sg13g2_inv_1 _12521_ (.Y(_06721_),
    .A(net4005));
 sg13g2_inv_1 _12522_ (.Y(_06722_),
    .A(\fpga_top.io_frc.frc_cmp_val[24] ));
 sg13g2_inv_2 _12523_ (.Y(_06723_),
    .A(net6165));
 sg13g2_inv_2 _12524_ (.Y(_06724_),
    .A(net4072));
 sg13g2_inv_1 _12525_ (.Y(_06725_),
    .A(\fpga_top.io_frc.frc_cmp_val[22] ));
 sg13g2_inv_2 _12526_ (.Y(_06726_),
    .A(net3824));
 sg13g2_inv_1 _12527_ (.Y(_06727_),
    .A(\fpga_top.io_frc.frc_cmp_val[21] ));
 sg13g2_inv_4 _12528_ (.A(net3756),
    .Y(_06728_));
 sg13g2_inv_2 _12529_ (.Y(_06729_),
    .A(net6273));
 sg13g2_inv_2 _12530_ (.Y(_06730_),
    .A(net4039));
 sg13g2_inv_4 _12531_ (.A(net3803),
    .Y(_06731_));
 sg13g2_inv_1 _12532_ (.Y(_06732_),
    .A(\fpga_top.io_frc.frc_cntr_val[18] ));
 sg13g2_inv_1 _12533_ (.Y(_06733_),
    .A(\fpga_top.io_frc.frc_cntr_val[63] ));
 sg13g2_inv_1 _12534_ (.Y(_06734_),
    .A(\fpga_top.io_frc.frc_cntr_val[62] ));
 sg13g2_inv_1 _12535_ (.Y(_06735_),
    .A(\fpga_top.io_frc.frc_cmp_val[62] ));
 sg13g2_inv_1 _12536_ (.Y(_06736_),
    .A(\fpga_top.io_frc.frc_cmp_val[61] ));
 sg13g2_inv_1 _12537_ (.Y(_06737_),
    .A(\fpga_top.io_frc.frc_cntr_val[60] ));
 sg13g2_inv_2 _12538_ (.Y(_06738_),
    .A(net2208));
 sg13g2_inv_1 _12539_ (.Y(_06739_),
    .A(\fpga_top.io_frc.frc_cntr_val[57] ));
 sg13g2_inv_1 _12540_ (.Y(_06740_),
    .A(\fpga_top.io_frc.frc_cntr_val[56] ));
 sg13g2_inv_1 _12541_ (.Y(_06741_),
    .A(\fpga_top.io_frc.frc_cmp_val[49] ));
 sg13g2_inv_1 _12542_ (.Y(_06742_),
    .A(\fpga_top.io_frc.frc_cntr_val[48] ));
 sg13g2_inv_1 _12543_ (.Y(_06743_),
    .A(\fpga_top.io_frc.frc_cmp_val[48] ));
 sg13g2_inv_1 _12544_ (.Y(_06744_),
    .A(\fpga_top.io_frc.frc_cntr_val[51] ));
 sg13g2_inv_1 _12545_ (.Y(_06745_),
    .A(\fpga_top.io_frc.frc_cmp_val[51] ));
 sg13g2_inv_2 _12546_ (.Y(_06746_),
    .A(net3645));
 sg13g2_inv_1 _12547_ (.Y(_06747_),
    .A(\fpga_top.io_frc.frc_cmp_val[50] ));
 sg13g2_inv_2 _12548_ (.Y(_06748_),
    .A(\fpga_top.io_frc.frc_cntr_val[55] ));
 sg13g2_inv_1 _12549_ (.Y(_06749_),
    .A(\fpga_top.io_frc.frc_cmp_val[55] ));
 sg13g2_inv_1 _12550_ (.Y(_06750_),
    .A(\fpga_top.io_frc.frc_cmp_val[54] ));
 sg13g2_inv_2 _12551_ (.Y(_06751_),
    .A(\fpga_top.io_frc.frc_cntr_val[53] ));
 sg13g2_inv_2 _12552_ (.Y(_06752_),
    .A(net2138));
 sg13g2_inv_1 _12553_ (.Y(_06753_),
    .A(\fpga_top.io_frc.frc_cmp_val[52] ));
 sg13g2_inv_1 _12554_ (.Y(_06754_),
    .A(\fpga_top.io_frc.frc_cntr_val[40] ));
 sg13g2_inv_2 _12555_ (.Y(_06755_),
    .A(net1958));
 sg13g2_inv_2 _12556_ (.Y(_06756_),
    .A(\fpga_top.io_frc.frc_cntr_val[46] ));
 sg13g2_inv_1 _12557_ (.Y(_06757_),
    .A(\fpga_top.io_frc.frc_cmp_val[39] ));
 sg13g2_inv_2 _12558_ (.Y(_06758_),
    .A(\fpga_top.io_frc.frc_cntr_val[38] ));
 sg13g2_inv_1 _12559_ (.Y(_06759_),
    .A(\fpga_top.io_frc.frc_cmp_val[38] ));
 sg13g2_inv_2 _12560_ (.Y(_06760_),
    .A(\fpga_top.io_frc.frc_cntr_val[37] ));
 sg13g2_inv_1 _12561_ (.Y(_06761_),
    .A(\fpga_top.io_frc.frc_cntr_val[36] ));
 sg13g2_inv_1 _12562_ (.Y(_06762_),
    .A(net3964));
 sg13g2_inv_1 _12563_ (.Y(_06763_),
    .A(net4024));
 sg13g2_inv_2 _12564_ (.Y(_06764_),
    .A(\fpga_top.io_frc.frc_cntr_val[34] ));
 sg13g2_inv_2 _12565_ (.Y(_06765_),
    .A(net2182));
 sg13g2_inv_1 _12566_ (.Y(_06766_),
    .A(\fpga_top.io_frc.frc_cmp_val[33] ));
 sg13g2_inv_2 _12567_ (.Y(_06767_),
    .A(\fpga_top.io_frc.frc_cntr_val[32] ));
 sg13g2_inv_1 _12568_ (.Y(_06768_),
    .A(\fpga_top.io_frc.frc_cmp_val[32] ));
 sg13g2_inv_1 _12569_ (.Y(_06769_),
    .A(net3839));
 sg13g2_inv_1 _12570_ (.Y(_06770_),
    .A(\fpga_top.dbg_bpoint_en[0] ));
 sg13g2_inv_2 _12571_ (.Y(_06771_),
    .A(net6353));
 sg13g2_inv_1 _12572_ (.Y(_06772_),
    .A(net4057));
 sg13g2_inv_4 _12573_ (.A(\fpga_top.cpu_top.execution.csr_array.frc_cntr_val_leq ),
    .Y(_06773_));
 sg13g2_inv_1 _12574_ (.Y(_06774_),
    .A(\fpga_top.cpu_top.pc_stage.frc_cntr_val_leq_lat ));
 sg13g2_inv_4 _12575_ (.A(net5588),
    .Y(_06775_));
 sg13g2_inv_1 _12576_ (.Y(_06776_),
    .A(\fpga_top.interrupter.int_status_int0 ));
 sg13g2_inv_1 _12577_ (.Y(_06777_),
    .A(net2835));
 sg13g2_inv_1 _12578_ (.Y(_06778_),
    .A(\fpga_top.io_spi_lite.sck_div[2] ));
 sg13g2_inv_1 _12579_ (.Y(_06779_),
    .A(\fpga_top.io_spi_lite.spi_sck_div[4] ));
 sg13g2_inv_1 _12580_ (.Y(_06780_),
    .A(\fpga_top.io_spi_lite.sck_div[5] ));
 sg13g2_inv_1 _12581_ (.Y(_06781_),
    .A(\fpga_top.io_spi_lite.spi_sck_div[6] ));
 sg13g2_inv_1 _12582_ (.Y(_06782_),
    .A(\fpga_top.io_spi_lite.sck_div[7] ));
 sg13g2_inv_1 _12583_ (.Y(_06783_),
    .A(\fpga_top.io_spi_lite.spi_sck_div[8] ));
 sg13g2_inv_1 _12584_ (.Y(_06784_),
    .A(\fpga_top.io_spi_lite.sck_div[9] ));
 sg13g2_inv_1 _12585_ (.Y(_06785_),
    .A(\fpga_top.io_spi_lite.spi_sck_div[9] ));
 sg13g2_inv_2 _12586_ (.Y(_06786_),
    .A(net6491));
 sg13g2_inv_2 _12587_ (.Y(_06787_),
    .A(net6536));
 sg13g2_inv_4 _12588_ (.A(net5833),
    .Y(_06788_));
 sg13g2_inv_4 _12589_ (.A(net5663),
    .Y(_06789_));
 sg13g2_inv_8 _12590_ (.Y(_06790_),
    .A(\fpga_top.cpu_start_adr[6] ));
 sg13g2_inv_4 _12591_ (.A(net5656),
    .Y(_06791_));
 sg13g2_inv_8 _12592_ (.Y(_06792_),
    .A(net5653));
 sg13g2_inv_8 _12593_ (.Y(_06793_),
    .A(net5651));
 sg13g2_inv_2 _12594_ (.Y(_06794_),
    .A(\fpga_top.cpu_start_adr[12] ));
 sg13g2_inv_1 _12595_ (.Y(_06795_),
    .A(\fpga_top.cpu_start_adr[13] ));
 sg13g2_inv_8 _12596_ (.Y(_06796_),
    .A(net5650));
 sg13g2_inv_1 _12597_ (.Y(_06797_),
    .A(\fpga_top.cpu_start_adr[15] ));
 sg13g2_inv_8 _12598_ (.Y(_06798_),
    .A(net5649));
 sg13g2_inv_8 _12599_ (.Y(_06799_),
    .A(net5648));
 sg13g2_inv_8 _12600_ (.Y(_06800_),
    .A(net5647));
 sg13g2_inv_8 _12601_ (.Y(_06801_),
    .A(\fpga_top.cpu_start_adr[19] ));
 sg13g2_inv_8 _12602_ (.Y(_06802_),
    .A(net5646));
 sg13g2_inv_8 _12603_ (.Y(_06803_),
    .A(net5643));
 sg13g2_inv_4 _12604_ (.A(net5642),
    .Y(_06804_));
 sg13g2_inv_8 _12605_ (.Y(_06805_),
    .A(\fpga_top.cpu_start_adr[24] ));
 sg13g2_inv_16 _12606_ (.A(net6560),
    .Y(_06806_));
 sg13g2_inv_8 _12607_ (.Y(_06807_),
    .A(\fpga_top.cpu_start_adr[26] ));
 sg13g2_inv_4 _12608_ (.A(net5638),
    .Y(_06808_));
 sg13g2_inv_8 _12609_ (.Y(_06809_),
    .A(net5637));
 sg13g2_inv_4 _12610_ (.A(net5635),
    .Y(_06810_));
 sg13g2_inv_4 _12611_ (.A(net2221),
    .Y(_06811_));
 sg13g2_inv_1 _12612_ (.Y(_06812_),
    .A(net8));
 sg13g2_inv_1 _12613_ (.Y(_06813_),
    .A(\fpga_top.qspi_if.dbg_2div_cec_lat ));
 sg13g2_inv_1 _12614_ (.Y(_06814_),
    .A(\fpga_top.qspi_if.wdata[0] ));
 sg13g2_inv_4 _12615_ (.A(net5701),
    .Y(_06815_));
 sg13g2_inv_1 _12616_ (.Y(_06816_),
    .A(\fpga_top.qspi_if.adr_rw[12] ));
 sg13g2_inv_1 _12617_ (.Y(_06817_),
    .A(\fpga_top.qspi_if.wrcmd0[0] ));
 sg13g2_inv_1 _12618_ (.Y(_06818_),
    .A(\fpga_top.qspi_if.rdcmd1[2] ));
 sg13g2_inv_1 _12619_ (.Y(_06819_),
    .A(\fpga_top.qspi_if.wrcmd1[2] ));
 sg13g2_inv_1 _12620_ (.Y(_06820_),
    .A(\fpga_top.qspi_if.wdata[1] ));
 sg13g2_inv_1 _12621_ (.Y(_06821_),
    .A(\fpga_top.qspi_if.wdata[5] ));
 sg13g2_inv_1 _12622_ (.Y(_06822_),
    .A(\fpga_top.qspi_if.wdata[29] ));
 sg13g2_inv_1 _12623_ (.Y(_06823_),
    .A(\fpga_top.qspi_if.wdata[6] ));
 sg13g2_inv_1 _12624_ (.Y(_06824_),
    .A(\fpga_top.qspi_if.wdata[30] ));
 sg13g2_inv_1 _12625_ (.Y(_06825_),
    .A(\fpga_top.qspi_if.wdata[7] ));
 sg13g2_inv_1 _12626_ (.Y(_06826_),
    .A(\fpga_top.qspi_if.wdata[31] ));
 sg13g2_inv_1 _12627_ (.Y(_06827_),
    .A(net6471));
 sg13g2_inv_1 _12628_ (.Y(_06828_),
    .A(\fpga_top.qspi_if.word_data[28] ));
 sg13g2_inv_1 _12629_ (.Y(_06829_),
    .A(net6151));
 sg13g2_inv_1 _12630_ (.Y(_06830_),
    .A(net3888));
 sg13g2_inv_2 _12631_ (.Y(_06831_),
    .A(net3838));
 sg13g2_inv_2 _12632_ (.Y(_06832_),
    .A(net1973));
 sg13g2_inv_2 _12633_ (.Y(_06833_),
    .A(net2123));
 sg13g2_inv_1 _12634_ (.Y(_06834_),
    .A(net2113));
 sg13g2_inv_1 _12635_ (.Y(_06835_),
    .A(net3973));
 sg13g2_inv_2 _12636_ (.Y(_06836_),
    .A(net2373));
 sg13g2_inv_1 _12637_ (.Y(_06837_),
    .A(net3142));
 sg13g2_inv_2 _12638_ (.Y(_06838_),
    .A(net3606));
 sg13g2_inv_1 _12639_ (.Y(_06839_),
    .A(net3965));
 sg13g2_inv_2 _12640_ (.Y(_06840_),
    .A(net3305));
 sg13g2_inv_1 _12641_ (.Y(_06841_),
    .A(net3988));
 sg13g2_inv_1 _12642_ (.Y(_06842_),
    .A(net6174));
 sg13g2_inv_2 _12643_ (.Y(_06843_),
    .A(net4022));
 sg13g2_inv_2 _12644_ (.Y(_06844_),
    .A(net4043));
 sg13g2_inv_1 _12645_ (.Y(_06845_),
    .A(net6111));
 sg13g2_inv_4 _12646_ (.A(net6147),
    .Y(_06846_));
 sg13g2_inv_1 _12647_ (.Y(_06847_),
    .A(net1385));
 sg13g2_inv_1 _12648_ (.Y(_06848_),
    .A(net5410));
 sg13g2_inv_1 _12649_ (.Y(_06849_),
    .A(net1631));
 sg13g2_inv_1 _12650_ (.Y(_06850_),
    .A(net1809));
 sg13g2_inv_1 _12651_ (.Y(_06851_),
    .A(net1830));
 sg13g2_inv_1 _12652_ (.Y(_06852_),
    .A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][2] ));
 sg13g2_inv_1 _12653_ (.Y(_06853_),
    .A(net1814));
 sg13g2_inv_1 _12654_ (.Y(_06854_),
    .A(net1956));
 sg13g2_inv_1 _12655_ (.Y(_06855_),
    .A(net1738));
 sg13g2_inv_1 _12656_ (.Y(_06856_),
    .A(net1853));
 sg13g2_inv_1 _12657_ (.Y(_06857_),
    .A(net3720));
 sg13g2_inv_1 _12658_ (.Y(_06858_),
    .A(net3718));
 sg13g2_inv_1 _12659_ (.Y(_06859_),
    .A(net2971));
 sg13g2_inv_1 _12660_ (.Y(_06860_),
    .A(net3811));
 sg13g2_inv_1 _12661_ (.Y(_06861_),
    .A(\fpga_top.uart_top.uart_logics.data_0[22] ));
 sg13g2_inv_1 _12662_ (.Y(_06862_),
    .A(\fpga_top.io_uart_out.uart_io_char[7] ));
 sg13g2_inv_2 _12663_ (.Y(_06863_),
    .A(net5465));
 sg13g2_inv_4 _12664_ (.A(net5452),
    .Y(_06864_));
 sg13g2_inv_1 _12665_ (.Y(_06865_),
    .A(uio_oe[4]));
 sg13g2_inv_2 _12666_ (.Y(_06866_),
    .A(net1686));
 sg13g2_inv_1 _12667_ (.Y(_06867_),
    .A(\fpga_top.io_uart_out.re_uart_rdflg_dly[4] ));
 sg13g2_inv_1 _12668_ (.Y(_06868_),
    .A(\fpga_top.io_led.re_gpio_value_dly[1] ));
 sg13g2_inv_1 _12669_ (.Y(_06869_),
    .A(net5710));
 sg13g2_inv_1 _12670_ (.Y(_06870_),
    .A(net5720));
 sg13g2_inv_8 _12671_ (.Y(_06871_),
    .A(net5745));
 sg13g2_inv_1 _12672_ (.Y(_06872_),
    .A(net5689));
 sg13g2_inv_8 _12673_ (.Y(_06873_),
    .A(net5696));
 sg13g2_inv_4 _12674_ (.A(net5387),
    .Y(_06874_));
 sg13g2_inv_2 _12675_ (.Y(_06875_),
    .A(\fpga_top.io_spi_lite.spi_mode[0] ));
 sg13g2_inv_1 _12676_ (.Y(_06876_),
    .A(net1705));
 sg13g2_inv_1 _12677_ (.Y(_06877_),
    .A(net1569));
 sg13g2_inv_1 _12678_ (.Y(_06878_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_sie ));
 sg13g2_inv_1 _12679_ (.Y(_06879_),
    .A(uio_out[5]));
 sg13g2_inv_1 _12680_ (.Y(_06880_),
    .A(\fpga_top.io_led.gpio_in_lat2[1] ));
 sg13g2_inv_1 _12681_ (.Y(_06881_),
    .A(net1575));
 sg13g2_inv_1 _12682_ (.Y(_06882_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[2] ));
 sg13g2_inv_1 _12683_ (.Y(_06883_),
    .A(net1857));
 sg13g2_inv_1 _12684_ (.Y(_06884_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[3] ));
 sg13g2_inv_1 _12685_ (.Y(_06885_),
    .A(net1626));
 sg13g2_inv_1 _12686_ (.Y(_06886_),
    .A(net1993));
 sg13g2_inv_2 _12687_ (.Y(_06887_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[4] ));
 sg13g2_inv_1 _12688_ (.Y(_06888_),
    .A(net1562));
 sg13g2_inv_1 _12689_ (.Y(_06889_),
    .A(net1740));
 sg13g2_inv_1 _12690_ (.Y(_06890_),
    .A(net2184));
 sg13g2_inv_1 _12691_ (.Y(_06891_),
    .A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][5] ));
 sg13g2_inv_1 _12692_ (.Y(_06892_),
    .A(net1566));
 sg13g2_inv_1 _12693_ (.Y(_06893_),
    .A(net1623));
 sg13g2_inv_2 _12694_ (.Y(_06894_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[7] ));
 sg13g2_inv_1 _12695_ (.Y(_06895_),
    .A(net1711));
 sg13g2_inv_1 _12696_ (.Y(_06896_),
    .A(net1947));
 sg13g2_inv_1 _12697_ (.Y(_06897_),
    .A(net1772));
 sg13g2_inv_1 _12698_ (.Y(_06898_),
    .A(net1946));
 sg13g2_inv_1 _12699_ (.Y(_06899_),
    .A(net1929));
 sg13g2_inv_2 _12700_ (.Y(_06900_),
    .A(net3890));
 sg13g2_inv_1 _12701_ (.Y(_06901_),
    .A(net2777));
 sg13g2_inv_2 _12702_ (.Y(_06902_),
    .A(net4014));
 sg13g2_inv_1 _12703_ (.Y(_06903_),
    .A(\fpga_top.io_uart_out.rx_write_error ));
 sg13g2_inv_1 _12704_ (.Y(_06904_),
    .A(net1786));
 sg13g2_inv_1 _12705_ (.Y(_06905_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[11] ));
 sg13g2_inv_1 _12706_ (.Y(_06906_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[12] ));
 sg13g2_inv_1 _12707_ (.Y(_06907_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[13] ));
 sg13g2_inv_1 _12708_ (.Y(_06908_),
    .A(net1549));
 sg13g2_inv_2 _12709_ (.Y(_06909_),
    .A(net4018));
 sg13g2_inv_1 _12710_ (.Y(_06910_),
    .A(\fpga_top.cpu_top.csr_mepc_ex[17] ));
 sg13g2_inv_2 _12711_ (.Y(_06911_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[17] ));
 sg13g2_inv_1 _12712_ (.Y(_06912_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[18] ));
 sg13g2_inv_1 _12713_ (.Y(_06913_),
    .A(net3829));
 sg13g2_inv_1 _12714_ (.Y(_06914_),
    .A(net1606));
 sg13g2_inv_1 _12715_ (.Y(_06915_),
    .A(net1801));
 sg13g2_inv_1 _12716_ (.Y(_06916_),
    .A(net1625));
 sg13g2_inv_2 _12717_ (.Y(_06917_),
    .A(net3843));
 sg13g2_inv_2 _12718_ (.Y(_06918_),
    .A(net3612));
 sg13g2_inv_1 _12719_ (.Y(_06919_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[27] ));
 sg13g2_inv_1 _12720_ (.Y(_06920_),
    .A(\fpga_top.cpu_top.csr_mepc_ex[30] ));
 sg13g2_inv_1 _12721_ (.Y(_06921_),
    .A(net1788));
 sg13g2_inv_1 _12722_ (.Y(_06922_),
    .A(\fpga_top.cpu_top.csr_mepc_ex[31] ));
 sg13g2_inv_2 _12723_ (.Y(_06923_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[31] ));
 sg13g2_inv_2 _12724_ (.Y(_06924_),
    .A(net6));
 sg13g2_inv_4 _12725_ (.A(net5436),
    .Y(_06925_));
 sg13g2_inv_1 _12726_ (.Y(_06926_),
    .A(\fpga_top.io_spi_lite.sel_sck[1] ));
 sg13g2_inv_1 _12727_ (.Y(_06927_),
    .A(\fpga_top.io_spi_lite.sel_sck[3] ));
 sg13g2_inv_2 _12728_ (.Y(_06928_),
    .A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[2] ));
 sg13g2_inv_1 _12729_ (.Y(_06929_),
    .A(net6597));
 sg13g2_inv_1 _12730_ (.Y(_06930_),
    .A(_00088_));
 sg13g2_inv_4 _12731_ (.A(_00091_),
    .Y(uo_out[1]));
 sg13g2_inv_4 _12732_ (.A(_00092_),
    .Y(uo_out[2]));
 sg13g2_inv_4 _12733_ (.A(_00093_),
    .Y(uo_out[3]));
 sg13g2_nor2b_1 _12734_ (.A(net1620),
    .B_N(net3682),
    .Y(_06931_));
 sg13g2_nand2b_1 _12735_ (.Y(_06932_),
    .B(net2105),
    .A_N(net1620));
 sg13g2_nor2b_2 _12736_ (.A(net6306),
    .B_N(net1807),
    .Y(_06933_));
 sg13g2_nand2b_1 _12737_ (.Y(_06934_),
    .B(\fpga_top.qspi_if.inner_state[0] ),
    .A_N(\fpga_top.qspi_if.inner_state[1] ));
 sg13g2_nor2b_1 _12738_ (.A(net1807),
    .B_N(net6306),
    .Y(_06935_));
 sg13g2_nand2b_2 _12739_ (.Y(_06936_),
    .B(\fpga_top.qspi_if.inner_state[1] ),
    .A_N(\fpga_top.qspi_if.inner_state[0] ));
 sg13g2_nor2_1 _12740_ (.A(_06933_),
    .B(net5346),
    .Y(_06937_));
 sg13g2_nand2_2 _12741_ (.Y(_06938_),
    .A(net5348),
    .B(_06936_));
 sg13g2_a21oi_1 _12742_ (.A1(net5353),
    .A2(_06938_),
    .Y(_06939_),
    .B1(_00125_));
 sg13g2_nor2_1 _12743_ (.A(net3079),
    .B(net6153),
    .Y(_06940_));
 sg13g2_a21oi_1 _12744_ (.A1(_06660_),
    .A2(\fpga_top.qspi_if.dbg_2div_trt ),
    .Y(_06941_),
    .B1(_06940_));
 sg13g2_nand2b_1 _12745_ (.Y(_06942_),
    .B(net5355),
    .A_N(\fpga_top.qspi_if.rst_cntr[0] ));
 sg13g2_nor4_2 _12746_ (.A(net3524),
    .B(net3589),
    .C(net3788),
    .Y(_06943_),
    .D(_06942_));
 sg13g2_or2_1 _12747_ (.X(_06944_),
    .B(_06942_),
    .A(net3524));
 sg13g2_a221oi_1 _12748_ (.B2(net1400),
    .C1(_06939_),
    .B1(_06943_),
    .A1(net5354),
    .Y(_00145_),
    .A2(_06941_));
 sg13g2_a21oi_1 _12749_ (.A1(\fpga_top.qspi_if.dbg_2div_cew_pre ),
    .A2(\fpga_top.qspi_if.dbg_2div_cew_lat ),
    .Y(_06945_),
    .B1(net3926));
 sg13g2_nand4_1 _12750_ (.B(net3975),
    .C(_06940_),
    .A(_06813_),
    .Y(_06946_),
    .D(_06945_));
 sg13g2_nor2b_2 _12751_ (.A(\fpga_top.qspi_if.word_adr[24] ),
    .B_N(\fpga_top.qspi_if.word_adr[25] ),
    .Y(_06947_));
 sg13g2_nand2b_2 _12752_ (.Y(_06948_),
    .B(_06947_),
    .A_N(_06946_));
 sg13g2_inv_4 _12753_ (.A(_06948_),
    .Y(_00134_));
 sg13g2_nor2b_2 _12754_ (.A(net6262),
    .B_N(net6529),
    .Y(_06949_));
 sg13g2_nand2b_2 _12755_ (.Y(_06950_),
    .B(_06949_),
    .A_N(_06946_));
 sg13g2_inv_2 _12756_ (.Y(_00133_),
    .A(_06950_));
 sg13g2_nor3_1 _12757_ (.A(\fpga_top.qspi_if.word_adr[24] ),
    .B(net6262),
    .C(_06946_),
    .Y(_00132_));
 sg13g2_nor2_1 _12758_ (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[3] ),
    .B(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ),
    .Y(_06951_));
 sg13g2_nor3_1 _12759_ (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ),
    .B(net6586),
    .C(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ),
    .Y(_06952_));
 sg13g2_nand2b_1 _12760_ (.Y(_06953_),
    .B(_06951_),
    .A_N(net6467));
 sg13g2_nor2_2 _12761_ (.A(net5632),
    .B(net5630),
    .Y(_06954_));
 sg13g2_nand2_2 _12762_ (.Y(_06955_),
    .A(_06952_),
    .B(_06954_));
 sg13g2_nor2b_1 _12763_ (.A(\fpga_top.uart_top.uart_rec_char.pdata[7] ),
    .B_N(\fpga_top.uart_top.uart_rec_char.pdata[5] ),
    .Y(_06956_));
 sg13g2_nand3_1 _12764_ (.B(\fpga_top.uart_top.uart_rec_char.pdata[6] ),
    .C(_06956_),
    .A(_06544_),
    .Y(_06957_));
 sg13g2_nand3_1 _12765_ (.B(\fpga_top.uart_top.uart_rec_char.data_en ),
    .C(_06956_),
    .A(\fpga_top.uart_top.uart_rec_char.pdata[6] ),
    .Y(_06958_));
 sg13g2_nor2_1 _12766_ (.A(\fpga_top.uart_top.uart_rec_char.pdata[4] ),
    .B(_06958_),
    .Y(_06959_));
 sg13g2_nand2_1 _12767_ (.Y(_06960_),
    .A(_06543_),
    .B(net5626));
 sg13g2_nor2_1 _12768_ (.A(net5628),
    .B(_06542_),
    .Y(_06961_));
 sg13g2_nor2b_1 _12769_ (.A(_06960_),
    .B_N(_06961_),
    .Y(_06962_));
 sg13g2_nand2_1 _12770_ (.Y(_06963_),
    .A(net5628),
    .B(\fpga_top.uart_top.uart_rec_char.pdata[0] ));
 sg13g2_inv_1 _12771_ (.Y(_06964_),
    .A(_06963_));
 sg13g2_nor3_1 _12772_ (.A(\fpga_top.uart_top.uart_rec_char.pdata[2] ),
    .B(net5626),
    .C(_06963_),
    .Y(_06965_));
 sg13g2_or3_1 _12773_ (.A(net5627),
    .B(net5625),
    .C(_06963_),
    .X(_06966_));
 sg13g2_nor2_2 _12774_ (.A(_06544_),
    .B(_06958_),
    .Y(_06967_));
 sg13g2_a22oi_1 _12775_ (.Y(_06968_),
    .B1(_06965_),
    .B2(_06967_),
    .A2(_06962_),
    .A1(_06959_));
 sg13g2_nor3_1 _12776_ (.A(_06543_),
    .B(net5626),
    .C(_06963_),
    .Y(_06969_));
 sg13g2_nor2b_1 _12777_ (.A(_06958_),
    .B_N(_06969_),
    .Y(_06970_));
 sg13g2_nand2_1 _12778_ (.Y(_06971_),
    .A(net5628),
    .B(_06542_));
 sg13g2_nor2_1 _12779_ (.A(_06960_),
    .B(_06971_),
    .Y(_06972_));
 sg13g2_or2_1 _12780_ (.X(_06973_),
    .B(_06971_),
    .A(_06960_));
 sg13g2_and2_1 _12781_ (.A(_06959_),
    .B(_06972_),
    .X(_06974_));
 sg13g2_nor3_1 _12782_ (.A(net5627),
    .B(net5625),
    .C(_06971_),
    .Y(_06975_));
 sg13g2_a21oi_1 _12783_ (.A1(_06967_),
    .A2(_06975_),
    .Y(_06976_),
    .B1(_06974_));
 sg13g2_nor2_1 _12784_ (.A(net5628),
    .B(\fpga_top.uart_top.uart_rec_char.pdata[0] ),
    .Y(_06977_));
 sg13g2_nand2_1 _12785_ (.Y(_06978_),
    .A(net5627),
    .B(_06977_));
 sg13g2_and4_1 _12786_ (.A(net5627),
    .B(net5625),
    .C(_06959_),
    .D(_06977_),
    .X(_06979_));
 sg13g2_nor2_1 _12787_ (.A(net5625),
    .B(_06978_),
    .Y(_06980_));
 sg13g2_a21oi_1 _12788_ (.A1(_06967_),
    .A2(_06980_),
    .Y(_06981_),
    .B1(_06979_));
 sg13g2_nand3_1 _12789_ (.B(_06976_),
    .C(_06981_),
    .A(_06968_),
    .Y(_06982_));
 sg13g2_nor2_1 _12790_ (.A(_06970_),
    .B(_06982_),
    .Y(_06983_));
 sg13g2_nand2b_1 _12791_ (.Y(_06984_),
    .B(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.cmd_status[3] ));
 sg13g2_nor2_1 _12792_ (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ),
    .B(_06984_),
    .Y(_06985_));
 sg13g2_or2_1 _12793_ (.X(_06986_),
    .B(_06984_),
    .A(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ));
 sg13g2_nand2_2 _12794_ (.Y(_06987_),
    .A(\fpga_top.uart_top.uart_rec_char.cmd_status[0] ),
    .B(net5631));
 sg13g2_nor2_1 _12795_ (.A(_06986_),
    .B(_06987_),
    .Y(_06988_));
 sg13g2_nor2b_2 _12796_ (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ),
    .B_N(\fpga_top.uart_top.uart_rec_char.cmd_status[3] ),
    .Y(_06989_));
 sg13g2_nand2_2 _12797_ (.Y(_06990_),
    .A(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ),
    .B(_06989_));
 sg13g2_nor2_1 _12798_ (.A(_06987_),
    .B(_06990_),
    .Y(_06991_));
 sg13g2_or2_1 _12799_ (.X(_06992_),
    .B(_06990_),
    .A(_06987_));
 sg13g2_nor3_1 _12800_ (.A(\fpga_top.uart_top.uart_rec_char.pdata[5] ),
    .B(\fpga_top.uart_top.uart_rec_char.pdata[6] ),
    .C(\fpga_top.uart_top.uart_rec_char.pdata[7] ),
    .Y(_06993_));
 sg13g2_nand3_1 _12801_ (.B(\fpga_top.uart_top.uart_rec_char.data_en ),
    .C(_06993_),
    .A(_06544_),
    .Y(_06994_));
 sg13g2_inv_1 _12802_ (.Y(_06995_),
    .A(_06994_));
 sg13g2_nor2_1 _12803_ (.A(_06966_),
    .B(_06994_),
    .Y(_06996_));
 sg13g2_nor2_1 _12804_ (.A(\fpga_top.uart_top.uart_logics.status_dump[1] ),
    .B(\fpga_top.uart_top.uart_logics.status_dump[0] ),
    .Y(_06997_));
 sg13g2_nor3_2 _12805_ (.A(\fpga_top.uart_top.uart_logics.status_dump[2] ),
    .B(net1851),
    .C(net6458),
    .Y(_06998_));
 sg13g2_nor2_1 _12806_ (.A(net5228),
    .B(_06998_),
    .Y(_06999_));
 sg13g2_o21ai_1 _12807_ (.B1(_06999_),
    .Y(_07000_),
    .A1(_06988_),
    .A2(net5235));
 sg13g2_nor2_1 _12808_ (.A(net5633),
    .B(net5227),
    .Y(_07001_));
 sg13g2_nand3_1 _12809_ (.B(net5630),
    .C(_06952_),
    .A(net5632),
    .Y(_07002_));
 sg13g2_inv_1 _12810_ (.Y(_07003_),
    .A(_07002_));
 sg13g2_nor2b_2 _12811_ (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ),
    .B_N(_06989_),
    .Y(_07004_));
 sg13g2_nand2b_2 _12812_ (.Y(_07005_),
    .B(_06989_),
    .A_N(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ));
 sg13g2_nor2_1 _12813_ (.A(_06987_),
    .B(_07005_),
    .Y(_07006_));
 sg13g2_nor3_1 _12814_ (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ),
    .B(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ),
    .C(_06987_),
    .Y(_07007_));
 sg13g2_nand2_2 _12815_ (.Y(_07008_),
    .A(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ),
    .B(_06951_));
 sg13g2_nor2_2 _12816_ (.A(_06987_),
    .B(_07008_),
    .Y(_07009_));
 sg13g2_o21ai_1 _12817_ (.B1(_07001_),
    .Y(_07010_),
    .A1(_07007_),
    .A2(_07009_));
 sg13g2_nand2_1 _12818_ (.Y(_07011_),
    .A(_07000_),
    .B(_07010_));
 sg13g2_nor2b_1 _12819_ (.A(net5630),
    .B_N(net5632),
    .Y(_07012_));
 sg13g2_nand2b_1 _12820_ (.Y(_07013_),
    .B(net5632),
    .A_N(net5630));
 sg13g2_nand2_1 _12821_ (.Y(_07014_),
    .A(_06986_),
    .B(_07008_));
 sg13g2_nand3_1 _12822_ (.B(_06989_),
    .C(_07012_),
    .A(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ),
    .Y(_07015_));
 sg13g2_o21ai_1 _12823_ (.B1(_07012_),
    .Y(_07016_),
    .A1(_06951_),
    .A2(_06985_));
 sg13g2_nand2_1 _12824_ (.Y(_07017_),
    .A(_07015_),
    .B(_07016_));
 sg13g2_nor2_2 _12825_ (.A(_07005_),
    .B(_07013_),
    .Y(_07018_));
 sg13g2_nor2_1 _12826_ (.A(_07017_),
    .B(_07018_),
    .Y(_07019_));
 sg13g2_or2_1 _12827_ (.X(_07020_),
    .B(_07018_),
    .A(_07017_));
 sg13g2_nor2b_1 _12828_ (.A(net5632),
    .B_N(net5630),
    .Y(_07021_));
 sg13g2_nand2b_2 _12829_ (.Y(_07022_),
    .B(net5631),
    .A_N(net5632));
 sg13g2_nor2_1 _12830_ (.A(_06986_),
    .B(_07022_),
    .Y(_07023_));
 sg13g2_a21oi_1 _12831_ (.A1(_06986_),
    .A2(_07005_),
    .Y(_07024_),
    .B1(_07022_));
 sg13g2_nor2_1 _12832_ (.A(_06546_),
    .B(net5227),
    .Y(_07025_));
 sg13g2_a221oi_1 _12833_ (.B2(_07025_),
    .C1(_07011_),
    .B1(_07024_),
    .A1(_07001_),
    .Y(_07026_),
    .A2(_07020_));
 sg13g2_o21ai_1 _12834_ (.B1(_07026_),
    .Y(\fpga_top.uart_top.uart_rec_char.next_cmd_status[0] ),
    .A1(_06955_),
    .A2(_06983_));
 sg13g2_inv_1 _12835_ (.Y(_07027_),
    .A(\fpga_top.uart_top.uart_rec_char.next_cmd_status[0] ));
 sg13g2_nand2b_2 _12836_ (.Y(_07028_),
    .B(\fpga_top.cpu_top.decoder.illegal_ops_inst[4] ),
    .A_N(\fpga_top.cpu_top.decoder.illegal_ops_inst[3] ));
 sg13g2_nand3b_1 _12837_ (.B(net5585),
    .C(\fpga_top.cpu_top.decoder.illegal_ops_inst[4] ),
    .Y(_07029_),
    .A_N(\fpga_top.cpu_top.decoder.illegal_ops_inst[3] ));
 sg13g2_nand3b_1 _12838_ (.B(net3864),
    .C(net3922),
    .Y(_07030_),
    .A_N(net3806));
 sg13g2_nand2b_1 _12839_ (.Y(_07031_),
    .B(_06550_),
    .A_N(net5344));
 sg13g2_nor3_2 _12840_ (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[5] ),
    .B(_07029_),
    .C(net5344),
    .Y(_07032_));
 sg13g2_or2_1 _12841_ (.X(_07033_),
    .B(_07031_),
    .A(_07029_));
 sg13g2_nor2_2 _12842_ (.A(net5569),
    .B(net5314),
    .Y(_07034_));
 sg13g2_a21oi_1 _12843_ (.A1(_06557_),
    .A2(net5313),
    .Y(_07035_),
    .B1(net5220));
 sg13g2_nor2_1 _12844_ (.A(net5582),
    .B(net5583),
    .Y(_07036_));
 sg13g2_nor3_2 _12845_ (.A(net5581),
    .B(net5583),
    .C(net5575),
    .Y(_07037_));
 sg13g2_or3_1 _12846_ (.A(net5581),
    .B(net5584),
    .C(net5577),
    .X(_07038_));
 sg13g2_nand4_1 _12847_ (.B(\fpga_top.cpu_top.decoder.illegal_ops_inst[6] ),
    .C(\fpga_top.cpu_top.decoder.illegal_ops_inst[0] ),
    .A(\fpga_top.cpu_top.decoder.illegal_ops_inst[5] ),
    .Y(_07039_),
    .D(\fpga_top.cpu_top.decoder.illegal_ops_inst[1] ));
 sg13g2_nand2b_1 _12848_ (.Y(_07040_),
    .B(net5585),
    .A_N(\fpga_top.cpu_top.decoder.illegal_ops_inst[4] ));
 sg13g2_nor4_2 _12849_ (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[3] ),
    .B(_07038_),
    .C(_07039_),
    .Y(_07041_),
    .D(_07040_));
 sg13g2_or4_1 _12850_ (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[3] ),
    .B(_07038_),
    .C(_07039_),
    .D(_07040_),
    .X(_07042_));
 sg13g2_nand2_1 _12851_ (.Y(_07043_),
    .A(net5756),
    .B(net5304));
 sg13g2_o21ai_1 _12852_ (.B1(_07043_),
    .Y(_07044_),
    .A1(_06643_),
    .A2(net5304));
 sg13g2_and2_1 _12853_ (.A(_07035_),
    .B(_07044_),
    .X(_07045_));
 sg13g2_xor2_1 _12854_ (.B(_07044_),
    .A(_07035_),
    .X(_07046_));
 sg13g2_a21oi_1 _12855_ (.A1(_06556_),
    .A2(net5312),
    .Y(_07047_),
    .B1(net5220));
 sg13g2_nand2_1 _12856_ (.Y(_07048_),
    .A(net5759),
    .B(net5305));
 sg13g2_o21ai_1 _12857_ (.B1(_07048_),
    .Y(_07049_),
    .A1(_06641_),
    .A2(net5305));
 sg13g2_nor2_1 _12858_ (.A(_07047_),
    .B(_07049_),
    .Y(_07050_));
 sg13g2_a21oi_1 _12859_ (.A1(_06555_),
    .A2(net5310),
    .Y(_07051_),
    .B1(_07034_));
 sg13g2_nand2_1 _12860_ (.Y(_07052_),
    .A(net5590),
    .B(net5299));
 sg13g2_o21ai_1 _12861_ (.B1(_07052_),
    .Y(_07053_),
    .A1(_06580_),
    .A2(net5299));
 sg13g2_nand2_1 _12862_ (.Y(_07054_),
    .A(_07051_),
    .B(_07053_));
 sg13g2_xor2_1 _12863_ (.B(_07053_),
    .A(_07051_),
    .X(_07055_));
 sg13g2_inv_1 _12864_ (.Y(_07056_),
    .A(_07055_));
 sg13g2_a21oi_1 _12865_ (.A1(_06554_),
    .A2(net5310),
    .Y(_07057_),
    .B1(net5220));
 sg13g2_nand2_1 _12866_ (.Y(_07058_),
    .A(net5763),
    .B(net5305));
 sg13g2_o21ai_1 _12867_ (.B1(_07058_),
    .Y(_07059_),
    .A1(_06636_),
    .A2(net5305));
 sg13g2_nor2_1 _12868_ (.A(_07057_),
    .B(_07059_),
    .Y(_07060_));
 sg13g2_nand2_1 _12869_ (.Y(_07061_),
    .A(net5801),
    .B(net5301));
 sg13g2_o21ai_1 _12870_ (.B1(_07061_),
    .Y(_07062_),
    .A1(_06592_),
    .A2(net5303));
 sg13g2_and3_1 _12871_ (.X(_07063_),
    .A(net5570),
    .B(net5222),
    .C(_07062_));
 sg13g2_a21o_1 _12872_ (.A2(net5222),
    .A1(net5570),
    .B1(_07062_),
    .X(_07064_));
 sg13g2_nand2b_1 _12873_ (.Y(_07065_),
    .B(_07064_),
    .A_N(_07063_));
 sg13g2_nor2_1 _12874_ (.A(_06554_),
    .B(net5307),
    .Y(_07066_));
 sg13g2_nor2_1 _12875_ (.A(net5805),
    .B(net5297),
    .Y(_07067_));
 sg13g2_a21oi_1 _12876_ (.A1(_06590_),
    .A2(net5297),
    .Y(_07068_),
    .B1(_07067_));
 sg13g2_nand2_1 _12877_ (.Y(_07069_),
    .A(_07066_),
    .B(_07068_));
 sg13g2_nor2_1 _12878_ (.A(_06549_),
    .B(net5307),
    .Y(_07070_));
 sg13g2_nand2_1 _12879_ (.Y(_07071_),
    .A(net5809),
    .B(net5301));
 sg13g2_o21ai_1 _12880_ (.B1(_07071_),
    .Y(_07072_),
    .A1(_06588_),
    .A2(net5301));
 sg13g2_and2_1 _12881_ (.A(_07070_),
    .B(_07072_),
    .X(_07073_));
 sg13g2_nand2_1 _12882_ (.Y(_07074_),
    .A(net5812),
    .B(net5301));
 sg13g2_o21ai_1 _12883_ (.B1(_07074_),
    .Y(_07075_),
    .A1(_06587_),
    .A2(net5301));
 sg13g2_nand3_1 _12884_ (.B(net5221),
    .C(_07075_),
    .A(\fpga_top.cpu_top.br_ofs[5] ),
    .Y(_07076_));
 sg13g2_a21o_1 _12885_ (.A2(net5221),
    .A1(\fpga_top.cpu_top.br_ofs[5] ),
    .B1(_07075_),
    .X(_07077_));
 sg13g2_nand3b_1 _12886_ (.B(\fpga_top.cpu_top.decoder.illegal_ops_inst[3] ),
    .C(net5585),
    .Y(_07078_),
    .A_N(\fpga_top.cpu_top.decoder.illegal_ops_inst[4] ));
 sg13g2_nor2_2 _12887_ (.A(_07039_),
    .B(_07078_),
    .Y(_07079_));
 sg13g2_or2_1 _12888_ (.X(_07080_),
    .B(_07078_),
    .A(_07039_));
 sg13g2_nor2_1 _12889_ (.A(net5303),
    .B(_07079_),
    .Y(_07081_));
 sg13g2_nand2_2 _12890_ (.Y(_07082_),
    .A(net5298),
    .B(net5295));
 sg13g2_o21ai_1 _12891_ (.B1(net5221),
    .Y(_07083_),
    .A1(\fpga_top.cpu_top.alui_shamt[4] ),
    .A2(net5219));
 sg13g2_a21oi_1 _12892_ (.A1(_06576_),
    .A2(net5219),
    .Y(_07084_),
    .B1(_07083_));
 sg13g2_mux2_1 _12893_ (.A0(net5815),
    .A1(net5597),
    .S(net5297),
    .X(_07085_));
 sg13g2_nand2_1 _12894_ (.Y(_07086_),
    .A(_07084_),
    .B(_07085_));
 sg13g2_o21ai_1 _12895_ (.B1(net5221),
    .Y(_07087_),
    .A1(\fpga_top.cpu_top.alui_shamt[3] ),
    .A2(net5219));
 sg13g2_a21oi_1 _12896_ (.A1(_06569_),
    .A2(net5219),
    .Y(_07088_),
    .B1(_07087_));
 sg13g2_nor2_1 _12897_ (.A(net5818),
    .B(net5297),
    .Y(_07089_));
 sg13g2_a21oi_1 _12898_ (.A1(_06584_),
    .A2(net5298),
    .Y(_07090_),
    .B1(_07089_));
 sg13g2_and2_1 _12899_ (.A(_07088_),
    .B(_07090_),
    .X(_07091_));
 sg13g2_nor3_1 _12900_ (.A(\fpga_top.cpu_top.br_ofs[2] ),
    .B(net5301),
    .C(_07079_),
    .Y(_07092_));
 sg13g2_a21oi_1 _12901_ (.A1(net5297),
    .A2(net5295),
    .Y(_07093_),
    .B1(\fpga_top.cpu_top.alui_shamt[2] ));
 sg13g2_nor3_1 _12902_ (.A(net5308),
    .B(_07092_),
    .C(_07093_),
    .Y(_07094_));
 sg13g2_nor2_1 _12903_ (.A(net5821),
    .B(net5298),
    .Y(_07095_));
 sg13g2_a21oi_1 _12904_ (.A1(net5386),
    .A2(net5298),
    .Y(_07096_),
    .B1(_07095_));
 sg13g2_and2_1 _12905_ (.A(_07094_),
    .B(_07096_),
    .X(_07097_));
 sg13g2_xor2_1 _12906_ (.B(_07096_),
    .A(_07094_),
    .X(_07098_));
 sg13g2_o21ai_1 _12907_ (.B1(_06559_),
    .Y(_07099_),
    .A1(net5301),
    .A2(_07079_));
 sg13g2_nand3_1 _12908_ (.B(net5297),
    .C(net5295),
    .A(_06560_),
    .Y(_07100_));
 sg13g2_nand3_1 _12909_ (.B(_07099_),
    .C(_07100_),
    .A(net5223),
    .Y(_07101_));
 sg13g2_nand3_1 _12910_ (.B(net5572),
    .C(net5825),
    .A(net5824),
    .Y(_07102_));
 sg13g2_a21oi_1 _12911_ (.A1(net5572),
    .A2(net5825),
    .Y(_07103_),
    .B1(net5824));
 sg13g2_nand2b_1 _12912_ (.Y(_07104_),
    .B(net5301),
    .A_N(_07103_));
 sg13g2_a21oi_1 _12913_ (.A1(_07101_),
    .A2(_07102_),
    .Y(_07105_),
    .B1(_07104_));
 sg13g2_a21o_1 _12914_ (.A2(_07105_),
    .A1(_07098_),
    .B1(_07097_),
    .X(_07106_));
 sg13g2_or2_1 _12915_ (.X(_07107_),
    .B(_07090_),
    .A(_07088_));
 sg13g2_nand2b_1 _12916_ (.Y(_07108_),
    .B(_07107_),
    .A_N(_07091_));
 sg13g2_a21o_2 _12917_ (.A2(_07107_),
    .A1(_07106_),
    .B1(_07091_),
    .X(_07109_));
 sg13g2_xor2_1 _12918_ (.B(_07085_),
    .A(_07084_),
    .X(_07110_));
 sg13g2_nand2_1 _12919_ (.Y(_07111_),
    .A(_07109_),
    .B(_07110_));
 sg13g2_nand2_1 _12920_ (.Y(_07112_),
    .A(_07086_),
    .B(_07111_));
 sg13g2_nand2_1 _12921_ (.Y(_07113_),
    .A(_07076_),
    .B(_07086_));
 sg13g2_a21o_1 _12922_ (.A2(_07110_),
    .A1(_07109_),
    .B1(_07113_),
    .X(_07114_));
 sg13g2_and2_1 _12923_ (.A(_07077_),
    .B(_07114_),
    .X(_07115_));
 sg13g2_xnor2_1 _12924_ (.Y(_07116_),
    .A(_07070_),
    .B(_07072_));
 sg13g2_inv_1 _12925_ (.Y(_07117_),
    .A(_07116_));
 sg13g2_a21oi_1 _12926_ (.A1(_07115_),
    .A2(_07117_),
    .Y(_07118_),
    .B1(_07073_));
 sg13g2_o21ai_1 _12927_ (.B1(_07073_),
    .Y(_07119_),
    .A1(_07066_),
    .A2(_07068_));
 sg13g2_xor2_1 _12928_ (.B(_07068_),
    .A(_07066_),
    .X(_07120_));
 sg13g2_nand4_1 _12929_ (.B(_07114_),
    .C(_07117_),
    .A(_07077_),
    .Y(_07121_),
    .D(_07120_));
 sg13g2_nand3_1 _12930_ (.B(_07119_),
    .C(_07121_),
    .A(_07069_),
    .Y(_07122_));
 sg13g2_nor2_1 _12931_ (.A(_06555_),
    .B(net5309),
    .Y(_07123_));
 sg13g2_nand2_1 _12932_ (.Y(_07124_),
    .A(net5595),
    .B(net5297));
 sg13g2_o21ai_1 _12933_ (.B1(_07124_),
    .Y(_07125_),
    .A1(_06566_),
    .A2(net5298));
 sg13g2_and2_1 _12934_ (.A(_07123_),
    .B(_07125_),
    .X(_07126_));
 sg13g2_xnor2_1 _12935_ (.Y(_07127_),
    .A(_07123_),
    .B(_07125_));
 sg13g2_inv_1 _12936_ (.Y(_07128_),
    .A(_07127_));
 sg13g2_nand3b_1 _12937_ (.B(_07122_),
    .C(_07128_),
    .Y(_07129_),
    .A_N(_07065_));
 sg13g2_nor2_1 _12938_ (.A(_06557_),
    .B(net5309),
    .Y(_07130_));
 sg13g2_nand2_1 _12939_ (.Y(_07131_),
    .A(net5798),
    .B(net5302));
 sg13g2_o21ai_1 _12940_ (.B1(_07131_),
    .Y(_07132_),
    .A1(_06594_),
    .A2(net5303));
 sg13g2_nand2_1 _12941_ (.Y(_07133_),
    .A(_07130_),
    .B(_07132_));
 sg13g2_nor2_1 _12942_ (.A(net5569),
    .B(net5300),
    .Y(_07134_));
 sg13g2_a21oi_1 _12943_ (.A1(_06564_),
    .A2(net5300),
    .Y(_07135_),
    .B1(_07134_));
 sg13g2_a21oi_1 _12944_ (.A1(_06563_),
    .A2(_07079_),
    .Y(_07136_),
    .B1(net5308));
 sg13g2_o21ai_1 _12945_ (.B1(_07136_),
    .Y(_07137_),
    .A1(_07079_),
    .A2(_07135_));
 sg13g2_nand2_1 _12946_ (.Y(_07138_),
    .A(_06597_),
    .B(net5297));
 sg13g2_o21ai_1 _12947_ (.B1(_07138_),
    .Y(_07139_),
    .A1(net5797),
    .A2(net5298));
 sg13g2_a21oi_1 _12948_ (.A1(_07137_),
    .A2(_07139_),
    .Y(_07140_),
    .B1(_07133_));
 sg13g2_or2_1 _12949_ (.X(_07141_),
    .B(_07139_),
    .A(_07137_));
 sg13g2_a21oi_1 _12950_ (.A1(_07064_),
    .A2(_07126_),
    .Y(_07142_),
    .B1(_07063_));
 sg13g2_nor2b_1 _12951_ (.A(_07140_),
    .B_N(_07141_),
    .Y(_07143_));
 sg13g2_xnor2_1 _12952_ (.Y(_07144_),
    .A(_07130_),
    .B(_07132_));
 sg13g2_xor2_1 _12953_ (.B(_07139_),
    .A(_07137_),
    .X(_07145_));
 sg13g2_nand2b_1 _12954_ (.Y(_07146_),
    .B(_07145_),
    .A_N(_07144_));
 sg13g2_o21ai_1 _12955_ (.B1(_07143_),
    .Y(_07147_),
    .A1(_07142_),
    .A2(_07146_));
 sg13g2_nor3_1 _12956_ (.A(_07065_),
    .B(_07127_),
    .C(_07146_),
    .Y(_07148_));
 sg13g2_a21oi_2 _12957_ (.B1(_07147_),
    .Y(_07149_),
    .A2(_07148_),
    .A1(_07122_));
 sg13g2_nor3_2 _12958_ (.A(net5569),
    .B(net5309),
    .C(_07079_),
    .Y(_07150_));
 sg13g2_a21oi_1 _12959_ (.A1(net5222),
    .A2(net5295),
    .Y(_07151_),
    .B1(net5576));
 sg13g2_nor2_1 _12960_ (.A(_07150_),
    .B(_07151_),
    .Y(_07152_));
 sg13g2_nand2_1 _12961_ (.Y(_07153_),
    .A(net5790),
    .B(net5302));
 sg13g2_o21ai_1 _12962_ (.B1(_07153_),
    .Y(_07154_),
    .A1(_06603_),
    .A2(net5302));
 sg13g2_nand2_1 _12963_ (.Y(_07155_),
    .A(_07152_),
    .B(_07154_));
 sg13g2_xor2_1 _12964_ (.B(_07154_),
    .A(_07152_),
    .X(_07156_));
 sg13g2_inv_1 _12965_ (.Y(_07157_),
    .A(_07156_));
 sg13g2_a21oi_1 _12966_ (.A1(net5222),
    .A2(net5295),
    .Y(_07158_),
    .B1(\fpga_top.cpu_top.csr_uimm[0] ));
 sg13g2_nor2_1 _12967_ (.A(_07150_),
    .B(_07158_),
    .Y(_07159_));
 sg13g2_nand2_1 _12968_ (.Y(_07160_),
    .A(net5789),
    .B(net5302));
 sg13g2_o21ai_1 _12969_ (.B1(_07160_),
    .Y(_07161_),
    .A1(_06605_),
    .A2(net5302));
 sg13g2_nor2_1 _12970_ (.A(_07159_),
    .B(_07161_),
    .Y(_07162_));
 sg13g2_xor2_1 _12971_ (.B(_07161_),
    .A(_07159_),
    .X(_07163_));
 sg13g2_and2_1 _12972_ (.A(_07156_),
    .B(_07163_),
    .X(_07164_));
 sg13g2_a21oi_1 _12973_ (.A1(net5222),
    .A2(net5295),
    .Y(_07165_),
    .B1(net5582));
 sg13g2_nor2_1 _12974_ (.A(_07150_),
    .B(_07165_),
    .Y(_07166_));
 sg13g2_nand2_1 _12975_ (.Y(_07167_),
    .A(net5792),
    .B(net5302));
 sg13g2_o21ai_1 _12976_ (.B1(_07167_),
    .Y(_07168_),
    .A1(_06601_),
    .A2(net5302));
 sg13g2_nand2_1 _12977_ (.Y(_07169_),
    .A(_07166_),
    .B(_07168_));
 sg13g2_nor2_1 _12978_ (.A(_07166_),
    .B(_07168_),
    .Y(_07170_));
 sg13g2_xor2_1 _12979_ (.B(_07168_),
    .A(_07166_),
    .X(_07171_));
 sg13g2_a21oi_1 _12980_ (.A1(net5223),
    .A2(net5295),
    .Y(_07172_),
    .B1(net5583));
 sg13g2_nor2_1 _12981_ (.A(_07150_),
    .B(_07172_),
    .Y(_07173_));
 sg13g2_nand2_1 _12982_ (.Y(_07174_),
    .A(net5795),
    .B(net5302));
 sg13g2_o21ai_1 _12983_ (.B1(_07174_),
    .Y(_07175_),
    .A1(_06599_),
    .A2(net5303));
 sg13g2_nand2_1 _12984_ (.Y(_07176_),
    .A(_07173_),
    .B(_07175_));
 sg13g2_xor2_1 _12985_ (.B(_07175_),
    .A(_07173_),
    .X(_07177_));
 sg13g2_inv_1 _12986_ (.Y(_07178_),
    .A(_07177_));
 sg13g2_nand3_1 _12987_ (.B(_07171_),
    .C(_07177_),
    .A(_07164_),
    .Y(_07179_));
 sg13g2_o21ai_1 _12988_ (.B1(_07169_),
    .Y(_07180_),
    .A1(_07170_),
    .A2(_07176_));
 sg13g2_nor2_1 _12989_ (.A(_07155_),
    .B(_07162_),
    .Y(_07181_));
 sg13g2_a221oi_1 _12990_ (.B2(_07180_),
    .C1(_07181_),
    .B1(_07164_),
    .A1(_07159_),
    .Y(_07182_),
    .A2(_07161_));
 sg13g2_o21ai_1 _12991_ (.B1(_07182_),
    .Y(_07183_),
    .A1(_07149_),
    .A2(_07179_));
 sg13g2_a21oi_1 _12992_ (.A1(_06548_),
    .A2(net5310),
    .Y(_07184_),
    .B1(net5220));
 sg13g2_nand2_1 _12993_ (.Y(_07185_),
    .A(net5591),
    .B(net5300));
 sg13g2_o21ai_1 _12994_ (.B1(_07185_),
    .Y(_07186_),
    .A1(_06579_),
    .A2(net5299));
 sg13g2_nand2_1 _12995_ (.Y(_07187_),
    .A(_07184_),
    .B(_07186_));
 sg13g2_xor2_1 _12996_ (.B(_07186_),
    .A(_07184_),
    .X(_07188_));
 sg13g2_inv_1 _12997_ (.Y(_07189_),
    .A(_07188_));
 sg13g2_a21oi_1 _12998_ (.A1(_06568_),
    .A2(net5310),
    .Y(_07190_),
    .B1(_07034_));
 sg13g2_nand2_1 _12999_ (.Y(_07191_),
    .A(net5773),
    .B(net5305));
 sg13g2_o21ai_1 _13000_ (.B1(_07191_),
    .Y(_07192_),
    .A1(_06626_),
    .A2(net5305));
 sg13g2_nor2_1 _13001_ (.A(_07190_),
    .B(_07192_),
    .Y(_07193_));
 sg13g2_xor2_1 _13002_ (.B(_07192_),
    .A(_07190_),
    .X(_07194_));
 sg13g2_and2_1 _13003_ (.A(_07188_),
    .B(_07194_),
    .X(_07195_));
 sg13g2_a21oi_1 _13004_ (.A1(_06559_),
    .A2(net5310),
    .Y(_07196_),
    .B1(net5220));
 sg13g2_nor2_1 _13005_ (.A(net5776),
    .B(net5299),
    .Y(_07197_));
 sg13g2_a21oi_1 _13006_ (.A1(_06623_),
    .A2(net5300),
    .Y(_07198_),
    .B1(_07197_));
 sg13g2_nand2_1 _13007_ (.Y(_07199_),
    .A(_07196_),
    .B(_07198_));
 sg13g2_nor2_1 _13008_ (.A(_07196_),
    .B(_07198_),
    .Y(_07200_));
 sg13g2_xnor2_1 _13009_ (.Y(_07201_),
    .A(_07196_),
    .B(_07198_));
 sg13g2_a21oi_1 _13010_ (.A1(_06563_),
    .A2(net5310),
    .Y(_07202_),
    .B1(net5220));
 sg13g2_nand2_1 _13011_ (.Y(_07203_),
    .A(net5777),
    .B(net5304));
 sg13g2_o21ai_1 _13012_ (.B1(_07203_),
    .Y(_07204_),
    .A1(_06620_),
    .A2(net5304));
 sg13g2_nand2_1 _13013_ (.Y(_07205_),
    .A(_07202_),
    .B(_07204_));
 sg13g2_xor2_1 _13014_ (.B(_07204_),
    .A(_07202_),
    .X(_07206_));
 sg13g2_inv_1 _13015_ (.Y(_07207_),
    .A(_07206_));
 sg13g2_nor2_1 _13016_ (.A(_07201_),
    .B(_07207_),
    .Y(_07208_));
 sg13g2_nand2_1 _13017_ (.Y(_07209_),
    .A(_07195_),
    .B(_07208_));
 sg13g2_a21oi_1 _13018_ (.A1(net5223),
    .A2(net5296),
    .Y(_07210_),
    .B1(\fpga_top.cpu_top.csr_uimm[4] ));
 sg13g2_nor2_2 _13019_ (.A(_07150_),
    .B(_07210_),
    .Y(_07211_));
 sg13g2_nand2_1 _13020_ (.Y(_07212_),
    .A(net5780),
    .B(net5306));
 sg13g2_o21ai_1 _13021_ (.B1(_07212_),
    .Y(_07213_),
    .A1(_06617_),
    .A2(net5306));
 sg13g2_nor2_1 _13022_ (.A(_07211_),
    .B(_07213_),
    .Y(_07214_));
 sg13g2_xor2_1 _13023_ (.B(_07213_),
    .A(_07211_),
    .X(_07215_));
 sg13g2_a21oi_1 _13024_ (.A1(net5225),
    .A2(net5296),
    .Y(_07216_),
    .B1(\fpga_top.cpu_top.csr_uimm[3] ));
 sg13g2_nor2_1 _13025_ (.A(_07150_),
    .B(_07216_),
    .Y(_07217_));
 sg13g2_nand2_1 _13026_ (.Y(_07218_),
    .A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[18] ),
    .B(net5306));
 sg13g2_o21ai_1 _13027_ (.B1(_07218_),
    .Y(_07219_),
    .A1(_06614_),
    .A2(net5306));
 sg13g2_nand2_1 _13028_ (.Y(_07220_),
    .A(_07217_),
    .B(_07219_));
 sg13g2_xor2_1 _13029_ (.B(_07219_),
    .A(_07217_),
    .X(_07221_));
 sg13g2_inv_1 _13030_ (.Y(_07222_),
    .A(_07221_));
 sg13g2_and2_1 _13031_ (.A(_07215_),
    .B(_07221_),
    .X(_07223_));
 sg13g2_a21oi_1 _13032_ (.A1(net5223),
    .A2(net5296),
    .Y(_07224_),
    .B1(\fpga_top.cpu_top.csr_uimm[1] ));
 sg13g2_nor2_1 _13033_ (.A(_07150_),
    .B(_07224_),
    .Y(_07225_));
 sg13g2_nand2_1 _13034_ (.Y(_07226_),
    .A(net5593),
    .B(net5299));
 sg13g2_o21ai_1 _13035_ (.B1(_07226_),
    .Y(_07227_),
    .A1(_06574_),
    .A2(net5299));
 sg13g2_and2_1 _13036_ (.A(_07225_),
    .B(_07227_),
    .X(_07228_));
 sg13g2_xor2_1 _13037_ (.B(_07227_),
    .A(_07225_),
    .X(_07229_));
 sg13g2_a21oi_1 _13038_ (.A1(net5225),
    .A2(net5296),
    .Y(_07230_),
    .B1(\fpga_top.cpu_top.csr_uimm[2] ));
 sg13g2_nor2_2 _13039_ (.A(_07150_),
    .B(_07230_),
    .Y(_07231_));
 sg13g2_nor2_1 _13040_ (.A(net5785),
    .B(net5299),
    .Y(_07232_));
 sg13g2_a21oi_2 _13041_ (.B1(_07232_),
    .Y(_07233_),
    .A2(net5299),
    .A1(_06611_));
 sg13g2_nor2_1 _13042_ (.A(_07231_),
    .B(_07233_),
    .Y(_07234_));
 sg13g2_xor2_1 _13043_ (.B(_07233_),
    .A(_07231_),
    .X(_07235_));
 sg13g2_and2_1 _13044_ (.A(_07229_),
    .B(_07235_),
    .X(_07236_));
 sg13g2_nand2_1 _13045_ (.Y(_07237_),
    .A(_07223_),
    .B(_07236_));
 sg13g2_inv_1 _13046_ (.Y(_07238_),
    .A(_07237_));
 sg13g2_nor2_1 _13047_ (.A(_07209_),
    .B(_07237_),
    .Y(_07239_));
 sg13g2_a21oi_1 _13048_ (.A1(_07231_),
    .A2(_07233_),
    .Y(_07240_),
    .B1(_07228_));
 sg13g2_nor2_1 _13049_ (.A(_07234_),
    .B(_07240_),
    .Y(_07241_));
 sg13g2_nor2_1 _13050_ (.A(_07214_),
    .B(_07220_),
    .Y(_07242_));
 sg13g2_a221oi_1 _13051_ (.B2(_07241_),
    .C1(_07242_),
    .B1(_07223_),
    .A1(_07211_),
    .Y(_07243_),
    .A2(_07213_));
 sg13g2_inv_1 _13052_ (.Y(_07244_),
    .A(_07243_));
 sg13g2_nor2_1 _13053_ (.A(_07187_),
    .B(_07193_),
    .Y(_07245_));
 sg13g2_o21ai_1 _13054_ (.B1(_07199_),
    .Y(_07246_),
    .A1(_07200_),
    .A2(_07205_));
 sg13g2_a221oi_1 _13055_ (.B2(_07246_),
    .C1(_07245_),
    .B1(_07195_),
    .A1(_07190_),
    .Y(_07247_),
    .A2(_07192_));
 sg13g2_o21ai_1 _13056_ (.B1(_07247_),
    .Y(_07248_),
    .A1(_07209_),
    .A2(_07243_));
 sg13g2_a21oi_2 _13057_ (.B1(_07248_),
    .Y(_07249_),
    .A2(_07239_),
    .A1(_07183_));
 sg13g2_a21oi_1 _13058_ (.A1(_06558_),
    .A2(net5313),
    .Y(_07250_),
    .B1(net5220));
 sg13g2_nand2_1 _13059_ (.Y(_07251_),
    .A(net5768),
    .B(net5304));
 sg13g2_o21ai_1 _13060_ (.B1(_07251_),
    .Y(_07252_),
    .A1(_06631_),
    .A2(net5304));
 sg13g2_nor2_1 _13061_ (.A(_07250_),
    .B(_07252_),
    .Y(_07253_));
 sg13g2_nand2_1 _13062_ (.Y(_07254_),
    .A(_07250_),
    .B(_07252_));
 sg13g2_nor2b_1 _13063_ (.A(_07253_),
    .B_N(_07254_),
    .Y(_07255_));
 sg13g2_a21oi_1 _13064_ (.A1(_06575_),
    .A2(net5313),
    .Y(_07256_),
    .B1(net5220));
 sg13g2_nand2_1 _13065_ (.Y(_07257_),
    .A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[24] ),
    .B(net5304));
 sg13g2_o21ai_1 _13066_ (.B1(_07257_),
    .Y(_07258_),
    .A1(_06629_),
    .A2(net5304));
 sg13g2_nand2_1 _13067_ (.Y(_07259_),
    .A(_07256_),
    .B(_07258_));
 sg13g2_xor2_1 _13068_ (.B(_07258_),
    .A(_07256_),
    .X(_07260_));
 sg13g2_inv_1 _13069_ (.Y(_07261_),
    .A(_07260_));
 sg13g2_nand2_1 _13070_ (.Y(_07262_),
    .A(_07255_),
    .B(_07260_));
 sg13g2_o21ai_1 _13071_ (.B1(_07254_),
    .Y(_07263_),
    .A1(_07253_),
    .A2(_07259_));
 sg13g2_inv_1 _13072_ (.Y(_07264_),
    .A(_07263_));
 sg13g2_o21ai_1 _13073_ (.B1(_07264_),
    .Y(_07265_),
    .A1(_07249_),
    .A2(_07262_));
 sg13g2_a21oi_1 _13074_ (.A1(_06549_),
    .A2(net5310),
    .Y(_07266_),
    .B1(_07034_));
 sg13g2_nand2_1 _13075_ (.Y(_07267_),
    .A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[26] ),
    .B(net5305));
 sg13g2_o21ai_1 _13076_ (.B1(_07267_),
    .Y(_07268_),
    .A1(_06634_),
    .A2(net5305));
 sg13g2_nand2_1 _13077_ (.Y(_07269_),
    .A(_07266_),
    .B(_07268_));
 sg13g2_xor2_1 _13078_ (.B(_07268_),
    .A(_07266_),
    .X(_07270_));
 sg13g2_nand2_1 _13079_ (.Y(_07271_),
    .A(_07265_),
    .B(_07270_));
 sg13g2_xor2_1 _13080_ (.B(_07059_),
    .A(_07057_),
    .X(_07272_));
 sg13g2_and2_1 _13081_ (.A(_07270_),
    .B(_07272_),
    .X(_07273_));
 sg13g2_nor2_1 _13082_ (.A(_07060_),
    .B(_07269_),
    .Y(_07274_));
 sg13g2_a221oi_1 _13083_ (.B2(_07273_),
    .C1(_07274_),
    .B1(_07265_),
    .A1(_07057_),
    .Y(_07275_),
    .A2(_07059_));
 sg13g2_o21ai_1 _13084_ (.B1(_07054_),
    .Y(_07276_),
    .A1(_07056_),
    .A2(_07275_));
 sg13g2_nand2_1 _13085_ (.Y(_07277_),
    .A(_07047_),
    .B(_07049_));
 sg13g2_o21ai_1 _13086_ (.B1(_07277_),
    .Y(_07278_),
    .A1(_07050_),
    .A2(_07054_));
 sg13g2_inv_1 _13087_ (.Y(_07279_),
    .A(_07278_));
 sg13g2_nor2b_1 _13088_ (.A(_07050_),
    .B_N(_07277_),
    .Y(_07280_));
 sg13g2_nand2_1 _13089_ (.Y(_07281_),
    .A(_07055_),
    .B(_07280_));
 sg13g2_o21ai_1 _13090_ (.B1(_07279_),
    .Y(_07282_),
    .A1(_07275_),
    .A2(_07281_));
 sg13g2_a21oi_1 _13091_ (.A1(_07046_),
    .A2(_07282_),
    .Y(_07283_),
    .B1(_07045_));
 sg13g2_nand2_1 _13092_ (.Y(_07284_),
    .A(net5754),
    .B(net5306));
 sg13g2_o21ai_1 _13093_ (.B1(_07284_),
    .Y(_07285_),
    .A1(_06646_),
    .A2(net5306));
 sg13g2_xnor2_1 _13094_ (.Y(_07286_),
    .A(net5569),
    .B(_07285_));
 sg13g2_xnor2_1 _13095_ (.Y(_07287_),
    .A(_07283_),
    .B(_07286_));
 sg13g2_nor2_1 _13096_ (.A(\fpga_top.cpu_top.br_ofs[7] ),
    .B(net5569),
    .Y(_07288_));
 sg13g2_nor4_1 _13097_ (.A(\fpga_top.cpu_top.br_ofs[7] ),
    .B(\fpga_top.cpu_top.br_ofs[8] ),
    .C(net5570),
    .D(\fpga_top.cpu_top.br_ofs[12] ),
    .Y(_07289_));
 sg13g2_nand3_1 _13098_ (.B(_06556_),
    .C(_07288_),
    .A(_06555_),
    .Y(_07290_));
 sg13g2_nor2_1 _13099_ (.A(_06557_),
    .B(_07290_),
    .Y(_07291_));
 sg13g2_nand2_2 _13100_ (.Y(_07292_),
    .A(\fpga_top.cpu_top.br_ofs[10] ),
    .B(_07289_));
 sg13g2_nor2_1 _13101_ (.A(_06550_),
    .B(net5344),
    .Y(_07293_));
 sg13g2_or2_1 _13102_ (.X(_07294_),
    .B(net5344),
    .A(_06550_));
 sg13g2_or2_1 _13103_ (.X(_07295_),
    .B(\fpga_top.cpu_top.br_ofs[5] ),
    .A(net5571));
 sg13g2_nor3_1 _13104_ (.A(net5585),
    .B(_07028_),
    .C(_07295_),
    .Y(_07296_));
 sg13g2_nor3_2 _13105_ (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[4] ),
    .B(net6282),
    .C(net5586),
    .Y(_07297_));
 sg13g2_nor2b_2 _13106_ (.A(net5344),
    .B_N(_07297_),
    .Y(_07298_));
 sg13g2_nand2b_2 _13107_ (.Y(_07299_),
    .B(_07297_),
    .A_N(net5344));
 sg13g2_nor4_2 _13108_ (.A(net5585),
    .B(\fpga_top.cpu_top.decoder.illegal_ops_inst[5] ),
    .C(_07028_),
    .Y(_07300_),
    .D(net5344));
 sg13g2_or4_1 _13109_ (.A(net5586),
    .B(\fpga_top.cpu_top.decoder.illegal_ops_inst[5] ),
    .C(_07028_),
    .D(_07030_),
    .X(_07301_));
 sg13g2_nor2b_1 _13110_ (.A(net5581),
    .B_N(net5583),
    .Y(_07302_));
 sg13g2_nand2_2 _13111_ (.Y(_07303_),
    .A(net5382),
    .B(net5583));
 sg13g2_a21oi_1 _13112_ (.A1(_07300_),
    .A2(_07303_),
    .Y(_07304_),
    .B1(net5294));
 sg13g2_o21ai_1 _13113_ (.B1(_07299_),
    .Y(_07305_),
    .A1(_07301_),
    .A2(net5342));
 sg13g2_and2_1 _13114_ (.A(\fpga_top.cpu_top.br_ofs[12] ),
    .B(_07305_),
    .X(_07306_));
 sg13g2_nand2_1 _13115_ (.Y(_07307_),
    .A(_06549_),
    .B(net5342));
 sg13g2_nor3_2 _13116_ (.A(net5571),
    .B(_07301_),
    .C(_07303_),
    .Y(_07308_));
 sg13g2_nand3_1 _13117_ (.B(_07300_),
    .C(net5342),
    .A(_06549_),
    .Y(_07309_));
 sg13g2_nor2_2 _13118_ (.A(net5206),
    .B(_07308_),
    .Y(_07310_));
 sg13g2_a21o_2 _13119_ (.A2(net5113),
    .A1(\fpga_top.bus_gather.d_write_data[30] ),
    .B1(net5116),
    .X(_07311_));
 sg13g2_nor4_1 _13120_ (.A(net5585),
    .B(_07028_),
    .C(_07294_),
    .D(_07295_),
    .Y(_07312_));
 sg13g2_and2_1 _13121_ (.A(_07291_),
    .B(_07312_),
    .X(_07313_));
 sg13g2_nand2_1 _13122_ (.Y(_07314_),
    .A(_07291_),
    .B(_07312_));
 sg13g2_xnor2_1 _13123_ (.Y(_07315_),
    .A(_07311_),
    .B(net5109));
 sg13g2_and2_1 _13124_ (.A(_06581_),
    .B(_07315_),
    .X(_07316_));
 sg13g2_a21o_2 _13125_ (.A2(net5113),
    .A1(\fpga_top.bus_gather.d_write_data[29] ),
    .B1(net5116),
    .X(_07317_));
 sg13g2_inv_1 _13126_ (.Y(_07318_),
    .A(_07317_));
 sg13g2_xnor2_1 _13127_ (.Y(_07319_),
    .A(net5110),
    .B(_07317_));
 sg13g2_inv_1 _13128_ (.Y(_07320_),
    .A(_07319_));
 sg13g2_a21o_2 _13129_ (.A2(net5112),
    .A1(\fpga_top.bus_gather.d_write_data[21] ),
    .B1(net5115),
    .X(_07321_));
 sg13g2_inv_1 _13130_ (.Y(_07322_),
    .A(_07321_));
 sg13g2_xnor2_1 _13131_ (.Y(_07323_),
    .A(net5109),
    .B(_07321_));
 sg13g2_nor2b_1 _13132_ (.A(_07323_),
    .B_N(net5775),
    .Y(_07324_));
 sg13g2_xnor2_1 _13133_ (.Y(_07325_),
    .A(net5775),
    .B(_07323_));
 sg13g2_a21o_2 _13134_ (.A2(net5112),
    .A1(\fpga_top.bus_gather.d_write_data[22] ),
    .B1(net5115),
    .X(_07326_));
 sg13g2_xnor2_1 _13135_ (.Y(_07327_),
    .A(net5106),
    .B(_07326_));
 sg13g2_xnor2_1 _13136_ (.Y(_07328_),
    .A(_06579_),
    .B(_07327_));
 sg13g2_and2_1 _13137_ (.A(_07325_),
    .B(_07328_),
    .X(_07329_));
 sg13g2_a21o_2 _13138_ (.A2(net5113),
    .A1(\fpga_top.bus_gather.d_write_data[19] ),
    .B1(net5116),
    .X(_07330_));
 sg13g2_inv_1 _13139_ (.Y(_07331_),
    .A(_07330_));
 sg13g2_xnor2_1 _13140_ (.Y(_07332_),
    .A(net5109),
    .B(_07330_));
 sg13g2_nor2b_1 _13141_ (.A(_07332_),
    .B_N(net5778),
    .Y(_07333_));
 sg13g2_xor2_1 _13142_ (.B(_07332_),
    .A(net5778),
    .X(_07334_));
 sg13g2_a21o_2 _13143_ (.A2(net5112),
    .A1(\fpga_top.bus_gather.d_write_data[20] ),
    .B1(net5115),
    .X(_07335_));
 sg13g2_xnor2_1 _13144_ (.Y(_07336_),
    .A(net5109),
    .B(_07335_));
 sg13g2_nor2_1 _13145_ (.A(_06578_),
    .B(_07336_),
    .Y(_07337_));
 sg13g2_xnor2_1 _13146_ (.Y(_07338_),
    .A(net5777),
    .B(_07336_));
 sg13g2_nor2b_1 _13147_ (.A(_07334_),
    .B_N(_07338_),
    .Y(_07339_));
 sg13g2_nand2_1 _13148_ (.Y(_07340_),
    .A(_07329_),
    .B(_07339_));
 sg13g2_o21ai_1 _13149_ (.B1(_07324_),
    .Y(_07341_),
    .A1(net5774),
    .A2(_07327_));
 sg13g2_inv_1 _13150_ (.Y(_07342_),
    .A(_07341_));
 sg13g2_nor2_1 _13151_ (.A(_07333_),
    .B(_07337_),
    .Y(_07343_));
 sg13g2_a21oi_1 _13152_ (.A1(_06578_),
    .A2(_07336_),
    .Y(_07344_),
    .B1(_07343_));
 sg13g2_a221oi_1 _13153_ (.B2(_07344_),
    .C1(_07342_),
    .B1(_07329_),
    .A1(net5774),
    .Y(_07345_),
    .A2(_07327_));
 sg13g2_a21o_2 _13154_ (.A2(net5111),
    .A1(\fpga_top.bus_gather.d_write_data[13] ),
    .B1(net5114),
    .X(_07346_));
 sg13g2_inv_1 _13155_ (.Y(_07347_),
    .A(_07346_));
 sg13g2_xnor2_1 _13156_ (.Y(_07348_),
    .A(net5108),
    .B(_07346_));
 sg13g2_nand2b_1 _13157_ (.Y(_07349_),
    .B(net5791),
    .A_N(_07348_));
 sg13g2_inv_1 _13158_ (.Y(_07350_),
    .A(_07349_));
 sg13g2_xnor2_1 _13159_ (.Y(_07351_),
    .A(net5791),
    .B(_07348_));
 sg13g2_xor2_1 _13160_ (.B(_07348_),
    .A(net5791),
    .X(_07352_));
 sg13g2_a21o_2 _13161_ (.A2(net5111),
    .A1(\fpga_top.bus_gather.d_write_data[14] ),
    .B1(net5114),
    .X(_07353_));
 sg13g2_xnor2_1 _13162_ (.Y(_07354_),
    .A(net5108),
    .B(_07353_));
 sg13g2_nand2_1 _13163_ (.Y(_07355_),
    .A(_06573_),
    .B(_07354_));
 sg13g2_nor2_1 _13164_ (.A(_06573_),
    .B(_07354_),
    .Y(_07356_));
 sg13g2_xnor2_1 _13165_ (.Y(_07357_),
    .A(_06573_),
    .B(_07354_));
 sg13g2_nor2_1 _13166_ (.A(_07352_),
    .B(_07357_),
    .Y(_07358_));
 sg13g2_a21o_2 _13167_ (.A2(_07310_),
    .A1(\fpga_top.bus_gather.d_write_data[11] ),
    .B1(net5114),
    .X(_07359_));
 sg13g2_xnor2_1 _13168_ (.Y(_07360_),
    .A(net5107),
    .B(_07359_));
 sg13g2_nor2_1 _13169_ (.A(_06572_),
    .B(_07360_),
    .Y(_07361_));
 sg13g2_xnor2_1 _13170_ (.Y(_07362_),
    .A(_06572_),
    .B(_07360_));
 sg13g2_a21oi_2 _13171_ (.B1(net5114),
    .Y(_07363_),
    .A2(net5111),
    .A1(\fpga_top.bus_gather.d_write_data[12] ));
 sg13g2_xnor2_1 _13172_ (.Y(_07364_),
    .A(net5108),
    .B(_07363_));
 sg13g2_and2_1 _13173_ (.A(net5794),
    .B(_07364_),
    .X(_07365_));
 sg13g2_or2_1 _13174_ (.X(_07366_),
    .B(_07364_),
    .A(net5794));
 sg13g2_xnor2_1 _13175_ (.Y(_07367_),
    .A(net5794),
    .B(_07364_));
 sg13g2_or2_1 _13176_ (.X(_07368_),
    .B(_07367_),
    .A(_07362_));
 sg13g2_a21o_1 _13177_ (.A2(_07366_),
    .A1(_07361_),
    .B1(_07365_),
    .X(_07369_));
 sg13g2_a21oi_1 _13178_ (.A1(_07361_),
    .A2(_07366_),
    .Y(_07370_),
    .B1(_07365_));
 sg13g2_nand3b_1 _13179_ (.B(_07297_),
    .C(_06550_),
    .Y(_07371_),
    .A_N(_07030_));
 sg13g2_a22oi_1 _13180_ (.Y(_07372_),
    .B1(_07300_),
    .B2(_07303_),
    .A2(net5294),
    .A1(_06550_));
 sg13g2_o21ai_1 _13181_ (.B1(_07371_),
    .Y(_07373_),
    .A1(_07301_),
    .A2(net5342));
 sg13g2_a21oi_1 _13182_ (.A1(net5205),
    .A2(_07372_),
    .Y(_07374_),
    .B1(\fpga_top.cpu_top.alui_shamt[2] ));
 sg13g2_nor3_1 _13183_ (.A(\fpga_top.bus_gather.d_write_data[2] ),
    .B(net5206),
    .C(_07308_),
    .Y(_07375_));
 sg13g2_nor2_1 _13184_ (.A(_06550_),
    .B(_07299_),
    .Y(_07376_));
 sg13g2_nand2_2 _13185_ (.Y(_07377_),
    .A(net6314),
    .B(net5294));
 sg13g2_nor2_1 _13186_ (.A(\fpga_top.cpu_top.br_ofs[2] ),
    .B(_07377_),
    .Y(_07378_));
 sg13g2_nor3_1 _13187_ (.A(_07374_),
    .B(_07375_),
    .C(_07378_),
    .Y(_07379_));
 sg13g2_or3_1 _13188_ (.A(_07374_),
    .B(_07375_),
    .C(_07378_),
    .X(_07380_));
 sg13g2_xnor2_1 _13189_ (.Y(_07381_),
    .A(net5104),
    .B(net5012));
 sg13g2_nor2_1 _13190_ (.A(net5819),
    .B(_07381_),
    .Y(_07382_));
 sg13g2_o21ai_1 _13191_ (.B1(\fpga_top.bus_gather.d_write_data[1] ),
    .Y(_07383_),
    .A1(_07301_),
    .A2(_07307_));
 sg13g2_nand4_1 _13192_ (.B(\fpga_top.cpu_top.alui_shamt[1] ),
    .C(_07300_),
    .A(_06549_),
    .Y(_07384_),
    .D(net5342));
 sg13g2_nand3_1 _13193_ (.B(_07383_),
    .C(_07384_),
    .A(_07377_),
    .Y(_07385_));
 sg13g2_a21oi_1 _13194_ (.A1(_06560_),
    .A2(_07376_),
    .Y(_07386_),
    .B1(_07373_));
 sg13g2_nor2_1 _13195_ (.A(_06559_),
    .B(_07372_),
    .Y(_07387_));
 sg13g2_a21oi_2 _13196_ (.B1(_07387_),
    .Y(_07388_),
    .A2(_07386_),
    .A1(_07385_));
 sg13g2_a21o_2 _13197_ (.A2(_07386_),
    .A1(_07385_),
    .B1(_07387_),
    .X(_07389_));
 sg13g2_xnor2_1 _13198_ (.Y(_07390_),
    .A(net5105),
    .B(net4997));
 sg13g2_nor2b_1 _13199_ (.A(_07390_),
    .B_N(net5822),
    .Y(_07391_));
 sg13g2_xnor2_1 _13200_ (.Y(_07392_),
    .A(net5822),
    .B(_07390_));
 sg13g2_a21oi_1 _13201_ (.A1(net5205),
    .A2(_07372_),
    .Y(_07393_),
    .B1(net5573));
 sg13g2_a221oi_1 _13202_ (.B2(_06564_),
    .C1(_07393_),
    .B1(_07376_),
    .A1(_06562_),
    .Y(_07394_),
    .A2(net5111));
 sg13g2_nor2b_2 _13203_ (.A(net5825),
    .B_N(net4977),
    .Y(_07395_));
 sg13g2_nor2_1 _13204_ (.A(net5107),
    .B(net4977),
    .Y(_07396_));
 sg13g2_nor2_1 _13205_ (.A(_07395_),
    .B(_07396_),
    .Y(_07397_));
 sg13g2_a21oi_1 _13206_ (.A1(_07392_),
    .A2(_07397_),
    .Y(_07398_),
    .B1(_07391_));
 sg13g2_a221oi_1 _13207_ (.B2(_07397_),
    .C1(_07391_),
    .B1(_07392_),
    .A1(net5819),
    .Y(_07399_),
    .A2(_07381_));
 sg13g2_nor3_1 _13208_ (.A(\fpga_top.bus_gather.d_write_data[3] ),
    .B(net5206),
    .C(_07308_),
    .Y(_07400_));
 sg13g2_nor2_1 _13209_ (.A(\fpga_top.cpu_top.br_ofs[3] ),
    .B(_07377_),
    .Y(_07401_));
 sg13g2_a21oi_1 _13210_ (.A1(_07309_),
    .A2(_07372_),
    .Y(_07402_),
    .B1(\fpga_top.cpu_top.alui_shamt[3] ));
 sg13g2_nor3_2 _13211_ (.A(_07400_),
    .B(_07401_),
    .C(_07402_),
    .Y(_07403_));
 sg13g2_or3_1 _13212_ (.A(_07400_),
    .B(_07401_),
    .C(_07402_),
    .X(_07404_));
 sg13g2_xnor2_1 _13213_ (.Y(_07405_),
    .A(net5105),
    .B(net4965));
 sg13g2_nand2_1 _13214_ (.Y(_07406_),
    .A(net5817),
    .B(_07405_));
 sg13g2_xnor2_1 _13215_ (.Y(_07407_),
    .A(net5817),
    .B(_07405_));
 sg13g2_or3_1 _13216_ (.A(_07382_),
    .B(_07399_),
    .C(_07407_),
    .X(_07408_));
 sg13g2_nor2_1 _13217_ (.A(\fpga_top.bus_gather.d_write_data[4] ),
    .B(_07308_),
    .Y(_07409_));
 sg13g2_o21ai_1 _13218_ (.B1(_07304_),
    .Y(_07410_),
    .A1(\fpga_top.cpu_top.alui_shamt[4] ),
    .A2(_07309_));
 sg13g2_nor2_1 _13219_ (.A(_07409_),
    .B(_07410_),
    .Y(_07411_));
 sg13g2_a22oi_1 _13220_ (.Y(_07412_),
    .B1(_07376_),
    .B2(\fpga_top.cpu_top.br_ofs[4] ),
    .A2(_07373_),
    .A1(\fpga_top.cpu_top.alui_shamt[4] ));
 sg13g2_nor2b_1 _13221_ (.A(_07411_),
    .B_N(_07412_),
    .Y(_07413_));
 sg13g2_o21ai_1 _13222_ (.B1(_07412_),
    .Y(_07414_),
    .A1(_07409_),
    .A2(_07410_));
 sg13g2_xnor2_1 _13223_ (.Y(_07415_),
    .A(net5105),
    .B(net4954));
 sg13g2_nand2_1 _13224_ (.Y(_07416_),
    .A(net5814),
    .B(_07415_));
 sg13g2_a22oi_1 _13225_ (.Y(_07417_),
    .B1(net5111),
    .B2(\fpga_top.bus_gather.d_write_data[6] ),
    .A2(net5206),
    .A1(net5571));
 sg13g2_xnor2_1 _13226_ (.Y(_07418_),
    .A(net5107),
    .B(_07417_));
 sg13g2_and2_1 _13227_ (.A(net5807),
    .B(_07418_),
    .X(_07419_));
 sg13g2_or2_1 _13228_ (.X(_07420_),
    .B(_07418_),
    .A(net5807));
 sg13g2_xor2_1 _13229_ (.B(_07418_),
    .A(net5807),
    .X(_07421_));
 sg13g2_nand3_1 _13230_ (.B(net5207),
    .C(net5205),
    .A(\fpga_top.bus_gather.d_write_data[5] ),
    .Y(_07422_));
 sg13g2_o21ai_1 _13231_ (.B1(_07422_),
    .Y(_07423_),
    .A1(_06558_),
    .A2(net5207));
 sg13g2_xnor2_1 _13232_ (.Y(_07424_),
    .A(net5107),
    .B(_07423_));
 sg13g2_nor2_1 _13233_ (.A(_06565_),
    .B(_07424_),
    .Y(_07425_));
 sg13g2_xnor2_1 _13234_ (.Y(_07426_),
    .A(net5810),
    .B(_07424_));
 sg13g2_or2_1 _13235_ (.X(_07427_),
    .B(_07415_),
    .A(net5814));
 sg13g2_and2_1 _13236_ (.A(_07426_),
    .B(_07427_),
    .X(_07428_));
 sg13g2_nand3_1 _13237_ (.B(_07426_),
    .C(_07427_),
    .A(_07421_),
    .Y(_07429_));
 sg13g2_nand4_1 _13238_ (.B(_07421_),
    .C(_07426_),
    .A(_07416_),
    .Y(_07430_),
    .D(_07427_));
 sg13g2_nand2_1 _13239_ (.Y(_07431_),
    .A(_07416_),
    .B(_07427_));
 sg13g2_nor4_2 _13240_ (.A(_07382_),
    .B(_07399_),
    .C(_07407_),
    .Y(_07432_),
    .D(_07430_));
 sg13g2_and2_1 _13241_ (.A(_07406_),
    .B(_07416_),
    .X(_07433_));
 sg13g2_o21ai_1 _13242_ (.B1(_07420_),
    .Y(_07434_),
    .A1(_07419_),
    .A2(_07425_));
 sg13g2_o21ai_1 _13243_ (.B1(_07434_),
    .Y(_07435_),
    .A1(_07429_),
    .A2(_07433_));
 sg13g2_nand2_2 _13244_ (.Y(_07436_),
    .A(net5570),
    .B(net5206));
 sg13g2_nand3_1 _13245_ (.B(net5207),
    .C(net5205),
    .A(\fpga_top.bus_gather.d_write_data[9] ),
    .Y(_07437_));
 sg13g2_nand2_2 _13246_ (.Y(_07438_),
    .A(_07436_),
    .B(_07437_));
 sg13g2_nand3_1 _13247_ (.B(_07436_),
    .C(_07437_),
    .A(net5104),
    .Y(_07439_));
 sg13g2_a21o_1 _13248_ (.A2(_07437_),
    .A1(_07436_),
    .B1(net5104),
    .X(_07440_));
 sg13g2_and3_1 _13249_ (.X(_07441_),
    .A(net5800),
    .B(_07439_),
    .C(_07440_));
 sg13g2_nand3_1 _13250_ (.B(_07439_),
    .C(_07440_),
    .A(net5800),
    .Y(_07442_));
 sg13g2_a21oi_1 _13251_ (.A1(_07439_),
    .A2(_07440_),
    .Y(_07443_),
    .B1(net5800));
 sg13g2_nor2_1 _13252_ (.A(_07441_),
    .B(_07443_),
    .Y(_07444_));
 sg13g2_nor2_1 _13253_ (.A(_06557_),
    .B(net5207),
    .Y(_07445_));
 sg13g2_nand2_1 _13254_ (.Y(_07446_),
    .A(\fpga_top.cpu_top.br_ofs[10] ),
    .B(net5206));
 sg13g2_nor3_1 _13255_ (.A(_06593_),
    .B(net5206),
    .C(_07308_),
    .Y(_07447_));
 sg13g2_nand3_1 _13256_ (.B(net5207),
    .C(net5205),
    .A(\fpga_top.bus_gather.d_write_data[10] ),
    .Y(_07448_));
 sg13g2_nand2_2 _13257_ (.Y(_07449_),
    .A(_07446_),
    .B(_07448_));
 sg13g2_a21oi_1 _13258_ (.A1(_07446_),
    .A2(_07448_),
    .Y(_07450_),
    .B1(net5107));
 sg13g2_o21ai_1 _13259_ (.B1(net5104),
    .Y(_07451_),
    .A1(_07445_),
    .A2(_07447_));
 sg13g2_nor3_1 _13260_ (.A(net5104),
    .B(_07445_),
    .C(_07447_),
    .Y(_07452_));
 sg13g2_nand3_1 _13261_ (.B(_07446_),
    .C(_07448_),
    .A(net5107),
    .Y(_07453_));
 sg13g2_a21oi_1 _13262_ (.A1(_07451_),
    .A2(_07453_),
    .Y(_07454_),
    .B1(_06571_));
 sg13g2_o21ai_1 _13263_ (.B1(net5798),
    .Y(_07455_),
    .A1(_07450_),
    .A2(_07452_));
 sg13g2_nor3_1 _13264_ (.A(net5798),
    .B(_07450_),
    .C(_07452_),
    .Y(_07456_));
 sg13g2_nor2_1 _13265_ (.A(_07454_),
    .B(_07456_),
    .Y(_07457_));
 sg13g2_nor4_1 _13266_ (.A(_07441_),
    .B(_07443_),
    .C(_07454_),
    .D(_07456_),
    .Y(_07458_));
 sg13g2_nand2_1 _13267_ (.Y(_07459_),
    .A(\fpga_top.cpu_top.br_ofs[8] ),
    .B(_07305_));
 sg13g2_nand3_1 _13268_ (.B(net5207),
    .C(net5205),
    .A(\fpga_top.bus_gather.d_write_data[8] ),
    .Y(_07460_));
 sg13g2_and2_1 _13269_ (.A(_07459_),
    .B(_07460_),
    .X(_07461_));
 sg13g2_a21oi_1 _13270_ (.A1(_07459_),
    .A2(_07460_),
    .Y(_07462_),
    .B1(net5107));
 sg13g2_and3_1 _13271_ (.X(_07463_),
    .A(net5107),
    .B(_07459_),
    .C(_07460_));
 sg13g2_nor3_1 _13272_ (.A(net5803),
    .B(_07462_),
    .C(_07463_),
    .Y(_07464_));
 sg13g2_o21ai_1 _13273_ (.B1(net5803),
    .Y(_07465_),
    .A1(_07462_),
    .A2(_07463_));
 sg13g2_nor2b_1 _13274_ (.A(_07464_),
    .B_N(_07465_),
    .Y(_07466_));
 sg13g2_nand2_1 _13275_ (.Y(_07467_),
    .A(\fpga_top.cpu_top.br_ofs[7] ),
    .B(net5206));
 sg13g2_nand3_1 _13276_ (.B(net5207),
    .C(net5205),
    .A(\fpga_top.bus_gather.d_write_data[7] ),
    .Y(_07468_));
 sg13g2_and2_1 _13277_ (.A(_07467_),
    .B(_07468_),
    .X(_07469_));
 sg13g2_inv_1 _13278_ (.Y(_07470_),
    .A(_07469_));
 sg13g2_nand3_1 _13279_ (.B(_07467_),
    .C(_07468_),
    .A(net5104),
    .Y(_07471_));
 sg13g2_a21oi_1 _13280_ (.A1(_07467_),
    .A2(_07468_),
    .Y(_07472_),
    .B1(net5104));
 sg13g2_xnor2_1 _13281_ (.Y(_07473_),
    .A(net5104),
    .B(_07469_));
 sg13g2_nand3b_1 _13282_ (.B(net5805),
    .C(_07471_),
    .Y(_07474_),
    .A_N(_07472_));
 sg13g2_xnor2_1 _13283_ (.Y(_07475_),
    .A(net5805),
    .B(_07473_));
 sg13g2_nand3_1 _13284_ (.B(_07466_),
    .C(_07475_),
    .A(_07458_),
    .Y(_07476_));
 sg13g2_inv_1 _13285_ (.Y(_07477_),
    .A(_07476_));
 sg13g2_o21ai_1 _13286_ (.B1(_07477_),
    .Y(_07478_),
    .A1(_07432_),
    .A2(_07435_));
 sg13g2_a21oi_1 _13287_ (.A1(_07465_),
    .A2(_07474_),
    .Y(_07479_),
    .B1(_07464_));
 sg13g2_a21o_1 _13288_ (.A2(_07474_),
    .A1(_07465_),
    .B1(_07464_),
    .X(_07480_));
 sg13g2_a21oi_1 _13289_ (.A1(_07442_),
    .A2(_07455_),
    .Y(_07481_),
    .B1(_07456_));
 sg13g2_a21oi_2 _13290_ (.B1(_07481_),
    .Y(_07482_),
    .A2(_07479_),
    .A1(_07458_));
 sg13g2_o21ai_1 _13291_ (.B1(_07370_),
    .Y(_07483_),
    .A1(_07368_),
    .A2(_07482_));
 sg13g2_a221oi_1 _13292_ (.B2(_07483_),
    .C1(_07356_),
    .B1(_07358_),
    .A1(_07350_),
    .Y(_07484_),
    .A2(_07355_));
 sg13g2_nor4_1 _13293_ (.A(_07352_),
    .B(_07357_),
    .C(_07368_),
    .D(_07476_),
    .Y(_07485_));
 sg13g2_o21ai_1 _13294_ (.B1(_07485_),
    .Y(_07486_),
    .A1(_07432_),
    .A2(_07435_));
 sg13g2_a21o_2 _13295_ (.A2(net5111),
    .A1(\fpga_top.bus_gather.d_write_data[15] ),
    .B1(net5114),
    .X(_07487_));
 sg13g2_inv_1 _13296_ (.Y(_07488_),
    .A(_07487_));
 sg13g2_xnor2_1 _13297_ (.Y(_07489_),
    .A(net5108),
    .B(_07487_));
 sg13g2_nor2b_1 _13298_ (.A(_07489_),
    .B_N(net5787),
    .Y(_07490_));
 sg13g2_xor2_1 _13299_ (.B(_07489_),
    .A(net5787),
    .X(_07491_));
 sg13g2_a21oi_1 _13300_ (.A1(_07484_),
    .A2(_07486_),
    .Y(_07492_),
    .B1(_07491_));
 sg13g2_a21o_2 _13301_ (.A2(net5113),
    .A1(\fpga_top.bus_gather.d_write_data[17] ),
    .B1(net5114),
    .X(_07493_));
 sg13g2_inv_1 _13302_ (.Y(_07494_),
    .A(_07493_));
 sg13g2_xnor2_1 _13303_ (.Y(_07495_),
    .A(net5106),
    .B(_07493_));
 sg13g2_and2_1 _13304_ (.A(net5783),
    .B(_07495_),
    .X(_07496_));
 sg13g2_xnor2_1 _13305_ (.Y(_07497_),
    .A(net5783),
    .B(_07495_));
 sg13g2_a21o_2 _13306_ (.A2(net5113),
    .A1(\fpga_top.bus_gather.d_write_data[18] ),
    .B1(net5114),
    .X(_07498_));
 sg13g2_inv_1 _13307_ (.Y(_07499_),
    .A(_07498_));
 sg13g2_xnor2_1 _13308_ (.Y(_07500_),
    .A(net5106),
    .B(_07498_));
 sg13g2_or2_1 _13309_ (.X(_07501_),
    .B(_07500_),
    .A(net5781));
 sg13g2_xor2_1 _13310_ (.B(_07500_),
    .A(net5781),
    .X(_07502_));
 sg13g2_nor2b_1 _13311_ (.A(_07497_),
    .B_N(_07502_),
    .Y(_07503_));
 sg13g2_a21o_2 _13312_ (.A2(net5111),
    .A1(\fpga_top.bus_gather.d_write_data[16] ),
    .B1(_07306_),
    .X(_07504_));
 sg13g2_inv_1 _13313_ (.Y(_07505_),
    .A(_07504_));
 sg13g2_xnor2_1 _13314_ (.Y(_07506_),
    .A(net5108),
    .B(_07504_));
 sg13g2_nand2_1 _13315_ (.Y(_07507_),
    .A(_06574_),
    .B(_07506_));
 sg13g2_nor2_1 _13316_ (.A(_06574_),
    .B(_07506_),
    .Y(_07508_));
 sg13g2_xnor2_1 _13317_ (.Y(_07509_),
    .A(net5786),
    .B(_07506_));
 sg13g2_nand3b_1 _13318_ (.B(_07503_),
    .C(_07509_),
    .Y(_07510_),
    .A_N(_07491_));
 sg13g2_a21o_2 _13319_ (.A2(_07486_),
    .A1(_07484_),
    .B1(_07510_),
    .X(_07511_));
 sg13g2_nor2_1 _13320_ (.A(_07490_),
    .B(_07508_),
    .Y(_07512_));
 sg13g2_inv_1 _13321_ (.Y(_07513_),
    .A(_07512_));
 sg13g2_nor2b_1 _13322_ (.A(_07512_),
    .B_N(_07503_),
    .Y(_07514_));
 sg13g2_a21o_1 _13323_ (.A2(_07500_),
    .A1(net5781),
    .B1(_07496_),
    .X(_07515_));
 sg13g2_a22oi_1 _13324_ (.Y(_07516_),
    .B1(_07515_),
    .B2(_07501_),
    .A2(_07514_),
    .A1(_07507_));
 sg13g2_and2_1 _13325_ (.A(_07345_),
    .B(_07516_),
    .X(_07517_));
 sg13g2_a22oi_1 _13326_ (.Y(_07518_),
    .B1(_07511_),
    .B2(_07517_),
    .A2(_07345_),
    .A1(_07340_));
 sg13g2_a21o_2 _13327_ (.A2(net5112),
    .A1(\fpga_top.bus_gather.d_write_data[23] ),
    .B1(net5115),
    .X(_07519_));
 sg13g2_inv_1 _13328_ (.Y(_07520_),
    .A(_07519_));
 sg13g2_xnor2_1 _13329_ (.Y(_07521_),
    .A(net5109),
    .B(_07519_));
 sg13g2_nor2b_1 _13330_ (.A(_07521_),
    .B_N(net5771),
    .Y(_07522_));
 sg13g2_xnor2_1 _13331_ (.Y(_07523_),
    .A(net5771),
    .B(_07521_));
 sg13g2_inv_1 _13332_ (.Y(_07524_),
    .A(_07523_));
 sg13g2_a221oi_1 _13333_ (.B2(_07517_),
    .C1(_07524_),
    .B1(_07511_),
    .A1(_07340_),
    .Y(_07525_),
    .A2(_07345_));
 sg13g2_a21o_2 _13334_ (.A2(net5112),
    .A1(\fpga_top.bus_gather.d_write_data[25] ),
    .B1(net5116),
    .X(_07526_));
 sg13g2_inv_1 _13335_ (.Y(_07527_),
    .A(_07526_));
 sg13g2_xnor2_1 _13336_ (.Y(_07528_),
    .A(net5109),
    .B(_07526_));
 sg13g2_nand2b_1 _13337_ (.Y(_07529_),
    .B(net5767),
    .A_N(_07528_));
 sg13g2_xnor2_1 _13338_ (.Y(_07530_),
    .A(net5767),
    .B(_07528_));
 sg13g2_inv_1 _13339_ (.Y(_07531_),
    .A(_07530_));
 sg13g2_a21o_2 _13340_ (.A2(net5113),
    .A1(\fpga_top.bus_gather.d_write_data[26] ),
    .B1(net5115),
    .X(_07532_));
 sg13g2_inv_1 _13341_ (.Y(_07533_),
    .A(_07532_));
 sg13g2_xnor2_1 _13342_ (.Y(_07534_),
    .A(net5106),
    .B(_07532_));
 sg13g2_nor2_1 _13343_ (.A(net5765),
    .B(_07534_),
    .Y(_07535_));
 sg13g2_xor2_1 _13344_ (.B(_07534_),
    .A(net5765),
    .X(_07536_));
 sg13g2_and2_1 _13345_ (.A(_07530_),
    .B(_07536_),
    .X(_07537_));
 sg13g2_a21oi_2 _13346_ (.B1(net5115),
    .Y(_07538_),
    .A2(net5112),
    .A1(\fpga_top.bus_gather.d_write_data[24] ));
 sg13g2_xnor2_1 _13347_ (.Y(_07539_),
    .A(net5110),
    .B(_07538_));
 sg13g2_or2_1 _13348_ (.X(_07540_),
    .B(_07539_),
    .A(net5770));
 sg13g2_xor2_1 _13349_ (.B(_07539_),
    .A(net5770),
    .X(_07541_));
 sg13g2_nand3_1 _13350_ (.B(_07537_),
    .C(_07541_),
    .A(_07523_),
    .Y(_07542_));
 sg13g2_a221oi_1 _13351_ (.B2(_07517_),
    .C1(_07542_),
    .B1(_07511_),
    .A1(_07340_),
    .Y(_07543_),
    .A2(_07345_));
 sg13g2_a21o_1 _13352_ (.A2(_07539_),
    .A1(net5770),
    .B1(_07522_),
    .X(_07544_));
 sg13g2_nand3_1 _13353_ (.B(_07540_),
    .C(_07544_),
    .A(_07537_),
    .Y(_07545_));
 sg13g2_o21ai_1 _13354_ (.B1(_07545_),
    .Y(_07546_),
    .A1(_07529_),
    .A2(_07535_));
 sg13g2_a21o_1 _13355_ (.A2(_07534_),
    .A1(net5765),
    .B1(_07546_),
    .X(_07547_));
 sg13g2_nor2_1 _13356_ (.A(_07543_),
    .B(_07547_),
    .Y(_07548_));
 sg13g2_a21o_2 _13357_ (.A2(net5112),
    .A1(\fpga_top.bus_gather.d_write_data[28] ),
    .B1(net5115),
    .X(_07549_));
 sg13g2_xnor2_1 _13358_ (.Y(_07550_),
    .A(net5109),
    .B(_07549_));
 sg13g2_inv_1 _13359_ (.Y(_07551_),
    .A(_07550_));
 sg13g2_xnor2_1 _13360_ (.Y(_07552_),
    .A(net5760),
    .B(_07550_));
 sg13g2_inv_1 _13361_ (.Y(_07553_),
    .A(_07552_));
 sg13g2_a21o_2 _13362_ (.A2(net5112),
    .A1(\fpga_top.bus_gather.d_write_data[27] ),
    .B1(net5115),
    .X(_07554_));
 sg13g2_inv_1 _13363_ (.Y(_07555_),
    .A(_07554_));
 sg13g2_xnor2_1 _13364_ (.Y(_07556_),
    .A(net5106),
    .B(_07554_));
 sg13g2_nand2_1 _13365_ (.Y(_07557_),
    .A(net5761),
    .B(_07556_));
 sg13g2_xnor2_1 _13366_ (.Y(_07558_),
    .A(net5761),
    .B(_07556_));
 sg13g2_nor2_1 _13367_ (.A(_07553_),
    .B(_07558_),
    .Y(_07559_));
 sg13g2_o21ai_1 _13368_ (.B1(_07559_),
    .Y(_07560_),
    .A1(_07543_),
    .A2(_07547_));
 sg13g2_a21oi_1 _13369_ (.A1(_06580_),
    .A2(_07550_),
    .Y(_07561_),
    .B1(_07557_));
 sg13g2_a21oi_1 _13370_ (.A1(net5760),
    .A2(_07551_),
    .Y(_07562_),
    .B1(_07561_));
 sg13g2_xor2_1 _13371_ (.B(_07319_),
    .A(net5758),
    .X(_07563_));
 sg13g2_a21oi_1 _13372_ (.A1(_07560_),
    .A2(_07562_),
    .Y(_07564_),
    .B1(_07563_));
 sg13g2_a21oi_2 _13373_ (.B1(_07564_),
    .Y(_07565_),
    .A2(_07320_),
    .A1(net5758));
 sg13g2_nand2b_1 _13374_ (.Y(_07566_),
    .B(net5756),
    .A_N(_07315_));
 sg13g2_o21ai_1 _13375_ (.B1(_07566_),
    .Y(_07567_),
    .A1(_07316_),
    .A2(_07565_));
 sg13g2_a21oi_2 _13376_ (.B1(net5114),
    .Y(_07568_),
    .A2(net5111),
    .A1(\fpga_top.bus_gather.d_write_data[31] ));
 sg13g2_inv_1 _13377_ (.Y(_07569_),
    .A(_07568_));
 sg13g2_xnor2_1 _13378_ (.Y(_07570_),
    .A(net5754),
    .B(_07568_));
 sg13g2_xnor2_1 _13379_ (.Y(_07571_),
    .A(net5109),
    .B(_07570_));
 sg13g2_nor2_2 _13380_ (.A(_07037_),
    .B(_07298_),
    .Y(_07572_));
 sg13g2_nand2_1 _13381_ (.Y(_07573_),
    .A(_07038_),
    .B(_07299_));
 sg13g2_xnor2_1 _13382_ (.Y(_07574_),
    .A(_07567_),
    .B(_07571_));
 sg13g2_nor3_2 _13383_ (.A(net5586),
    .B(_07028_),
    .C(_07039_),
    .Y(_07575_));
 sg13g2_or3_1 _13384_ (.A(net5586),
    .B(_07028_),
    .C(_07039_),
    .X(_07576_));
 sg13g2_nor4_2 _13385_ (.A(net5585),
    .B(_07028_),
    .C(_07037_),
    .Y(_07577_),
    .D(_07039_));
 sg13g2_nand2_2 _13386_ (.Y(_07578_),
    .A(_07038_),
    .B(_07575_));
 sg13g2_nor2_1 _13387_ (.A(net5574),
    .B(net5294),
    .Y(_07579_));
 sg13g2_nor4_2 _13388_ (.A(net5574),
    .B(net5294),
    .C(_07303_),
    .Y(_07580_),
    .D(net4860));
 sg13g2_nand3_1 _13389_ (.B(net4954),
    .C(_07579_),
    .A(net5342),
    .Y(_07581_));
 sg13g2_mux2_1 _13390_ (.A0(net5800),
    .A1(net5804),
    .S(net4978),
    .X(_07582_));
 sg13g2_mux2_1 _13391_ (.A0(net5797),
    .A1(net5798),
    .S(net4978),
    .X(_07583_));
 sg13g2_mux2_1 _13392_ (.A0(_07582_),
    .A1(_07583_),
    .S(net4996),
    .X(_07584_));
 sg13g2_mux2_1 _13393_ (.A0(net5791),
    .A1(net5794),
    .S(net4979),
    .X(_07585_));
 sg13g2_nor2_1 _13394_ (.A(net5788),
    .B(net4981),
    .Y(_07586_));
 sg13g2_a21oi_1 _13395_ (.A1(_06573_),
    .A2(net4981),
    .Y(_07587_),
    .B1(_07586_));
 sg13g2_mux2_1 _13396_ (.A0(_07585_),
    .A1(_07587_),
    .S(net4996),
    .X(_07588_));
 sg13g2_mux2_1 _13397_ (.A0(_07584_),
    .A1(_07588_),
    .S(net5004),
    .X(_07589_));
 sg13g2_nor2_1 _13398_ (.A(net5822),
    .B(net4975),
    .Y(_07590_));
 sg13g2_mux4_1 _13399_ (.S0(net4975),
    .A0(net5822),
    .A1(net5825),
    .A2(net5816),
    .A3(net5820),
    .S1(net4995),
    .X(_07591_));
 sg13g2_mux2_1 _13400_ (.A0(net5806),
    .A1(net5807),
    .S(net4978),
    .X(_07592_));
 sg13g2_mux4_1 _13401_ (.S0(net4996),
    .A0(net5810),
    .A1(net5805),
    .A2(net5813),
    .A3(net5807),
    .S1(net4978),
    .X(_07593_));
 sg13g2_mux2_1 _13402_ (.A0(_07591_),
    .A1(_07593_),
    .S(net5003),
    .X(_07594_));
 sg13g2_mux2_1 _13403_ (.A0(_07589_),
    .A1(_07594_),
    .S(net4967),
    .X(_07595_));
 sg13g2_nor3_2 _13404_ (.A(_06582_),
    .B(net4992),
    .C(net4986),
    .Y(_07596_));
 sg13g2_nand2_1 _13405_ (.Y(_07597_),
    .A(net5007),
    .B(_07596_));
 sg13g2_nand3_1 _13406_ (.B(net4958),
    .C(_07596_),
    .A(net5007),
    .Y(_07598_));
 sg13g2_nand2_1 _13407_ (.Y(_07599_),
    .A(_07292_),
    .B(_07598_));
 sg13g2_nor2_1 _13408_ (.A(net5754),
    .B(_07292_),
    .Y(_07600_));
 sg13g2_nor2_2 _13409_ (.A(net5208),
    .B(net4858),
    .Y(_07601_));
 sg13g2_nand2_1 _13410_ (.Y(_07602_),
    .A(net5574),
    .B(net5342));
 sg13g2_nor2_2 _13411_ (.A(net5294),
    .B(_07602_),
    .Y(_07603_));
 sg13g2_nand2b_2 _13412_ (.Y(_07604_),
    .B(_07299_),
    .A_N(_07602_));
 sg13g2_nor3_1 _13413_ (.A(_07600_),
    .B(_07601_),
    .C(_07604_),
    .Y(_07605_));
 sg13g2_nor2_2 _13414_ (.A(net5382),
    .B(net5583),
    .Y(_07606_));
 sg13g2_nand2_2 _13415_ (.Y(_07607_),
    .A(net5574),
    .B(_07606_));
 sg13g2_nor3_2 _13416_ (.A(net5382),
    .B(_06552_),
    .C(net5379),
    .Y(_07608_));
 sg13g2_nand3_1 _13417_ (.B(net5583),
    .C(net5574),
    .A(net5582),
    .Y(_07609_));
 sg13g2_o21ai_1 _13418_ (.B1(_07607_),
    .Y(_07610_),
    .A1(_07568_),
    .A2(_07609_));
 sg13g2_o21ai_1 _13419_ (.B1(net5200),
    .Y(_07611_),
    .A1(_07568_),
    .A2(_07607_));
 sg13g2_nor2_1 _13420_ (.A(net5294),
    .B(_07609_),
    .Y(_07612_));
 sg13g2_nor2_2 _13421_ (.A(net5294),
    .B(_07607_),
    .Y(_07613_));
 sg13g2_a21o_1 _13422_ (.A2(_07610_),
    .A1(net5754),
    .B1(_07611_),
    .X(_07614_));
 sg13g2_nor4_2 _13423_ (.A(net5582),
    .B(net5584),
    .C(net5380),
    .Y(_07615_),
    .D(_07298_));
 sg13g2_nand3_1 _13424_ (.B(_07036_),
    .C(_07299_),
    .A(net5574),
    .Y(_07616_));
 sg13g2_a221oi_1 _13425_ (.B2(_07570_),
    .C1(_07614_),
    .B1(net5186),
    .A1(_07599_),
    .Y(_07617_),
    .A2(_07605_));
 sg13g2_mux2_1 _13426_ (.A0(net5766),
    .A1(net5769),
    .S(net4985),
    .X(_07618_));
 sg13g2_mux2_1 _13427_ (.A0(net5761),
    .A1(net5764),
    .S(net4984),
    .X(_07619_));
 sg13g2_mux2_1 _13428_ (.A0(_07618_),
    .A1(_07619_),
    .S(net4998),
    .X(_07620_));
 sg13g2_nor2_1 _13429_ (.A(net5757),
    .B(net4985),
    .Y(_07621_));
 sg13g2_a21oi_1 _13430_ (.A1(_06580_),
    .A2(net4985),
    .Y(_07622_),
    .B1(_07621_));
 sg13g2_nand2_1 _13431_ (.Y(_07623_),
    .A(net4992),
    .B(_07622_));
 sg13g2_nor2_1 _13432_ (.A(net5015),
    .B(_07596_),
    .Y(_07624_));
 sg13g2_nand3_1 _13433_ (.B(net5001),
    .C(net4986),
    .A(net5756),
    .Y(_07625_));
 sg13g2_nand3_1 _13434_ (.B(_07624_),
    .C(_07625_),
    .A(_07623_),
    .Y(_07626_));
 sg13g2_o21ai_1 _13435_ (.B1(_07626_),
    .Y(_07627_),
    .A1(net5007),
    .A2(_07620_));
 sg13g2_nor4_1 _13436_ (.A(net5575),
    .B(_07298_),
    .C(_07303_),
    .D(net4954),
    .Y(_07628_));
 sg13g2_nand3_1 _13437_ (.B(net4860),
    .C(_07579_),
    .A(net5342),
    .Y(_07629_));
 sg13g2_nor2_1 _13438_ (.A(net5783),
    .B(net4983),
    .Y(_07630_));
 sg13g2_a21oi_1 _13439_ (.A1(_06574_),
    .A2(net4983),
    .Y(_07631_),
    .B1(_07630_));
 sg13g2_mux2_1 _13440_ (.A0(net5778),
    .A1(net5781),
    .S(net4983),
    .X(_07632_));
 sg13g2_mux2_1 _13441_ (.A0(_07631_),
    .A1(_07632_),
    .S(net5002),
    .X(_07633_));
 sg13g2_nand2_1 _13442_ (.Y(_07634_),
    .A(_06578_),
    .B(net4986));
 sg13g2_o21ai_1 _13443_ (.B1(_07634_),
    .Y(_07635_),
    .A1(net5775),
    .A2(net4986));
 sg13g2_nor2_1 _13444_ (.A(net5771),
    .B(net4985),
    .Y(_07636_));
 sg13g2_a21oi_1 _13445_ (.A1(_06579_),
    .A2(net4985),
    .Y(_07637_),
    .B1(_07636_));
 sg13g2_nand2_1 _13446_ (.Y(_07638_),
    .A(net4998),
    .B(_07637_));
 sg13g2_o21ai_1 _13447_ (.B1(_07638_),
    .Y(_07639_),
    .A1(net4998),
    .A2(_07635_));
 sg13g2_mux2_1 _13448_ (.A0(_07633_),
    .A1(_07639_),
    .S(net5006),
    .X(_07640_));
 sg13g2_o21ai_1 _13449_ (.B1(net4853),
    .Y(_07641_),
    .A1(net4956),
    .A2(_07640_));
 sg13g2_a21oi_1 _13450_ (.A1(net4956),
    .A2(_07627_),
    .Y(_07642_),
    .B1(_07641_));
 sg13g2_a21oi_1 _13451_ (.A1(net4786),
    .A2(_07595_),
    .Y(_07643_),
    .B1(_07642_));
 sg13g2_a21oi_1 _13452_ (.A1(_07617_),
    .A2(_07643_),
    .Y(_07644_),
    .B1(net5292));
 sg13g2_o21ai_1 _13453_ (.B1(_07644_),
    .Y(_07645_),
    .A1(net5204),
    .A2(_07574_));
 sg13g2_nand2_1 _13454_ (.Y(_07646_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[31] ),
    .B(net5292));
 sg13g2_a21oi_1 _13455_ (.A1(_07645_),
    .A2(_07646_),
    .Y(_07647_),
    .B1(net5314));
 sg13g2_o21ai_1 _13456_ (.B1(net5218),
    .Y(_07648_),
    .A1(net5225),
    .A2(_07287_));
 sg13g2_nor2_2 _13457_ (.A(_07029_),
    .B(_07294_),
    .Y(_07649_));
 sg13g2_or3_1 _13458_ (.A(_06550_),
    .B(_07029_),
    .C(net5344),
    .X(_07650_));
 sg13g2_nand3_1 _13459_ (.B(\fpga_top.bus_gather.i_read_adr[3] ),
    .C(net5597),
    .A(\fpga_top.bus_gather.i_read_adr[2] ),
    .Y(_07651_));
 sg13g2_and4_1 _13460_ (.A(\fpga_top.bus_gather.i_read_adr[2] ),
    .B(\fpga_top.bus_gather.i_read_adr[3] ),
    .C(net5597),
    .D(\fpga_top.bus_gather.i_read_adr[5] ),
    .X(_07652_));
 sg13g2_nand3_1 _13461_ (.B(\fpga_top.bus_gather.i_read_adr[7] ),
    .C(_07652_),
    .A(net5596),
    .Y(_07653_));
 sg13g2_nand4_1 _13462_ (.B(\fpga_top.bus_gather.i_read_adr[7] ),
    .C(net5595),
    .A(net5596),
    .Y(_07654_),
    .D(_07652_));
 sg13g2_nor2_1 _13463_ (.A(_06592_),
    .B(_07654_),
    .Y(_07655_));
 sg13g2_nand3_1 _13464_ (.B(\fpga_top.bus_gather.i_read_adr[11] ),
    .C(_07655_),
    .A(\fpga_top.bus_gather.i_read_adr[10] ),
    .Y(_07656_));
 sg13g2_nor2_1 _13465_ (.A(_06599_),
    .B(_07656_),
    .Y(_07657_));
 sg13g2_nand2_1 _13466_ (.Y(_07658_),
    .A(\fpga_top.bus_gather.i_read_adr[13] ),
    .B(_07657_));
 sg13g2_nand3_1 _13467_ (.B(\fpga_top.bus_gather.i_read_adr[14] ),
    .C(_07657_),
    .A(\fpga_top.bus_gather.i_read_adr[13] ),
    .Y(_07659_));
 sg13g2_nor2_1 _13468_ (.A(_06605_),
    .B(_07659_),
    .Y(_07660_));
 sg13g2_nand3_1 _13469_ (.B(\fpga_top.bus_gather.i_read_adr[17] ),
    .C(_07660_),
    .A(net5593),
    .Y(_07661_));
 sg13g2_nor2_2 _13470_ (.A(_06614_),
    .B(_07661_),
    .Y(_07662_));
 sg13g2_nand3_1 _13471_ (.B(\fpga_top.bus_gather.i_read_adr[20] ),
    .C(_07662_),
    .A(\fpga_top.bus_gather.i_read_adr[19] ),
    .Y(_07663_));
 sg13g2_nor2_1 _13472_ (.A(_06623_),
    .B(_07663_),
    .Y(_07664_));
 sg13g2_nand3_1 _13473_ (.B(\fpga_top.bus_gather.i_read_adr[23] ),
    .C(_07664_),
    .A(net5591),
    .Y(_07665_));
 sg13g2_nor2_1 _13474_ (.A(_06629_),
    .B(_07665_),
    .Y(_07666_));
 sg13g2_nand3_1 _13475_ (.B(\fpga_top.bus_gather.i_read_adr[26] ),
    .C(_07666_),
    .A(\fpga_top.bus_gather.i_read_adr[25] ),
    .Y(_07667_));
 sg13g2_nor2_1 _13476_ (.A(_06636_),
    .B(_07667_),
    .Y(_07668_));
 sg13g2_nand3_1 _13477_ (.B(\fpga_top.bus_gather.i_read_adr[29] ),
    .C(_07668_),
    .A(net5590),
    .Y(_07669_));
 sg13g2_or2_1 _13478_ (.X(_07670_),
    .B(_07669_),
    .A(_06643_));
 sg13g2_xnor2_1 _13479_ (.Y(_07671_),
    .A(_06646_),
    .B(_07670_));
 sg13g2_a21oi_1 _13480_ (.A1(net5214),
    .A2(_07671_),
    .Y(_07672_),
    .B1(net5182));
 sg13g2_o21ai_1 _13481_ (.B1(_07672_),
    .Y(_07673_),
    .A1(_07647_),
    .A2(_07648_));
 sg13g2_nand2_2 _13482_ (.Y(_07674_),
    .A(net5569),
    .B(net5177));
 sg13g2_nand2_2 _13483_ (.Y(_07675_),
    .A(_07673_),
    .B(_07674_));
 sg13g2_xnor2_1 _13484_ (.Y(_07676_),
    .A(_07046_),
    .B(_07282_));
 sg13g2_o21ai_1 _13485_ (.B1(net5209),
    .Y(_07677_),
    .A1(_06582_),
    .A2(net4959));
 sg13g2_nor2_1 _13486_ (.A(net5755),
    .B(net5009),
    .Y(_07678_));
 sg13g2_nor2_1 _13487_ (.A(_06582_),
    .B(net4999),
    .Y(_07679_));
 sg13g2_mux2_1 _13488_ (.A0(net5756),
    .A1(net5755),
    .S(net4982),
    .X(_07680_));
 sg13g2_a21o_1 _13489_ (.A2(_07680_),
    .A1(net4999),
    .B1(_07679_),
    .X(_07681_));
 sg13g2_inv_1 _13490_ (.Y(_07682_),
    .A(_07681_));
 sg13g2_mux2_1 _13491_ (.A0(net5754),
    .A1(_07681_),
    .S(net5008),
    .X(_07683_));
 sg13g2_a21oi_1 _13492_ (.A1(net4959),
    .A2(_07683_),
    .Y(_07684_),
    .B1(_07677_));
 sg13g2_inv_1 _13493_ (.Y(_07685_),
    .A(_07684_));
 sg13g2_a21oi_1 _13494_ (.A1(net4952),
    .A2(_07600_),
    .Y(_07686_),
    .B1(net5190));
 sg13g2_nor2b_2 _13495_ (.A(_07601_),
    .B_N(_07686_),
    .Y(_07687_));
 sg13g2_o21ai_1 _13496_ (.B1(_07686_),
    .Y(_07688_),
    .A1(net5208),
    .A2(net4858));
 sg13g2_nor2_2 _13497_ (.A(net5208),
    .B(net4959),
    .Y(_07689_));
 sg13g2_nand3_1 _13498_ (.B(net4999),
    .C(_07680_),
    .A(net5008),
    .Y(_07690_));
 sg13g2_o21ai_1 _13499_ (.B1(_07292_),
    .Y(_07691_),
    .A1(net4971),
    .A2(_07690_));
 sg13g2_nand2_1 _13500_ (.Y(_07692_),
    .A(net4756),
    .B(_07691_));
 sg13g2_a21oi_1 _13501_ (.A1(net4858),
    .A2(_07684_),
    .Y(_07693_),
    .B1(_07692_));
 sg13g2_nand2b_1 _13502_ (.Y(_07694_),
    .B(net4978),
    .A_N(net5806));
 sg13g2_o21ai_1 _13503_ (.B1(_07694_),
    .Y(_07695_),
    .A1(net5803),
    .A2(net4978));
 sg13g2_nor2_1 _13504_ (.A(net5798),
    .B(net4975),
    .Y(_07696_));
 sg13g2_a21oi_1 _13505_ (.A1(_06567_),
    .A2(net4975),
    .Y(_07697_),
    .B1(_07696_));
 sg13g2_nor2_1 _13506_ (.A(net4990),
    .B(_07697_),
    .Y(_07698_));
 sg13g2_a21oi_1 _13507_ (.A1(net4991),
    .A2(_07695_),
    .Y(_07699_),
    .B1(_07698_));
 sg13g2_nor2_1 _13508_ (.A(net5794),
    .B(net4976),
    .Y(_07700_));
 sg13g2_a21oi_1 _13509_ (.A1(_06572_),
    .A2(net4976),
    .Y(_07701_),
    .B1(_07700_));
 sg13g2_mux2_1 _13510_ (.A0(net5790),
    .A1(net5791),
    .S(net4980),
    .X(_07702_));
 sg13g2_mux2_1 _13511_ (.A0(_07701_),
    .A1(_07702_),
    .S(net4995),
    .X(_07703_));
 sg13g2_mux2_1 _13512_ (.A0(_07699_),
    .A1(_07703_),
    .S(net5003),
    .X(_07704_));
 sg13g2_nor2b_2 _13513_ (.A(net4977),
    .B_N(net5825),
    .Y(_07705_));
 sg13g2_nand2b_2 _13514_ (.Y(_07706_),
    .B(net5825),
    .A_N(net4976));
 sg13g2_mux2_1 _13515_ (.A0(net5820),
    .A1(net5823),
    .S(net4975),
    .X(_07707_));
 sg13g2_nand2_1 _13516_ (.Y(_07708_),
    .A(net4990),
    .B(_07706_));
 sg13g2_o21ai_1 _13517_ (.B1(_07708_),
    .Y(_07709_),
    .A1(net4990),
    .A2(_07707_));
 sg13g2_mux2_1 _13518_ (.A0(net5813),
    .A1(net5816),
    .S(net4975),
    .X(_07710_));
 sg13g2_mux2_1 _13519_ (.A0(net5808),
    .A1(net5810),
    .S(net4975),
    .X(_07711_));
 sg13g2_mux2_1 _13520_ (.A0(_07710_),
    .A1(_07711_),
    .S(net4995),
    .X(_07712_));
 sg13g2_nand2_1 _13521_ (.Y(_07713_),
    .A(net5003),
    .B(_07712_));
 sg13g2_o21ai_1 _13522_ (.B1(_07713_),
    .Y(_07714_),
    .A1(net5003),
    .A2(_07709_));
 sg13g2_mux2_1 _13523_ (.A0(_07704_),
    .A1(_07714_),
    .S(net4967),
    .X(_07715_));
 sg13g2_nand3_1 _13524_ (.B(_07311_),
    .C(net5288),
    .A(net5756),
    .Y(_07716_));
 sg13g2_o21ai_1 _13525_ (.B1(net5103),
    .Y(_07717_),
    .A1(net5756),
    .A2(_07311_));
 sg13g2_xnor2_1 _13526_ (.Y(_07718_),
    .A(_06581_),
    .B(_07311_));
 sg13g2_a22oi_1 _13527_ (.Y(_07719_),
    .B1(_07718_),
    .B2(net5186),
    .A2(_07715_),
    .A1(net4786));
 sg13g2_nand4_1 _13528_ (.B(_07716_),
    .C(_07717_),
    .A(net5202),
    .Y(_07720_),
    .D(_07719_));
 sg13g2_mux2_1 _13529_ (.A0(net5769),
    .A1(net5772),
    .S(net4984),
    .X(_07721_));
 sg13g2_mux2_1 _13530_ (.A0(net5764),
    .A1(net5766),
    .S(net4984),
    .X(_07722_));
 sg13g2_mux2_1 _13531_ (.A0(_07721_),
    .A1(_07722_),
    .S(net4998),
    .X(_07723_));
 sg13g2_nor2b_1 _13532_ (.A(net5762),
    .B_N(net4984),
    .Y(_07724_));
 sg13g2_nor2_1 _13533_ (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[28] ),
    .B(net4984),
    .Y(_07725_));
 sg13g2_mux2_1 _13534_ (.A0(net5786),
    .A1(net5787),
    .S(net4979),
    .X(_07726_));
 sg13g2_mux2_1 _13535_ (.A0(net5782),
    .A1(net5783),
    .S(net4982),
    .X(_07727_));
 sg13g2_mux2_1 _13536_ (.A0(_07726_),
    .A1(_07727_),
    .S(net5002),
    .X(_07728_));
 sg13g2_mux2_1 _13537_ (.A0(net5777),
    .A1(net5779),
    .S(net4983),
    .X(_07729_));
 sg13g2_mux2_1 _13538_ (.A0(net5774),
    .A1(net5775),
    .S(net4984),
    .X(_07730_));
 sg13g2_mux2_1 _13539_ (.A0(_07729_),
    .A1(_07730_),
    .S(net4998),
    .X(_07731_));
 sg13g2_mux2_1 _13540_ (.A0(_07728_),
    .A1(_07731_),
    .S(net5006),
    .X(_07732_));
 sg13g2_mux4_1 _13541_ (.S0(net5001),
    .A0(net5760),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[30] ),
    .A2(net5762),
    .A3(net5757),
    .S1(net4984),
    .X(_07733_));
 sg13g2_nand2_1 _13542_ (.Y(_07734_),
    .A(net5015),
    .B(_07723_));
 sg13g2_a21oi_1 _13543_ (.A1(net5007),
    .A2(_07733_),
    .Y(_07735_),
    .B1(net4969));
 sg13g2_o21ai_1 _13544_ (.B1(net4853),
    .Y(_07736_),
    .A1(net4958),
    .A2(_07732_));
 sg13g2_a21oi_1 _13545_ (.A1(_07734_),
    .A2(_07735_),
    .Y(_07737_),
    .B1(_07736_));
 sg13g2_or3_1 _13546_ (.A(_07693_),
    .B(_07720_),
    .C(_07737_),
    .X(_07738_));
 sg13g2_nor2b_1 _13547_ (.A(_07316_),
    .B_N(_07566_),
    .Y(_07739_));
 sg13g2_xnor2_1 _13548_ (.Y(_07740_),
    .A(_07565_),
    .B(_07739_));
 sg13g2_o21ai_1 _13549_ (.B1(_07738_),
    .Y(_07741_),
    .A1(net5202),
    .A2(_07740_));
 sg13g2_o21ai_1 _13550_ (.B1(net5226),
    .Y(_07742_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[30] ),
    .A2(net5194));
 sg13g2_a21oi_1 _13551_ (.A1(net5194),
    .A2(_07741_),
    .Y(_07743_),
    .B1(_07742_));
 sg13g2_o21ai_1 _13552_ (.B1(net5217),
    .Y(_07744_),
    .A1(net5226),
    .A2(_07676_));
 sg13g2_or2_1 _13553_ (.X(_07745_),
    .B(_07744_),
    .A(_07743_));
 sg13g2_xnor2_1 _13554_ (.Y(_07746_),
    .A(_06643_),
    .B(_07669_));
 sg13g2_a21oi_1 _13555_ (.A1(net5210),
    .A2(_07746_),
    .Y(_07747_),
    .B1(net5178));
 sg13g2_nand2_1 _13556_ (.Y(_07748_),
    .A(_07745_),
    .B(_07747_));
 sg13g2_nand2_1 _13557_ (.Y(_07749_),
    .A(\fpga_top.cpu_top.br_ofs[10] ),
    .B(net5177));
 sg13g2_a22oi_1 _13558_ (.Y(_07750_),
    .B1(_07745_),
    .B2(_07747_),
    .A2(net5177),
    .A1(\fpga_top.cpu_top.br_ofs[10] ));
 sg13g2_xnor2_1 _13559_ (.Y(_07751_),
    .A(_06644_),
    .B(_07750_));
 sg13g2_xor2_1 _13560_ (.B(_07280_),
    .A(_07276_),
    .X(_07752_));
 sg13g2_and3_1 _13561_ (.X(_07753_),
    .A(_07560_),
    .B(_07562_),
    .C(_07563_));
 sg13g2_o21ai_1 _13562_ (.B1(net5197),
    .Y(_07754_),
    .A1(_07564_),
    .A2(_07753_));
 sg13g2_mux2_1 _13563_ (.A0(net5757),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[30] ),
    .S(net4987),
    .X(_07755_));
 sg13g2_a21oi_1 _13564_ (.A1(net4999),
    .A2(_07755_),
    .Y(_07756_),
    .B1(_07679_));
 sg13g2_a21oi_1 _13565_ (.A1(net5008),
    .A2(_07756_),
    .Y(_07757_),
    .B1(_07678_));
 sg13g2_a21oi_1 _13566_ (.A1(net4961),
    .A2(_07757_),
    .Y(_07758_),
    .B1(_07677_));
 sg13g2_nor3_1 _13567_ (.A(_06582_),
    .B(net4998),
    .C(net4987),
    .Y(_07759_));
 sg13g2_a21oi_1 _13568_ (.A1(net4999),
    .A2(_07755_),
    .Y(_07760_),
    .B1(_07759_));
 sg13g2_nor2_1 _13569_ (.A(net5018),
    .B(_07760_),
    .Y(_07761_));
 sg13g2_a21oi_1 _13570_ (.A1(net4961),
    .A2(_07761_),
    .Y(_07762_),
    .B1(net5208));
 sg13g2_nand2b_1 _13571_ (.Y(_07763_),
    .B(net4756),
    .A_N(_07762_));
 sg13g2_a21oi_1 _13572_ (.A1(net4858),
    .A2(_07758_),
    .Y(_07764_),
    .B1(_07763_));
 sg13g2_mux2_1 _13573_ (.A0(_07582_),
    .A1(_07592_),
    .S(net4990),
    .X(_07765_));
 sg13g2_mux2_1 _13574_ (.A0(_07583_),
    .A1(_07585_),
    .S(net4995),
    .X(_07766_));
 sg13g2_mux2_1 _13575_ (.A0(_07765_),
    .A1(_07766_),
    .S(net5005),
    .X(_07767_));
 sg13g2_nor2_1 _13576_ (.A(net4966),
    .B(_07767_),
    .Y(_07768_));
 sg13g2_or3_1 _13577_ (.A(net4990),
    .B(_07395_),
    .C(_07590_),
    .X(_07769_));
 sg13g2_nor2_1 _13578_ (.A(net5003),
    .B(_07769_),
    .Y(_07770_));
 sg13g2_mux4_1 _13579_ (.S0(net4996),
    .A0(net5816),
    .A1(net5810),
    .A2(net5820),
    .A3(net5813),
    .S1(net4978),
    .X(_07771_));
 sg13g2_a21oi_1 _13580_ (.A1(net5003),
    .A2(_07771_),
    .Y(_07772_),
    .B1(_07770_));
 sg13g2_a21oi_2 _13581_ (.B1(_07768_),
    .Y(_07773_),
    .A2(_07772_),
    .A1(net4966));
 sg13g2_nand3_1 _13582_ (.B(_07317_),
    .C(net5288),
    .A(net5757),
    .Y(_07774_));
 sg13g2_o21ai_1 _13583_ (.B1(net5101),
    .Y(_07775_),
    .A1(net5757),
    .A2(_07317_));
 sg13g2_xor2_1 _13584_ (.B(_07317_),
    .A(net5757),
    .X(_07776_));
 sg13g2_a22oi_1 _13585_ (.Y(_07777_),
    .B1(_07776_),
    .B2(net5185),
    .A2(_07773_),
    .A1(_07580_));
 sg13g2_nand4_1 _13586_ (.B(_07774_),
    .C(_07775_),
    .A(net5202),
    .Y(_07778_),
    .D(_07777_));
 sg13g2_mux2_1 _13587_ (.A0(_07587_),
    .A1(_07631_),
    .S(net5002),
    .X(_07779_));
 sg13g2_nand2_1 _13588_ (.Y(_07780_),
    .A(net4994),
    .B(_07632_));
 sg13g2_o21ai_1 _13589_ (.B1(_07780_),
    .Y(_07781_),
    .A1(net4994),
    .A2(_07635_));
 sg13g2_mux2_1 _13590_ (.A0(_07779_),
    .A1(_07781_),
    .S(net5006),
    .X(_07782_));
 sg13g2_nor2_1 _13591_ (.A(net4958),
    .B(_07782_),
    .Y(_07783_));
 sg13g2_mux2_1 _13592_ (.A0(_07618_),
    .A1(_07637_),
    .S(net4992),
    .X(_07784_));
 sg13g2_nor2_1 _13593_ (.A(net4998),
    .B(_07619_),
    .Y(_07785_));
 sg13g2_o21ai_1 _13594_ (.B1(net5007),
    .Y(_07786_),
    .A1(net4993),
    .A2(_07622_));
 sg13g2_o21ai_1 _13595_ (.B1(net4958),
    .Y(_07787_),
    .A1(_07785_),
    .A2(_07786_));
 sg13g2_a21oi_1 _13596_ (.A1(net5015),
    .A2(_07784_),
    .Y(_07788_),
    .B1(_07787_));
 sg13g2_nor3_1 _13597_ (.A(net4784),
    .B(_07783_),
    .C(_07788_),
    .Y(_07789_));
 sg13g2_nor3_1 _13598_ (.A(_07764_),
    .B(_07778_),
    .C(_07789_),
    .Y(_07790_));
 sg13g2_nor2_1 _13599_ (.A(net5291),
    .B(_07790_),
    .Y(_07791_));
 sg13g2_a22oi_1 _13600_ (.Y(_07792_),
    .B1(_07754_),
    .B2(_07791_),
    .A2(net5290),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[29] ));
 sg13g2_o21ai_1 _13601_ (.B1(net5217),
    .Y(_07793_),
    .A1(net5311),
    .A2(_07792_));
 sg13g2_a21o_2 _13602_ (.A2(_07752_),
    .A1(net5311),
    .B1(_07793_),
    .X(_07794_));
 sg13g2_a21o_1 _13603_ (.A2(_07668_),
    .A1(\fpga_top.bus_gather.i_read_adr[28] ),
    .B1(\fpga_top.bus_gather.i_read_adr[29] ),
    .X(_07795_));
 sg13g2_nand2_2 _13604_ (.Y(_07796_),
    .A(_07669_),
    .B(_07795_));
 sg13g2_a21oi_1 _13605_ (.A1(net5214),
    .A2(_07796_),
    .Y(_07797_),
    .B1(net5180));
 sg13g2_a22oi_1 _13606_ (.Y(_07798_),
    .B1(_07794_),
    .B2(_07797_),
    .A2(net5180),
    .A1(net5570));
 sg13g2_nand2_1 _13607_ (.Y(_07799_),
    .A(_06548_),
    .B(net5181));
 sg13g2_nand2b_1 _13608_ (.Y(_07800_),
    .B(net5290),
    .A_N(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[22] ));
 sg13g2_a21o_1 _13609_ (.A2(_07516_),
    .A1(_07511_),
    .B1(_07334_),
    .X(_07801_));
 sg13g2_a22oi_1 _13610_ (.Y(_07802_),
    .B1(_07343_),
    .B2(_07801_),
    .A2(_07336_),
    .A1(_06578_));
 sg13g2_a21oi_1 _13611_ (.A1(_07325_),
    .A2(_07802_),
    .Y(_07803_),
    .B1(_07324_));
 sg13g2_xor2_1 _13612_ (.B(_07803_),
    .A(_07328_),
    .X(_07804_));
 sg13g2_nor2_2 _13613_ (.A(_07292_),
    .B(net4959),
    .Y(_07805_));
 sg13g2_nand2b_1 _13614_ (.Y(_07806_),
    .B(_07805_),
    .A_N(_07683_));
 sg13g2_mux2_1 _13615_ (.A0(net5769),
    .A1(net5766),
    .S(net4987),
    .X(_07807_));
 sg13g2_mux2_1 _13616_ (.A0(net5774),
    .A1(net5772),
    .S(net4987),
    .X(_07808_));
 sg13g2_mux2_1 _13617_ (.A0(_07807_),
    .A1(_07808_),
    .S(net4999),
    .X(_07809_));
 sg13g2_mux2_1 _13618_ (.A0(net5760),
    .A1(net5757),
    .S(net4987),
    .X(_07810_));
 sg13g2_mux2_1 _13619_ (.A0(net5764),
    .A1(net5761),
    .S(net4987),
    .X(_07811_));
 sg13g2_mux2_1 _13620_ (.A0(_07810_),
    .A1(_07811_),
    .S(net4999),
    .X(_07812_));
 sg13g2_mux2_1 _13621_ (.A0(_07809_),
    .A1(_07812_),
    .S(net5017),
    .X(_07813_));
 sg13g2_nand2_1 _13622_ (.Y(_07814_),
    .A(_07689_),
    .B(_07690_));
 sg13g2_o21ai_1 _13623_ (.B1(_07814_),
    .Y(_07815_),
    .A1(net4972),
    .A2(_07813_));
 sg13g2_nand2b_2 _13624_ (.Y(_07816_),
    .B(_07806_),
    .A_N(_07815_));
 sg13g2_a21oi_2 _13625_ (.B1(_07688_),
    .Y(_07817_),
    .A2(_07816_),
    .A1(net4858));
 sg13g2_mux2_1 _13626_ (.A0(_07704_),
    .A1(_07732_),
    .S(net4956),
    .X(_07818_));
 sg13g2_xnor2_1 _13627_ (.Y(_07819_),
    .A(_06579_),
    .B(_07326_));
 sg13g2_o21ai_1 _13628_ (.B1(net5101),
    .Y(_07820_),
    .A1(net5774),
    .A2(_07326_));
 sg13g2_nand3_1 _13629_ (.B(_07326_),
    .C(net5188),
    .A(net5774),
    .Y(_07821_));
 sg13g2_nand3_1 _13630_ (.B(_07820_),
    .C(_07821_),
    .A(net5195),
    .Y(_07822_));
 sg13g2_a21oi_1 _13631_ (.A1(net5186),
    .A2(_07819_),
    .Y(_07823_),
    .B1(_07822_));
 sg13g2_nand2_1 _13632_ (.Y(_07824_),
    .A(net4963),
    .B(_07714_));
 sg13g2_o21ai_1 _13633_ (.B1(_07823_),
    .Y(_07825_),
    .A1(_07581_),
    .A2(_07824_));
 sg13g2_a21oi_1 _13634_ (.A1(net4854),
    .A2(_07818_),
    .Y(_07826_),
    .B1(_07825_));
 sg13g2_o21ai_1 _13635_ (.B1(_07826_),
    .Y(_07827_),
    .A1(net5202),
    .A2(_07804_));
 sg13g2_o21ai_1 _13636_ (.B1(_07800_),
    .Y(_07828_),
    .A1(_07817_),
    .A2(_07827_));
 sg13g2_a21oi_1 _13637_ (.A1(_07183_),
    .A2(_07238_),
    .Y(_07829_),
    .B1(_07244_));
 sg13g2_a21o_1 _13638_ (.A2(_07238_),
    .A1(_07183_),
    .B1(_07244_),
    .X(_07830_));
 sg13g2_a21oi_1 _13639_ (.A1(_07208_),
    .A2(_07830_),
    .Y(_07831_),
    .B1(_07246_));
 sg13g2_xnor2_1 _13640_ (.Y(_07832_),
    .A(_07188_),
    .B(_07831_));
 sg13g2_o21ai_1 _13641_ (.B1(net5217),
    .Y(_07833_),
    .A1(net5226),
    .A2(_07832_));
 sg13g2_a21oi_1 _13642_ (.A1(net5226),
    .A2(_07828_),
    .Y(_07834_),
    .B1(_07833_));
 sg13g2_xnor2_1 _13643_ (.Y(_07835_),
    .A(net5591),
    .B(_07664_));
 sg13g2_o21ai_1 _13644_ (.B1(net5286),
    .Y(_07836_),
    .A1(net5217),
    .A2(_07835_));
 sg13g2_o21ai_1 _13645_ (.B1(_07799_),
    .Y(_07837_),
    .A1(_07834_),
    .A2(_07836_));
 sg13g2_xor2_1 _13646_ (.B(_07837_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[22] ),
    .X(_07838_));
 sg13g2_xnor2_1 _13647_ (.Y(_07839_),
    .A(_07325_),
    .B(_07802_));
 sg13g2_nor2b_1 _13648_ (.A(_07757_),
    .B_N(_07805_),
    .Y(_07840_));
 sg13g2_mux4_1 _13649_ (.S0(net4988),
    .A0(net5776),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[22] ),
    .A2(net5772),
    .A3(net5769),
    .S1(net4992),
    .X(_07841_));
 sg13g2_mux4_1 _13650_ (.S0(net4984),
    .A0(net5766),
    .A1(net5764),
    .A2(net5762),
    .A3(\fpga_top.cpu_top.execution.csr_array.rs1_sel[28] ),
    .S1(net4992),
    .X(_07842_));
 sg13g2_mux2_1 _13651_ (.A0(_07841_),
    .A1(_07842_),
    .S(net5016),
    .X(_07843_));
 sg13g2_nor2_1 _13652_ (.A(net4972),
    .B(_07843_),
    .Y(_07844_));
 sg13g2_nor2b_1 _13653_ (.A(_07761_),
    .B_N(_07689_),
    .Y(_07845_));
 sg13g2_nor3_1 _13654_ (.A(_07840_),
    .B(_07844_),
    .C(_07845_),
    .Y(_07846_));
 sg13g2_o21ai_1 _13655_ (.B1(_07687_),
    .Y(_07847_),
    .A1(net4952),
    .A2(_07846_));
 sg13g2_nor2_1 _13656_ (.A(net4956),
    .B(_07767_),
    .Y(_07848_));
 sg13g2_o21ai_1 _13657_ (.B1(net4854),
    .Y(_07849_),
    .A1(net4969),
    .A2(_07782_));
 sg13g2_nor2_1 _13658_ (.A(_07848_),
    .B(_07849_),
    .Y(_07850_));
 sg13g2_nor2_2 _13659_ (.A(net4968),
    .B(_07772_),
    .Y(_07851_));
 sg13g2_xor2_1 _13660_ (.B(_07321_),
    .A(net5775),
    .X(_07852_));
 sg13g2_o21ai_1 _13661_ (.B1(net5101),
    .Y(_07853_),
    .A1(net5775),
    .A2(_07321_));
 sg13g2_nand3_1 _13662_ (.B(_07321_),
    .C(net5188),
    .A(net5775),
    .Y(_07854_));
 sg13g2_a22oi_1 _13663_ (.Y(_07855_),
    .B1(_07852_),
    .B2(net5185),
    .A2(_07851_),
    .A1(net4786));
 sg13g2_nand4_1 _13664_ (.B(_07853_),
    .C(_07854_),
    .A(net5203),
    .Y(_07856_),
    .D(_07855_));
 sg13g2_nor2_1 _13665_ (.A(_07850_),
    .B(_07856_),
    .Y(_07857_));
 sg13g2_a221oi_1 _13666_ (.B2(_07857_),
    .C1(net5291),
    .B1(_07847_),
    .A1(net5196),
    .Y(_07858_),
    .A2(_07839_));
 sg13g2_a21o_1 _13667_ (.A2(net5289),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[21] ),
    .B1(net5311),
    .X(_07859_));
 sg13g2_o21ai_1 _13668_ (.B1(_07205_),
    .Y(_07860_),
    .A1(_07207_),
    .A2(_07829_));
 sg13g2_xor2_1 _13669_ (.B(_07860_),
    .A(_07201_),
    .X(_07861_));
 sg13g2_a21oi_1 _13670_ (.A1(net5312),
    .A2(_07861_),
    .Y(_07862_),
    .B1(net5215));
 sg13g2_o21ai_1 _13671_ (.B1(_07862_),
    .Y(_07863_),
    .A1(_07858_),
    .A2(_07859_));
 sg13g2_xnor2_1 _13672_ (.Y(_07864_),
    .A(_06623_),
    .B(_07663_));
 sg13g2_inv_1 _13673_ (.Y(_07865_),
    .A(_07864_));
 sg13g2_a21oi_1 _13674_ (.A1(net5215),
    .A2(_07865_),
    .Y(_07866_),
    .B1(net5182));
 sg13g2_a22oi_1 _13675_ (.Y(_07867_),
    .B1(_07863_),
    .B2(_07866_),
    .A2(net5181),
    .A1(_06559_));
 sg13g2_nor2_1 _13676_ (.A(_07522_),
    .B(_07525_),
    .Y(_07868_));
 sg13g2_xor2_1 _13677_ (.B(_07868_),
    .A(_07541_),
    .X(_07869_));
 sg13g2_mux2_1 _13678_ (.A0(_07680_),
    .A1(_07810_),
    .S(net4999),
    .X(_07870_));
 sg13g2_mux2_1 _13679_ (.A0(_07807_),
    .A1(_07811_),
    .S(net4994),
    .X(_07871_));
 sg13g2_mux2_1 _13680_ (.A0(_07870_),
    .A1(_07871_),
    .S(net5005),
    .X(_07872_));
 sg13g2_a22oi_1 _13681_ (.Y(_07873_),
    .B1(_07872_),
    .B2(net4955),
    .A2(_07805_),
    .A1(net5754));
 sg13g2_a21oi_1 _13682_ (.A1(net4858),
    .A2(_07873_),
    .Y(_07874_),
    .B1(_07688_));
 sg13g2_mux2_1 _13683_ (.A0(_07727_),
    .A1(_07729_),
    .S(net5002),
    .X(_07875_));
 sg13g2_inv_1 _13684_ (.Y(_07876_),
    .A(_07875_));
 sg13g2_mux2_1 _13685_ (.A0(_07721_),
    .A1(_07730_),
    .S(net4992),
    .X(_07877_));
 sg13g2_a21oi_1 _13686_ (.A1(net5016),
    .A2(_07876_),
    .Y(_07878_),
    .B1(net4969));
 sg13g2_o21ai_1 _13687_ (.B1(_07878_),
    .Y(_07879_),
    .A1(net5016),
    .A2(_07877_));
 sg13g2_mux2_1 _13688_ (.A0(_07697_),
    .A1(_07701_),
    .S(net4995),
    .X(_07880_));
 sg13g2_mux2_1 _13689_ (.A0(_07702_),
    .A1(_07726_),
    .S(net4995),
    .X(_07881_));
 sg13g2_mux2_1 _13690_ (.A0(_07880_),
    .A1(_07881_),
    .S(net5003),
    .X(_07882_));
 sg13g2_nand2_1 _13691_ (.Y(_07883_),
    .A(net4966),
    .B(_07882_));
 sg13g2_a21oi_1 _13692_ (.A1(_07879_),
    .A2(_07883_),
    .Y(_07884_),
    .B1(net4784));
 sg13g2_mux2_1 _13693_ (.A0(_07707_),
    .A1(_07710_),
    .S(net4995),
    .X(_07885_));
 sg13g2_mux4_1 _13694_ (.S0(net4997),
    .A0(net5808),
    .A1(net5803),
    .A2(net5810),
    .A3(net5805),
    .S1(net4975),
    .X(_07886_));
 sg13g2_mux2_1 _13695_ (.A0(_07885_),
    .A1(_07886_),
    .S(net5004),
    .X(_07887_));
 sg13g2_nand3_1 _13696_ (.B(net4997),
    .C(_07705_),
    .A(net5004),
    .Y(_07888_));
 sg13g2_nand2_1 _13697_ (.Y(_07889_),
    .A(net4964),
    .B(_07888_));
 sg13g2_o21ai_1 _13698_ (.B1(_07889_),
    .Y(_07890_),
    .A1(net4964),
    .A2(_07887_));
 sg13g2_nor2_1 _13699_ (.A(_07581_),
    .B(_07890_),
    .Y(_07891_));
 sg13g2_nand2b_1 _13700_ (.Y(_07892_),
    .B(_07538_),
    .A_N(net5769));
 sg13g2_nor2b_1 _13701_ (.A(_07538_),
    .B_N(net5770),
    .Y(_07893_));
 sg13g2_xor2_1 _13702_ (.B(_07538_),
    .A(net5769),
    .X(_07894_));
 sg13g2_a22oi_1 _13703_ (.Y(_07895_),
    .B1(_07893_),
    .B2(net5188),
    .A2(_07892_),
    .A1(net5101));
 sg13g2_o21ai_1 _13704_ (.B1(_07895_),
    .Y(_07896_),
    .A1(_07616_),
    .A2(_07894_));
 sg13g2_nor4_1 _13705_ (.A(_07874_),
    .B(_07884_),
    .C(_07891_),
    .D(_07896_),
    .Y(_07897_));
 sg13g2_o21ai_1 _13706_ (.B1(_07897_),
    .Y(_07898_),
    .A1(net5202),
    .A2(_07869_));
 sg13g2_nand2_1 _13707_ (.Y(_07899_),
    .A(net5194),
    .B(_07898_));
 sg13g2_a21oi_1 _13708_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[24] ),
    .A2(net5290),
    .Y(_07900_),
    .B1(net5313));
 sg13g2_xnor2_1 _13709_ (.Y(_07901_),
    .A(_07249_),
    .B(_07261_));
 sg13g2_a221oi_1 _13710_ (.B2(net5313),
    .C1(net5215),
    .B1(_07901_),
    .A1(_07899_),
    .Y(_07902_),
    .A2(_07900_));
 sg13g2_xnor2_1 _13711_ (.Y(_07903_),
    .A(_06629_),
    .B(_07665_));
 sg13g2_o21ai_1 _13712_ (.B1(net5287),
    .Y(_07904_),
    .A1(net5218),
    .A2(_07903_));
 sg13g2_nor2_1 _13713_ (.A(_07902_),
    .B(_07904_),
    .Y(_07905_));
 sg13g2_nand2_1 _13714_ (.Y(_07906_),
    .A(_06575_),
    .B(net5180));
 sg13g2_nor2b_2 _13715_ (.A(_07905_),
    .B_N(_07906_),
    .Y(_07907_));
 sg13g2_o21ai_1 _13716_ (.B1(_07906_),
    .Y(_07908_),
    .A1(_07902_),
    .A2(_07904_));
 sg13g2_a21oi_1 _13717_ (.A1(_07478_),
    .A2(_07482_),
    .Y(_07909_),
    .B1(_07362_));
 sg13g2_nor2_1 _13718_ (.A(_07361_),
    .B(_07909_),
    .Y(_07910_));
 sg13g2_a21oi_1 _13719_ (.A1(_07478_),
    .A2(_07482_),
    .Y(_07911_),
    .B1(_07368_));
 sg13g2_o21ai_1 _13720_ (.B1(_07351_),
    .Y(_07912_),
    .A1(_07369_),
    .A2(_07911_));
 sg13g2_and3_1 _13721_ (.X(_07913_),
    .A(_07349_),
    .B(_07357_),
    .C(_07912_));
 sg13g2_a21oi_1 _13722_ (.A1(_07349_),
    .A2(_07912_),
    .Y(_07914_),
    .B1(_07357_));
 sg13g2_nor3_1 _13723_ (.A(net5201),
    .B(_07913_),
    .C(_07914_),
    .Y(_07915_));
 sg13g2_mux2_1 _13724_ (.A0(net5777),
    .A1(net5776),
    .S(net4987),
    .X(_07916_));
 sg13g2_mux2_1 _13725_ (.A0(net5782),
    .A1(net5778),
    .S(net4982),
    .X(_07917_));
 sg13g2_mux2_1 _13726_ (.A0(_07916_),
    .A1(_07917_),
    .S(net5000),
    .X(_07918_));
 sg13g2_mux2_1 _13727_ (.A0(net5786),
    .A1(net5784),
    .S(net4982),
    .X(_07919_));
 sg13g2_mux2_1 _13728_ (.A0(net5790),
    .A1(net5787),
    .S(net4983),
    .X(_07920_));
 sg13g2_mux2_1 _13729_ (.A0(_07919_),
    .A1(_07920_),
    .S(net5000),
    .X(_07921_));
 sg13g2_mux2_1 _13730_ (.A0(_07918_),
    .A1(_07921_),
    .S(net5008),
    .X(_07922_));
 sg13g2_nor2_1 _13731_ (.A(net4960),
    .B(_07813_),
    .Y(_07923_));
 sg13g2_nor2_1 _13732_ (.A(net4950),
    .B(_07923_),
    .Y(_07924_));
 sg13g2_o21ai_1 _13733_ (.B1(_07924_),
    .Y(_07925_),
    .A1(net4971),
    .A2(_07922_));
 sg13g2_nand3_1 _13734_ (.B(_07685_),
    .C(_07691_),
    .A(net4950),
    .Y(_07926_));
 sg13g2_a21oi_2 _13735_ (.B1(net5190),
    .Y(_07927_),
    .A2(_07926_),
    .A1(_07925_));
 sg13g2_and2_1 _13736_ (.A(net4853),
    .B(_07715_),
    .X(_07928_));
 sg13g2_xnor2_1 _13737_ (.Y(_07929_),
    .A(_06573_),
    .B(_07353_));
 sg13g2_nand2_1 _13738_ (.Y(_07930_),
    .A(net5184),
    .B(_07929_));
 sg13g2_nand3_1 _13739_ (.B(_07353_),
    .C(net5189),
    .A(net5790),
    .Y(_07931_));
 sg13g2_o21ai_1 _13740_ (.B1(net5100),
    .Y(_07932_),
    .A1(net5790),
    .A2(_07353_));
 sg13g2_nand4_1 _13741_ (.B(_07930_),
    .C(_07931_),
    .A(net5195),
    .Y(_07933_),
    .D(_07932_));
 sg13g2_nor4_2 _13742_ (.A(_07915_),
    .B(_07927_),
    .C(_07928_),
    .Y(_07934_),
    .D(_07933_));
 sg13g2_nor2_1 _13743_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[14] ),
    .B(net5194),
    .Y(_07935_));
 sg13g2_o21ai_1 _13744_ (.B1(net5225),
    .Y(_07936_),
    .A1(_07934_),
    .A2(_07935_));
 sg13g2_nor2_1 _13745_ (.A(_07149_),
    .B(_07178_),
    .Y(_07937_));
 sg13g2_a21oi_1 _13746_ (.A1(_07171_),
    .A2(_07937_),
    .Y(_07938_),
    .B1(_07180_));
 sg13g2_xnor2_1 _13747_ (.Y(_07939_),
    .A(_07157_),
    .B(_07938_));
 sg13g2_a21oi_1 _13748_ (.A1(net5309),
    .A2(_07939_),
    .Y(_07940_),
    .B1(net5214));
 sg13g2_xnor2_1 _13749_ (.Y(_07941_),
    .A(_06603_),
    .B(_07658_));
 sg13g2_o21ai_1 _13750_ (.B1(net5286),
    .Y(_07942_),
    .A1(net5219),
    .A2(_07941_));
 sg13g2_a21oi_1 _13751_ (.A1(_07936_),
    .A2(_07940_),
    .Y(_07943_),
    .B1(_07942_));
 sg13g2_a21oi_2 _13752_ (.B1(_07943_),
    .Y(_07944_),
    .A2(net5180),
    .A1(net5380));
 sg13g2_xnor2_1 _13753_ (.Y(_07945_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[14] ),
    .B(_07944_));
 sg13g2_and2_1 _13754_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[13] ),
    .B(net5292),
    .X(_07946_));
 sg13g2_or3_1 _13755_ (.A(_07351_),
    .B(_07369_),
    .C(_07911_),
    .X(_07947_));
 sg13g2_nand2_1 _13756_ (.Y(_07948_),
    .A(_07912_),
    .B(_07947_));
 sg13g2_or2_1 _13757_ (.X(_07949_),
    .B(_07762_),
    .A(_07758_));
 sg13g2_mux4_1 _13758_ (.S0(net4988),
    .A0(net5793),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[14] ),
    .A2(net5788),
    .A3(\fpga_top.cpu_top.execution.csr_array.rs1_sel[16] ),
    .S1(net4993),
    .X(_07950_));
 sg13g2_mux4_1 _13759_ (.S0(net4988),
    .A0(net5784),
    .A1(net5782),
    .A2(net5779),
    .A3(net5777),
    .S1(net4993),
    .X(_07951_));
 sg13g2_mux2_1 _13760_ (.A0(_07950_),
    .A1(_07951_),
    .S(net5018),
    .X(_07952_));
 sg13g2_nand2_1 _13761_ (.Y(_07953_),
    .A(net4961),
    .B(_07952_));
 sg13g2_a21oi_1 _13762_ (.A1(net4970),
    .A2(_07843_),
    .Y(_07954_),
    .B1(net4950));
 sg13g2_a221oi_1 _13763_ (.B2(_07954_),
    .C1(net5190),
    .B1(_07953_),
    .A1(net4951),
    .Y(_07955_),
    .A2(_07949_));
 sg13g2_xor2_1 _13764_ (.B(_07346_),
    .A(net5791),
    .X(_07956_));
 sg13g2_nand3_1 _13765_ (.B(_07346_),
    .C(net5288),
    .A(net5791),
    .Y(_07957_));
 sg13g2_o21ai_1 _13766_ (.B1(net5100),
    .Y(_07958_),
    .A1(net5792),
    .A2(_07346_));
 sg13g2_a22oi_1 _13767_ (.Y(_07959_),
    .B1(_07956_),
    .B2(net5184),
    .A2(_07773_),
    .A1(net4855));
 sg13g2_nand4_1 _13768_ (.B(_07957_),
    .C(_07958_),
    .A(net5201),
    .Y(_07960_),
    .D(_07959_));
 sg13g2_o21ai_1 _13769_ (.B1(net5195),
    .Y(_07961_),
    .A1(_07955_),
    .A2(_07960_));
 sg13g2_a21oi_1 _13770_ (.A1(net5197),
    .A2(_07948_),
    .Y(_07962_),
    .B1(_07961_));
 sg13g2_o21ai_1 _13771_ (.B1(net5225),
    .Y(_07963_),
    .A1(_07946_),
    .A2(_07962_));
 sg13g2_o21ai_1 _13772_ (.B1(_07176_),
    .Y(_07964_),
    .A1(_07149_),
    .A2(_07178_));
 sg13g2_xnor2_1 _13773_ (.Y(_07965_),
    .A(_07171_),
    .B(_07964_));
 sg13g2_nor2_1 _13774_ (.A(net5225),
    .B(_07965_),
    .Y(_07966_));
 sg13g2_nor2_1 _13775_ (.A(net5214),
    .B(_07966_),
    .Y(_07967_));
 sg13g2_xnor2_1 _13776_ (.Y(_07968_),
    .A(\fpga_top.bus_gather.i_read_adr[13] ),
    .B(_07657_));
 sg13g2_a221oi_1 _13777_ (.B2(net5214),
    .C1(net5180),
    .B1(_07968_),
    .A1(_07963_),
    .Y(_07969_),
    .A2(_07967_));
 sg13g2_a21o_2 _13778_ (.A2(net5177),
    .A1(net5581),
    .B1(_07969_),
    .X(_07970_));
 sg13g2_and2_1 _13779_ (.A(net5017),
    .B(_07809_),
    .X(_07971_));
 sg13g2_a21oi_1 _13780_ (.A1(net5008),
    .A2(_07918_),
    .Y(_07972_),
    .B1(_07971_));
 sg13g2_nand2_1 _13781_ (.Y(_07973_),
    .A(net4971),
    .B(_07972_));
 sg13g2_mux2_1 _13782_ (.A0(net5795),
    .A1(net5792),
    .S(net4982),
    .X(_07974_));
 sg13g2_mux2_1 _13783_ (.A0(net5799),
    .A1(net5797),
    .S(net4983),
    .X(_07975_));
 sg13g2_mux2_1 _13784_ (.A0(_07974_),
    .A1(_07975_),
    .S(net5000),
    .X(_07976_));
 sg13g2_mux2_1 _13785_ (.A0(_07921_),
    .A1(_07976_),
    .S(net5009),
    .X(_07977_));
 sg13g2_o21ai_1 _13786_ (.B1(_07973_),
    .Y(_07978_),
    .A1(net4971),
    .A2(_07977_));
 sg13g2_nor2_1 _13787_ (.A(net5017),
    .B(_07812_),
    .Y(_07979_));
 sg13g2_a21oi_1 _13788_ (.A1(net5017),
    .A2(_07682_),
    .Y(_07980_),
    .B1(_07979_));
 sg13g2_a21oi_1 _13789_ (.A1(net4960),
    .A2(_07980_),
    .Y(_07981_),
    .B1(_07677_));
 sg13g2_a21oi_1 _13790_ (.A1(net5000),
    .A2(_07680_),
    .Y(_07982_),
    .B1(net5008));
 sg13g2_nor2_1 _13791_ (.A(_07979_),
    .B(_07982_),
    .Y(_07983_));
 sg13g2_a21oi_1 _13792_ (.A1(net4959),
    .A2(_07983_),
    .Y(_07984_),
    .B1(net5208));
 sg13g2_nor2_1 _13793_ (.A(_07981_),
    .B(_07984_),
    .Y(_07985_));
 sg13g2_a21oi_1 _13794_ (.A1(net4857),
    .A2(_07978_),
    .Y(_07986_),
    .B1(net5190));
 sg13g2_o21ai_1 _13795_ (.B1(_07986_),
    .Y(_07987_),
    .A1(net4857),
    .A2(_07985_));
 sg13g2_xnor2_1 _13796_ (.Y(_07988_),
    .A(_06571_),
    .B(_07449_));
 sg13g2_nand2_1 _13797_ (.Y(_07989_),
    .A(net5183),
    .B(_07988_));
 sg13g2_o21ai_1 _13798_ (.B1(net5099),
    .Y(_07990_),
    .A1(net5798),
    .A2(_07449_));
 sg13g2_nand3_1 _13799_ (.B(_07449_),
    .C(net5187),
    .A(net5798),
    .Y(_07991_));
 sg13g2_nand4_1 _13800_ (.B(_07989_),
    .C(_07990_),
    .A(net5200),
    .Y(_07992_),
    .D(_07991_));
 sg13g2_mux2_1 _13801_ (.A0(_07699_),
    .A1(_07712_),
    .S(net5012),
    .X(_07993_));
 sg13g2_or2_1 _13802_ (.X(_07994_),
    .B(_07709_),
    .A(net5012));
 sg13g2_nand2_1 _13803_ (.Y(_07995_),
    .A(net4967),
    .B(_07994_));
 sg13g2_o21ai_1 _13804_ (.B1(_07995_),
    .Y(_07996_),
    .A1(net4967),
    .A2(_07993_));
 sg13g2_o21ai_1 _13805_ (.B1(_07987_),
    .Y(_07997_),
    .A1(net4785),
    .A2(_07996_));
 sg13g2_o21ai_1 _13806_ (.B1(_07475_),
    .Y(_07998_),
    .A1(_07432_),
    .A2(_07435_));
 sg13g2_o21ai_1 _13807_ (.B1(_07480_),
    .Y(_07999_),
    .A1(_07464_),
    .A2(_07998_));
 sg13g2_a21oi_1 _13808_ (.A1(_07444_),
    .A2(_07999_),
    .Y(_08000_),
    .B1(_07441_));
 sg13g2_a21oi_1 _13809_ (.A1(_07457_),
    .A2(_08000_),
    .Y(_08001_),
    .B1(net5199));
 sg13g2_o21ai_1 _13810_ (.B1(_08001_),
    .Y(_08002_),
    .A1(_07457_),
    .A2(_08000_));
 sg13g2_o21ai_1 _13811_ (.B1(_08002_),
    .Y(_08003_),
    .A1(_07992_),
    .A2(_07997_));
 sg13g2_o21ai_1 _13812_ (.B1(net5223),
    .Y(_08004_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[10] ),
    .A2(net5194));
 sg13g2_a21oi_1 _13813_ (.A1(net5192),
    .A2(_08003_),
    .Y(_08005_),
    .B1(_08004_));
 sg13g2_a21o_1 _13814_ (.A2(_07142_),
    .A1(_07129_),
    .B1(_07144_),
    .X(_08006_));
 sg13g2_nand3_1 _13815_ (.B(_07142_),
    .C(_07144_),
    .A(_07129_),
    .Y(_08007_));
 sg13g2_and2_1 _13816_ (.A(_08006_),
    .B(_08007_),
    .X(_08008_));
 sg13g2_a21o_1 _13817_ (.A2(_08008_),
    .A1(net5309),
    .B1(net5213),
    .X(_08009_));
 sg13g2_xnor2_1 _13818_ (.Y(_08010_),
    .A(\fpga_top.bus_gather.i_read_adr[10] ),
    .B(_07655_));
 sg13g2_a21oi_1 _13819_ (.A1(net5213),
    .A2(_08010_),
    .Y(_08011_),
    .B1(net5179));
 sg13g2_o21ai_1 _13820_ (.B1(_08011_),
    .Y(_08012_),
    .A1(_08005_),
    .A2(_08009_));
 sg13g2_xnor2_1 _13821_ (.Y(_08013_),
    .A(_06595_),
    .B(_08012_));
 sg13g2_nor2_1 _13822_ (.A(_07490_),
    .B(_07492_),
    .Y(_08014_));
 sg13g2_xnor2_1 _13823_ (.Y(_08015_),
    .A(_07509_),
    .B(_08014_));
 sg13g2_mux2_1 _13824_ (.A0(_07808_),
    .A1(_07916_),
    .S(net5000),
    .X(_08016_));
 sg13g2_mux2_1 _13825_ (.A0(_07917_),
    .A1(_07919_),
    .S(net5002),
    .X(_08017_));
 sg13g2_mux2_1 _13826_ (.A0(_08016_),
    .A1(_08017_),
    .S(net5005),
    .X(_08018_));
 sg13g2_mux2_1 _13827_ (.A0(_07872_),
    .A1(_08018_),
    .S(net4957),
    .X(_08019_));
 sg13g2_nand2b_1 _13828_ (.Y(_08020_),
    .B(net4856),
    .A_N(_08019_));
 sg13g2_nor2_1 _13829_ (.A(net4963),
    .B(_07887_),
    .Y(_08021_));
 sg13g2_o21ai_1 _13830_ (.B1(net4853),
    .Y(_08022_),
    .A1(net4967),
    .A2(_07882_));
 sg13g2_nor2_1 _13831_ (.A(net4964),
    .B(_07888_),
    .Y(_08023_));
 sg13g2_xnor2_1 _13832_ (.Y(_08024_),
    .A(_06574_),
    .B(_07504_));
 sg13g2_nand3_1 _13833_ (.B(_07504_),
    .C(net5189),
    .A(net5786),
    .Y(_08025_));
 sg13g2_o21ai_1 _13834_ (.B1(net5100),
    .Y(_08026_),
    .A1(net5786),
    .A2(_07504_));
 sg13g2_nand3_1 _13835_ (.B(_08025_),
    .C(_08026_),
    .A(net5195),
    .Y(_08027_));
 sg13g2_a221oi_1 _13836_ (.B2(net5184),
    .C1(_08027_),
    .B1(_08024_),
    .A1(net4786),
    .Y(_08028_),
    .A2(_08023_));
 sg13g2_o21ai_1 _13837_ (.B1(_08028_),
    .Y(_08029_),
    .A1(_08021_),
    .A2(_08022_));
 sg13g2_a221oi_1 _13838_ (.B2(net4756),
    .C1(_08029_),
    .B1(_08020_),
    .A1(net5196),
    .Y(_08030_),
    .A2(_08015_));
 sg13g2_a21oi_1 _13839_ (.A1(_06607_),
    .A2(net5292),
    .Y(_08031_),
    .B1(_08030_));
 sg13g2_xnor2_1 _13840_ (.Y(_08032_),
    .A(_07183_),
    .B(_07229_));
 sg13g2_a21oi_1 _13841_ (.A1(net5314),
    .A2(_08032_),
    .Y(_08033_),
    .B1(net5214));
 sg13g2_o21ai_1 _13842_ (.B1(_08033_),
    .Y(_08034_),
    .A1(net5314),
    .A2(_08031_));
 sg13g2_xnor2_1 _13843_ (.Y(_08035_),
    .A(net5593),
    .B(_07660_));
 sg13g2_inv_1 _13844_ (.Y(_08036_),
    .A(_08035_));
 sg13g2_a21oi_1 _13845_ (.A1(net5214),
    .A2(_08036_),
    .Y(_08037_),
    .B1(net5182));
 sg13g2_a22oi_1 _13846_ (.Y(_08038_),
    .B1(_08034_),
    .B2(_08037_),
    .A2(net5182),
    .A1(_06608_));
 sg13g2_xnor2_1 _13847_ (.Y(_08039_),
    .A(_06609_),
    .B(_08038_));
 sg13g2_or3_1 _13848_ (.A(_07432_),
    .B(_07435_),
    .C(_07475_),
    .X(_08040_));
 sg13g2_and2_1 _13849_ (.A(_07998_),
    .B(_08040_),
    .X(_08041_));
 sg13g2_mux4_1 _13850_ (.S0(net4985),
    .A0(net5772),
    .A1(net5769),
    .A2(net5766),
    .A3(net5764),
    .S1(net4992),
    .X(_08042_));
 sg13g2_mux4_1 _13851_ (.S0(net4985),
    .A0(net5762),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[28] ),
    .A2(net5758),
    .A3(\fpga_top.cpu_top.execution.csr_array.rs1_sel[30] ),
    .S1(net4993),
    .X(_08043_));
 sg13g2_mux2_1 _13852_ (.A0(_08042_),
    .A1(_08043_),
    .S(net5016),
    .X(_08044_));
 sg13g2_nor2_1 _13853_ (.A(net4970),
    .B(_08044_),
    .Y(_08045_));
 sg13g2_a221oi_1 _13854_ (.B2(_07597_),
    .C1(_08045_),
    .B1(_07689_),
    .A1(net4970),
    .Y(_08046_),
    .A2(_07600_));
 sg13g2_mux4_1 _13855_ (.S0(net4988),
    .A0(net5788),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[16] ),
    .A2(net5784),
    .A3(net5782),
    .S1(net4993),
    .X(_08047_));
 sg13g2_mux4_1 _13856_ (.S0(net4988),
    .A0(net5779),
    .A1(net5777),
    .A2(net5776),
    .A3(\fpga_top.cpu_top.execution.csr_array.rs1_sel[22] ),
    .S1(net4992),
    .X(_08048_));
 sg13g2_mux2_1 _13857_ (.A0(_08047_),
    .A1(_08048_),
    .S(net5018),
    .X(_08049_));
 sg13g2_mux4_1 _13858_ (.S0(net4988),
    .A0(net5806),
    .A1(net5804),
    .A2(net5802),
    .A3(net5799),
    .S1(net4993),
    .X(_08050_));
 sg13g2_nor2_1 _13859_ (.A(net5018),
    .B(_08050_),
    .Y(_08051_));
 sg13g2_mux4_1 _13860_ (.S0(net4988),
    .A0(net5797),
    .A1(net5796),
    .A2(net5793),
    .A3(\fpga_top.cpu_top.execution.csr_array.rs1_sel[14] ),
    .S1(net4993),
    .X(_08052_));
 sg13g2_o21ai_1 _13861_ (.B1(net4961),
    .Y(_08053_),
    .A1(net5009),
    .A2(_08052_));
 sg13g2_o21ai_1 _13862_ (.B1(net4857),
    .Y(_08054_),
    .A1(_08051_),
    .A2(_08053_));
 sg13g2_a21o_1 _13863_ (.A2(_08049_),
    .A1(net4972),
    .B1(_08054_),
    .X(_08055_));
 sg13g2_o21ai_1 _13864_ (.B1(_08055_),
    .Y(_08056_),
    .A1(net4858),
    .A2(_08046_));
 sg13g2_nand2_1 _13865_ (.Y(_08057_),
    .A(net4963),
    .B(_07594_));
 sg13g2_inv_2 _13866_ (.Y(_08058_),
    .A(_08057_));
 sg13g2_xnor2_1 _13867_ (.Y(_08059_),
    .A(net5805),
    .B(_07469_));
 sg13g2_nand3_1 _13868_ (.B(_07470_),
    .C(net5187),
    .A(net5805),
    .Y(_08060_));
 sg13g2_o21ai_1 _13869_ (.B1(net5099),
    .Y(_08061_),
    .A1(net5806),
    .A2(_07470_));
 sg13g2_nand3_1 _13870_ (.B(_08060_),
    .C(_08061_),
    .A(net5198),
    .Y(_08062_));
 sg13g2_a221oi_1 _13871_ (.B2(net5183),
    .C1(_08062_),
    .B1(_08059_),
    .A1(net4855),
    .Y(_08063_),
    .A2(_08058_));
 sg13g2_o21ai_1 _13872_ (.B1(_08063_),
    .Y(_08064_),
    .A1(net5190),
    .A2(_08056_));
 sg13g2_o21ai_1 _13873_ (.B1(_08064_),
    .Y(_08065_),
    .A1(net5198),
    .A2(_08041_));
 sg13g2_o21ai_1 _13874_ (.B1(net5221),
    .Y(_08066_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[7] ),
    .A2(net5191));
 sg13g2_a21o_1 _13875_ (.A2(_08065_),
    .A1(net5191),
    .B1(_08066_),
    .X(_08067_));
 sg13g2_xnor2_1 _13876_ (.Y(_08068_),
    .A(_07118_),
    .B(_07120_));
 sg13g2_a21oi_1 _13877_ (.A1(net5307),
    .A2(_08068_),
    .Y(_08069_),
    .B1(net5210));
 sg13g2_a21o_1 _13878_ (.A2(_07652_),
    .A1(net5596),
    .B1(\fpga_top.bus_gather.i_read_adr[7] ),
    .X(_08070_));
 sg13g2_nand2_2 _13879_ (.Y(_08071_),
    .A(_07653_),
    .B(_08070_));
 sg13g2_a22oi_1 _13880_ (.Y(_08072_),
    .B1(_08071_),
    .B2(net5210),
    .A2(_08069_),
    .A1(_08067_));
 sg13g2_nand2_2 _13881_ (.Y(_08073_),
    .A(net5286),
    .B(_08072_));
 sg13g2_xnor2_1 _13882_ (.Y(_08074_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[7] ),
    .B(_08073_));
 sg13g2_nand2_1 _13883_ (.Y(_08075_),
    .A(_07406_),
    .B(_07408_));
 sg13g2_nand3_1 _13884_ (.B(_07408_),
    .C(_07416_),
    .A(_07406_),
    .Y(_08076_));
 sg13g2_a21oi_1 _13885_ (.A1(_07427_),
    .A2(_08076_),
    .Y(_08077_),
    .B1(_07426_));
 sg13g2_a21oi_1 _13886_ (.A1(_07428_),
    .A2(_08076_),
    .Y(_08078_),
    .B1(_08077_));
 sg13g2_mux4_1 _13887_ (.S0(net4982),
    .A0(net5811),
    .A1(net5808),
    .A2(net5806),
    .A3(net5804),
    .S1(net4994),
    .X(_08079_));
 sg13g2_inv_1 _13888_ (.Y(_08080_),
    .A(_08079_));
 sg13g2_mux4_1 _13889_ (.S0(net4987),
    .A0(net5802),
    .A1(net5799),
    .A2(\fpga_top.cpu_top.execution.csr_array.rs1_sel[11] ),
    .A3(net5796),
    .S1(net4994),
    .X(_08081_));
 sg13g2_nor2_1 _13890_ (.A(net5009),
    .B(_08081_),
    .Y(_08082_));
 sg13g2_o21ai_1 _13891_ (.B1(net4960),
    .Y(_08083_),
    .A1(net5017),
    .A2(_08079_));
 sg13g2_a21oi_1 _13892_ (.A1(net4972),
    .A2(_07952_),
    .Y(_08084_),
    .B1(net4951));
 sg13g2_o21ai_1 _13893_ (.B1(_08084_),
    .Y(_08085_),
    .A1(_08082_),
    .A2(_08083_));
 sg13g2_o21ai_1 _13894_ (.B1(_08085_),
    .Y(_08086_),
    .A1(net4857),
    .A2(_07846_));
 sg13g2_o21ai_1 _13895_ (.B1(net5100),
    .Y(_08087_),
    .A1(net5810),
    .A2(_07423_));
 sg13g2_nand3_1 _13896_ (.B(_07423_),
    .C(net5288),
    .A(net5810),
    .Y(_08088_));
 sg13g2_nand3_1 _13897_ (.B(_08087_),
    .C(_08088_),
    .A(net5198),
    .Y(_08089_));
 sg13g2_xnor2_1 _13898_ (.Y(_08090_),
    .A(_06565_),
    .B(_07423_));
 sg13g2_a221oi_1 _13899_ (.B2(net5183),
    .C1(_08089_),
    .B1(_08090_),
    .A1(net4855),
    .Y(_08091_),
    .A2(_07851_));
 sg13g2_o21ai_1 _13900_ (.B1(_08091_),
    .Y(_08092_),
    .A1(net5190),
    .A2(_08086_));
 sg13g2_o21ai_1 _13901_ (.B1(_08092_),
    .Y(_08093_),
    .A1(net5198),
    .A2(_08078_));
 sg13g2_o21ai_1 _13902_ (.B1(net5221),
    .Y(_08094_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[5] ),
    .A2(net5192));
 sg13g2_a21oi_1 _13903_ (.A1(net5191),
    .A2(_08093_),
    .Y(_08095_),
    .B1(_08094_));
 sg13g2_nand2_1 _13904_ (.Y(_08096_),
    .A(_07076_),
    .B(_07077_));
 sg13g2_xnor2_1 _13905_ (.Y(_08097_),
    .A(_07112_),
    .B(_08096_));
 sg13g2_a21o_1 _13906_ (.A2(_08097_),
    .A1(net5307),
    .B1(net5210),
    .X(_08098_));
 sg13g2_xnor2_1 _13907_ (.Y(_08099_),
    .A(_06587_),
    .B(_07651_));
 sg13g2_a21oi_1 _13908_ (.A1(net5210),
    .A2(_08099_),
    .Y(_08100_),
    .B1(net5177));
 sg13g2_o21ai_1 _13909_ (.B1(_08100_),
    .Y(_08101_),
    .A1(_08095_),
    .A2(_08098_));
 sg13g2_xnor2_1 _13910_ (.Y(_08102_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[5] ),
    .B(_08101_));
 sg13g2_nor2_1 _13911_ (.A(_08074_),
    .B(_08102_),
    .Y(_08103_));
 sg13g2_nor2_1 _13912_ (.A(net4955),
    .B(_08018_),
    .Y(_08104_));
 sg13g2_mux2_1 _13913_ (.A0(net5804),
    .A1(net5802),
    .S(net4982),
    .X(_08105_));
 sg13g2_mux2_1 _13914_ (.A0(_07975_),
    .A1(_08105_),
    .S(net5000),
    .X(_08106_));
 sg13g2_mux2_1 _13915_ (.A0(_07920_),
    .A1(_07974_),
    .S(net5002),
    .X(_08107_));
 sg13g2_mux2_1 _13916_ (.A0(_08106_),
    .A1(_08107_),
    .S(net5013),
    .X(_08108_));
 sg13g2_nor2_1 _13917_ (.A(net4968),
    .B(_08108_),
    .Y(_08109_));
 sg13g2_o21ai_1 _13918_ (.B1(net4856),
    .Y(_08110_),
    .A1(_08104_),
    .A2(_08109_));
 sg13g2_a21oi_1 _13919_ (.A1(net4950),
    .A2(_07873_),
    .Y(_08111_),
    .B1(net5190));
 sg13g2_nand2_2 _13920_ (.Y(_08112_),
    .A(_08110_),
    .B(_08111_));
 sg13g2_nand2_1 _13921_ (.Y(_08113_),
    .A(_06566_),
    .B(_07461_));
 sg13g2_xnor2_1 _13922_ (.Y(_08114_),
    .A(net5803),
    .B(_07461_));
 sg13g2_nor3_1 _13923_ (.A(_06566_),
    .B(_07461_),
    .C(_07609_),
    .Y(_08115_));
 sg13g2_or2_1 _13924_ (.X(_08116_),
    .B(_07890_),
    .A(net4784));
 sg13g2_a221oi_1 _13925_ (.B2(net5183),
    .C1(_08115_),
    .B1(_08114_),
    .A1(net5099),
    .Y(_08117_),
    .A2(_08113_));
 sg13g2_nand4_1 _13926_ (.B(_08112_),
    .C(_08116_),
    .A(net5199),
    .Y(_08118_),
    .D(_08117_));
 sg13g2_nand2_1 _13927_ (.Y(_08119_),
    .A(_07474_),
    .B(_07998_));
 sg13g2_xor2_1 _13928_ (.B(_08119_),
    .A(_07466_),
    .X(_08120_));
 sg13g2_o21ai_1 _13929_ (.B1(_08118_),
    .Y(_08121_),
    .A1(net5198),
    .A2(_08120_));
 sg13g2_o21ai_1 _13930_ (.B1(net5224),
    .Y(_08122_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[8] ),
    .A2(net5192));
 sg13g2_a21oi_1 _13931_ (.A1(net5191),
    .A2(_08121_),
    .Y(_08123_),
    .B1(_08122_));
 sg13g2_xnor2_1 _13932_ (.Y(_08124_),
    .A(_07122_),
    .B(_07127_));
 sg13g2_a21o_1 _13933_ (.A2(_08124_),
    .A1(net5307),
    .B1(net5211),
    .X(_08125_));
 sg13g2_xor2_1 _13934_ (.B(_07653_),
    .A(net5595),
    .X(_08126_));
 sg13g2_a21oi_1 _13935_ (.A1(net5210),
    .A2(_08126_),
    .Y(_08127_),
    .B1(net5178));
 sg13g2_o21ai_1 _13936_ (.B1(_08127_),
    .Y(_08128_),
    .A1(_08123_),
    .A2(_08125_));
 sg13g2_inv_2 _13937_ (.Y(_08129_),
    .A(_08128_));
 sg13g2_nand2_1 _13938_ (.Y(_08130_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[8] ),
    .B(_08128_));
 sg13g2_nand2_1 _13939_ (.Y(_08131_),
    .A(net5386),
    .B(net5212));
 sg13g2_mux4_1 _13940_ (.S0(net4980),
    .A0(net5820),
    .A1(net5816),
    .A2(net5813),
    .A3(net5811),
    .S1(net4991),
    .X(_08132_));
 sg13g2_nand2b_1 _13941_ (.Y(_08133_),
    .B(net5005),
    .A_N(_08132_));
 sg13g2_mux4_1 _13942_ (.S0(net4982),
    .A0(net5808),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[7] ),
    .A2(net5803),
    .A3(net5801),
    .S1(net4994),
    .X(_08134_));
 sg13g2_o21ai_1 _13943_ (.B1(_08133_),
    .Y(_08135_),
    .A1(net5005),
    .A2(_08134_));
 sg13g2_o21ai_1 _13944_ (.B1(net4857),
    .Y(_08136_),
    .A1(net4955),
    .A2(_07977_));
 sg13g2_a21oi_1 _13945_ (.A1(net4957),
    .A2(_08135_),
    .Y(_08137_),
    .B1(_08136_));
 sg13g2_and3_1 _13946_ (.X(_08138_),
    .A(_07292_),
    .B(net4960),
    .C(_07972_));
 sg13g2_nor2b_1 _13947_ (.A(_07983_),
    .B_N(_07689_),
    .Y(_08139_));
 sg13g2_mux4_1 _13948_ (.S0(net4960),
    .A0(_07681_),
    .A1(_07809_),
    .A2(_07812_),
    .A3(_07918_),
    .S1(net5008),
    .X(_08140_));
 sg13g2_o21ai_1 _13949_ (.B1(net4950),
    .Y(_08141_),
    .A1(_07292_),
    .A2(_08140_));
 sg13g2_nor3_1 _13950_ (.A(_08138_),
    .B(_08139_),
    .C(_08141_),
    .Y(_08142_));
 sg13g2_o21ai_1 _13951_ (.B1(_07603_),
    .Y(_08143_),
    .A1(_08137_),
    .A2(_08142_));
 sg13g2_xnor2_1 _13952_ (.Y(_08144_),
    .A(net5819),
    .B(_07381_));
 sg13g2_o21ai_1 _13953_ (.B1(net5197),
    .Y(_08145_),
    .A1(_07398_),
    .A2(_08144_));
 sg13g2_a21oi_1 _13954_ (.A1(_07398_),
    .A2(_08144_),
    .Y(_08146_),
    .B1(_08145_));
 sg13g2_nor3_1 _13955_ (.A(net4964),
    .B(net4784),
    .C(_07994_),
    .Y(_08147_));
 sg13g2_xnor2_1 _13956_ (.Y(_08148_),
    .A(net5819),
    .B(net5012));
 sg13g2_nor2_1 _13957_ (.A(_07616_),
    .B(_08148_),
    .Y(_08149_));
 sg13g2_nand3_1 _13958_ (.B(net5012),
    .C(net5187),
    .A(net5819),
    .Y(_08150_));
 sg13g2_o21ai_1 _13959_ (.B1(net5099),
    .Y(_08151_),
    .A1(net5819),
    .A2(net5012));
 sg13g2_nand3_1 _13960_ (.B(_08150_),
    .C(_08151_),
    .A(net5193),
    .Y(_08152_));
 sg13g2_nor4_1 _13961_ (.A(_08146_),
    .B(_08147_),
    .C(_08149_),
    .D(_08152_),
    .Y(_08153_));
 sg13g2_a22oi_1 _13962_ (.Y(_08154_),
    .B1(_08143_),
    .B2(_08153_),
    .A2(net5293),
    .A1(_06583_));
 sg13g2_xnor2_1 _13963_ (.Y(_08155_),
    .A(_07098_),
    .B(_07105_));
 sg13g2_a21oi_1 _13964_ (.A1(net5309),
    .A2(_08155_),
    .Y(_08156_),
    .B1(net5212));
 sg13g2_o21ai_1 _13965_ (.B1(_08156_),
    .Y(_08157_),
    .A1(net5308),
    .A2(_08154_));
 sg13g2_a21o_2 _13966_ (.A2(_08157_),
    .A1(_08131_),
    .B1(net5178),
    .X(_08158_));
 sg13g2_inv_2 _13967_ (.Y(_08159_),
    .A(_08158_));
 sg13g2_xor2_1 _13968_ (.B(_08158_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[2] ),
    .X(_08160_));
 sg13g2_mux2_1 _13969_ (.A0(_08042_),
    .A1(_08048_),
    .S(net5007),
    .X(_08161_));
 sg13g2_mux2_1 _13970_ (.A0(net5755),
    .A1(_08043_),
    .S(net5010),
    .X(_08162_));
 sg13g2_mux2_1 _13971_ (.A0(_08161_),
    .A1(_08162_),
    .S(net4970),
    .X(_08163_));
 sg13g2_nand3_1 _13972_ (.B(net4951),
    .C(_08163_),
    .A(net5208),
    .Y(_08164_));
 sg13g2_and2_1 _13973_ (.A(net5018),
    .B(_08047_),
    .X(_08165_));
 sg13g2_a21oi_1 _13974_ (.A1(net5009),
    .A2(_08052_),
    .Y(_08166_),
    .B1(_08165_));
 sg13g2_mux4_1 _13975_ (.S0(net4978),
    .A0(net5816),
    .A1(net5814),
    .A2(net5811),
    .A3(net5808),
    .S1(net4994),
    .X(_08167_));
 sg13g2_mux4_1 _13976_ (.S0(net4962),
    .A0(_08047_),
    .A1(_08050_),
    .A2(_08052_),
    .A3(_08167_),
    .S1(net5009),
    .X(_08168_));
 sg13g2_mux2_1 _13977_ (.A0(_07596_),
    .A1(_08043_),
    .S(net5010),
    .X(_08169_));
 sg13g2_mux2_1 _13978_ (.A0(_08161_),
    .A1(_08169_),
    .S(net4970),
    .X(_08170_));
 sg13g2_a22oi_1 _13979_ (.Y(_08171_),
    .B1(_08170_),
    .B2(_07601_),
    .A2(_08168_),
    .A1(net4859));
 sg13g2_a21oi_2 _13980_ (.B1(net5190),
    .Y(_08172_),
    .A2(_08171_),
    .A1(_08164_));
 sg13g2_nand2_2 _13981_ (.Y(_08173_),
    .A(net5004),
    .B(_07591_));
 sg13g2_nor3_1 _13982_ (.A(net4965),
    .B(net4784),
    .C(_08173_),
    .Y(_08174_));
 sg13g2_o21ai_1 _13983_ (.B1(net5099),
    .Y(_08175_),
    .A1(net5816),
    .A2(net4965));
 sg13g2_xnor2_1 _13984_ (.Y(_08176_),
    .A(net5817),
    .B(net4965));
 sg13g2_nor2_1 _13985_ (.A(_07616_),
    .B(_08176_),
    .Y(_08177_));
 sg13g2_o21ai_1 _13986_ (.B1(_07407_),
    .Y(_08178_),
    .A1(_07382_),
    .A2(_07399_));
 sg13g2_nand3_1 _13987_ (.B(net4964),
    .C(net5187),
    .A(net5816),
    .Y(_08179_));
 sg13g2_nand3_1 _13988_ (.B(_08175_),
    .C(_08179_),
    .A(net5201),
    .Y(_08180_));
 sg13g2_nor4_1 _13989_ (.A(_08172_),
    .B(_08174_),
    .C(_08177_),
    .D(_08180_),
    .Y(_08181_));
 sg13g2_a21oi_1 _13990_ (.A1(_07408_),
    .A2(_08178_),
    .Y(_08182_),
    .B1(net5198));
 sg13g2_nor2_1 _13991_ (.A(_08181_),
    .B(_08182_),
    .Y(_08183_));
 sg13g2_nor2_1 _13992_ (.A(net5293),
    .B(_08183_),
    .Y(_08184_));
 sg13g2_o21ai_1 _13993_ (.B1(net5224),
    .Y(_08185_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[3] ),
    .A2(net5191));
 sg13g2_xnor2_1 _13994_ (.Y(_08186_),
    .A(_07106_),
    .B(_07108_));
 sg13g2_a21oi_1 _13995_ (.A1(net5307),
    .A2(_08186_),
    .Y(_08187_),
    .B1(net5212));
 sg13g2_o21ai_1 _13996_ (.B1(_08187_),
    .Y(_08188_),
    .A1(_08184_),
    .A2(_08185_));
 sg13g2_xnor2_1 _13997_ (.Y(_08189_),
    .A(\fpga_top.bus_gather.i_read_adr[2] ),
    .B(\fpga_top.bus_gather.i_read_adr[3] ));
 sg13g2_a21oi_1 _13998_ (.A1(net5211),
    .A2(_08189_),
    .Y(_08190_),
    .B1(net5177));
 sg13g2_nand2_2 _13999_ (.Y(_08191_),
    .A(_08188_),
    .B(_08190_));
 sg13g2_inv_2 _14000_ (.Y(_08192_),
    .A(_08191_));
 sg13g2_xnor2_1 _14001_ (.Y(_08193_),
    .A(_07431_),
    .B(_08075_));
 sg13g2_a21oi_1 _14002_ (.A1(net5755),
    .A2(net5209),
    .Y(_08194_),
    .B1(net5005));
 sg13g2_nor2_1 _14003_ (.A(net5017),
    .B(_07870_),
    .Y(_08195_));
 sg13g2_nor2_1 _14004_ (.A(_08194_),
    .B(_08195_),
    .Y(_08196_));
 sg13g2_mux2_1 _14005_ (.A0(_07871_),
    .A1(_08016_),
    .S(net5005),
    .X(_08197_));
 sg13g2_mux2_1 _14006_ (.A0(_08196_),
    .A1(_08197_),
    .S(net4957),
    .X(_08198_));
 sg13g2_mux2_1 _14007_ (.A0(_08017_),
    .A1(_08107_),
    .S(net5011),
    .X(_08199_));
 sg13g2_nor2_1 _14008_ (.A(net5006),
    .B(_08106_),
    .Y(_08200_));
 sg13g2_mux4_1 _14009_ (.S0(net4979),
    .A0(net5813),
    .A1(net5811),
    .A2(net5808),
    .A3(\fpga_top.cpu_top.execution.csr_array.rs1_sel[7] ),
    .S1(net4991),
    .X(_08201_));
 sg13g2_o21ai_1 _14010_ (.B1(net4955),
    .Y(_08202_),
    .A1(net5013),
    .A2(_08201_));
 sg13g2_o21ai_1 _14011_ (.B1(net4859),
    .Y(_08203_),
    .A1(_08200_),
    .A2(_08202_));
 sg13g2_a21oi_1 _14012_ (.A1(net4968),
    .A2(_08199_),
    .Y(_08204_),
    .B1(_08203_));
 sg13g2_o21ai_1 _14013_ (.B1(_07603_),
    .Y(_08205_),
    .A1(net4856),
    .A2(_08198_));
 sg13g2_o21ai_1 _14014_ (.B1(net5012),
    .Y(_08206_),
    .A1(net4990),
    .A2(_07706_));
 sg13g2_o21ai_1 _14015_ (.B1(_08206_),
    .Y(_08207_),
    .A1(net5020),
    .A2(_07885_));
 sg13g2_nor2_1 _14016_ (.A(net4967),
    .B(_08207_),
    .Y(_08208_));
 sg13g2_xor2_1 _14017_ (.B(net4954),
    .A(net5814),
    .X(_08209_));
 sg13g2_o21ai_1 _14018_ (.B1(net5103),
    .Y(_08210_),
    .A1(net5813),
    .A2(net4953));
 sg13g2_nand3_1 _14019_ (.B(net4953),
    .C(net5188),
    .A(net5813),
    .Y(_08211_));
 sg13g2_nand3_1 _14020_ (.B(_08210_),
    .C(_08211_),
    .A(net5195),
    .Y(_08212_));
 sg13g2_a221oi_1 _14021_ (.B2(net5186),
    .C1(_08212_),
    .B1(_08209_),
    .A1(net4853),
    .Y(_08213_),
    .A2(_08208_));
 sg13g2_o21ai_1 _14022_ (.B1(_08213_),
    .Y(_08214_),
    .A1(_08204_),
    .A2(_08205_));
 sg13g2_a21oi_2 _14023_ (.B1(_08214_),
    .Y(_08215_),
    .A2(_08193_),
    .A1(net5197));
 sg13g2_o21ai_1 _14024_ (.B1(net5221),
    .Y(_08216_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[4] ),
    .A2(net5191));
 sg13g2_or2_1 _14025_ (.X(_08217_),
    .B(_08216_),
    .A(_08215_));
 sg13g2_xor2_1 _14026_ (.B(_07110_),
    .A(_07109_),
    .X(_08218_));
 sg13g2_a21oi_1 _14027_ (.A1(net5307),
    .A2(_08218_),
    .Y(_08219_),
    .B1(net5211));
 sg13g2_a21o_1 _14028_ (.A2(\fpga_top.bus_gather.i_read_adr[3] ),
    .A1(\fpga_top.bus_gather.i_read_adr[2] ),
    .B1(net5598),
    .X(_08220_));
 sg13g2_nand2_2 _14029_ (.Y(_08221_),
    .A(_07651_),
    .B(_08220_));
 sg13g2_a221oi_1 _14030_ (.B2(net5211),
    .C1(net5178),
    .B1(_08221_),
    .A1(_08217_),
    .Y(_08222_),
    .A2(_08219_));
 sg13g2_xnor2_1 _14031_ (.Y(_08223_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[4] ),
    .B(_08222_));
 sg13g2_xor2_1 _14032_ (.B(_08191_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[3] ),
    .X(_08224_));
 sg13g2_and4_1 _14033_ (.A(_08130_),
    .B(_08160_),
    .C(_08223_),
    .D(_08224_),
    .X(_08225_));
 sg13g2_nor2_1 _14034_ (.A(net5014),
    .B(_08134_),
    .Y(_08226_));
 sg13g2_o21ai_1 _14035_ (.B1(net4960),
    .Y(_08227_),
    .A1(net5008),
    .A2(_07976_));
 sg13g2_o21ai_1 _14036_ (.B1(net4857),
    .Y(_08228_),
    .A1(_08226_),
    .A2(_08227_));
 sg13g2_a21oi_1 _14037_ (.A1(net4971),
    .A2(_07922_),
    .Y(_08229_),
    .B1(_08228_));
 sg13g2_a21oi_2 _14038_ (.B1(_08229_),
    .Y(_08230_),
    .A2(_07816_),
    .A1(net4950));
 sg13g2_nor2b_1 _14039_ (.A(_07417_),
    .B_N(net5807),
    .Y(_08231_));
 sg13g2_nor2b_1 _14040_ (.A(net5807),
    .B_N(_07417_),
    .Y(_08232_));
 sg13g2_o21ai_1 _14041_ (.B1(net5198),
    .Y(_08233_),
    .A1(_07607_),
    .A2(_08232_));
 sg13g2_nor2_1 _14042_ (.A(_08231_),
    .B(_08232_),
    .Y(_08234_));
 sg13g2_a221oi_1 _14043_ (.B2(net5183),
    .C1(_08233_),
    .B1(_08234_),
    .A1(net5187),
    .Y(_08235_),
    .A2(_08231_));
 sg13g2_o21ai_1 _14044_ (.B1(_08235_),
    .Y(_08236_),
    .A1(net4785),
    .A2(_07824_));
 sg13g2_a21o_2 _14045_ (.A2(_08230_),
    .A1(_07603_),
    .B1(_08236_),
    .X(_08237_));
 sg13g2_a21oi_1 _14046_ (.A1(_07428_),
    .A2(_08076_),
    .Y(_08238_),
    .B1(_07425_));
 sg13g2_xnor2_1 _14047_ (.Y(_08239_),
    .A(_07421_),
    .B(_08238_));
 sg13g2_o21ai_1 _14048_ (.B1(_08237_),
    .Y(_08240_),
    .A1(net5199),
    .A2(_08239_));
 sg13g2_o21ai_1 _14049_ (.B1(net5221),
    .Y(_08241_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[6] ),
    .A2(net5191));
 sg13g2_a21oi_1 _14050_ (.A1(net5191),
    .A2(_08240_),
    .Y(_08242_),
    .B1(_08241_));
 sg13g2_xnor2_1 _14051_ (.Y(_08243_),
    .A(_07115_),
    .B(_07116_));
 sg13g2_a21o_1 _14052_ (.A2(_08243_),
    .A1(net5307),
    .B1(net5210),
    .X(_08244_));
 sg13g2_xnor2_1 _14053_ (.Y(_08245_),
    .A(net5596),
    .B(_07652_));
 sg13g2_a21oi_1 _14054_ (.A1(net5210),
    .A2(_08245_),
    .Y(_08246_),
    .B1(net5177));
 sg13g2_o21ai_1 _14055_ (.B1(_08246_),
    .Y(_08247_),
    .A1(_08242_),
    .A2(_08244_));
 sg13g2_a22oi_1 _14056_ (.Y(_08248_),
    .B1(_08247_),
    .B2(\fpga_top.uart_top.uart_rec_char.bpoint[6] ),
    .A2(_08129_),
    .A1(_06591_));
 sg13g2_a21oi_1 _14057_ (.A1(_07133_),
    .A2(_08006_),
    .Y(_08249_),
    .B1(_07145_));
 sg13g2_and3_1 _14058_ (.X(_08250_),
    .A(_07133_),
    .B(_07145_),
    .C(_08006_));
 sg13g2_nor2_1 _14059_ (.A(_08249_),
    .B(_08250_),
    .Y(_08251_));
 sg13g2_o21ai_1 _14060_ (.B1(net5308),
    .Y(_08252_),
    .A1(_08249_),
    .A2(_08250_));
 sg13g2_nand3_1 _14061_ (.B(_07478_),
    .C(_07482_),
    .A(_07362_),
    .Y(_08253_));
 sg13g2_nor2_1 _14062_ (.A(net5199),
    .B(_07909_),
    .Y(_08254_));
 sg13g2_nor2_1 _14063_ (.A(net4961),
    .B(_08161_),
    .Y(_08255_));
 sg13g2_a21oi_1 _14064_ (.A1(net4961),
    .A2(_08166_),
    .Y(_08256_),
    .B1(_08255_));
 sg13g2_a21oi_1 _14065_ (.A1(net4962),
    .A2(_08162_),
    .Y(_08257_),
    .B1(_07677_));
 sg13g2_a21oi_1 _14066_ (.A1(net4958),
    .A2(_08169_),
    .Y(_08258_),
    .B1(net5209));
 sg13g2_nor2_1 _14067_ (.A(_08257_),
    .B(_08258_),
    .Y(_08259_));
 sg13g2_mux2_1 _14068_ (.A0(_08256_),
    .A1(_08259_),
    .S(net4951),
    .X(_08260_));
 sg13g2_mux2_1 _14069_ (.A0(_07584_),
    .A1(_07593_),
    .S(net5013),
    .X(_08261_));
 sg13g2_nor2_1 _14070_ (.A(net4966),
    .B(_08261_),
    .Y(_08262_));
 sg13g2_a21oi_1 _14071_ (.A1(net4966),
    .A2(_08173_),
    .Y(_08263_),
    .B1(_08262_));
 sg13g2_nand3_1 _14072_ (.B(_07359_),
    .C(net5187),
    .A(net5797),
    .Y(_08264_));
 sg13g2_xnor2_1 _14073_ (.Y(_08265_),
    .A(_06572_),
    .B(_07359_));
 sg13g2_nand2_1 _14074_ (.Y(_08266_),
    .A(net5183),
    .B(_08265_));
 sg13g2_o21ai_1 _14075_ (.B1(net5099),
    .Y(_08267_),
    .A1(net5797),
    .A2(_07359_));
 sg13g2_nand3_1 _14076_ (.B(_08266_),
    .C(_08267_),
    .A(_08264_),
    .Y(_08268_));
 sg13g2_a221oi_1 _14077_ (.B2(net4855),
    .C1(_08268_),
    .B1(_08263_),
    .A1(_07603_),
    .Y(_08269_),
    .A2(_08260_));
 sg13g2_nand2_1 _14078_ (.Y(_08270_),
    .A(_07578_),
    .B(_08269_));
 sg13g2_a21o_2 _14079_ (.A2(_08254_),
    .A1(_08253_),
    .B1(_08270_),
    .X(_08271_));
 sg13g2_a21oi_1 _14080_ (.A1(_06596_),
    .A2(net5293),
    .Y(_08272_),
    .B1(net5308));
 sg13g2_a21oi_2 _14081_ (.B1(net5212),
    .Y(_08273_),
    .A2(_08272_),
    .A1(_08271_));
 sg13g2_a21o_1 _14082_ (.A2(_07655_),
    .A1(\fpga_top.bus_gather.i_read_adr[10] ),
    .B1(\fpga_top.bus_gather.i_read_adr[11] ),
    .X(_08274_));
 sg13g2_nand2_2 _14083_ (.Y(_08275_),
    .A(_07656_),
    .B(_08274_));
 sg13g2_nand3_1 _14084_ (.B(net5295),
    .C(net5286),
    .A(net5298),
    .Y(_08276_));
 sg13g2_a21o_1 _14085_ (.A2(_08275_),
    .A1(net5211),
    .B1(net5179),
    .X(_08277_));
 sg13g2_a21oi_2 _14086_ (.B1(_08277_),
    .Y(_08278_),
    .A2(_08273_),
    .A1(_08252_));
 sg13g2_a21o_2 _14087_ (.A2(_08273_),
    .A1(_08252_),
    .B1(_08277_),
    .X(_08279_));
 sg13g2_xnor2_1 _14088_ (.Y(_08280_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[11] ),
    .B(_08279_));
 sg13g2_xor2_1 _14089_ (.B(_07999_),
    .A(_07444_),
    .X(_08281_));
 sg13g2_mux2_1 _14090_ (.A0(_07841_),
    .A1(_07951_),
    .S(net5009),
    .X(_08282_));
 sg13g2_nor2_1 _14091_ (.A(net4959),
    .B(_08282_),
    .Y(_08283_));
 sg13g2_mux2_1 _14092_ (.A0(_07950_),
    .A1(_08081_),
    .S(net5010),
    .X(_08284_));
 sg13g2_o21ai_1 _14093_ (.B1(net4857),
    .Y(_08285_),
    .A1(net4971),
    .A2(_08284_));
 sg13g2_nor2_1 _14094_ (.A(_08283_),
    .B(_08285_),
    .Y(_08286_));
 sg13g2_nor2_1 _14095_ (.A(net5015),
    .B(_07842_),
    .Y(_08287_));
 sg13g2_a21oi_1 _14096_ (.A1(net5017),
    .A2(_07756_),
    .Y(_08288_),
    .B1(_08287_));
 sg13g2_a21oi_1 _14097_ (.A1(net4959),
    .A2(_08288_),
    .Y(_08289_),
    .B1(_07677_));
 sg13g2_a21oi_1 _14098_ (.A1(net5017),
    .A2(_07760_),
    .Y(_08290_),
    .B1(_08287_));
 sg13g2_nor2_1 _14099_ (.A(net5208),
    .B(_08290_),
    .Y(_08291_));
 sg13g2_nor3_1 _14100_ (.A(_07689_),
    .B(_08289_),
    .C(_08291_),
    .Y(_08292_));
 sg13g2_nor4_1 _14101_ (.A(net4857),
    .B(_07689_),
    .C(_08289_),
    .D(_08291_),
    .Y(_08293_));
 sg13g2_o21ai_1 _14102_ (.B1(_07603_),
    .Y(_08294_),
    .A1(_08286_),
    .A2(_08293_));
 sg13g2_mux2_1 _14103_ (.A0(_07765_),
    .A1(_07771_),
    .S(net5013),
    .X(_08295_));
 sg13g2_o21ai_1 _14104_ (.B1(net4968),
    .Y(_08296_),
    .A1(net5013),
    .A2(_07769_));
 sg13g2_o21ai_1 _14105_ (.B1(_08296_),
    .Y(_08297_),
    .A1(net4968),
    .A2(_08295_));
 sg13g2_or2_1 _14106_ (.X(_08298_),
    .B(_08297_),
    .A(net4784));
 sg13g2_nand3_1 _14107_ (.B(_07438_),
    .C(net5288),
    .A(net5800),
    .Y(_08299_));
 sg13g2_xnor2_1 _14108_ (.Y(_08300_),
    .A(_06567_),
    .B(_07438_));
 sg13g2_o21ai_1 _14109_ (.B1(net5099),
    .Y(_08301_),
    .A1(net5800),
    .A2(_07438_));
 sg13g2_nand3_1 _14110_ (.B(_08299_),
    .C(_08301_),
    .A(net5199),
    .Y(_08302_));
 sg13g2_a21oi_1 _14111_ (.A1(net5183),
    .A2(_08300_),
    .Y(_08303_),
    .B1(_08302_));
 sg13g2_nand3_1 _14112_ (.B(_08298_),
    .C(_08303_),
    .A(_08294_),
    .Y(_08304_));
 sg13g2_o21ai_1 _14113_ (.B1(_08304_),
    .Y(_08305_),
    .A1(net5200),
    .A2(_08281_));
 sg13g2_o21ai_1 _14114_ (.B1(net5223),
    .Y(_08306_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[9] ),
    .A2(net5192));
 sg13g2_a21oi_1 _14115_ (.A1(net5192),
    .A2(_08305_),
    .Y(_08307_),
    .B1(_08306_));
 sg13g2_a21oi_1 _14116_ (.A1(_07122_),
    .A2(_07128_),
    .Y(_08308_),
    .B1(_07126_));
 sg13g2_xnor2_1 _14117_ (.Y(_08309_),
    .A(_07065_),
    .B(_08308_));
 sg13g2_o21ai_1 _14118_ (.B1(net5219),
    .Y(_08310_),
    .A1(net5222),
    .A2(_08309_));
 sg13g2_xnor2_1 _14119_ (.Y(_08311_),
    .A(_06592_),
    .B(_07654_));
 sg13g2_a21oi_1 _14120_ (.A1(net5213),
    .A2(_08311_),
    .Y(_08312_),
    .B1(net5179));
 sg13g2_o21ai_1 _14121_ (.B1(_08312_),
    .Y(_08313_),
    .A1(_08307_),
    .A2(_08310_));
 sg13g2_and2_1 _14122_ (.A(\fpga_top.uart_top.uart_rec_char.bpoint[9] ),
    .B(_08313_),
    .X(_08314_));
 sg13g2_nor2_1 _14123_ (.A(\fpga_top.uart_top.uart_rec_char.bpoint[9] ),
    .B(_08313_),
    .Y(_08315_));
 sg13g2_nor2_1 _14124_ (.A(\fpga_top.uart_top.uart_rec_char.bpoint[6] ),
    .B(_08247_),
    .Y(_08316_));
 sg13g2_nor4_1 _14125_ (.A(_08280_),
    .B(_08314_),
    .C(_08315_),
    .D(_08316_),
    .Y(_08317_));
 sg13g2_nand4_1 _14126_ (.B(_08225_),
    .C(_08248_),
    .A(_08103_),
    .Y(_08318_),
    .D(_08317_));
 sg13g2_nor2_1 _14127_ (.A(_06552_),
    .B(net5286),
    .Y(_08319_));
 sg13g2_xnor2_1 _14128_ (.Y(_08320_),
    .A(_07367_),
    .B(_07910_));
 sg13g2_nand2_1 _14129_ (.Y(_08321_),
    .A(net5197),
    .B(_08320_));
 sg13g2_nor2_1 _14130_ (.A(net4974),
    .B(_08199_),
    .Y(_08322_));
 sg13g2_o21ai_1 _14131_ (.B1(net4856),
    .Y(_08323_),
    .A1(net4955),
    .A2(_08197_));
 sg13g2_nor2_1 _14132_ (.A(_08322_),
    .B(_08323_),
    .Y(_08324_));
 sg13g2_a22oi_1 _14133_ (.Y(_08325_),
    .B1(_08196_),
    .B2(net4959),
    .A2(_07805_),
    .A1(net5755));
 sg13g2_nor2_1 _14134_ (.A(net4856),
    .B(_08325_),
    .Y(_08326_));
 sg13g2_o21ai_1 _14135_ (.B1(_07603_),
    .Y(_08327_),
    .A1(_08324_),
    .A2(_08326_));
 sg13g2_mux2_1 _14136_ (.A0(_07880_),
    .A1(_07886_),
    .S(net5020),
    .X(_08328_));
 sg13g2_nor2_1 _14137_ (.A(net4964),
    .B(_08328_),
    .Y(_08329_));
 sg13g2_a21oi_2 _14138_ (.B1(_08329_),
    .Y(_08330_),
    .A2(_08207_),
    .A1(net4964));
 sg13g2_nand2b_1 _14139_ (.Y(_08331_),
    .B(_07363_),
    .A_N(net5794));
 sg13g2_nor2b_1 _14140_ (.A(_07363_),
    .B_N(net5794),
    .Y(_08332_));
 sg13g2_a221oi_1 _14141_ (.B2(net5189),
    .C1(net5197),
    .B1(_08332_),
    .A1(_07613_),
    .Y(_08333_),
    .A2(_08331_));
 sg13g2_xnor2_1 _14142_ (.Y(_08334_),
    .A(net5794),
    .B(_07363_));
 sg13g2_a22oi_1 _14143_ (.Y(_08335_),
    .B1(_08334_),
    .B2(net5184),
    .A2(_08330_),
    .A1(net4855));
 sg13g2_nand3_1 _14144_ (.B(_08333_),
    .C(_08335_),
    .A(_08327_),
    .Y(_08336_));
 sg13g2_o21ai_1 _14145_ (.B1(net5222),
    .Y(_08337_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[12] ),
    .A2(net5192));
 sg13g2_a21oi_1 _14146_ (.A1(_08321_),
    .A2(_08336_),
    .Y(_08338_),
    .B1(net5293));
 sg13g2_xnor2_1 _14147_ (.Y(_08339_),
    .A(_07149_),
    .B(_07178_));
 sg13g2_nor2_1 _14148_ (.A(net5222),
    .B(_08339_),
    .Y(_08340_));
 sg13g2_nor2_1 _14149_ (.A(net5213),
    .B(_08340_),
    .Y(_08341_));
 sg13g2_o21ai_1 _14150_ (.B1(_08341_),
    .Y(_08342_),
    .A1(_08337_),
    .A2(_08338_));
 sg13g2_xnor2_1 _14151_ (.Y(_08343_),
    .A(_06599_),
    .B(_07656_));
 sg13g2_a21oi_1 _14152_ (.A1(net5213),
    .A2(_08343_),
    .Y(_08344_),
    .B1(net5179));
 sg13g2_a21o_2 _14153_ (.A2(_08344_),
    .A1(_08342_),
    .B1(_08319_),
    .X(_08345_));
 sg13g2_xor2_1 _14154_ (.B(_08345_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[12] ),
    .X(_08346_));
 sg13g2_nand2_1 _14155_ (.Y(_08347_),
    .A(\fpga_top.cpu_top.csr_uimm[2] ),
    .B(net5180));
 sg13g2_o21ai_1 _14156_ (.B1(_07507_),
    .Y(_08348_),
    .A1(_07492_),
    .A2(_07513_));
 sg13g2_nor2_1 _14157_ (.A(_07497_),
    .B(_08348_),
    .Y(_08349_));
 sg13g2_xor2_1 _14158_ (.B(_08348_),
    .A(_07497_),
    .X(_08350_));
 sg13g2_nand2b_1 _14159_ (.Y(_08351_),
    .B(_07805_),
    .A_N(_08288_));
 sg13g2_o21ai_1 _14160_ (.B1(_08351_),
    .Y(_08352_),
    .A1(net4971),
    .A2(_08282_));
 sg13g2_a21oi_2 _14161_ (.B1(_08352_),
    .Y(_08353_),
    .A2(_08291_),
    .A1(net4971));
 sg13g2_o21ai_1 _14162_ (.B1(net4756),
    .Y(_08354_),
    .A1(net4953),
    .A2(_08353_));
 sg13g2_nor2_1 _14163_ (.A(net4955),
    .B(_08295_),
    .Y(_08355_));
 sg13g2_mux2_1 _14164_ (.A0(_07766_),
    .A1(_07779_),
    .S(net5006),
    .X(_08356_));
 sg13g2_nor2_1 _14165_ (.A(net4784),
    .B(_08355_),
    .Y(_08357_));
 sg13g2_o21ai_1 _14166_ (.B1(_08357_),
    .Y(_08358_),
    .A1(net4967),
    .A2(_08356_));
 sg13g2_xnor2_1 _14167_ (.Y(_08359_),
    .A(net5783),
    .B(_07493_));
 sg13g2_or2_1 _14168_ (.X(_08360_),
    .B(_08359_),
    .A(_07616_));
 sg13g2_o21ai_1 _14169_ (.B1(net5100),
    .Y(_08361_),
    .A1(net5783),
    .A2(_07493_));
 sg13g2_nand3_1 _14170_ (.B(_07493_),
    .C(net5288),
    .A(net5783),
    .Y(_08362_));
 sg13g2_nand4_1 _14171_ (.B(_08360_),
    .C(_08361_),
    .A(net5204),
    .Y(_08363_),
    .D(_08362_));
 sg13g2_nor3_1 _14172_ (.A(net5012),
    .B(net4964),
    .C(_07769_),
    .Y(_08364_));
 sg13g2_a21oi_1 _14173_ (.A1(net4786),
    .A2(_08364_),
    .Y(_08365_),
    .B1(_08363_));
 sg13g2_nand3_1 _14174_ (.B(_08358_),
    .C(_08365_),
    .A(_08354_),
    .Y(_08366_));
 sg13g2_o21ai_1 _14175_ (.B1(_08366_),
    .Y(_08367_),
    .A1(net5204),
    .A2(_08350_));
 sg13g2_o21ai_1 _14176_ (.B1(net5226),
    .Y(_08368_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[17] ),
    .A2(net5195));
 sg13g2_a21oi_1 _14177_ (.A1(net5194),
    .A2(_08367_),
    .Y(_08369_),
    .B1(_08368_));
 sg13g2_a21oi_1 _14178_ (.A1(_07183_),
    .A2(_07229_),
    .Y(_08370_),
    .B1(_07228_));
 sg13g2_xor2_1 _14179_ (.B(_08370_),
    .A(_07235_),
    .X(_08371_));
 sg13g2_o21ai_1 _14180_ (.B1(net5218),
    .Y(_08372_),
    .A1(net5225),
    .A2(_08371_));
 sg13g2_nor2_1 _14181_ (.A(_08369_),
    .B(_08372_),
    .Y(_08373_));
 sg13g2_a21o_1 _14182_ (.A2(_07660_),
    .A1(net5594),
    .B1(\fpga_top.bus_gather.i_read_adr[17] ),
    .X(_08374_));
 sg13g2_and2_1 _14183_ (.A(_07661_),
    .B(_08374_),
    .X(_08375_));
 sg13g2_o21ai_1 _14184_ (.B1(net5286),
    .Y(_08376_),
    .A1(net5218),
    .A2(_08375_));
 sg13g2_o21ai_1 _14185_ (.B1(_08347_),
    .Y(_08377_),
    .A1(_08373_),
    .A2(_08376_));
 sg13g2_xnor2_1 _14186_ (.Y(_08378_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[17] ),
    .B(_08377_));
 sg13g2_a21oi_1 _14187_ (.A1(_07183_),
    .A2(_07236_),
    .Y(_08379_),
    .B1(_07241_));
 sg13g2_o21ai_1 _14188_ (.B1(_07220_),
    .Y(_08380_),
    .A1(_07222_),
    .A2(_08379_));
 sg13g2_xor2_1 _14189_ (.B(_08380_),
    .A(_07215_),
    .X(_08381_));
 sg13g2_nand3_1 _14190_ (.B(_07511_),
    .C(_07516_),
    .A(_07334_),
    .Y(_08382_));
 sg13g2_a21oi_1 _14191_ (.A1(_07801_),
    .A2(_08382_),
    .Y(_08383_),
    .B1(net5202));
 sg13g2_nor2_1 _14192_ (.A(net5208),
    .B(_08170_),
    .Y(_08384_));
 sg13g2_nor3_1 _14193_ (.A(_07292_),
    .B(net4951),
    .C(_08163_),
    .Y(_08385_));
 sg13g2_nor3_1 _14194_ (.A(_07688_),
    .B(_08384_),
    .C(_08385_),
    .Y(_08386_));
 sg13g2_nor2_1 _14195_ (.A(net4956),
    .B(_08261_),
    .Y(_08387_));
 sg13g2_mux2_1 _14196_ (.A0(_07588_),
    .A1(_07633_),
    .S(net5006),
    .X(_08388_));
 sg13g2_o21ai_1 _14197_ (.B1(net4854),
    .Y(_08389_),
    .A1(net4969),
    .A2(_08388_));
 sg13g2_nor3_1 _14198_ (.A(net4966),
    .B(_07581_),
    .C(_08173_),
    .Y(_08390_));
 sg13g2_xor2_1 _14199_ (.B(_07330_),
    .A(net5778),
    .X(_08391_));
 sg13g2_nand2_1 _14200_ (.Y(_08392_),
    .A(net5185),
    .B(_08391_));
 sg13g2_nand3_1 _14201_ (.B(_07330_),
    .C(_07608_),
    .A(net5778),
    .Y(_08393_));
 sg13g2_o21ai_1 _14202_ (.B1(net5101),
    .Y(_08394_),
    .A1(net5778),
    .A2(_07330_));
 sg13g2_o21ai_1 _14203_ (.B1(net5204),
    .Y(_08395_),
    .A1(_08387_),
    .A2(_08389_));
 sg13g2_nand3_1 _14204_ (.B(_08393_),
    .C(_08394_),
    .A(_08392_),
    .Y(_08396_));
 sg13g2_nor4_1 _14205_ (.A(_08386_),
    .B(_08390_),
    .C(_08395_),
    .D(_08396_),
    .Y(_08397_));
 sg13g2_or3_1 _14206_ (.A(net5290),
    .B(_08383_),
    .C(_08397_),
    .X(_08398_));
 sg13g2_a21oi_1 _14207_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[19] ),
    .A2(net5289),
    .Y(_08399_),
    .B1(net5311));
 sg13g2_a21oi_1 _14208_ (.A1(_08398_),
    .A2(_08399_),
    .Y(_08400_),
    .B1(net5216));
 sg13g2_o21ai_1 _14209_ (.B1(_08400_),
    .Y(_08401_),
    .A1(net5226),
    .A2(_08381_));
 sg13g2_xnor2_1 _14210_ (.Y(_08402_),
    .A(\fpga_top.bus_gather.i_read_adr[19] ),
    .B(_07662_));
 sg13g2_nor2_1 _14211_ (.A(net5218),
    .B(_08402_),
    .Y(_08403_));
 sg13g2_nor2_1 _14212_ (.A(net5182),
    .B(_08403_),
    .Y(_08404_));
 sg13g2_a22oi_1 _14213_ (.Y(_08405_),
    .B1(_08401_),
    .B2(_08404_),
    .A2(net5182),
    .A1(_06618_));
 sg13g2_nor2b_1 _14214_ (.A(_07333_),
    .B_N(_07801_),
    .Y(_08406_));
 sg13g2_xnor2_1 _14215_ (.Y(_08407_),
    .A(_07338_),
    .B(_08406_));
 sg13g2_nand2_1 _14216_ (.Y(_08408_),
    .A(net5013),
    .B(_07881_));
 sg13g2_o21ai_1 _14217_ (.B1(_08408_),
    .Y(_08409_),
    .A1(net5014),
    .A2(_07876_));
 sg13g2_mux2_1 _14218_ (.A0(_08328_),
    .A1(_08409_),
    .S(net4956),
    .X(_08410_));
 sg13g2_xnor2_1 _14219_ (.Y(_08411_),
    .A(_06578_),
    .B(_07335_));
 sg13g2_nand3_1 _14220_ (.B(_07335_),
    .C(net5188),
    .A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[20] ),
    .Y(_08412_));
 sg13g2_o21ai_1 _14221_ (.B1(net5101),
    .Y(_08413_),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[20] ),
    .A2(_07335_));
 sg13g2_nand2_1 _14222_ (.Y(_08414_),
    .A(_08412_),
    .B(_08413_));
 sg13g2_o21ai_1 _14223_ (.B1(net4756),
    .Y(_08415_),
    .A1(net4953),
    .A2(_08198_));
 sg13g2_a221oi_1 _14224_ (.B2(net4853),
    .C1(_08414_),
    .B1(_08410_),
    .A1(net4786),
    .Y(_08416_),
    .A2(_08208_));
 sg13g2_nand2_1 _14225_ (.Y(_08417_),
    .A(_08415_),
    .B(_08416_));
 sg13g2_a221oi_1 _14226_ (.B2(net5185),
    .C1(_08417_),
    .B1(_08411_),
    .A1(net5196),
    .Y(_08418_),
    .A2(_08407_));
 sg13g2_a21oi_1 _14227_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[20] ),
    .A2(net5289),
    .Y(_08419_),
    .B1(net5311));
 sg13g2_o21ai_1 _14228_ (.B1(_08419_),
    .Y(_08420_),
    .A1(net5290),
    .A2(_08418_));
 sg13g2_xnor2_1 _14229_ (.Y(_08421_),
    .A(_07207_),
    .B(_07829_));
 sg13g2_a21oi_1 _14230_ (.A1(net5310),
    .A2(_08421_),
    .Y(_08422_),
    .B1(net5215));
 sg13g2_a21o_1 _14231_ (.A2(_07662_),
    .A1(\fpga_top.bus_gather.i_read_adr[19] ),
    .B1(\fpga_top.bus_gather.i_read_adr[20] ),
    .X(_08423_));
 sg13g2_nand2_1 _14232_ (.Y(_08424_),
    .A(_07663_),
    .B(_08423_));
 sg13g2_o21ai_1 _14233_ (.B1(net5287),
    .Y(_08425_),
    .A1(net5217),
    .A2(_08424_));
 sg13g2_a21o_2 _14234_ (.A2(_08422_),
    .A1(_08420_),
    .B1(_08425_),
    .X(_08426_));
 sg13g2_o21ai_1 _14235_ (.B1(_08426_),
    .Y(_08427_),
    .A1(net5572),
    .A2(net5286));
 sg13g2_inv_2 _14236_ (.Y(_08428_),
    .A(_08427_));
 sg13g2_xnor2_1 _14237_ (.Y(_08429_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[20] ),
    .B(_08427_));
 sg13g2_nand2_1 _14238_ (.Y(_08430_),
    .A(\fpga_top.cpu_top.br_ofs[7] ),
    .B(net5179));
 sg13g2_nand2_1 _14239_ (.Y(_08431_),
    .A(_07269_),
    .B(_07271_));
 sg13g2_xor2_1 _14240_ (.B(_08431_),
    .A(_07272_),
    .X(_08432_));
 sg13g2_or2_1 _14241_ (.X(_08433_),
    .B(_07558_),
    .A(_07548_));
 sg13g2_xnor2_1 _14242_ (.Y(_08434_),
    .A(_07548_),
    .B(_07558_));
 sg13g2_o21ai_1 _14243_ (.B1(net4756),
    .Y(_08435_),
    .A1(net4952),
    .A2(_08259_));
 sg13g2_nor2_1 _14244_ (.A(net5007),
    .B(_07639_),
    .Y(_08436_));
 sg13g2_o21ai_1 _14245_ (.B1(net4958),
    .Y(_08437_),
    .A1(net5015),
    .A2(_07620_));
 sg13g2_nand2_1 _14246_ (.Y(_08438_),
    .A(net4969),
    .B(_08388_));
 sg13g2_o21ai_1 _14247_ (.B1(_08438_),
    .Y(_08439_),
    .A1(_08436_),
    .A2(_08437_));
 sg13g2_xor2_1 _14248_ (.B(_07554_),
    .A(net5761),
    .X(_08440_));
 sg13g2_nand2_1 _14249_ (.Y(_08441_),
    .A(net5185),
    .B(_08440_));
 sg13g2_nand3_1 _14250_ (.B(_07554_),
    .C(net5288),
    .A(net5761),
    .Y(_08442_));
 sg13g2_o21ai_1 _14251_ (.B1(net5101),
    .Y(_08443_),
    .A1(net5761),
    .A2(_07554_));
 sg13g2_nand4_1 _14252_ (.B(_08441_),
    .C(_08442_),
    .A(net5203),
    .Y(_08444_),
    .D(_08443_));
 sg13g2_a221oi_1 _14253_ (.B2(net4854),
    .C1(_08444_),
    .B1(_08439_),
    .A1(net4786),
    .Y(_08445_),
    .A2(_08263_));
 sg13g2_a221oi_1 _14254_ (.B2(_08445_),
    .C1(net5291),
    .B1(_08435_),
    .A1(net5196),
    .Y(_08446_),
    .A2(_08434_));
 sg13g2_a21oi_1 _14255_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[27] ),
    .A2(net5289),
    .Y(_08447_),
    .B1(_08446_));
 sg13g2_o21ai_1 _14256_ (.B1(net5217),
    .Y(_08448_),
    .A1(net5311),
    .A2(_08447_));
 sg13g2_a21oi_1 _14257_ (.A1(net5311),
    .A2(_08432_),
    .Y(_08449_),
    .B1(_08448_));
 sg13g2_xnor2_1 _14258_ (.Y(_08450_),
    .A(_06636_),
    .B(_07667_));
 sg13g2_a21o_1 _14259_ (.A2(_08450_),
    .A1(net5214),
    .B1(net5181),
    .X(_08451_));
 sg13g2_o21ai_1 _14260_ (.B1(_08430_),
    .Y(_08452_),
    .A1(_08449_),
    .A2(_08451_));
 sg13g2_xnor2_1 _14261_ (.Y(_08453_),
    .A(_06637_),
    .B(_08452_));
 sg13g2_o21ai_1 _14262_ (.B1(_07187_),
    .Y(_08454_),
    .A1(_07189_),
    .A2(_07831_));
 sg13g2_xor2_1 _14263_ (.B(_08454_),
    .A(_07194_),
    .X(_08455_));
 sg13g2_xnor2_1 _14264_ (.Y(_08456_),
    .A(_07518_),
    .B(_07523_));
 sg13g2_o21ai_1 _14265_ (.B1(_07687_),
    .Y(_08457_),
    .A1(net4952),
    .A2(_08046_));
 sg13g2_nor2_1 _14266_ (.A(net4956),
    .B(_07589_),
    .Y(_08458_));
 sg13g2_nor2_1 _14267_ (.A(net4785),
    .B(_08458_),
    .Y(_08459_));
 sg13g2_o21ai_1 _14268_ (.B1(_08459_),
    .Y(_08460_),
    .A1(net4969),
    .A2(_07640_));
 sg13g2_xor2_1 _14269_ (.B(_07519_),
    .A(net5771),
    .X(_08461_));
 sg13g2_nand3_1 _14270_ (.B(_07519_),
    .C(_07608_),
    .A(net5771),
    .Y(_08462_));
 sg13g2_o21ai_1 _14271_ (.B1(net5102),
    .Y(_08463_),
    .A1(net5771),
    .A2(_07519_));
 sg13g2_nand3_1 _14272_ (.B(_08462_),
    .C(_08463_),
    .A(net5203),
    .Y(_08464_));
 sg13g2_a221oi_1 _14273_ (.B2(net5185),
    .C1(_08464_),
    .B1(_08461_),
    .A1(_07580_),
    .Y(_08465_),
    .A2(_08058_));
 sg13g2_and2_1 _14274_ (.A(_08460_),
    .B(_08465_),
    .X(_08466_));
 sg13g2_a221oi_1 _14275_ (.B2(_08466_),
    .C1(net5291),
    .B1(_08457_),
    .A1(net5196),
    .Y(_08467_),
    .A2(_08456_));
 sg13g2_a21oi_1 _14276_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[23] ),
    .A2(net5289),
    .Y(_08468_),
    .B1(_08467_));
 sg13g2_a21oi_1 _14277_ (.A1(net5226),
    .A2(_08468_),
    .Y(_08469_),
    .B1(net5216));
 sg13g2_o21ai_1 _14278_ (.B1(_08469_),
    .Y(_08470_),
    .A1(net5226),
    .A2(_08455_));
 sg13g2_a21o_1 _14279_ (.A2(_07664_),
    .A1(net5591),
    .B1(\fpga_top.bus_gather.i_read_adr[23] ),
    .X(_08471_));
 sg13g2_nand2_1 _14280_ (.Y(_08472_),
    .A(_07665_),
    .B(_08471_));
 sg13g2_inv_1 _14281_ (.Y(_08473_),
    .A(_08472_));
 sg13g2_a21oi_1 _14282_ (.A1(net5215),
    .A2(_08473_),
    .Y(_08474_),
    .B1(net5181));
 sg13g2_a22oi_1 _14283_ (.Y(_08475_),
    .B1(_08470_),
    .B2(_08474_),
    .A2(net5181),
    .A1(_06568_));
 sg13g2_xnor2_1 _14284_ (.Y(_08476_),
    .A(_06627_),
    .B(_08475_));
 sg13g2_o21ai_1 _14285_ (.B1(_07540_),
    .Y(_08477_),
    .A1(_07525_),
    .A2(_07544_));
 sg13g2_xnor2_1 _14286_ (.Y(_08478_),
    .A(_07530_),
    .B(_08477_));
 sg13g2_o21ai_1 _14287_ (.B1(net4756),
    .Y(_08479_),
    .A1(net4952),
    .A2(_08292_));
 sg13g2_nor2_1 _14288_ (.A(net5016),
    .B(_07784_),
    .Y(_08480_));
 sg13g2_o21ai_1 _14289_ (.B1(net4956),
    .Y(_08481_),
    .A1(net5006),
    .A2(_07781_));
 sg13g2_nand2_1 _14290_ (.Y(_08482_),
    .A(net4966),
    .B(_08356_));
 sg13g2_o21ai_1 _14291_ (.B1(_08482_),
    .Y(_08483_),
    .A1(_08480_),
    .A2(_08481_));
 sg13g2_xor2_1 _14292_ (.B(_07526_),
    .A(net5766),
    .X(_08484_));
 sg13g2_nand3_1 _14293_ (.B(_07526_),
    .C(net5188),
    .A(net5766),
    .Y(_08485_));
 sg13g2_o21ai_1 _14294_ (.B1(net5102),
    .Y(_08486_),
    .A1(net5766),
    .A2(_07526_));
 sg13g2_nand3_1 _14295_ (.B(_08485_),
    .C(_08486_),
    .A(net5203),
    .Y(_08487_));
 sg13g2_a21oi_1 _14296_ (.A1(net5186),
    .A2(_08484_),
    .Y(_08488_),
    .B1(_08487_));
 sg13g2_o21ai_1 _14297_ (.B1(_08488_),
    .Y(_08489_),
    .A1(_07581_),
    .A2(_08297_));
 sg13g2_a21oi_1 _14298_ (.A1(net4854),
    .A2(_08483_),
    .Y(_08490_),
    .B1(_08489_));
 sg13g2_a21oi_1 _14299_ (.A1(_08479_),
    .A2(_08490_),
    .Y(_08491_),
    .B1(net5291));
 sg13g2_o21ai_1 _14300_ (.B1(_08491_),
    .Y(_08492_),
    .A1(net5202),
    .A2(_08478_));
 sg13g2_a21oi_1 _14301_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[25] ),
    .A2(net5290),
    .Y(_08493_),
    .B1(net5313));
 sg13g2_o21ai_1 _14302_ (.B1(_07259_),
    .Y(_08494_),
    .A1(_07249_),
    .A2(_07261_));
 sg13g2_xnor2_1 _14303_ (.Y(_08495_),
    .A(_07255_),
    .B(_08494_));
 sg13g2_a22oi_1 _14304_ (.Y(_08496_),
    .B1(_08495_),
    .B2(net5313),
    .A2(_08493_),
    .A1(_08492_));
 sg13g2_xnor2_1 _14305_ (.Y(_08497_),
    .A(\fpga_top.bus_gather.i_read_adr[25] ),
    .B(_07666_));
 sg13g2_o21ai_1 _14306_ (.B1(net5287),
    .Y(_08498_),
    .A1(net5217),
    .A2(_08497_));
 sg13g2_a21oi_1 _14307_ (.A1(net5217),
    .A2(_08496_),
    .Y(_08499_),
    .B1(_08498_));
 sg13g2_a21oi_2 _14308_ (.B1(_08499_),
    .Y(_08500_),
    .A2(net5181),
    .A1(_06558_));
 sg13g2_xnor2_1 _14309_ (.Y(_08501_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[25] ),
    .B(_08500_));
 sg13g2_nor2_1 _14310_ (.A(\fpga_top.cpu_top.csr_uimm[3] ),
    .B(net5287),
    .Y(_08502_));
 sg13g2_o21ai_1 _14311_ (.B1(_07502_),
    .Y(_08503_),
    .A1(_07496_),
    .A2(_08349_));
 sg13g2_or3_1 _14312_ (.A(_07496_),
    .B(_07502_),
    .C(_08349_),
    .X(_08504_));
 sg13g2_nand3_1 _14313_ (.B(_08503_),
    .C(_08504_),
    .A(net5196),
    .Y(_08505_));
 sg13g2_nor3_1 _14314_ (.A(_07292_),
    .B(net4950),
    .C(_08140_),
    .Y(_08506_));
 sg13g2_nor4_2 _14315_ (.A(_07688_),
    .B(_08138_),
    .C(_08139_),
    .Y(_08507_),
    .D(_08506_));
 sg13g2_mux2_1 _14316_ (.A0(_07703_),
    .A1(_07728_),
    .S(net5005),
    .X(_08508_));
 sg13g2_nor2_1 _14317_ (.A(net4955),
    .B(_07993_),
    .Y(_08509_));
 sg13g2_o21ai_1 _14318_ (.B1(net4853),
    .Y(_08510_),
    .A1(net4966),
    .A2(_08508_));
 sg13g2_nor2_1 _14319_ (.A(_08509_),
    .B(_08510_),
    .Y(_08511_));
 sg13g2_nor3_1 _14320_ (.A(net4967),
    .B(_07581_),
    .C(_07994_),
    .Y(_08512_));
 sg13g2_xor2_1 _14321_ (.B(_07498_),
    .A(net5781),
    .X(_08513_));
 sg13g2_nand2_1 _14322_ (.Y(_08514_),
    .A(net5186),
    .B(_08513_));
 sg13g2_o21ai_1 _14323_ (.B1(net5103),
    .Y(_08515_),
    .A1(net5781),
    .A2(_07498_));
 sg13g2_nand3_1 _14324_ (.B(_07498_),
    .C(net5188),
    .A(net5781),
    .Y(_08516_));
 sg13g2_nand4_1 _14325_ (.B(_08514_),
    .C(_08515_),
    .A(net5195),
    .Y(_08517_),
    .D(_08516_));
 sg13g2_nor4_1 _14326_ (.A(_08507_),
    .B(_08511_),
    .C(_08512_),
    .D(_08517_),
    .Y(_08518_));
 sg13g2_a22oi_1 _14327_ (.Y(_08519_),
    .B1(_08505_),
    .B2(_08518_),
    .A2(net5292),
    .A1(_06613_));
 sg13g2_xnor2_1 _14328_ (.Y(_08520_),
    .A(_07222_),
    .B(_08379_));
 sg13g2_a21oi_1 _14329_ (.A1(net5314),
    .A2(_08520_),
    .Y(_08521_),
    .B1(net5215));
 sg13g2_o21ai_1 _14330_ (.B1(_08521_),
    .Y(_08522_),
    .A1(net5314),
    .A2(_08519_));
 sg13g2_xnor2_1 _14331_ (.Y(_08523_),
    .A(_06614_),
    .B(_07661_));
 sg13g2_inv_1 _14332_ (.Y(_08524_),
    .A(_08523_));
 sg13g2_a21oi_1 _14333_ (.A1(net5216),
    .A2(_08524_),
    .Y(_08525_),
    .B1(net5181));
 sg13g2_a21o_2 _14334_ (.A2(_08525_),
    .A1(_08522_),
    .B1(_08502_),
    .X(_08526_));
 sg13g2_xnor2_1 _14335_ (.Y(_08527_),
    .A(_06615_),
    .B(_08526_));
 sg13g2_nand2_1 _14336_ (.Y(_08528_),
    .A(\fpga_top.cpu_top.csr_uimm[0] ),
    .B(net5180));
 sg13g2_o21ai_1 _14337_ (.B1(_07155_),
    .Y(_08529_),
    .A1(_07157_),
    .A2(_07938_));
 sg13g2_xor2_1 _14338_ (.B(_08529_),
    .A(_07163_),
    .X(_08530_));
 sg13g2_and3_1 _14339_ (.X(_08531_),
    .A(_07484_),
    .B(_07486_),
    .C(_07491_));
 sg13g2_o21ai_1 _14340_ (.B1(net5196),
    .Y(_08532_),
    .A1(_07492_),
    .A2(_08531_));
 sg13g2_mux2_1 _14341_ (.A0(_08044_),
    .A1(_08049_),
    .S(net4962),
    .X(_08533_));
 sg13g2_o21ai_1 _14342_ (.B1(_07686_),
    .Y(_08534_),
    .A1(net4952),
    .A2(_08533_));
 sg13g2_a21oi_2 _14343_ (.B1(_08534_),
    .Y(_08535_),
    .A2(_07601_),
    .A1(_07598_));
 sg13g2_nand3_1 _14344_ (.B(_07487_),
    .C(net5187),
    .A(net5787),
    .Y(_08536_));
 sg13g2_o21ai_1 _14345_ (.B1(net5100),
    .Y(_08537_),
    .A1(net5787),
    .A2(_07487_));
 sg13g2_xor2_1 _14346_ (.B(_07487_),
    .A(net5787),
    .X(_08538_));
 sg13g2_a22oi_1 _14347_ (.Y(_08539_),
    .B1(_08538_),
    .B2(net5184),
    .A2(net4853),
    .A1(_07595_));
 sg13g2_nand4_1 _14348_ (.B(_08536_),
    .C(_08537_),
    .A(net5201),
    .Y(_08540_),
    .D(_08539_));
 sg13g2_or2_1 _14349_ (.X(_08541_),
    .B(_08540_),
    .A(_08535_));
 sg13g2_a21oi_1 _14350_ (.A1(_08532_),
    .A2(_08541_),
    .Y(_08542_),
    .B1(net5292));
 sg13g2_o21ai_1 _14351_ (.B1(net5225),
    .Y(_08543_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[15] ),
    .A2(net5194));
 sg13g2_o21ai_1 _14352_ (.B1(net5218),
    .Y(_08544_),
    .A1(_08542_),
    .A2(_08543_));
 sg13g2_a21oi_1 _14353_ (.A1(net5309),
    .A2(_08530_),
    .Y(_08545_),
    .B1(_08544_));
 sg13g2_xnor2_1 _14354_ (.Y(_08546_),
    .A(_06605_),
    .B(_07659_));
 sg13g2_a21o_1 _14355_ (.A2(_08546_),
    .A1(net5213),
    .B1(net5180),
    .X(_08547_));
 sg13g2_o21ai_1 _14356_ (.B1(_08528_),
    .Y(_08548_),
    .A1(_08545_),
    .A2(_08547_));
 sg13g2_xor2_1 _14357_ (.B(_08548_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[15] ),
    .X(_08549_));
 sg13g2_nand2_1 _14358_ (.Y(_08550_),
    .A(\fpga_top.cpu_top.br_ofs[8] ),
    .B(net5179));
 sg13g2_and3_1 _14359_ (.X(_08551_),
    .A(_07552_),
    .B(_07557_),
    .C(_08433_));
 sg13g2_a21oi_1 _14360_ (.A1(_07557_),
    .A2(_08433_),
    .Y(_08552_),
    .B1(_07552_));
 sg13g2_nor3_1 _14361_ (.A(net5203),
    .B(_08551_),
    .C(_08552_),
    .Y(_08553_));
 sg13g2_a21oi_1 _14362_ (.A1(net4858),
    .A2(_08325_),
    .Y(_08554_),
    .B1(_07688_));
 sg13g2_o21ai_1 _14363_ (.B1(net5001),
    .Y(_08555_),
    .A1(_07724_),
    .A2(_07725_));
 sg13g2_o21ai_1 _14364_ (.B1(_08555_),
    .Y(_08556_),
    .A1(net4998),
    .A2(_07722_));
 sg13g2_a21oi_1 _14365_ (.A1(net5015),
    .A2(_07877_),
    .Y(_08557_),
    .B1(net4969));
 sg13g2_o21ai_1 _14366_ (.B1(_08557_),
    .Y(_08558_),
    .A1(net5015),
    .A2(_08556_));
 sg13g2_o21ai_1 _14367_ (.B1(_08558_),
    .Y(_08559_),
    .A1(net4958),
    .A2(_08409_));
 sg13g2_nor2_1 _14368_ (.A(net4785),
    .B(_08559_),
    .Y(_08560_));
 sg13g2_nand3_1 _14369_ (.B(_07549_),
    .C(net5188),
    .A(net5760),
    .Y(_08561_));
 sg13g2_o21ai_1 _14370_ (.B1(net5101),
    .Y(_08562_),
    .A1(net5760),
    .A2(_07549_));
 sg13g2_xnor2_1 _14371_ (.Y(_08563_),
    .A(_06580_),
    .B(_07549_));
 sg13g2_a22oi_1 _14372_ (.Y(_08564_),
    .B1(_08563_),
    .B2(net5185),
    .A2(_08330_),
    .A1(net4786));
 sg13g2_nand4_1 _14373_ (.B(_08561_),
    .C(_08562_),
    .A(net5202),
    .Y(_08565_),
    .D(_08564_));
 sg13g2_nor3_1 _14374_ (.A(_08554_),
    .B(_08560_),
    .C(_08565_),
    .Y(_08566_));
 sg13g2_o21ai_1 _14375_ (.B1(net5194),
    .Y(_08567_),
    .A1(_08553_),
    .A2(_08566_));
 sg13g2_a21oi_1 _14376_ (.A1(_06638_),
    .A2(net5289),
    .Y(_08568_),
    .B1(net5312));
 sg13g2_xnor2_1 _14377_ (.Y(_08569_),
    .A(_07055_),
    .B(_07275_));
 sg13g2_a221oi_1 _14378_ (.B2(net5311),
    .C1(net5216),
    .B1(_08569_),
    .A1(_08567_),
    .Y(_08570_),
    .A2(_08568_));
 sg13g2_xor2_1 _14379_ (.B(_07668_),
    .A(net5590),
    .X(_08571_));
 sg13g2_inv_1 _14380_ (.Y(_08572_),
    .A(_08571_));
 sg13g2_o21ai_1 _14381_ (.B1(net5286),
    .Y(_08573_),
    .A1(net5218),
    .A2(_08571_));
 sg13g2_o21ai_1 _14382_ (.B1(_08550_),
    .Y(_08574_),
    .A1(_08570_),
    .A2(_08573_));
 sg13g2_xor2_1 _14383_ (.B(_08574_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[28] ),
    .X(_08575_));
 sg13g2_o21ai_1 _14384_ (.B1(_07529_),
    .Y(_08576_),
    .A1(_07531_),
    .A2(_08477_));
 sg13g2_xnor2_1 _14385_ (.Y(_08577_),
    .A(_07536_),
    .B(_08576_));
 sg13g2_o21ai_1 _14386_ (.B1(net4756),
    .Y(_08578_),
    .A1(net4952),
    .A2(_07985_));
 sg13g2_nor2_1 _14387_ (.A(net5015),
    .B(_07723_),
    .Y(_08579_));
 sg13g2_o21ai_1 _14388_ (.B1(net4958),
    .Y(_08580_),
    .A1(net5007),
    .A2(_07731_));
 sg13g2_nand2_1 _14389_ (.Y(_08581_),
    .A(net4969),
    .B(_08508_));
 sg13g2_o21ai_1 _14390_ (.B1(_08581_),
    .Y(_08582_),
    .A1(_08579_),
    .A2(_08580_));
 sg13g2_xor2_1 _14391_ (.B(_07532_),
    .A(net5764),
    .X(_08583_));
 sg13g2_nand3_1 _14392_ (.B(_07532_),
    .C(net5189),
    .A(net5764),
    .Y(_08584_));
 sg13g2_o21ai_1 _14393_ (.B1(net5102),
    .Y(_08585_),
    .A1(net5764),
    .A2(_07532_));
 sg13g2_nand3_1 _14394_ (.B(_08584_),
    .C(_08585_),
    .A(net5203),
    .Y(_08586_));
 sg13g2_a21oi_1 _14395_ (.A1(net5185),
    .A2(_08583_),
    .Y(_08587_),
    .B1(_08586_));
 sg13g2_o21ai_1 _14396_ (.B1(_08587_),
    .Y(_08588_),
    .A1(_07581_),
    .A2(_07996_));
 sg13g2_a21oi_1 _14397_ (.A1(net4854),
    .A2(_08582_),
    .Y(_08589_),
    .B1(_08588_));
 sg13g2_a22oi_1 _14398_ (.Y(_08590_),
    .B1(_08578_),
    .B2(_08589_),
    .A2(_08577_),
    .A1(net5196));
 sg13g2_a21oi_1 _14399_ (.A1(_06632_),
    .A2(net5289),
    .Y(_08591_),
    .B1(net5314));
 sg13g2_o21ai_1 _14400_ (.B1(_08591_),
    .Y(_08592_),
    .A1(net5289),
    .A2(_08590_));
 sg13g2_xor2_1 _14401_ (.B(_07270_),
    .A(_07265_),
    .X(_08593_));
 sg13g2_a21oi_1 _14402_ (.A1(net5312),
    .A2(_08593_),
    .Y(_08594_),
    .B1(net5215));
 sg13g2_a21o_1 _14403_ (.A2(_07666_),
    .A1(\fpga_top.bus_gather.i_read_adr[25] ),
    .B1(\fpga_top.bus_gather.i_read_adr[26] ),
    .X(_08595_));
 sg13g2_nand2_2 _14404_ (.Y(_08596_),
    .A(_07667_),
    .B(_08595_));
 sg13g2_a221oi_1 _14405_ (.B2(net5215),
    .C1(net5181),
    .B1(_08596_),
    .A1(_08592_),
    .Y(_08597_),
    .A2(_08594_));
 sg13g2_a21o_1 _14406_ (.A2(net5177),
    .A1(\fpga_top.cpu_top.br_ofs[6] ),
    .B1(_08597_),
    .X(_08598_));
 sg13g2_xnor2_1 _14407_ (.Y(_08599_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[26] ),
    .B(_08598_));
 sg13g2_xnor2_1 _14408_ (.Y(_08600_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[21] ),
    .B(_07867_));
 sg13g2_xor2_1 _14409_ (.B(_07970_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[13] ),
    .X(_08601_));
 sg13g2_xnor2_1 _14410_ (.Y(_08602_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[19] ),
    .B(_08405_));
 sg13g2_xor2_1 _14411_ (.B(_07908_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[24] ),
    .X(_08603_));
 sg13g2_nor2_1 _14412_ (.A(\fpga_top.uart_top.uart_rec_char.bpoint[29] ),
    .B(_07798_),
    .Y(_08604_));
 sg13g2_nor4_1 _14413_ (.A(_08039_),
    .B(_08318_),
    .C(_08346_),
    .D(_08601_),
    .Y(_08605_));
 sg13g2_nand4_1 _14414_ (.B(_08378_),
    .C(_08527_),
    .A(_08013_),
    .Y(_08606_),
    .D(_08605_));
 sg13g2_nor4_1 _14415_ (.A(_08429_),
    .B(_08549_),
    .C(_08604_),
    .D(_08606_),
    .Y(_08607_));
 sg13g2_nand3_1 _14416_ (.B(_08602_),
    .C(_08603_),
    .A(_07945_),
    .Y(_08608_));
 sg13g2_nand2_1 _14417_ (.Y(_08609_),
    .A(_08501_),
    .B(_08600_));
 sg13g2_nor4_1 _14418_ (.A(_08453_),
    .B(_08476_),
    .C(_08608_),
    .D(_08609_),
    .Y(_08610_));
 sg13g2_a21oi_1 _14419_ (.A1(\fpga_top.uart_top.uart_rec_char.bpoint[29] ),
    .A2(_07798_),
    .Y(_08611_),
    .B1(_08575_));
 sg13g2_nand4_1 _14420_ (.B(_08607_),
    .C(_08610_),
    .A(_07838_),
    .Y(_08612_),
    .D(_08611_));
 sg13g2_nand2_2 _14421_ (.Y(_08613_),
    .A(_07751_),
    .B(_08599_));
 sg13g2_xor2_1 _14422_ (.B(_07675_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint[31] ),
    .X(_08614_));
 sg13g2_nand3_1 _14423_ (.B(\fpga_top.uart_top.uart_rec_char.bpoint_ld ),
    .C(\fpga_top.uart_top.uart_rec_char.bpoint_en ),
    .A(\fpga_top.cmd_ld_ma ),
    .Y(_08615_));
 sg13g2_or4_1 _14424_ (.A(_08612_),
    .B(_08613_),
    .C(_08614_),
    .D(_08615_),
    .X(_08616_));
 sg13g2_nand3b_1 _14425_ (.B(\fpga_top.uart_top.uart_rec_char.bpoint_en ),
    .C(\fpga_top.cmd_st_ma ),
    .Y(_08617_),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint_ld ));
 sg13g2_nor4_2 _14426_ (.A(_08612_),
    .B(_08613_),
    .C(_08614_),
    .Y(_08618_),
    .D(_08617_));
 sg13g2_or4_1 _14427_ (.A(_08612_),
    .B(_08613_),
    .C(_08614_),
    .D(_08617_),
    .X(_08619_));
 sg13g2_nand2_1 _14428_ (.Y(_08620_),
    .A(net5386),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[2] ));
 sg13g2_nand2_1 _14429_ (.Y(_08621_),
    .A(_06599_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[12] ));
 sg13g2_nand2b_1 _14430_ (.Y(_08622_),
    .B(\fpga_top.bus_gather.i_read_adr[25] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[25] ));
 sg13g2_nor2_1 _14431_ (.A(_06587_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[5] ),
    .Y(_08623_));
 sg13g2_nand2_1 _14432_ (.Y(_08624_),
    .A(_06605_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[15] ));
 sg13g2_nor2_1 _14433_ (.A(_06629_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[24] ),
    .Y(_08625_));
 sg13g2_nand2_1 _14434_ (.Y(_08626_),
    .A(_06643_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[30] ));
 sg13g2_nor2_1 _14435_ (.A(net5595),
    .B(_06591_),
    .Y(_08627_));
 sg13g2_xnor2_1 _14436_ (.Y(_08628_),
    .A(\fpga_top.bus_gather.i_read_adr[21] ),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[21] ));
 sg13g2_nand2_1 _14437_ (.Y(_08629_),
    .A(_06590_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[7] ));
 sg13g2_nand2b_1 _14438_ (.Y(_08630_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[28] ),
    .A_N(net5590));
 sg13g2_xor2_1 _14439_ (.B(\fpga_top.uart_top.uart_rec_char.bpoint[13] ),
    .A(\fpga_top.bus_gather.i_read_adr[13] ),
    .X(_08631_));
 sg13g2_xor2_1 _14440_ (.B(\fpga_top.uart_top.uart_rec_char.bpoint[14] ),
    .A(\fpga_top.bus_gather.i_read_adr[14] ),
    .X(_08632_));
 sg13g2_nand2b_1 _14441_ (.Y(_08633_),
    .B(\fpga_top.bus_gather.i_read_adr[12] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[12] ));
 sg13g2_nand2b_1 _14442_ (.Y(_08634_),
    .B(net5597),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[4] ));
 sg13g2_nand2_1 _14443_ (.Y(_08635_),
    .A(_06631_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[25] ));
 sg13g2_xor2_1 _14444_ (.B(\fpga_top.uart_top.uart_rec_char.bpoint[19] ),
    .A(\fpga_top.bus_gather.i_read_adr[19] ),
    .X(_08636_));
 sg13g2_nor2_1 _14445_ (.A(net5386),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[2] ),
    .Y(_08637_));
 sg13g2_nand2b_1 _14446_ (.Y(_08638_),
    .B(net5591),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[22] ));
 sg13g2_nand2_1 _14447_ (.Y(_08639_),
    .A(net5595),
    .B(_06591_));
 sg13g2_nand2b_1 _14448_ (.Y(_08640_),
    .B(\fpga_top.bus_gather.i_read_adr[7] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[7] ));
 sg13g2_nand2_1 _14449_ (.Y(_08641_),
    .A(_06636_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[27] ));
 sg13g2_nand2b_1 _14450_ (.Y(_08642_),
    .B(\fpga_top.bus_gather.i_read_adr[3] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[3] ));
 sg13g2_nand2b_1 _14451_ (.Y(_08643_),
    .B(\fpga_top.bus_gather.i_read_adr[17] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[17] ));
 sg13g2_nand2b_1 _14452_ (.Y(_08644_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[4] ),
    .A_N(net5597));
 sg13g2_nand2b_1 _14453_ (.Y(_08645_),
    .B(\fpga_top.bus_gather.i_read_adr[31] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[31] ));
 sg13g2_nand2b_1 _14454_ (.Y(_08646_),
    .B(\fpga_top.bus_gather.i_read_adr[15] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[15] ));
 sg13g2_nand2b_1 _14455_ (.Y(_08647_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[22] ),
    .A_N(net5591));
 sg13g2_nand2_1 _14456_ (.Y(_08648_),
    .A(_06611_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[17] ));
 sg13g2_nand2_1 _14457_ (.Y(_08649_),
    .A(_06646_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[31] ));
 sg13g2_nand2b_1 _14458_ (.Y(_08650_),
    .B(net5590),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[28] ));
 sg13g2_nor2_1 _14459_ (.A(\fpga_top.bus_gather.i_read_adr[18] ),
    .B(_06615_),
    .Y(_08651_));
 sg13g2_nand2_1 _14460_ (.Y(_08652_),
    .A(_06584_),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[3] ));
 sg13g2_nand2b_1 _14461_ (.Y(_08653_),
    .B(\fpga_top.bus_gather.i_read_adr[29] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.bpoint[29] ));
 sg13g2_xnor2_1 _14462_ (.Y(_08654_),
    .A(\fpga_top.bus_gather.i_read_adr[9] ),
    .B(\fpga_top.uart_top.uart_rec_char.bpoint[9] ));
 sg13g2_nand4_1 _14463_ (.B(_08622_),
    .C(_08629_),
    .A(_08620_),
    .Y(_08655_),
    .D(_08654_));
 sg13g2_a22oi_1 _14464_ (.Y(_08656_),
    .B1(\fpga_top.bus_gather.i_read_adr[27] ),
    .B2(_06637_),
    .A2(\fpga_top.uart_top.uart_rec_char.bpoint[6] ),
    .A1(_06588_));
 sg13g2_nand4_1 _14465_ (.B(_08649_),
    .C(_08652_),
    .A(_08630_),
    .Y(_08657_),
    .D(_08656_));
 sg13g2_a221oi_1 _14466_ (.B2(\fpga_top.uart_top.uart_rec_char.bpoint[29] ),
    .C1(_08625_),
    .B1(_06641_),
    .A1(\fpga_top.bus_gather.i_read_adr[20] ),
    .Y(_08658_),
    .A2(_06621_));
 sg13g2_nand4_1 _14467_ (.B(_08624_),
    .C(_08626_),
    .A(_08621_),
    .Y(_08659_),
    .D(_08658_));
 sg13g2_a22oi_1 _14468_ (.Y(_08660_),
    .B1(_06626_),
    .B2(\fpga_top.uart_top.uart_rec_char.bpoint[23] ),
    .A2(_06615_),
    .A1(\fpga_top.bus_gather.i_read_adr[18] ));
 sg13g2_nand4_1 _14469_ (.B(_08648_),
    .C(_08653_),
    .A(_08638_),
    .Y(_08661_),
    .D(_08660_));
 sg13g2_a221oi_1 _14470_ (.B2(_06627_),
    .C1(_08661_),
    .B1(\fpga_top.bus_gather.i_read_adr[23] ),
    .A1(net5593),
    .Y(_08662_),
    .A2(_06609_));
 sg13g2_nand4_1 _14471_ (.B(_08639_),
    .C(_08640_),
    .A(_08634_),
    .Y(_08663_),
    .D(_08647_));
 sg13g2_nor4_1 _14472_ (.A(_08636_),
    .B(_08637_),
    .C(_08651_),
    .D(_08663_),
    .Y(_08664_));
 sg13g2_nand3_1 _14473_ (.B(_08662_),
    .C(_08664_),
    .A(_08646_),
    .Y(_08665_));
 sg13g2_nor4_1 _14474_ (.A(_08655_),
    .B(_08657_),
    .C(_08659_),
    .D(_08665_),
    .Y(_08666_));
 sg13g2_o21ai_1 _14475_ (.B1(_08643_),
    .Y(_08667_),
    .A1(_06597_),
    .A2(\fpga_top.uart_top.uart_rec_char.bpoint[11] ));
 sg13g2_o21ai_1 _14476_ (.B1(_08633_),
    .Y(_08668_),
    .A1(net5593),
    .A2(_06609_));
 sg13g2_xor2_1 _14477_ (.B(\fpga_top.uart_top.uart_rec_char.bpoint[26] ),
    .A(\fpga_top.bus_gather.i_read_adr[26] ),
    .X(_08669_));
 sg13g2_nor2_1 _14478_ (.A(_08632_),
    .B(_08669_),
    .Y(_08670_));
 sg13g2_a22oi_1 _14479_ (.Y(_08671_),
    .B1(_06597_),
    .B2(\fpga_top.uart_top.uart_rec_char.bpoint[11] ),
    .A2(_06595_),
    .A1(\fpga_top.bus_gather.i_read_adr[10] ));
 sg13g2_nand4_1 _14480_ (.B(_08645_),
    .C(_08670_),
    .A(\fpga_top.uart_top.uart_rec_char.bpoint_en ),
    .Y(_08672_),
    .D(_08671_));
 sg13g2_nor4_1 _14481_ (.A(_08631_),
    .B(_08667_),
    .C(_08668_),
    .D(_08672_),
    .Y(_08673_));
 sg13g2_nand3_1 _14482_ (.B(_08641_),
    .C(_08650_),
    .A(_08628_),
    .Y(_08674_));
 sg13g2_nand3_1 _14483_ (.B(_08642_),
    .C(_08644_),
    .A(_08635_),
    .Y(_08675_));
 sg13g2_nor3_1 _14484_ (.A(_08627_),
    .B(_08674_),
    .C(_08675_),
    .Y(_08676_));
 sg13g2_a221oi_1 _14485_ (.B2(_06644_),
    .C1(_08623_),
    .B1(\fpga_top.bus_gather.i_read_adr[30] ),
    .A1(_06594_),
    .Y(_08677_),
    .A2(\fpga_top.uart_top.uart_rec_char.bpoint[10] ));
 sg13g2_a22oi_1 _14486_ (.Y(_08678_),
    .B1(_06629_),
    .B2(\fpga_top.uart_top.uart_rec_char.bpoint[24] ),
    .A2(_06589_),
    .A1(net5596));
 sg13g2_nand2_1 _14487_ (.Y(_08679_),
    .A(_08677_),
    .B(_08678_));
 sg13g2_a221oi_1 _14488_ (.B2(\fpga_top.uart_top.uart_rec_char.bpoint[20] ),
    .C1(_08679_),
    .B1(_06620_),
    .A1(_06587_),
    .Y(_08680_),
    .A2(\fpga_top.uart_top.uart_rec_char.bpoint[5] ));
 sg13g2_and4_1 _14489_ (.A(_08666_),
    .B(_08673_),
    .C(_08676_),
    .D(_08680_),
    .X(_08681_));
 sg13g2_nand4_1 _14490_ (.B(_08673_),
    .C(_08676_),
    .A(_08666_),
    .Y(_08682_),
    .D(_08680_));
 sg13g2_nand3_1 _14491_ (.B(_08619_),
    .C(_08682_),
    .A(_08616_),
    .Y(_08683_));
 sg13g2_a21oi_1 _14492_ (.A1(net5426),
    .A2(_08683_),
    .Y(_08684_),
    .B1(net5227));
 sg13g2_nor2_1 _14493_ (.A(_06953_),
    .B(_07022_),
    .Y(_08685_));
 sg13g2_inv_1 _14494_ (.Y(_08686_),
    .A(_08685_));
 sg13g2_a221oi_1 _14495_ (.B2(net5426),
    .C1(_08686_),
    .B1(_08683_),
    .A1(_06965_),
    .Y(_08687_),
    .A2(_06995_));
 sg13g2_nor2_2 _14496_ (.A(_07008_),
    .B(_07022_),
    .Y(_08688_));
 sg13g2_and2_1 _14497_ (.A(_07001_),
    .B(_08688_),
    .X(_08689_));
 sg13g2_nor4_1 _14498_ (.A(net5628),
    .B(\fpga_top.uart_top.uart_rec_char.pdata[0] ),
    .C(net5627),
    .D(net5625),
    .Y(_08690_));
 sg13g2_a21oi_1 _14499_ (.A1(_06967_),
    .A2(_08690_),
    .Y(_08691_),
    .B1(_06974_));
 sg13g2_a21oi_1 _14500_ (.A1(_06967_),
    .A2(_06969_),
    .Y(_08692_),
    .B1(_06979_));
 sg13g2_a21oi_1 _14501_ (.A1(_08691_),
    .A2(_08692_),
    .Y(_08693_),
    .B1(_06955_));
 sg13g2_o21ai_1 _14502_ (.B1(_07021_),
    .Y(_08694_),
    .A1(_06985_),
    .A2(_06989_));
 sg13g2_nand2_1 _14503_ (.Y(_08695_),
    .A(net5633),
    .B(_07017_));
 sg13g2_a21oi_1 _14504_ (.A1(_08694_),
    .A2(_08695_),
    .Y(_08696_),
    .B1(net5227));
 sg13g2_or4_1 _14505_ (.A(_07011_),
    .B(_08689_),
    .C(_08693_),
    .D(_08696_),
    .X(_08697_));
 sg13g2_nor2_1 _14506_ (.A(_08687_),
    .B(_08697_),
    .Y(_08698_));
 sg13g2_inv_1 _14507_ (.Y(\fpga_top.uart_top.uart_rec_char.next_cmd_status[1] ),
    .A(_08698_));
 sg13g2_nand3_1 _14508_ (.B(net5625),
    .C(_06961_),
    .A(net5627),
    .Y(_08699_));
 sg13g2_nor3_1 _14509_ (.A(\fpga_top.uart_top.uart_rec_char.pdata[4] ),
    .B(_06958_),
    .C(_08699_),
    .Y(_08700_));
 sg13g2_nand3_1 _14510_ (.B(_06959_),
    .C(_06961_),
    .A(net5625),
    .Y(_08701_));
 sg13g2_a21oi_1 _14511_ (.A1(_06976_),
    .A2(_08701_),
    .Y(_08702_),
    .B1(_06955_));
 sg13g2_nor3_1 _14512_ (.A(net5632),
    .B(net5630),
    .C(_06984_),
    .Y(_08703_));
 sg13g2_nand2_1 _14513_ (.Y(_08704_),
    .A(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ),
    .B(_08703_));
 sg13g2_nor3_1 _14514_ (.A(net5633),
    .B(net5227),
    .C(_08704_),
    .Y(_08705_));
 sg13g2_o21ai_1 _14515_ (.B1(_07015_),
    .Y(_08706_),
    .A1(_06990_),
    .A2(_07022_));
 sg13g2_nand2b_1 _14516_ (.Y(_08707_),
    .B(_06998_),
    .A_N(_06987_));
 sg13g2_nor3_1 _14517_ (.A(net6539),
    .B(net5631),
    .C(_06990_),
    .Y(_08708_));
 sg13g2_nor2_1 _14518_ (.A(net5235),
    .B(_08708_),
    .Y(_08709_));
 sg13g2_nor2b_1 _14519_ (.A(_08709_),
    .B_N(_06999_),
    .Y(_08710_));
 sg13g2_a221oi_1 _14520_ (.B2(_06985_),
    .C1(_08706_),
    .B1(_08707_),
    .A1(net5633),
    .Y(_08711_),
    .A2(_07007_));
 sg13g2_nor2_1 _14521_ (.A(net5227),
    .B(_08711_),
    .Y(_08712_));
 sg13g2_or4_1 _14522_ (.A(_08702_),
    .B(_08705_),
    .C(_08710_),
    .D(_08712_),
    .X(\fpga_top.uart_top.uart_rec_char.next_cmd_status[2] ));
 sg13g2_nand3_1 _14523_ (.B(_06954_),
    .C(_07004_),
    .A(net5624),
    .Y(_08713_));
 sg13g2_nand2_1 _14524_ (.Y(_08714_),
    .A(net5633),
    .B(_08688_));
 sg13g2_a221oi_1 _14525_ (.B2(_06546_),
    .C1(_08706_),
    .B1(_07018_),
    .A1(net5630),
    .Y(_08715_),
    .A2(_07004_));
 sg13g2_and3_1 _14526_ (.X(_08716_),
    .A(_08713_),
    .B(_08714_),
    .C(_08715_));
 sg13g2_a21oi_1 _14527_ (.A1(_06968_),
    .A2(_08691_),
    .Y(_08717_),
    .B1(_06955_));
 sg13g2_nor2_1 _14528_ (.A(_08710_),
    .B(_08717_),
    .Y(_08718_));
 sg13g2_o21ai_1 _14529_ (.B1(_08718_),
    .Y(\fpga_top.uart_top.uart_rec_char.next_cmd_status[3] ),
    .A1(net5227),
    .A2(_08716_));
 sg13g2_a21oi_1 _14530_ (.A1(_06967_),
    .A2(_06972_),
    .Y(_08719_),
    .B1(_08700_));
 sg13g2_a21oi_1 _14531_ (.A1(_06981_),
    .A2(_08719_),
    .Y(_08720_),
    .B1(_06955_));
 sg13g2_nor3_1 _14532_ (.A(net5630),
    .B(net5228),
    .C(_07008_),
    .Y(_08721_));
 sg13g2_o21ai_1 _14533_ (.B1(_07001_),
    .Y(_08722_),
    .A1(_07009_),
    .A2(_08688_));
 sg13g2_nor3_1 _14534_ (.A(_08705_),
    .B(_08720_),
    .C(_08721_),
    .Y(_08723_));
 sg13g2_nand2_1 _14535_ (.Y(\fpga_top.uart_top.uart_rec_char.next_cmd_status[4] ),
    .A(_08722_),
    .B(_08723_));
 sg13g2_nor2b_1 _14536_ (.A(\fpga_top.uart_top.uart_logics.status_dump[1] ),
    .B_N(\fpga_top.uart_top.uart_logics.status_dump[0] ),
    .Y(_08724_));
 sg13g2_nor2b_2 _14537_ (.A(net6573),
    .B_N(_08724_),
    .Y(\fpga_top.uart_top.uart_logics.radr_enable ));
 sg13g2_nor3_2 _14538_ (.A(net3944),
    .B(net3911),
    .C(net4067),
    .Y(_08725_));
 sg13g2_nor2b_2 _14539_ (.A(net1489),
    .B_N(_08725_),
    .Y(_08726_));
 sg13g2_nand2b_2 _14540_ (.Y(_08727_),
    .B(_08725_),
    .A_N(net1489));
 sg13g2_nand2_2 _14541_ (.Y(_08728_),
    .A(net3978),
    .B(_08726_));
 sg13g2_nor2_1 _14542_ (.A(net5351),
    .B(_08728_),
    .Y(_08729_));
 sg13g2_nand3_1 _14543_ (.B(net5353),
    .C(_08726_),
    .A(net3978),
    .Y(_08730_));
 sg13g2_nand2_1 _14544_ (.Y(_08731_),
    .A(_06988_),
    .B(net5228));
 sg13g2_nor2b_1 _14545_ (.A(\fpga_top.uart_top.uart_logics.status_dump[2] ),
    .B_N(net1851),
    .Y(_08732_));
 sg13g2_and4_1 _14546_ (.A(net6458),
    .B(net5098),
    .C(_08731_),
    .D(_08732_),
    .X(_08733_));
 sg13g2_inv_1 _14547_ (.Y(_08734_),
    .A(_08733_));
 sg13g2_nand2_1 _14548_ (.Y(_08735_),
    .A(net5228),
    .B(_08708_));
 sg13g2_nor2b_1 _14549_ (.A(net6458),
    .B_N(_08732_),
    .Y(_08736_));
 sg13g2_nand2_1 _14550_ (.Y(_08737_),
    .A(_08735_),
    .B(_08736_));
 sg13g2_o21ai_1 _14551_ (.B1(net5228),
    .Y(_08738_),
    .A1(_06988_),
    .A2(_08708_));
 sg13g2_nor2_1 _14552_ (.A(net5423),
    .B(\fpga_top.uart_top.uart_send_char.send_cntr[2] ),
    .Y(_08739_));
 sg13g2_nor3_2 _14553_ (.A(net5423),
    .B(net5422),
    .C(\fpga_top.uart_top.uart_send_char.send_cntr[2] ),
    .Y(_08740_));
 sg13g2_nor2b_2 _14554_ (.A(net6117),
    .B_N(\fpga_top.uart_top.uart_send_char.send_cntr[4] ),
    .Y(_08741_));
 sg13g2_nand2b_2 _14555_ (.Y(_08742_),
    .B(net6318),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[3] ));
 sg13g2_or3_1 _14556_ (.A(net5424),
    .B(net5423),
    .C(_08742_),
    .X(_08743_));
 sg13g2_nor3_1 _14557_ (.A(net5424),
    .B(net5423),
    .C(net6297),
    .Y(_08744_));
 sg13g2_nand2_1 _14558_ (.Y(_08745_),
    .A(_06501_),
    .B(_08740_));
 sg13g2_nor2_1 _14559_ (.A(net5340),
    .B(_08745_),
    .Y(_08746_));
 sg13g2_nand3_1 _14560_ (.B(_08740_),
    .C(net5341),
    .A(_06501_),
    .Y(_08747_));
 sg13g2_and2_1 _14561_ (.A(\fpga_top.uart_top.uart_logics.status_dump[2] ),
    .B(_06997_),
    .X(_08748_));
 sg13g2_nor2b_1 _14562_ (.A(net1851),
    .B_N(\fpga_top.uart_top.uart_logics.status_dump[2] ),
    .Y(\fpga_top.uart_top.uart_logics.rdata_snd_wait ));
 sg13g2_nand3_1 _14563_ (.B(_08747_),
    .C(net1852),
    .A(_08738_),
    .Y(_08749_));
 sg13g2_o21ai_1 _14564_ (.B1(net5634),
    .Y(_08750_),
    .A1(_07006_),
    .A2(_07023_));
 sg13g2_nand2b_2 _14565_ (.Y(_08751_),
    .B(\fpga_top.uart_top.uart_rec_char.next_cmd_status[0] ),
    .A_N(\fpga_top.uart_top.uart_rec_char.next_cmd_status[4] ));
 sg13g2_nand2_1 _14566_ (.Y(_08752_),
    .A(\fpga_top.uart_top.uart_rec_char.next_cmd_status[2] ),
    .B(\fpga_top.uart_top.uart_rec_char.next_cmd_status[3] ));
 sg13g2_nor4_2 _14567_ (.A(_06955_),
    .B(_08698_),
    .C(_08751_),
    .Y(_08753_),
    .D(_08752_));
 sg13g2_nand3_1 _14568_ (.B(_08750_),
    .C(_08753_),
    .A(net6459),
    .Y(_08754_));
 sg13g2_nand4_1 _14569_ (.B(_08737_),
    .C(_08749_),
    .A(_08734_),
    .Y(\fpga_top.uart_top.uart_logics.next_status_dump[2] ),
    .D(_08754_));
 sg13g2_nand2_1 _14570_ (.Y(_08755_),
    .A(net2500),
    .B(_06540_));
 sg13g2_a22oi_1 _14571_ (.Y(_08756_),
    .B1(_06541_),
    .B2(net5613),
    .A2(\fpga_top.bus_gather.u_read_adr[31] ),
    .A1(_06539_));
 sg13g2_nand2_1 _14572_ (.Y(_08757_),
    .A(_06534_),
    .B(\fpga_top.uart_top.uart_logics.cmd_read_end[29] ));
 sg13g2_a22oi_1 _14573_ (.Y(_08758_),
    .B1(\fpga_top.bus_gather.u_read_adr[28] ),
    .B2(_06536_),
    .A2(_06535_),
    .A1(\fpga_top.bus_gather.u_read_adr[29] ));
 sg13g2_a22oi_1 _14574_ (.Y(_08759_),
    .B1(\fpga_top.bus_gather.u_read_adr[26] ),
    .B2(_06538_),
    .A2(_06537_),
    .A1(\fpga_top.bus_gather.u_read_adr[27] ));
 sg13g2_nand2b_1 _14575_ (.Y(_08760_),
    .B(\fpga_top.uart_top.uart_logics.cmd_read_end[28] ),
    .A_N(\fpga_top.bus_gather.u_read_adr[28] ));
 sg13g2_o21ai_1 _14576_ (.B1(_08760_),
    .Y(_08761_),
    .A1(\fpga_top.bus_gather.u_read_adr[27] ),
    .A2(_06537_));
 sg13g2_o21ai_1 _14577_ (.B1(_08758_),
    .Y(_08762_),
    .A1(_08759_),
    .A2(_08761_));
 sg13g2_nand2_1 _14578_ (.Y(_08763_),
    .A(_06516_),
    .B(\fpga_top.bus_gather.u_read_adr[16] ));
 sg13g2_o21ai_1 _14579_ (.B1(_08763_),
    .Y(_08764_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[17] ),
    .A2(_06515_));
 sg13g2_nand2_1 _14580_ (.Y(_08765_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[17] ),
    .B(_06515_));
 sg13g2_nor2b_1 _14581_ (.A(\fpga_top.bus_gather.u_read_adr[15] ),
    .B_N(\fpga_top.uart_top.uart_logics.cmd_read_end[15] ),
    .Y(_08766_));
 sg13g2_o21ai_1 _14582_ (.B1(_08765_),
    .Y(_08767_),
    .A1(_06516_),
    .A2(\fpga_top.bus_gather.u_read_adr[16] ));
 sg13g2_nor3_1 _14583_ (.A(_08764_),
    .B(_08766_),
    .C(_08767_),
    .Y(_08768_));
 sg13g2_nand2b_1 _14584_ (.Y(_08769_),
    .B(\fpga_top.bus_gather.u_read_adr[15] ),
    .A_N(\fpga_top.uart_top.uart_logics.cmd_read_end[15] ));
 sg13g2_o21ai_1 _14585_ (.B1(_08769_),
    .Y(_08770_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[14] ),
    .A2(_06518_));
 sg13g2_nand2_1 _14586_ (.Y(_08771_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[7] ),
    .B(_06513_));
 sg13g2_nor2_1 _14587_ (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[6] ),
    .B(_06514_),
    .Y(_08772_));
 sg13g2_nand2b_1 _14588_ (.Y(_08773_),
    .B(net5615),
    .A_N(\fpga_top.uart_top.uart_logics.cmd_read_end[3] ));
 sg13g2_nand3_1 _14589_ (.B(_06504_),
    .C(_08773_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[2] ),
    .Y(_08774_));
 sg13g2_a22oi_1 _14590_ (.Y(_08775_),
    .B1(\fpga_top.uart_top.uart_logics.cmd_read_end[4] ),
    .B2(_06508_),
    .A2(_06505_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[3] ));
 sg13g2_nor2_1 _14591_ (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[4] ),
    .B(_06508_),
    .Y(_08776_));
 sg13g2_a221oi_1 _14592_ (.B2(_08775_),
    .C1(_08776_),
    .B1(_08774_),
    .A1(_06506_),
    .Y(_08777_),
    .A2(\fpga_top.bus_gather.u_read_adr[5] ));
 sg13g2_a221oi_1 _14593_ (.B2(_06514_),
    .C1(_08777_),
    .B1(\fpga_top.uart_top.uart_logics.cmd_read_end[6] ),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[5] ),
    .Y(_08778_),
    .A2(_06507_));
 sg13g2_o21ai_1 _14594_ (.B1(_08771_),
    .Y(_08779_),
    .A1(_08772_),
    .A2(_08778_));
 sg13g2_a22oi_1 _14595_ (.Y(_08780_),
    .B1(_06512_),
    .B2(\fpga_top.bus_gather.u_read_adr[7] ),
    .A2(\fpga_top.bus_gather.u_read_adr[8] ),
    .A1(_06510_));
 sg13g2_a22oi_1 _14596_ (.Y(_08781_),
    .B1(_08779_),
    .B2(_08780_),
    .A2(_06509_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[9] ));
 sg13g2_o21ai_1 _14597_ (.B1(_08781_),
    .Y(_08782_),
    .A1(_06510_),
    .A2(\fpga_top.bus_gather.u_read_adr[8] ));
 sg13g2_o21ai_1 _14598_ (.B1(_08782_),
    .Y(_08783_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[9] ),
    .A2(_06509_));
 sg13g2_nand2_1 _14599_ (.Y(_08784_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[10] ),
    .B(_06523_));
 sg13g2_nand2b_1 _14600_ (.Y(_08785_),
    .B(\fpga_top.bus_gather.u_read_adr[10] ),
    .A_N(\fpga_top.uart_top.uart_logics.cmd_read_end[10] ));
 sg13g2_o21ai_1 _14601_ (.B1(_08785_),
    .Y(_08786_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[11] ),
    .A2(_06522_));
 sg13g2_a21oi_1 _14602_ (.A1(_08783_),
    .A2(_08784_),
    .Y(_08787_),
    .B1(_08786_));
 sg13g2_a221oi_1 _14603_ (.B2(_06522_),
    .C1(_08787_),
    .B1(\fpga_top.uart_top.uart_logics.cmd_read_end[11] ),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[12] ),
    .Y(_08788_),
    .A2(_06521_));
 sg13g2_a21oi_1 _14604_ (.A1(_06519_),
    .A2(\fpga_top.bus_gather.u_read_adr[13] ),
    .Y(_08789_),
    .B1(_08788_));
 sg13g2_o21ai_1 _14605_ (.B1(_08789_),
    .Y(_08790_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[12] ),
    .A2(_06521_));
 sg13g2_a22oi_1 _14606_ (.Y(_08791_),
    .B1(\fpga_top.uart_top.uart_logics.cmd_read_end[13] ),
    .B2(_06520_),
    .A2(_06518_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[14] ));
 sg13g2_a21o_1 _14607_ (.A2(_08791_),
    .A1(_08790_),
    .B1(_08770_),
    .X(_08792_));
 sg13g2_a22oi_1 _14608_ (.Y(_08793_),
    .B1(_08768_),
    .B2(_08792_),
    .A2(_08765_),
    .A1(_08764_));
 sg13g2_a22oi_1 _14609_ (.Y(_08794_),
    .B1(_06533_),
    .B2(\fpga_top.bus_gather.u_read_adr[22] ),
    .A2(net5614),
    .A1(_06524_));
 sg13g2_nor2_1 _14610_ (.A(_06533_),
    .B(\fpga_top.bus_gather.u_read_adr[22] ),
    .Y(_08795_));
 sg13g2_nor2_1 _14611_ (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[25] ),
    .B(_06530_),
    .Y(_08796_));
 sg13g2_nor2_1 _14612_ (.A(_06524_),
    .B(net5614),
    .Y(_08797_));
 sg13g2_nand2b_1 _14613_ (.Y(_08798_),
    .B(\fpga_top.uart_top.uart_logics.cmd_read_end[20] ),
    .A_N(\fpga_top.bus_gather.u_read_adr[20] ));
 sg13g2_a22oi_1 _14614_ (.Y(_08799_),
    .B1(_06528_),
    .B2(\fpga_top.bus_gather.u_read_adr[18] ),
    .A2(\fpga_top.bus_gather.u_read_adr[19] ),
    .A1(_06526_));
 sg13g2_a22oi_1 _14615_ (.Y(_08800_),
    .B1(\fpga_top.uart_top.uart_logics.cmd_read_end[23] ),
    .B2(_06532_),
    .A2(_06531_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[24] ));
 sg13g2_nand2_1 _14616_ (.Y(_08801_),
    .A(\fpga_top.uart_top.uart_logics.cmd_read_end[25] ),
    .B(_06530_));
 sg13g2_nor2_1 _14617_ (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[24] ),
    .B(_06531_),
    .Y(_08802_));
 sg13g2_nand3b_1 _14618_ (.B(_08800_),
    .C(_08801_),
    .Y(_08803_),
    .A_N(_08802_));
 sg13g2_nor2_1 _14619_ (.A(_06526_),
    .B(\fpga_top.bus_gather.u_read_adr[19] ),
    .Y(_08804_));
 sg13g2_a21o_1 _14620_ (.A2(_06529_),
    .A1(\fpga_top.uart_top.uart_logics.cmd_read_end[18] ),
    .B1(_08804_),
    .X(_08805_));
 sg13g2_nand2b_1 _14621_ (.Y(_08806_),
    .B(\fpga_top.bus_gather.u_read_adr[20] ),
    .A_N(\fpga_top.uart_top.uart_logics.cmd_read_end[20] ));
 sg13g2_nand2b_1 _14622_ (.Y(_08807_),
    .B(\fpga_top.bus_gather.u_read_adr[23] ),
    .A_N(\fpga_top.uart_top.uart_logics.cmd_read_end[23] ));
 sg13g2_nand3b_1 _14623_ (.B(_08798_),
    .C(_08806_),
    .Y(_08808_),
    .A_N(_08797_));
 sg13g2_nor4_1 _14624_ (.A(_08795_),
    .B(_08803_),
    .C(_08805_),
    .D(_08808_),
    .Y(_08809_));
 sg13g2_nor2b_1 _14625_ (.A(_08796_),
    .B_N(_08807_),
    .Y(_08810_));
 sg13g2_nand4_1 _14626_ (.B(_08799_),
    .C(_08809_),
    .A(_08794_),
    .Y(_08811_),
    .D(_08810_));
 sg13g2_nor2_1 _14627_ (.A(_08793_),
    .B(_08811_),
    .Y(_08812_));
 sg13g2_o21ai_1 _14628_ (.B1(_08794_),
    .Y(_08813_),
    .A1(_08797_),
    .A2(_08806_));
 sg13g2_nor3_1 _14629_ (.A(_08799_),
    .B(_08804_),
    .C(_08808_),
    .Y(_08814_));
 sg13g2_nor2_1 _14630_ (.A(_08813_),
    .B(_08814_),
    .Y(_08815_));
 sg13g2_o21ai_1 _14631_ (.B1(_08807_),
    .Y(_08816_),
    .A1(_08795_),
    .A2(_08815_));
 sg13g2_nand2b_1 _14632_ (.Y(_08817_),
    .B(_08816_),
    .A_N(_08803_));
 sg13g2_a21oi_1 _14633_ (.A1(_08801_),
    .A2(_08802_),
    .Y(_08818_),
    .B1(_08796_));
 sg13g2_nand3b_1 _14634_ (.B(_08817_),
    .C(_08818_),
    .Y(_08819_),
    .A_N(_08812_));
 sg13g2_nand2b_1 _14635_ (.Y(_08820_),
    .B(\fpga_top.uart_top.uart_logics.cmd_read_end[26] ),
    .A_N(\fpga_top.bus_gather.u_read_adr[26] ));
 sg13g2_nand4_1 _14636_ (.B(_08758_),
    .C(_08759_),
    .A(_08757_),
    .Y(_08821_),
    .D(_08820_));
 sg13g2_nor2_1 _14637_ (.A(_08761_),
    .B(_08821_),
    .Y(_08822_));
 sg13g2_a22oi_1 _14638_ (.Y(_08823_),
    .B1(_08819_),
    .B2(_08822_),
    .A2(_08762_),
    .A1(_08757_));
 sg13g2_nor2_1 _14639_ (.A(_06541_),
    .B(net5613),
    .Y(_08824_));
 sg13g2_o21ai_1 _14640_ (.B1(_08756_),
    .Y(_08825_),
    .A1(_08823_),
    .A2(_08824_));
 sg13g2_a21oi_2 _14641_ (.B1(net1641),
    .Y(_08826_),
    .A2(_08825_),
    .A1(_08755_));
 sg13g2_nand4_1 _14642_ (.B(_08746_),
    .C(_08748_),
    .A(_08738_),
    .Y(_08827_),
    .D(_08826_));
 sg13g2_nand4_1 _14643_ (.B(_08730_),
    .C(_08731_),
    .A(net6458),
    .Y(_08828_),
    .D(_08732_));
 sg13g2_nand2_1 _14644_ (.Y(_08829_),
    .A(net5285),
    .B(_08735_));
 sg13g2_nand3_1 _14645_ (.B(net6459),
    .C(_07023_),
    .A(net5634),
    .Y(_08830_));
 sg13g2_nand4_1 _14646_ (.B(_08828_),
    .C(_08829_),
    .A(_08827_),
    .Y(\fpga_top.uart_top.uart_logics.next_status_dump[1] ),
    .D(_08830_));
 sg13g2_nand2b_1 _14647_ (.Y(_08831_),
    .B(_08750_),
    .A_N(_08753_));
 sg13g2_a21o_1 _14648_ (.A2(_08826_),
    .A1(net5229),
    .B1(_08747_),
    .X(_08832_));
 sg13g2_nand4_1 _14649_ (.B(_08724_),
    .C(_08738_),
    .A(\fpga_top.uart_top.uart_logics.status_dump[2] ),
    .Y(_08833_),
    .D(_08832_));
 sg13g2_nand4_1 _14650_ (.B(_08827_),
    .C(_08828_),
    .A(_08737_),
    .Y(_08834_),
    .D(_08833_));
 sg13g2_a21o_1 _14651_ (.A2(_08831_),
    .A1(net6459),
    .B1(_08834_),
    .X(\fpga_top.uart_top.uart_logics.next_status_dump[0] ));
 sg13g2_nor2_2 _14652_ (.A(net6192),
    .B(net3827),
    .Y(_08835_));
 sg13g2_inv_4 _14653_ (.A(_08835_),
    .Y(\fpga_top.io_spi_lite.cs_all_status ));
 sg13g2_o21ai_1 _14654_ (.B1(_07027_),
    .Y(_08836_),
    .A1(_08687_),
    .A2(_08697_));
 sg13g2_nor3_1 _14655_ (.A(net6468),
    .B(_07013_),
    .C(_08836_),
    .Y(\fpga_top.uart_top.uart_rec_char.g_crlf ));
 sg13g2_a21oi_2 _14656_ (.B1(_07750_),
    .Y(_08837_),
    .A2(_07674_),
    .A1(_07673_));
 sg13g2_and2_1 _14657_ (.A(net6369),
    .B(_08837_),
    .X(\fpga_top.cpu_top.data_rw_mem.dma_io_radr_en ));
 sg13g2_nor2b_1 _14658_ (.A(net6542),
    .B_N(net6427),
    .Y(_08838_));
 sg13g2_nor2_1 _14659_ (.A(net6427),
    .B(net3934),
    .Y(_08839_));
 sg13g2_nor3_2 _14660_ (.A(\fpga_top.cpu_top.data_rw_mem.data_state[1] ),
    .B(net6427),
    .C(net3934),
    .Y(_08840_));
 sg13g2_o21ai_1 _14661_ (.B1(_08838_),
    .Y(_08841_),
    .A1(net3934),
    .A2(net5174));
 sg13g2_inv_1 _14662_ (.Y(_08842_),
    .A(_08841_));
 sg13g2_a21oi_2 _14663_ (.B1(_08842_),
    .Y(_08843_),
    .A2(net6428),
    .A1(net6369));
 sg13g2_inv_1 _14664_ (.Y(\fpga_top.cpu_top.data_rw_mem.next_data_state[0] ),
    .A(net6429));
 sg13g2_nor2_1 _14665_ (.A(_08838_),
    .B(_08839_),
    .Y(_08844_));
 sg13g2_nand2b_2 _14666_ (.Y(_08845_),
    .B(net6577),
    .A_N(_08837_));
 sg13g2_nand3_1 _14667_ (.B(\fpga_top.cmd_st_ma ),
    .C(_07606_),
    .A(net5379),
    .Y(_08846_));
 sg13g2_or2_1 _14668_ (.X(_08847_),
    .B(_08846_),
    .A(\fpga_top.cmd_ld_ma ));
 sg13g2_o21ai_1 _14669_ (.B1(_08847_),
    .Y(_08848_),
    .A1(_06647_),
    .A2(_08837_));
 sg13g2_nand2b_2 _14670_ (.Y(_08849_),
    .B(net6369),
    .A_N(_08837_));
 sg13g2_nand3_1 _14671_ (.B(_08848_),
    .C(_08849_),
    .A(net6428),
    .Y(_08850_));
 sg13g2_nor2_1 _14672_ (.A(net5683),
    .B(net6195),
    .Y(_08851_));
 sg13g2_nor3_1 _14673_ (.A(net5682),
    .B(net5683),
    .C(\fpga_top.qspi_if.wdata_ofs[1] ),
    .Y(_08852_));
 sg13g2_nand2b_1 _14674_ (.Y(_08853_),
    .B(_08851_),
    .A_N(net5682));
 sg13g2_nand2_1 _14675_ (.Y(_08854_),
    .A(net5629),
    .B(net5354));
 sg13g2_nor2_2 _14676_ (.A(_08853_),
    .B(_08854_),
    .Y(_08855_));
 sg13g2_nand3_1 _14677_ (.B(net5354),
    .C(net5339),
    .A(net5629),
    .Y(_08856_));
 sg13g2_and2_1 _14678_ (.A(\fpga_top.cpu_top.data_rw_mem.data_state[1] ),
    .B(_08839_),
    .X(_08857_));
 sg13g2_a21oi_1 _14679_ (.A1(_08856_),
    .A2(_08857_),
    .Y(_08858_),
    .B1(net3934));
 sg13g2_a21o_2 _14680_ (.A2(_08858_),
    .A1(_08850_),
    .B1(_08844_),
    .X(_08859_));
 sg13g2_inv_1 _14681_ (.Y(\fpga_top.cpu_top.data_rw_mem.next_data_state[1] ),
    .A(net6543));
 sg13g2_or2_1 _14682_ (.X(_08860_),
    .B(\fpga_top.qspi_if.rwait_cntr[1] ),
    .A(\fpga_top.qspi_if.rwait_cntr[0] ));
 sg13g2_or2_1 _14683_ (.X(_08861_),
    .B(_08860_),
    .A(net6473));
 sg13g2_nor2_2 _14684_ (.A(net2398),
    .B(_08861_),
    .Y(_08862_));
 sg13g2_nand2_1 _14685_ (.Y(_08863_),
    .A(net3762),
    .B(_08862_));
 sg13g2_o21ai_1 _14686_ (.B1(net3762),
    .Y(_08864_),
    .A1(net5350),
    .A2(_08863_));
 sg13g2_nor2_2 _14687_ (.A(net5681),
    .B(net6157),
    .Y(_08865_));
 sg13g2_nand3b_1 _14688_ (.B(_08865_),
    .C(net6481),
    .Y(_08866_),
    .A_N(net5680));
 sg13g2_or2_1 _14689_ (.X(_08867_),
    .B(_08866_),
    .A(net5348));
 sg13g2_o21ai_1 _14690_ (.B1(_08864_),
    .Y(_00023_),
    .A1(net5350),
    .A2(_08867_));
 sg13g2_nor2b_1 _14691_ (.A(net1378),
    .B_N(net5624),
    .Y(_00084_));
 sg13g2_o21ai_1 _14692_ (.B1(net5629),
    .Y(_08868_),
    .A1(net5351),
    .A2(_08853_));
 sg13g2_nand2_1 _14693_ (.Y(_08869_),
    .A(net5353),
    .B(net5346));
 sg13g2_o21ai_1 _14694_ (.B1(_08868_),
    .Y(_00014_),
    .A1(_08866_),
    .A2(_08869_));
 sg13g2_nand2_1 _14695_ (.Y(_08870_),
    .A(\fpga_top.qspi_if.qspi_state[11] ),
    .B(_08727_));
 sg13g2_o21ai_1 _14696_ (.B1(net3978),
    .Y(_08871_),
    .A1(net5350),
    .A2(_08727_));
 sg13g2_o21ai_1 _14697_ (.B1(net3979),
    .Y(_00015_),
    .A1(net5350),
    .A2(_08863_));
 sg13g2_nor2_1 _14698_ (.A(net1897),
    .B(net2176),
    .Y(_08872_));
 sg13g2_nor4_1 _14699_ (.A(net1390),
    .B(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[0] ),
    .C(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[3] ),
    .D(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[2] ),
    .Y(_08873_));
 sg13g2_inv_2 _14700_ (.Y(\fpga_top.uart_top.rx_fifo_dvalid ),
    .A(net5338));
 sg13g2_nor3_2 _14701_ (.A(_06546_),
    .B(_06990_),
    .C(_07022_),
    .Y(_08874_));
 sg13g2_and3_2 _14702_ (.X(_08875_),
    .A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[30] ),
    .B(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[31] ),
    .C(_08874_));
 sg13g2_and3_1 _14703_ (.X(_08876_),
    .A(\fpga_top.dma_io_wadr_u[14] ),
    .B(\fpga_top.dma_io_wadr_u[15] ),
    .C(net5083));
 sg13g2_a221oi_1 _14704_ (.B2(_07749_),
    .C1(_08846_),
    .B1(_07748_),
    .A1(_07673_),
    .Y(_08877_),
    .A2(_07674_));
 sg13g2_nand2_1 _14705_ (.Y(_08878_),
    .A(_07944_),
    .B(_08548_));
 sg13g2_nor2_1 _14706_ (.A(net5084),
    .B(_08878_),
    .Y(_08879_));
 sg13g2_a21o_2 _14707_ (.A2(_08879_),
    .A1(_08877_),
    .B1(_08876_),
    .X(_08880_));
 sg13g2_nand2_1 _14708_ (.Y(_08881_),
    .A(net4035),
    .B(\fpga_top.cpu_top.csr_wadr_mon[11] ));
 sg13g2_nand2_2 _14709_ (.Y(_08882_),
    .A(net5083),
    .B(_08881_));
 sg13g2_nand2_2 _14710_ (.Y(_08883_),
    .A(_07970_),
    .B(_08345_));
 sg13g2_nand2b_2 _14711_ (.Y(_08884_),
    .B(_08883_),
    .A_N(net5080));
 sg13g2_and2_1 _14712_ (.A(_08882_),
    .B(_08884_),
    .X(_08885_));
 sg13g2_and2_1 _14713_ (.A(_08880_),
    .B(_08885_),
    .X(_08886_));
 sg13g2_nand2_1 _14714_ (.Y(_08887_),
    .A(\fpga_top.cpu_top.csr_wadr_mon[8] ),
    .B(net5081));
 sg13g2_o21ai_1 _14715_ (.B1(_08887_),
    .Y(_08888_),
    .A1(_08012_),
    .A2(net5081));
 sg13g2_inv_1 _14716_ (.Y(_08889_),
    .A(_08888_));
 sg13g2_nor2_1 _14717_ (.A(_08279_),
    .B(net5082),
    .Y(_08890_));
 sg13g2_a21oi_2 _14718_ (.B1(_08890_),
    .Y(_08891_),
    .A2(net5082),
    .A1(\fpga_top.cpu_top.csr_wadr_mon[9] ));
 sg13g2_inv_2 _14719_ (.Y(_08892_),
    .A(_08891_));
 sg13g2_nand4_1 _14720_ (.B(_08885_),
    .C(_08889_),
    .A(_08880_),
    .Y(_08893_),
    .D(_08892_));
 sg13g2_nand2_1 _14721_ (.Y(_08894_),
    .A(net5665),
    .B(net5086));
 sg13g2_o21ai_1 _14722_ (.B1(_08894_),
    .Y(_08895_),
    .A1(_08158_),
    .A2(net5082));
 sg13g2_nand2_1 _14723_ (.Y(_08896_),
    .A(\fpga_top.cpu_top.csr_wadr_mon[1] ),
    .B(net5086));
 sg13g2_o21ai_1 _14724_ (.B1(_08896_),
    .Y(_08897_),
    .A1(_08191_),
    .A2(net5082));
 sg13g2_or2_1 _14725_ (.X(_08898_),
    .B(_08897_),
    .A(_08895_));
 sg13g2_nand2_1 _14726_ (.Y(_08899_),
    .A(\fpga_top.cpu_top.csr_wadr_mon[3] ),
    .B(net5085));
 sg13g2_o21ai_1 _14727_ (.B1(_08899_),
    .Y(_08900_),
    .A1(_08101_),
    .A2(net5081));
 sg13g2_mux2_1 _14728_ (.A0(_08222_),
    .A1(\fpga_top.cpu_top.csr_wadr_mon[2] ),
    .S(net5081),
    .X(_08901_));
 sg13g2_nand2b_2 _14729_ (.Y(_08902_),
    .B(_08901_),
    .A_N(_08900_));
 sg13g2_nor3_1 _14730_ (.A(\fpga_top.cpu_top.csr_wadr_mon[4] ),
    .B(\fpga_top.cpu_top.csr_wadr_mon[5] ),
    .C(\fpga_top.cpu_top.csr_wadr_mon[6] ),
    .Y(_08903_));
 sg13g2_nand2_1 _14731_ (.Y(_08904_),
    .A(net5081),
    .B(_08903_));
 sg13g2_nand3_1 _14732_ (.B(_08128_),
    .C(_08247_),
    .A(_08073_),
    .Y(_08905_));
 sg13g2_o21ai_1 _14733_ (.B1(_08904_),
    .Y(_08906_),
    .A1(net5082),
    .A2(_08905_));
 sg13g2_nor2_1 _14734_ (.A(_08313_),
    .B(net5081),
    .Y(_08907_));
 sg13g2_a21oi_2 _14735_ (.B1(_08907_),
    .Y(_08908_),
    .A2(net5081),
    .A1(\fpga_top.cpu_top.csr_wadr_mon[7] ));
 sg13g2_and2_1 _14736_ (.A(_08906_),
    .B(_08908_),
    .X(_08909_));
 sg13g2_nand2b_2 _14737_ (.Y(_08910_),
    .B(_08909_),
    .A_N(_08902_));
 sg13g2_or2_1 _14738_ (.X(_08911_),
    .B(_08910_),
    .A(_08898_));
 sg13g2_nor2_2 _14739_ (.A(_08893_),
    .B(_08911_),
    .Y(_08912_));
 sg13g2_nor2b_1 _14740_ (.A(net5087),
    .B_N(\fpga_top.bus_gather.d_write_data[2] ),
    .Y(_08913_));
 sg13g2_a21oi_1 _14741_ (.A1(net5664),
    .A2(net5086),
    .Y(_08914_),
    .B1(_08913_));
 sg13g2_a21o_2 _14742_ (.A2(net5085),
    .A1(net5664),
    .B1(_08913_),
    .X(_08915_));
 sg13g2_nor3_1 _14743_ (.A(_08893_),
    .B(_08911_),
    .C(_08915_),
    .Y(\fpga_top.io_frc.frc_cntr_val_rst_pre ));
 sg13g2_o21ai_1 _14744_ (.B1(\fpga_top.cpu_top.csr_rmie ),
    .Y(_08916_),
    .A1(\fpga_top.interrupter.int_status_int0 ),
    .A2(\fpga_top.interrupter.int_status_rx ));
 sg13g2_inv_2 _14745_ (.Y(\fpga_top.cpu_top.execution.csr_array.g_interrupt ),
    .A(_08916_));
 sg13g2_and2_1 _14746_ (.A(\fpga_top.qspi_if.dbg_2div_trt ),
    .B(net6153),
    .X(_08917_));
 sg13g2_mux2_1 _14747_ (.A0(net3926),
    .A1(net6154),
    .S(net5353),
    .X(_00017_));
 sg13g2_nor2b_1 _14748_ (.A(_06943_),
    .B_N(net1534),
    .Y(_00016_));
 sg13g2_nor2_1 _14749_ (.A(net6602),
    .B(net6420),
    .Y(_08918_));
 sg13g2_nand2_2 _14750_ (.Y(_08919_),
    .A(_06938_),
    .B(_08918_));
 sg13g2_nor2_1 _14751_ (.A(\fpga_top.qspi_if.cmd_ofs[2] ),
    .B(_08919_),
    .Y(_08920_));
 sg13g2_or2_1 _14752_ (.X(_08921_),
    .B(_08919_),
    .A(\fpga_top.qspi_if.cmd_ofs[2] ));
 sg13g2_o21ai_1 _14753_ (.B1(net3898),
    .Y(_08922_),
    .A1(net5350),
    .A2(_08921_));
 sg13g2_nor2_1 _14754_ (.A(_00125_),
    .B(_06937_),
    .Y(_08923_));
 sg13g2_nand2b_1 _14755_ (.Y(_08924_),
    .B(_06938_),
    .A_N(net3975));
 sg13g2_o21ai_1 _14756_ (.B1(_08922_),
    .Y(_00021_),
    .A1(net5350),
    .A2(_08924_));
 sg13g2_nor2_1 _14757_ (.A(net1375),
    .B(net5351),
    .Y(_08925_));
 sg13g2_o21ai_1 _14758_ (.B1(_08925_),
    .Y(_08926_),
    .A1(\fpga_top.qspi_if.dbg_2div_read_half_end ),
    .A2(_08728_));
 sg13g2_o21ai_1 _14759_ (.B1(_08926_),
    .Y(_08927_),
    .A1(\fpga_top.qspi_if.qspi_state[4] ),
    .A2(net5353));
 sg13g2_o21ai_1 _14760_ (.B1(_08927_),
    .Y(_00019_),
    .A1(net3326),
    .A2(_08856_));
 sg13g2_nor2b_1 _14761_ (.A(_06943_),
    .B_N(net1400),
    .Y(_08928_));
 sg13g2_inv_1 _14762_ (.Y(_08929_),
    .A(_08928_));
 sg13g2_a21o_1 _14763_ (.A2(_06943_),
    .A1(net1534),
    .B1(_08928_),
    .X(_00022_));
 sg13g2_and2_1 _14764_ (.A(net3326),
    .B(_08855_),
    .X(_08930_));
 sg13g2_a21oi_1 _14765_ (.A1(net1375),
    .A2(net5351),
    .Y(_08931_),
    .B1(_08930_));
 sg13g2_o21ai_1 _14766_ (.B1(_08931_),
    .Y(_00020_),
    .A1(_06671_),
    .A2(_08730_));
 sg13g2_nor3_1 _14767_ (.A(net5350),
    .B(_06937_),
    .C(_08866_),
    .Y(_08932_));
 sg13g2_nand3_1 _14768_ (.B(net5353),
    .C(_08920_),
    .A(net3898),
    .Y(_08933_));
 sg13g2_o21ai_1 _14769_ (.B1(net3899),
    .Y(_00018_),
    .A1(net5378),
    .A2(_08932_));
 sg13g2_nor2_2 _14770_ (.A(\fpga_top.cpu_top.data_rw_mem.dma_io_radr_en ),
    .B(_08877_),
    .Y(_08934_));
 sg13g2_nor2b_1 _14771_ (.A(_08934_),
    .B_N(_08840_),
    .Y(_08935_));
 sg13g2_a21o_1 _14772_ (.A2(_08838_),
    .A1(net3934),
    .B1(_08935_),
    .X(\fpga_top.cpu_top.data_rw_mem.next_data_state[2] ));
 sg13g2_nand2b_1 _14773_ (.Y(_08936_),
    .B(\fpga_top.io_spi_lite.spi_sck_div[4] ),
    .A_N(\fpga_top.io_spi_lite.sck_div[4] ));
 sg13g2_nand2b_1 _14774_ (.Y(_08937_),
    .B(\fpga_top.io_spi_lite.sck_div[5] ),
    .A_N(\fpga_top.io_spi_lite.spi_sck_div[5] ));
 sg13g2_nand2b_1 _14775_ (.Y(_08938_),
    .B(\fpga_top.io_spi_lite.spi_sck_div[6] ),
    .A_N(\fpga_top.io_spi_lite.sck_div[6] ));
 sg13g2_o21ai_1 _14776_ (.B1(_08937_),
    .Y(_08939_),
    .A1(_06778_),
    .A2(\fpga_top.io_spi_lite.spi_sck_div[2] ));
 sg13g2_o21ai_1 _14777_ (.B1(_08936_),
    .Y(_08940_),
    .A1(\fpga_top.io_spi_lite.sck_div[8] ),
    .A2(_06783_));
 sg13g2_xor2_1 _14778_ (.B(\fpga_top.io_spi_lite.spi_sck_div[1] ),
    .A(\fpga_top.io_spi_lite.sck_div[1] ),
    .X(_08941_));
 sg13g2_a221oi_1 _14779_ (.B2(_06783_),
    .C1(_08941_),
    .B1(\fpga_top.io_spi_lite.sck_div[8] ),
    .A1(\fpga_top.io_spi_lite.sck_div[6] ),
    .Y(_08942_),
    .A2(_06781_));
 sg13g2_o21ai_1 _14780_ (.B1(_08942_),
    .Y(_08943_),
    .A1(_06782_),
    .A2(net1621));
 sg13g2_xor2_1 _14781_ (.B(\fpga_top.io_spi_lite.spi_sck_div[3] ),
    .A(\fpga_top.io_spi_lite.sck_div[3] ),
    .X(_08944_));
 sg13g2_a221oi_1 _14782_ (.B2(\fpga_top.io_spi_lite.spi_sck_div[9] ),
    .C1(_08944_),
    .B1(_06784_),
    .A1(_06780_),
    .Y(_08945_),
    .A2(\fpga_top.io_spi_lite.spi_sck_div[5] ));
 sg13g2_xor2_1 _14783_ (.B(\fpga_top.io_spi_lite.spi_sck_div[0] ),
    .A(\fpga_top.io_spi_lite.sck_div[0] ),
    .X(_08946_));
 sg13g2_a221oi_1 _14784_ (.B2(\fpga_top.io_spi_lite.spi_sck_div[7] ),
    .C1(_08946_),
    .B1(_06782_),
    .A1(_06778_),
    .Y(_08947_),
    .A2(\fpga_top.io_spi_lite.spi_sck_div[2] ));
 sg13g2_a22oi_1 _14785_ (.Y(_08948_),
    .B1(\fpga_top.io_spi_lite.sck_div[9] ),
    .B2(_06785_),
    .A2(_06779_),
    .A1(\fpga_top.io_spi_lite.sck_div[4] ));
 sg13g2_nand4_1 _14786_ (.B(_08945_),
    .C(_08947_),
    .A(_08938_),
    .Y(_08949_),
    .D(_08948_));
 sg13g2_nor4_1 _14787_ (.A(_08939_),
    .B(_08940_),
    .C(_08943_),
    .D(_08949_),
    .Y(_08950_));
 sg13g2_nor2_1 _14788_ (.A(net1404),
    .B(net5075),
    .Y(_00028_));
 sg13g2_xnor2_1 _14789_ (.Y(_08951_),
    .A(net1404),
    .B(net3797));
 sg13g2_nor2_1 _14790_ (.A(net5075),
    .B(_08951_),
    .Y(_00029_));
 sg13g2_a21oi_1 _14791_ (.A1(net1404),
    .A2(\fpga_top.io_spi_lite.sck_div[1] ),
    .Y(_08952_),
    .B1(net1899));
 sg13g2_and3_1 _14792_ (.X(_08953_),
    .A(net1404),
    .B(net3797),
    .C(net1899));
 sg13g2_nor3_1 _14793_ (.A(net5076),
    .B(net1900),
    .C(_08953_),
    .Y(_00030_));
 sg13g2_nor2_1 _14794_ (.A(net4001),
    .B(_08953_),
    .Y(_08954_));
 sg13g2_and2_1 _14795_ (.A(net4001),
    .B(_08953_),
    .X(_08955_));
 sg13g2_nor3_1 _14796_ (.A(net5076),
    .B(_08954_),
    .C(_08955_),
    .Y(_00031_));
 sg13g2_nor2_1 _14797_ (.A(net3871),
    .B(_08955_),
    .Y(_08956_));
 sg13g2_and2_1 _14798_ (.A(net3871),
    .B(_08955_),
    .X(_08957_));
 sg13g2_nor3_1 _14799_ (.A(net5075),
    .B(net3872),
    .C(_08957_),
    .Y(_00032_));
 sg13g2_nor2_1 _14800_ (.A(net3874),
    .B(_08957_),
    .Y(_08958_));
 sg13g2_and2_1 _14801_ (.A(net3874),
    .B(_08957_),
    .X(_08959_));
 sg13g2_nor3_1 _14802_ (.A(net5075),
    .B(net3875),
    .C(_08959_),
    .Y(_00033_));
 sg13g2_nor2_1 _14803_ (.A(net3878),
    .B(_08959_),
    .Y(_08960_));
 sg13g2_and2_1 _14804_ (.A(net3878),
    .B(_08959_),
    .X(_08961_));
 sg13g2_nor3_1 _14805_ (.A(net5075),
    .B(_08960_),
    .C(_08961_),
    .Y(_00034_));
 sg13g2_nor2_1 _14806_ (.A(net3725),
    .B(_08961_),
    .Y(_08962_));
 sg13g2_and2_1 _14807_ (.A(net3725),
    .B(_08961_),
    .X(_08963_));
 sg13g2_nor3_1 _14808_ (.A(net5075),
    .B(net3726),
    .C(_08963_),
    .Y(_00035_));
 sg13g2_nor2_1 _14809_ (.A(net3893),
    .B(_08963_),
    .Y(_08964_));
 sg13g2_and2_1 _14810_ (.A(net3893),
    .B(_08963_),
    .X(_08965_));
 sg13g2_nor3_1 _14811_ (.A(net5075),
    .B(_08964_),
    .C(_08965_),
    .Y(_00036_));
 sg13g2_a21oi_1 _14812_ (.A1(net6084),
    .A2(_08965_),
    .Y(_08966_),
    .B1(net5075));
 sg13g2_o21ai_1 _14813_ (.B1(_08966_),
    .Y(_08967_),
    .A1(net6084),
    .A2(_08965_));
 sg13g2_inv_1 _14814_ (.Y(_00037_),
    .A(_08967_));
 sg13g2_nand2_1 _14815_ (.Y(_08968_),
    .A(net1975),
    .B(net1703));
 sg13g2_nor2b_1 _14816_ (.A(\fpga_top.io_spi_lite.org_sck ),
    .B_N(\fpga_top.io_spi_lite.org_sck_dly ),
    .Y(_08969_));
 sg13g2_nand2b_1 _14817_ (.Y(_08970_),
    .B(\fpga_top.io_spi_lite.org_sck ),
    .A_N(\fpga_top.io_spi_lite.org_sck_dly ));
 sg13g2_nand2_1 _14818_ (.Y(_08971_),
    .A(\fpga_top.io_spi_lite.spi_mode[1] ),
    .B(_08970_));
 sg13g2_o21ai_1 _14819_ (.B1(_08971_),
    .Y(_08972_),
    .A1(\fpga_top.io_spi_lite.spi_mode[1] ),
    .A2(_08969_));
 sg13g2_nor2_2 _14820_ (.A(_08968_),
    .B(_08972_),
    .Y(_08973_));
 sg13g2_and2_1 _14821_ (.A(net1915),
    .B(_08973_),
    .X(_08974_));
 sg13g2_nand2_2 _14822_ (.Y(_08975_),
    .A(net1915),
    .B(_08973_));
 sg13g2_xnor2_1 _14823_ (.Y(\fpga_top.io_spi_lite.mosi_fifo.radr_early[0] ),
    .A(net1892),
    .B(_08975_));
 sg13g2_nand3_1 _14824_ (.B(net1587),
    .C(_08974_),
    .A(\fpga_top.io_spi_lite.mosi_fifo.radr[0] ),
    .Y(_08976_));
 sg13g2_a21o_1 _14825_ (.A2(_08974_),
    .A1(net1892),
    .B1(net1587),
    .X(_08977_));
 sg13g2_and2_1 _14826_ (.A(net1588),
    .B(_08977_),
    .X(\fpga_top.io_spi_lite.mosi_fifo.radr_early[1] ));
 sg13g2_xnor2_1 _14827_ (.Y(\fpga_top.io_spi_lite.mosi_fifo.radr_early[2] ),
    .A(net1572),
    .B(_08976_));
 sg13g2_xor2_1 _14828_ (.B(net1861),
    .A(net5831),
    .X(\fpga_top.io_spi_lite.miso_fifo.radr_early[0] ));
 sg13g2_nor2b_2 _14829_ (.A(_08908_),
    .B_N(_08906_),
    .Y(_08978_));
 sg13g2_inv_1 _14830_ (.Y(_08979_),
    .A(_08978_));
 sg13g2_nand2_1 _14831_ (.Y(_08980_),
    .A(net5652),
    .B(net5087));
 sg13g2_o21ai_1 _14832_ (.B1(_08980_),
    .Y(_08981_),
    .A1(_06593_),
    .A2(net5087));
 sg13g2_or2_1 _14833_ (.X(_08982_),
    .B(_08901_),
    .A(_08900_));
 sg13g2_nand2_1 _14834_ (.Y(_08983_),
    .A(_08895_),
    .B(_08897_));
 sg13g2_nor2_1 _14835_ (.A(_08982_),
    .B(_08983_),
    .Y(_08984_));
 sg13g2_nand3_1 _14836_ (.B(_08889_),
    .C(_08891_),
    .A(_08886_),
    .Y(_08985_));
 sg13g2_inv_1 _14837_ (.Y(_08986_),
    .A(_08985_));
 sg13g2_nand4_1 _14838_ (.B(_08981_),
    .C(_08984_),
    .A(_08978_),
    .Y(_08987_),
    .D(_08986_));
 sg13g2_and3_1 _14839_ (.X(_08988_),
    .A(_08880_),
    .B(_08882_),
    .C(_08884_));
 sg13g2_nand3_1 _14840_ (.B(_08891_),
    .C(_08988_),
    .A(_08889_),
    .Y(_08989_));
 sg13g2_and2_1 _14841_ (.A(\fpga_top.io_spi_lite.miso_fifo.radr_early[0] ),
    .B(_08987_),
    .X(_00038_));
 sg13g2_nand3_1 _14842_ (.B(net1861),
    .C(net6442),
    .A(net5832),
    .Y(_08990_));
 sg13g2_a21o_1 _14843_ (.A2(net1861),
    .A1(net5832),
    .B1(net6442),
    .X(_08991_));
 sg13g2_and2_1 _14844_ (.A(_08990_),
    .B(_08991_),
    .X(\fpga_top.io_spi_lite.miso_fifo.radr_early[1] ));
 sg13g2_and2_1 _14845_ (.A(_08987_),
    .B(\fpga_top.io_spi_lite.miso_fifo.radr_early[1] ),
    .X(_00039_));
 sg13g2_xnor2_1 _14846_ (.Y(\fpga_top.io_spi_lite.miso_fifo.radr_early[2] ),
    .A(net1991),
    .B(_08990_));
 sg13g2_and2_1 _14847_ (.A(_08987_),
    .B(net1992),
    .X(_00040_));
 sg13g2_mux2_1 _14848_ (.A0(_00087_),
    .A1(_00086_),
    .S(\fpga_top.qspi_if.wredge[0] ),
    .X(_08992_));
 sg13g2_nand2b_1 _14849_ (.Y(_08993_),
    .B(_08992_),
    .A_N(_00094_));
 sg13g2_o21ai_1 _14850_ (.B1(_00094_),
    .Y(_08994_),
    .A1(\fpga_top.qspi_if.wredge[0] ),
    .A2(_00089_));
 sg13g2_a21oi_1 _14851_ (.A1(\fpga_top.qspi_if.wredge[0] ),
    .A2(_06930_),
    .Y(_08995_),
    .B1(_08994_));
 sg13g2_nand3b_1 _14852_ (.B(\fpga_top.qspi_if.wredge[2] ),
    .C(_08993_),
    .Y(_08996_),
    .A_N(_08995_));
 sg13g2_mux4_1 _14853_ (.S0(\fpga_top.qspi_if.wredge[0] ),
    .A0(_00107_),
    .A1(_00095_),
    .A2(_00123_),
    .A3(_00115_),
    .S1(_00094_),
    .X(_08997_));
 sg13g2_o21ai_1 _14854_ (.B1(_08996_),
    .Y(\fpga_top.qspi_if.sck ),
    .A1(\fpga_top.qspi_if.wredge[2] ),
    .A2(_08997_));
 sg13g2_a22oi_1 _14855_ (.Y(_08998_),
    .B1(net5346),
    .B2(net3773),
    .A2(_06933_),
    .A1(net3690));
 sg13g2_nor2_1 _14856_ (.A(net3976),
    .B(_08998_),
    .Y(\fpga_top.qspi_if.dbg_2div_cec_pre ));
 sg13g2_and2_1 _14857_ (.A(\fpga_top.qspi_if.rdwrch[0] ),
    .B(_06950_),
    .X(_08999_));
 sg13g2_a21oi_2 _14858_ (.B1(_08999_),
    .Y(_09000_),
    .A2(_00133_),
    .A1(\fpga_top.qspi_if.rdwrch[2] ));
 sg13g2_a21o_2 _14859_ (.A2(_00133_),
    .A1(\fpga_top.qspi_if.rdwrch[2] ),
    .B1(_08999_),
    .X(_09001_));
 sg13g2_o21ai_1 _14860_ (.B1(net5349),
    .Y(_09002_),
    .A1(\fpga_top.qspi_if.rdcmd0[2] ),
    .A2(net4949));
 sg13g2_a21oi_1 _14861_ (.A1(_06818_),
    .A2(net4949),
    .Y(_09003_),
    .B1(_09002_));
 sg13g2_mux2_1 _14862_ (.A0(\fpga_top.qspi_if.rdwrch[3] ),
    .A1(\fpga_top.qspi_if.rdwrch[1] ),
    .S(_06950_),
    .X(_09004_));
 sg13g2_o21ai_1 _14863_ (.B1(net5345),
    .Y(_09005_),
    .A1(\fpga_top.qspi_if.wrcmd0[2] ),
    .A2(net5074));
 sg13g2_a21oi_1 _14864_ (.A1(_06819_),
    .A2(_09004_),
    .Y(_09006_),
    .B1(_09005_));
 sg13g2_nor2_1 _14865_ (.A(_09003_),
    .B(_09006_),
    .Y(_09007_));
 sg13g2_nor2_1 _14866_ (.A(\fpga_top.qspi_if.cmd_ofs[0] ),
    .B(_09007_),
    .Y(_09008_));
 sg13g2_mux2_1 _14867_ (.A0(_00099_),
    .A1(_00096_),
    .S(net5074),
    .X(_09009_));
 sg13g2_mux2_1 _14868_ (.A0(_00110_),
    .A1(_00104_),
    .S(_09001_),
    .X(_09010_));
 sg13g2_a221oi_1 _14869_ (.B2(net5349),
    .C1(_06675_),
    .B1(_09010_),
    .A1(net5346),
    .Y(_09011_),
    .A2(_09009_));
 sg13g2_o21ai_1 _14870_ (.B1(_06948_),
    .Y(_09012_),
    .A1(_09008_),
    .A2(_09011_));
 sg13g2_a21oi_1 _14871_ (.A1(net5684),
    .A2(_06819_),
    .Y(_09013_),
    .B1(_06936_));
 sg13g2_o21ai_1 _14872_ (.B1(_09013_),
    .Y(_09014_),
    .A1(net5685),
    .A2(\fpga_top.qspi_if.wrcmd0[2] ));
 sg13g2_a21oi_1 _14873_ (.A1(net5687),
    .A2(_06818_),
    .Y(_09015_),
    .B1(net5348));
 sg13g2_o21ai_1 _14874_ (.B1(_09015_),
    .Y(_09016_),
    .A1(net5687),
    .A2(\fpga_top.qspi_if.rdcmd0[2] ));
 sg13g2_a21oi_1 _14875_ (.A1(_09014_),
    .A2(_09016_),
    .Y(_09017_),
    .B1(\fpga_top.qspi_if.cmd_ofs[0] ));
 sg13g2_mux2_1 _14876_ (.A0(_00099_),
    .A1(_00096_),
    .S(net5685),
    .X(_09018_));
 sg13g2_mux2_1 _14877_ (.A0(_00110_),
    .A1(_00104_),
    .S(net5687),
    .X(_09019_));
 sg13g2_a221oi_1 _14878_ (.B2(net5349),
    .C1(_06675_),
    .B1(_09019_),
    .A1(net5346),
    .Y(_09020_),
    .A2(_09018_));
 sg13g2_o21ai_1 _14879_ (.B1(_00134_),
    .Y(_09021_),
    .A1(_09017_),
    .A2(_09020_));
 sg13g2_nand3_1 _14880_ (.B(_09012_),
    .C(_09021_),
    .A(\fpga_top.qspi_if.cmd_ofs[1] ),
    .Y(_09022_));
 sg13g2_nand2_1 _14881_ (.Y(_09023_),
    .A(_00109_),
    .B(_09000_));
 sg13g2_a21oi_1 _14882_ (.A1(_00103_),
    .A2(net4949),
    .Y(_09024_),
    .B1(net5347));
 sg13g2_mux2_1 _14883_ (.A0(\fpga_top.qspi_if.wrcmd0[1] ),
    .A1(\fpga_top.qspi_if.wrcmd1[1] ),
    .S(net5074),
    .X(_09025_));
 sg13g2_a22oi_1 _14884_ (.Y(_09026_),
    .B1(_09025_),
    .B2(net5345),
    .A2(_09024_),
    .A1(_09023_));
 sg13g2_nor2_1 _14885_ (.A(_00134_),
    .B(_09026_),
    .Y(_09027_));
 sg13g2_nand2b_1 _14886_ (.Y(_09028_),
    .B(\fpga_top.qspi_if.cmd_ofs[0] ),
    .A_N(\fpga_top.qspi_if.cmd_ofs[1] ));
 sg13g2_mux2_1 _14887_ (.A0(\fpga_top.qspi_if.wrcmd0[1] ),
    .A1(\fpga_top.qspi_if.wrcmd1[1] ),
    .S(net5684),
    .X(_09029_));
 sg13g2_nor2b_1 _14888_ (.A(net5686),
    .B_N(_00109_),
    .Y(_09030_));
 sg13g2_a21oi_1 _14889_ (.A1(_00103_),
    .A2(net5686),
    .Y(_09031_),
    .B1(_09030_));
 sg13g2_a22oi_1 _14890_ (.Y(_09032_),
    .B1(_09031_),
    .B2(net5349),
    .A2(_09029_),
    .A1(net5345));
 sg13g2_nor2_1 _14891_ (.A(_06948_),
    .B(_09032_),
    .Y(_09033_));
 sg13g2_nor3_1 _14892_ (.A(_09027_),
    .B(_09028_),
    .C(_09033_),
    .Y(_09034_));
 sg13g2_o21ai_1 _14893_ (.B1(net5345),
    .Y(_09035_),
    .A1(_06817_),
    .A2(net5074));
 sg13g2_a21oi_1 _14894_ (.A1(\fpga_top.qspi_if.wrcmd1[0] ),
    .A2(net5074),
    .Y(_09036_),
    .B1(_09035_));
 sg13g2_o21ai_1 _14895_ (.B1(net5349),
    .Y(_09037_),
    .A1(_00102_),
    .A2(_09000_));
 sg13g2_a21oi_1 _14896_ (.A1(_06499_),
    .A2(_09000_),
    .Y(_09038_),
    .B1(_09037_));
 sg13g2_nor3_1 _14897_ (.A(_00134_),
    .B(_09036_),
    .C(_09038_),
    .Y(_09039_));
 sg13g2_nor2b_1 _14898_ (.A(net5684),
    .B_N(\fpga_top.qspi_if.wrcmd0[0] ),
    .Y(_09040_));
 sg13g2_a21oi_1 _14899_ (.A1(\fpga_top.qspi_if.wrcmd1[0] ),
    .A2(net5685),
    .Y(_09041_),
    .B1(_09040_));
 sg13g2_mux2_1 _14900_ (.A0(_00108_),
    .A1(_00102_),
    .S(net5686),
    .X(_09042_));
 sg13g2_a221oi_1 _14901_ (.B2(net5349),
    .C1(_06948_),
    .B1(_09042_),
    .A1(net5345),
    .Y(_09043_),
    .A2(_09041_));
 sg13g2_nor4_1 _14902_ (.A(\fpga_top.qspi_if.cmd_ofs[0] ),
    .B(\fpga_top.qspi_if.cmd_ofs[1] ),
    .C(_09039_),
    .D(_09043_),
    .Y(_09044_));
 sg13g2_nor3_1 _14903_ (.A(\fpga_top.qspi_if.cmd_ofs[2] ),
    .B(_09034_),
    .C(_09044_),
    .Y(_09045_));
 sg13g2_nand2_1 _14904_ (.Y(_09046_),
    .A(_00106_),
    .B(_09001_));
 sg13g2_a21oi_1 _14905_ (.A1(_00112_),
    .A2(_09000_),
    .Y(_09047_),
    .B1(net5347));
 sg13g2_mux2_1 _14906_ (.A0(\fpga_top.qspi_if.wrcmd0[6] ),
    .A1(\fpga_top.qspi_if.wrcmd1[6] ),
    .S(net5074),
    .X(_09048_));
 sg13g2_a22oi_1 _14907_ (.Y(_09049_),
    .B1(_09048_),
    .B2(net5345),
    .A2(_09047_),
    .A1(_09046_));
 sg13g2_mux2_1 _14908_ (.A0(\fpga_top.qspi_if.wrcmd0[6] ),
    .A1(\fpga_top.qspi_if.wrcmd1[6] ),
    .S(net5684),
    .X(_09050_));
 sg13g2_nor2b_1 _14909_ (.A(net5688),
    .B_N(_00112_),
    .Y(_09051_));
 sg13g2_a21oi_1 _14910_ (.A1(_00106_),
    .A2(net5686),
    .Y(_09052_),
    .B1(_09051_));
 sg13g2_a22oi_1 _14911_ (.Y(_09053_),
    .B1(_09052_),
    .B2(net5349),
    .A2(_09050_),
    .A1(net5345));
 sg13g2_a21oi_1 _14912_ (.A1(\fpga_top.qspi_if.rdcmd1[7] ),
    .A2(net4949),
    .Y(_09054_),
    .B1(net5347));
 sg13g2_o21ai_1 _14913_ (.B1(_09054_),
    .Y(_09055_),
    .A1(_00113_),
    .A2(net4949));
 sg13g2_mux2_1 _14914_ (.A0(\fpga_top.qspi_if.wrcmd0[7] ),
    .A1(\fpga_top.qspi_if.wrcmd1[7] ),
    .S(net5074),
    .X(_09056_));
 sg13g2_o21ai_1 _14915_ (.B1(_09055_),
    .Y(_09057_),
    .A1(_06936_),
    .A2(_09056_));
 sg13g2_mux2_1 _14916_ (.A0(\fpga_top.qspi_if.wrcmd0[7] ),
    .A1(\fpga_top.qspi_if.wrcmd1[7] ),
    .S(net5684),
    .X(_09058_));
 sg13g2_a21oi_1 _14917_ (.A1(net5686),
    .A2(\fpga_top.qspi_if.rdcmd1[7] ),
    .Y(_09059_),
    .B1(net5347));
 sg13g2_o21ai_1 _14918_ (.B1(_09059_),
    .Y(_09060_),
    .A1(_00113_),
    .A2(net5686));
 sg13g2_o21ai_1 _14919_ (.B1(_09060_),
    .Y(_09061_),
    .A1(_06936_),
    .A2(_09058_));
 sg13g2_mux4_1 _14920_ (.S0(_00134_),
    .A0(_09049_),
    .A1(_09053_),
    .A2(_09057_),
    .A3(_09061_),
    .S1(\fpga_top.qspi_if.cmd_ofs[0] ),
    .X(_09062_));
 sg13g2_mux2_1 _14921_ (.A0(_00100_),
    .A1(_00097_),
    .S(net5074),
    .X(_09063_));
 sg13g2_nand2_1 _14922_ (.Y(_09064_),
    .A(\fpga_top.qspi_if.rdcmd0[4] ),
    .B(_09000_));
 sg13g2_a21oi_1 _14923_ (.A1(\fpga_top.qspi_if.rdcmd1[4] ),
    .A2(net4949),
    .Y(_09065_),
    .B1(net5348));
 sg13g2_a221oi_1 _14924_ (.B2(_09065_),
    .C1(_00134_),
    .B1(_09064_),
    .A1(net5347),
    .Y(_09066_),
    .A2(_09063_));
 sg13g2_mux2_1 _14925_ (.A0(_00100_),
    .A1(_00097_),
    .S(net5684),
    .X(_09067_));
 sg13g2_nand2b_1 _14926_ (.Y(_09068_),
    .B(\fpga_top.qspi_if.rdcmd0[4] ),
    .A_N(net5687));
 sg13g2_a21oi_1 _14927_ (.A1(net5687),
    .A2(\fpga_top.qspi_if.rdcmd1[4] ),
    .Y(_09069_),
    .B1(net5347));
 sg13g2_a22oi_1 _14928_ (.Y(_09070_),
    .B1(_09068_),
    .B2(_09069_),
    .A2(_09067_),
    .A1(net5347));
 sg13g2_a21o_1 _14929_ (.A2(_09070_),
    .A1(_00134_),
    .B1(_08919_),
    .X(_09071_));
 sg13g2_a21oi_1 _14930_ (.A1(_00105_),
    .A2(net4949),
    .Y(_09072_),
    .B1(net5347));
 sg13g2_o21ai_1 _14931_ (.B1(_09072_),
    .Y(_09073_),
    .A1(_06498_),
    .A2(net4949));
 sg13g2_mux2_1 _14932_ (.A0(_00101_),
    .A1(_00098_),
    .S(_09004_),
    .X(_09074_));
 sg13g2_o21ai_1 _14933_ (.B1(_09073_),
    .Y(_09075_),
    .A1(_06936_),
    .A2(_09074_));
 sg13g2_nor2b_1 _14934_ (.A(net5684),
    .B_N(_00101_),
    .Y(_09076_));
 sg13g2_a21oi_1 _14935_ (.A1(_00098_),
    .A2(net5684),
    .Y(_09077_),
    .B1(_09076_));
 sg13g2_nor2_1 _14936_ (.A(_06498_),
    .B(net5686),
    .Y(_09078_));
 sg13g2_a21oi_1 _14937_ (.A1(_00105_),
    .A2(net5686),
    .Y(_09079_),
    .B1(_09078_));
 sg13g2_a22oi_1 _14938_ (.Y(_09080_),
    .B1(_09079_),
    .B2(net5349),
    .A2(_09077_),
    .A1(net5345));
 sg13g2_a21oi_1 _14939_ (.A1(_06948_),
    .A2(_09075_),
    .Y(_09081_),
    .B1(_09028_));
 sg13g2_o21ai_1 _14940_ (.B1(_09081_),
    .Y(_09082_),
    .A1(_06948_),
    .A2(_09080_));
 sg13g2_o21ai_1 _14941_ (.B1(\fpga_top.qspi_if.cmd_ofs[2] ),
    .Y(_09083_),
    .A1(_09066_),
    .A2(_09071_));
 sg13g2_a21oi_1 _14942_ (.A1(\fpga_top.qspi_if.cmd_ofs[1] ),
    .A2(_09062_),
    .Y(_09084_),
    .B1(_09083_));
 sg13g2_nand2_1 _14943_ (.Y(_09085_),
    .A(net6570),
    .B(_08920_));
 sg13g2_nand2_1 _14944_ (.Y(_09086_),
    .A(\fpga_top.qspi_if.qspi_state[3] ),
    .B(_08867_));
 sg13g2_nor3_1 _14945_ (.A(net3978),
    .B(net5629),
    .C(net1375),
    .Y(_09087_));
 sg13g2_nand4_1 _14946_ (.B(_09085_),
    .C(_09086_),
    .A(_08863_),
    .Y(_09088_),
    .D(_09087_));
 sg13g2_nor2_1 _14947_ (.A(_06937_),
    .B(_08866_),
    .Y(_09089_));
 sg13g2_nor4_1 _14948_ (.A(net3762),
    .B(net3926),
    .C(_08923_),
    .D(_09089_),
    .Y(_09090_));
 sg13g2_a21oi_1 _14949_ (.A1(net6570),
    .A2(_08921_),
    .Y(_09091_),
    .B1(_00022_));
 sg13g2_nand4_1 _14950_ (.B(_08870_),
    .C(_09090_),
    .A(_08868_),
    .Y(_09092_),
    .D(_09091_));
 sg13g2_nor2b_1 _14951_ (.A(_09088_),
    .B_N(_09092_),
    .Y(_09093_));
 sg13g2_inv_1 _14952_ (.Y(_09094_),
    .A(_09093_));
 sg13g2_nor4_1 _14953_ (.A(net1534),
    .B(\fpga_top.qspi_if.qspi_state[2] ),
    .C(\fpga_top.qspi_if.dbg_2div_cew_pre ),
    .D(_08917_),
    .Y(_09095_));
 sg13g2_nand4_1 _14954_ (.B(_08856_),
    .C(_08929_),
    .A(_08728_),
    .Y(_09096_),
    .D(_09095_));
 sg13g2_nor3_1 _14955_ (.A(net3762),
    .B(\fpga_top.qspi_if.qspi_state[2] ),
    .C(_08917_),
    .Y(_09097_));
 sg13g2_o21ai_1 _14956_ (.B1(net6616),
    .Y(_09098_),
    .A1(\fpga_top.qspi_if.dbg_2div_read_half_end ),
    .A2(_08727_));
 sg13g2_nand3_1 _14957_ (.B(net3927),
    .C(_09098_),
    .A(_08867_),
    .Y(_09099_));
 sg13g2_nor2_1 _14958_ (.A(_09096_),
    .B(_09099_),
    .Y(_09100_));
 sg13g2_nand2_1 _14959_ (.Y(_09101_),
    .A(_09093_),
    .B(_09100_));
 sg13g2_nand2b_2 _14960_ (.Y(_09102_),
    .B(_09101_),
    .A_N(net3898));
 sg13g2_a22oi_1 _14961_ (.Y(_09103_),
    .B1(_09082_),
    .B2(_09084_),
    .A2(_09045_),
    .A1(_09022_));
 sg13g2_nor2b_2 _14962_ (.A(net5682),
    .B_N(\fpga_top.qspi_if.wdata_ofs[1] ),
    .Y(_09104_));
 sg13g2_and2_1 _14963_ (.A(net5682),
    .B(_08851_),
    .X(_09105_));
 sg13g2_nand2_1 _14964_ (.Y(_09106_),
    .A(net5683),
    .B(net6195));
 sg13g2_nand3_1 _14965_ (.B(net5683),
    .C(\fpga_top.qspi_if.wdata_ofs[1] ),
    .A(net5682),
    .Y(_09107_));
 sg13g2_a21oi_1 _14966_ (.A1(_06814_),
    .A2(_09107_),
    .Y(_09108_),
    .B1(_09105_));
 sg13g2_o21ai_1 _14967_ (.B1(_09108_),
    .Y(_09109_),
    .A1(\fpga_top.qspi_if.wdata[4] ),
    .A2(_09107_));
 sg13g2_nor2b_2 _14968_ (.A(\fpga_top.qspi_if.wdata_ofs[1] ),
    .B_N(net5683),
    .Y(_09110_));
 sg13g2_nand2_2 _14969_ (.Y(_09111_),
    .A(net5682),
    .B(_09110_));
 sg13g2_a22oi_1 _14970_ (.Y(_09112_),
    .B1(_09110_),
    .B2(net5682),
    .A2(_09105_),
    .A1(\fpga_top.qspi_if.wdata[8] ));
 sg13g2_o21ai_1 _14971_ (.B1(net5699),
    .Y(_09113_),
    .A1(\fpga_top.qspi_if.wdata[12] ),
    .A2(_09111_));
 sg13g2_a21oi_1 _14972_ (.A1(_09109_),
    .A2(_09112_),
    .Y(_09114_),
    .B1(_09113_));
 sg13g2_nor2_1 _14973_ (.A(_09104_),
    .B(_09114_),
    .Y(_09115_));
 sg13g2_nand2_2 _14974_ (.Y(_09116_),
    .A(net5683),
    .B(_09104_));
 sg13g2_nor2b_1 _14975_ (.A(net5701),
    .B_N(\fpga_top.qspi_if.word_hw ),
    .Y(_09117_));
 sg13g2_nand2_2 _14976_ (.Y(_09118_),
    .A(\fpga_top.qspi_if.word_hw ),
    .B(_06815_));
 sg13g2_a221oi_1 _14977_ (.B2(net5332),
    .C1(_09116_),
    .B1(\fpga_top.qspi_if.wdata[4] ),
    .A1(net5699),
    .Y(_09119_),
    .A2(\fpga_top.qspi_if.wdata[20] ));
 sg13g2_nand2b_2 _14978_ (.Y(_09120_),
    .B(_09104_),
    .A_N(\fpga_top.qspi_if.wdata_ofs[0] ));
 sg13g2_a221oi_1 _14979_ (.B2(\fpga_top.qspi_if.wdata[0] ),
    .C1(_09120_),
    .B1(net5332),
    .A1(net5699),
    .Y(_09121_),
    .A2(\fpga_top.qspi_if.wdata[16] ));
 sg13g2_nor4_1 _14980_ (.A(net5339),
    .B(_09115_),
    .C(_09119_),
    .D(_09121_),
    .Y(_09122_));
 sg13g2_nor2b_2 _14981_ (.A(\fpga_top.qspi_if.wdata_ofs[2] ),
    .B_N(_09110_),
    .Y(_09123_));
 sg13g2_o21ai_1 _14982_ (.B1(net5339),
    .Y(_09124_),
    .A1(\fpga_top.qspi_if.wdata[24] ),
    .A2(_06815_));
 sg13g2_nor2_1 _14983_ (.A(\fpga_top.qspi_if.word_hw ),
    .B(net5701),
    .Y(_09125_));
 sg13g2_or2_1 _14984_ (.X(_09126_),
    .B(net5700),
    .A(\fpga_top.qspi_if.word_hw ));
 sg13g2_nor2_1 _14985_ (.A(\fpga_top.qspi_if.wdata[0] ),
    .B(_09126_),
    .Y(_09127_));
 sg13g2_nor2_1 _14986_ (.A(\fpga_top.qspi_if.wdata[8] ),
    .B(_09118_),
    .Y(_09128_));
 sg13g2_nor3_1 _14987_ (.A(_09124_),
    .B(_09127_),
    .C(_09128_),
    .Y(_09129_));
 sg13g2_or3_1 _14988_ (.A(_09122_),
    .B(_09123_),
    .C(_09129_),
    .X(_09130_));
 sg13g2_nor2_1 _14989_ (.A(net4053),
    .B(_09126_),
    .Y(_09131_));
 sg13g2_nand2b_1 _14990_ (.Y(_09132_),
    .B(net5332),
    .A_N(net6551));
 sg13g2_o21ai_1 _14991_ (.B1(_09132_),
    .Y(_09133_),
    .A1(_06815_),
    .A2(net4070));
 sg13g2_o21ai_1 _14992_ (.B1(_09123_),
    .Y(_09134_),
    .A1(_09131_),
    .A2(_09133_));
 sg13g2_nand4_1 _14993_ (.B(net5377),
    .C(_09130_),
    .A(net5629),
    .Y(_09135_),
    .D(_09134_));
 sg13g2_and2_1 _14994_ (.A(net5680),
    .B(_08865_),
    .X(_09136_));
 sg13g2_nor2b_2 _14995_ (.A(net5680),
    .B_N(\fpga_top.qspi_if.adr_ofs[1] ),
    .Y(_09137_));
 sg13g2_nand2_2 _14996_ (.Y(_09138_),
    .A(net5681),
    .B(_09137_));
 sg13g2_nor2b_2 _14997_ (.A(\fpga_top.qspi_if.adr_ofs[1] ),
    .B_N(net5681),
    .Y(_09139_));
 sg13g2_nor2b_2 _14998_ (.A(net5680),
    .B_N(_09139_),
    .Y(_09140_));
 sg13g2_nand2b_1 _14999_ (.Y(_09141_),
    .B(_09139_),
    .A_N(net5680));
 sg13g2_o21ai_1 _15000_ (.B1(\fpga_top.qspi_if.adr_rw[0] ),
    .Y(_09142_),
    .A1(\fpga_top.qspi_if.adr_ofs[2] ),
    .A2(_08865_));
 sg13g2_nand2b_2 _15001_ (.Y(_09143_),
    .B(_09137_),
    .A_N(net5681));
 sg13g2_inv_1 _15002_ (.Y(_09144_),
    .A(_09143_));
 sg13g2_and2_1 _15003_ (.A(net5680),
    .B(_09139_),
    .X(_09145_));
 sg13g2_nand2_1 _15004_ (.Y(_09146_),
    .A(\fpga_top.qspi_if.adr_ofs[2] ),
    .B(_09139_));
 sg13g2_o21ai_1 _15005_ (.B1(_09142_),
    .Y(_09147_),
    .A1(_06816_),
    .A2(_09138_));
 sg13g2_a221oi_1 _15006_ (.B2(\fpga_top.qspi_if.adr_rw[8] ),
    .C1(_09147_),
    .B1(_09144_),
    .A1(\fpga_top.qspi_if.adr_rw[4] ),
    .Y(_09148_),
    .A2(_09140_));
 sg13g2_o21ai_1 _15007_ (.B1(_09146_),
    .Y(_09149_),
    .A1(_09136_),
    .A2(_09148_));
 sg13g2_a21oi_1 _15008_ (.A1(net6261),
    .A2(_09136_),
    .Y(_09150_),
    .B1(_09149_));
 sg13g2_o21ai_1 _15009_ (.B1(net6481),
    .Y(_09151_),
    .A1(net6397),
    .A2(_09146_));
 sg13g2_nor2_2 _15010_ (.A(_09150_),
    .B(_09151_),
    .Y(_09152_));
 sg13g2_nor2_1 _15011_ (.A(_09102_),
    .B(_09152_),
    .Y(_09153_));
 sg13g2_a22oi_1 _15012_ (.Y(\fpga_top.qspi_if.sio_out_pre[0] ),
    .B1(_09135_),
    .B2(_09153_),
    .A2(_09103_),
    .A1(_09102_));
 sg13g2_a21oi_1 _15013_ (.A1(_06820_),
    .A2(_09107_),
    .Y(_09154_),
    .B1(_09105_));
 sg13g2_o21ai_1 _15014_ (.B1(_09154_),
    .Y(_09155_),
    .A1(\fpga_top.qspi_if.wdata[5] ),
    .A2(_09107_));
 sg13g2_a22oi_1 _15015_ (.Y(_09156_),
    .B1(_09110_),
    .B2(\fpga_top.qspi_if.wdata_ofs[2] ),
    .A2(_09105_),
    .A1(\fpga_top.qspi_if.wdata[9] ));
 sg13g2_o21ai_1 _15016_ (.B1(net5699),
    .Y(_09157_),
    .A1(\fpga_top.qspi_if.wdata[13] ),
    .A2(_09111_));
 sg13g2_a21oi_1 _15017_ (.A1(_09155_),
    .A2(_09156_),
    .Y(_09158_),
    .B1(_09157_));
 sg13g2_a221oi_1 _15018_ (.B2(net5332),
    .C1(_09116_),
    .B1(\fpga_top.qspi_if.wdata[5] ),
    .A1(net5709),
    .Y(_09159_),
    .A2(\fpga_top.qspi_if.wdata[21] ));
 sg13g2_a221oi_1 _15019_ (.B2(\fpga_top.qspi_if.wdata[1] ),
    .C1(_09120_),
    .B1(net5332),
    .A1(net5699),
    .Y(_09160_),
    .A2(\fpga_top.qspi_if.wdata[17] ));
 sg13g2_nor3_1 _15020_ (.A(net5339),
    .B(_09159_),
    .C(_09160_),
    .Y(_09161_));
 sg13g2_o21ai_1 _15021_ (.B1(_09161_),
    .Y(_09162_),
    .A1(_09104_),
    .A2(_09158_));
 sg13g2_o21ai_1 _15022_ (.B1(net5339),
    .Y(_09163_),
    .A1(_06815_),
    .A2(\fpga_top.qspi_if.wdata[25] ));
 sg13g2_nor2_1 _15023_ (.A(\fpga_top.qspi_if.wdata[1] ),
    .B(_09126_),
    .Y(_09164_));
 sg13g2_nor2_1 _15024_ (.A(\fpga_top.qspi_if.wdata[9] ),
    .B(_09118_),
    .Y(_09165_));
 sg13g2_nor3_1 _15025_ (.A(_09163_),
    .B(_09164_),
    .C(_09165_),
    .Y(_09166_));
 sg13g2_nor2_1 _15026_ (.A(_09123_),
    .B(_09166_),
    .Y(_09167_));
 sg13g2_a22oi_1 _15027_ (.Y(_09168_),
    .B1(net5331),
    .B2(_06821_),
    .A2(_06822_),
    .A1(net5699));
 sg13g2_o21ai_1 _15028_ (.B1(_09168_),
    .Y(_09169_),
    .A1(net6235),
    .A2(_09118_));
 sg13g2_a22oi_1 _15029_ (.Y(_09170_),
    .B1(_09169_),
    .B2(_09123_),
    .A2(_09167_),
    .A1(_09162_));
 sg13g2_nand2_1 _15030_ (.Y(_09171_),
    .A(net6338),
    .B(_09170_));
 sg13g2_nor2_1 _15031_ (.A(\fpga_top.qspi_if.adr_rw[5] ),
    .B(_09141_),
    .Y(_09172_));
 sg13g2_o21ai_1 _15032_ (.B1(_09143_),
    .Y(_09173_),
    .A1(\fpga_top.qspi_if.adr_rw[1] ),
    .A2(_09140_));
 sg13g2_o21ai_1 _15033_ (.B1(_09137_),
    .Y(_09174_),
    .A1(net5681),
    .A2(\fpga_top.qspi_if.adr_rw[9] ));
 sg13g2_o21ai_1 _15034_ (.B1(_09174_),
    .Y(_09175_),
    .A1(_09172_),
    .A2(_09173_));
 sg13g2_nor2_1 _15035_ (.A(\fpga_top.qspi_if.adr_rw[13] ),
    .B(_09138_),
    .Y(_09176_));
 sg13g2_nor2_1 _15036_ (.A(_09136_),
    .B(_09176_),
    .Y(_09177_));
 sg13g2_a22oi_1 _15037_ (.Y(_09178_),
    .B1(_09175_),
    .B2(_09177_),
    .A2(_09136_),
    .A1(\fpga_top.qspi_if.adr_rw[17] ));
 sg13g2_or2_1 _15038_ (.X(_09179_),
    .B(_09178_),
    .A(_09145_));
 sg13g2_a21oi_1 _15039_ (.A1(\fpga_top.qspi_if.adr_rw[21] ),
    .A2(_09145_),
    .Y(_09180_),
    .B1(net5377));
 sg13g2_a221oi_1 _15040_ (.B2(_09180_),
    .C1(_09102_),
    .B1(_09179_),
    .A1(net5377),
    .Y(\fpga_top.qspi_if.sio_out_pre[1] ),
    .A2(_09171_));
 sg13g2_nand2b_1 _15041_ (.Y(_09181_),
    .B(_09107_),
    .A_N(\fpga_top.qspi_if.wdata[2] ));
 sg13g2_nor2_1 _15042_ (.A(\fpga_top.qspi_if.wdata[6] ),
    .B(_09107_),
    .Y(_09182_));
 sg13g2_nor2_1 _15043_ (.A(_09105_),
    .B(_09182_),
    .Y(_09183_));
 sg13g2_a22oi_1 _15044_ (.Y(_09184_),
    .B1(_09181_),
    .B2(_09183_),
    .A2(_09105_),
    .A1(\fpga_top.qspi_if.wdata[10] ));
 sg13g2_o21ai_1 _15045_ (.B1(net5700),
    .Y(_09185_),
    .A1(\fpga_top.qspi_if.wdata[14] ),
    .A2(_09111_));
 sg13g2_a21oi_1 _15046_ (.A1(_09111_),
    .A2(_09184_),
    .Y(_09186_),
    .B1(_09185_));
 sg13g2_a221oi_1 _15047_ (.B2(net5332),
    .C1(_09116_),
    .B1(\fpga_top.qspi_if.wdata[6] ),
    .A1(net5700),
    .Y(_09187_),
    .A2(\fpga_top.qspi_if.wdata[22] ));
 sg13g2_a221oi_1 _15048_ (.B2(\fpga_top.qspi_if.wdata[2] ),
    .C1(_09120_),
    .B1(net5332),
    .A1(net5700),
    .Y(_09188_),
    .A2(\fpga_top.qspi_if.wdata[18] ));
 sg13g2_nor3_1 _15049_ (.A(net5339),
    .B(_09187_),
    .C(_09188_),
    .Y(_09189_));
 sg13g2_o21ai_1 _15050_ (.B1(_09189_),
    .Y(_09190_),
    .A1(_09104_),
    .A2(_09186_));
 sg13g2_o21ai_1 _15051_ (.B1(net5339),
    .Y(_09191_),
    .A1(_06815_),
    .A2(\fpga_top.qspi_if.wdata[26] ));
 sg13g2_nor2_1 _15052_ (.A(\fpga_top.qspi_if.wdata[2] ),
    .B(_09126_),
    .Y(_09192_));
 sg13g2_nor2_1 _15053_ (.A(\fpga_top.qspi_if.wdata[10] ),
    .B(_09118_),
    .Y(_09193_));
 sg13g2_nor3_1 _15054_ (.A(_09191_),
    .B(_09192_),
    .C(_09193_),
    .Y(_09194_));
 sg13g2_nor2_1 _15055_ (.A(_09123_),
    .B(_09194_),
    .Y(_09195_));
 sg13g2_a22oi_1 _15056_ (.Y(_09196_),
    .B1(net5331),
    .B2(_06823_),
    .A2(_06824_),
    .A1(net5699));
 sg13g2_o21ai_1 _15057_ (.B1(_09196_),
    .Y(_09197_),
    .A1(\fpga_top.qspi_if.wdata[14] ),
    .A2(_09118_));
 sg13g2_a22oi_1 _15058_ (.Y(_09198_),
    .B1(_09197_),
    .B2(_09123_),
    .A2(_09195_),
    .A1(_09190_));
 sg13g2_nand2_1 _15059_ (.Y(_09199_),
    .A(net6338),
    .B(_09198_));
 sg13g2_nor2_1 _15060_ (.A(\fpga_top.qspi_if.adr_rw[6] ),
    .B(_09141_),
    .Y(_09200_));
 sg13g2_o21ai_1 _15061_ (.B1(_09143_),
    .Y(_09201_),
    .A1(\fpga_top.qspi_if.adr_rw[2] ),
    .A2(_09140_));
 sg13g2_o21ai_1 _15062_ (.B1(_09137_),
    .Y(_09202_),
    .A1(\fpga_top.qspi_if.adr_ofs[0] ),
    .A2(\fpga_top.qspi_if.adr_rw[10] ));
 sg13g2_o21ai_1 _15063_ (.B1(_09202_),
    .Y(_09203_),
    .A1(_09200_),
    .A2(_09201_));
 sg13g2_nor2_1 _15064_ (.A(\fpga_top.qspi_if.adr_rw[14] ),
    .B(_09138_),
    .Y(_09204_));
 sg13g2_nor2_1 _15065_ (.A(_09136_),
    .B(_09204_),
    .Y(_09205_));
 sg13g2_a22oi_1 _15066_ (.Y(_09206_),
    .B1(_09203_),
    .B2(_09205_),
    .A2(_09136_),
    .A1(net6436));
 sg13g2_or2_1 _15067_ (.X(_09207_),
    .B(_09206_),
    .A(_09145_));
 sg13g2_a21oi_1 _15068_ (.A1(net6485),
    .A2(_09145_),
    .Y(_09208_),
    .B1(net5377));
 sg13g2_a221oi_1 _15069_ (.B2(_09208_),
    .C1(_09102_),
    .B1(_09207_),
    .A1(net5377),
    .Y(\fpga_top.qspi_if.sio_out_pre[2] ),
    .A2(_09199_));
 sg13g2_nand2b_1 _15070_ (.Y(_09209_),
    .B(_09107_),
    .A_N(\fpga_top.qspi_if.wdata[3] ));
 sg13g2_nor2_1 _15071_ (.A(\fpga_top.qspi_if.wdata[7] ),
    .B(_09107_),
    .Y(_09210_));
 sg13g2_nor2_1 _15072_ (.A(_09105_),
    .B(_09210_),
    .Y(_09211_));
 sg13g2_a22oi_1 _15073_ (.Y(_09212_),
    .B1(_09209_),
    .B2(_09211_),
    .A2(_09105_),
    .A1(\fpga_top.qspi_if.wdata[11] ));
 sg13g2_o21ai_1 _15074_ (.B1(net5700),
    .Y(_09213_),
    .A1(\fpga_top.qspi_if.wdata[15] ),
    .A2(_09111_));
 sg13g2_a21oi_1 _15075_ (.A1(_09111_),
    .A2(_09212_),
    .Y(_09214_),
    .B1(_09213_));
 sg13g2_a221oi_1 _15076_ (.B2(net5335),
    .C1(_09116_),
    .B1(\fpga_top.qspi_if.wdata[7] ),
    .A1(net5700),
    .Y(_09215_),
    .A2(\fpga_top.qspi_if.wdata[23] ));
 sg13g2_a221oi_1 _15077_ (.B2(\fpga_top.qspi_if.wdata[3] ),
    .C1(_09120_),
    .B1(net5332),
    .A1(net5700),
    .Y(_09216_),
    .A2(\fpga_top.qspi_if.wdata[19] ));
 sg13g2_nor3_1 _15078_ (.A(net5339),
    .B(_09215_),
    .C(_09216_),
    .Y(_09217_));
 sg13g2_o21ai_1 _15079_ (.B1(_09217_),
    .Y(_09218_),
    .A1(_09104_),
    .A2(_09214_));
 sg13g2_o21ai_1 _15080_ (.B1(_08852_),
    .Y(_09219_),
    .A1(_06815_),
    .A2(\fpga_top.qspi_if.wdata[27] ));
 sg13g2_nor2_1 _15081_ (.A(\fpga_top.qspi_if.wdata[3] ),
    .B(_09126_),
    .Y(_09220_));
 sg13g2_nor2_1 _15082_ (.A(\fpga_top.qspi_if.wdata[11] ),
    .B(_09118_),
    .Y(_09221_));
 sg13g2_nor3_1 _15083_ (.A(_09219_),
    .B(_09220_),
    .C(_09221_),
    .Y(_09222_));
 sg13g2_nor2_1 _15084_ (.A(_09123_),
    .B(_09222_),
    .Y(_09223_));
 sg13g2_a22oi_1 _15085_ (.Y(_09224_),
    .B1(net5330),
    .B2(_06825_),
    .A2(_06826_),
    .A1(net5700));
 sg13g2_o21ai_1 _15086_ (.B1(_09224_),
    .Y(_09225_),
    .A1(\fpga_top.qspi_if.wdata[15] ),
    .A2(_09118_));
 sg13g2_a22oi_1 _15087_ (.Y(_09226_),
    .B1(_09225_),
    .B2(_09123_),
    .A2(_09223_),
    .A1(_09218_));
 sg13g2_nand2_1 _15088_ (.Y(_09227_),
    .A(net6338),
    .B(_09226_));
 sg13g2_nand2_1 _15089_ (.Y(_09228_),
    .A(net6448),
    .B(_09136_));
 sg13g2_nor2_1 _15090_ (.A(\fpga_top.qspi_if.adr_rw[3] ),
    .B(_09140_),
    .Y(_09229_));
 sg13g2_o21ai_1 _15091_ (.B1(_09143_),
    .Y(_09230_),
    .A1(\fpga_top.qspi_if.adr_rw[7] ),
    .A2(_09141_));
 sg13g2_o21ai_1 _15092_ (.B1(_09137_),
    .Y(_09231_),
    .A1(\fpga_top.qspi_if.adr_ofs[0] ),
    .A2(\fpga_top.qspi_if.adr_rw[11] ));
 sg13g2_o21ai_1 _15093_ (.B1(_09231_),
    .Y(_09232_),
    .A1(_09229_),
    .A2(_09230_));
 sg13g2_o21ai_1 _15094_ (.B1(_09232_),
    .Y(_09233_),
    .A1(\fpga_top.qspi_if.adr_rw[15] ),
    .A2(_09138_));
 sg13g2_o21ai_1 _15095_ (.B1(_09228_),
    .Y(_09234_),
    .A1(_09136_),
    .A2(_09233_));
 sg13g2_nand2_1 _15096_ (.Y(_09235_),
    .A(_09146_),
    .B(_09234_));
 sg13g2_a21oi_1 _15097_ (.A1(net6513),
    .A2(_09145_),
    .Y(_09236_),
    .B1(net5378));
 sg13g2_a221oi_1 _15098_ (.B2(_09236_),
    .C1(_09102_),
    .B1(_09235_),
    .A1(net5377),
    .Y(\fpga_top.qspi_if.sio_out_pre[3] ),
    .A2(_09227_));
 sg13g2_nand2b_1 _15099_ (.Y(_09237_),
    .B(\fpga_top.qspi_if.sck_cntr[2] ),
    .A_N(\fpga_top.qspi_if.sck_div[2] ));
 sg13g2_xnor2_1 _15100_ (.Y(_09238_),
    .A(net6594),
    .B(\fpga_top.qspi_if.sck_div[9] ));
 sg13g2_nand2b_1 _15101_ (.Y(_09239_),
    .B(\fpga_top.qspi_if.sck_div[7] ),
    .A_N(\fpga_top.qspi_if.sck_cntr[7] ));
 sg13g2_nand2b_1 _15102_ (.Y(_09240_),
    .B(\fpga_top.qspi_if.sck_cntr[4] ),
    .A_N(\fpga_top.qspi_if.sck_div[4] ));
 sg13g2_nand2b_1 _15103_ (.Y(_09241_),
    .B(\fpga_top.qspi_if.sck_cntr[8] ),
    .A_N(\fpga_top.qspi_if.sck_div[8] ));
 sg13g2_xnor2_1 _15104_ (.Y(_09242_),
    .A(\fpga_top.qspi_if.sck_cntr[1] ),
    .B(\fpga_top.qspi_if.sck_div[1] ));
 sg13g2_a22oi_1 _15105_ (.Y(_09243_),
    .B1(\fpga_top.qspi_if.sck_cntr[5] ),
    .B2(_06655_),
    .A2(\fpga_top.qspi_if.sck_div[3] ),
    .A1(_06652_));
 sg13g2_o21ai_1 _15106_ (.B1(_09239_),
    .Y(_09244_),
    .A1(\fpga_top.qspi_if.sck_cntr[5] ),
    .A2(_06655_));
 sg13g2_a22oi_1 _15107_ (.Y(_09245_),
    .B1(_06651_),
    .B2(\fpga_top.qspi_if.sck_div[2] ),
    .A2(\fpga_top.qspi_if.sck_cntr[0] ),
    .A1(_00114_));
 sg13g2_a22oi_1 _15108_ (.Y(_09246_),
    .B1(_06656_),
    .B2(\fpga_top.qspi_if.sck_div[6] ),
    .A2(_06653_),
    .A1(\fpga_top.qspi_if.sck_cntr[3] ));
 sg13g2_nand4_1 _15109_ (.B(_09241_),
    .C(_09242_),
    .A(_09237_),
    .Y(_09247_),
    .D(_09246_));
 sg13g2_a221oi_1 _15110_ (.B2(\fpga_top.qspi_if.sck_div[8] ),
    .C1(_09247_),
    .B1(_06659_),
    .A1(_06654_),
    .Y(_09248_),
    .A2(\fpga_top.qspi_if.sck_div[4] ));
 sg13g2_o21ai_1 _15111_ (.B1(_09240_),
    .Y(_09249_),
    .A1(_00114_),
    .A2(\fpga_top.qspi_if.sck_cntr[0] ));
 sg13g2_a22oi_1 _15112_ (.Y(_09250_),
    .B1(\fpga_top.qspi_if.sck_cntr[7] ),
    .B2(_06658_),
    .A2(_06657_),
    .A1(\fpga_top.qspi_if.sck_cntr[6] ));
 sg13g2_nand2_1 _15113_ (.Y(_09251_),
    .A(_09245_),
    .B(_09250_));
 sg13g2_nor3_1 _15114_ (.A(_09244_),
    .B(_09249_),
    .C(_09251_),
    .Y(_09252_));
 sg13g2_and4_1 _15115_ (.A(_09238_),
    .B(_09243_),
    .C(_09248_),
    .D(_09252_),
    .X(_09253_));
 sg13g2_nor2_1 _15116_ (.A(net1485),
    .B(net4947),
    .Y(_00042_));
 sg13g2_xnor2_1 _15117_ (.Y(_09254_),
    .A(net1485),
    .B(net3953));
 sg13g2_nor2_1 _15118_ (.A(net4947),
    .B(_09254_),
    .Y(_00043_));
 sg13g2_nand3_1 _15119_ (.B(net3953),
    .C(net6355),
    .A(net1485),
    .Y(_09255_));
 sg13g2_a21o_1 _15120_ (.A2(net3953),
    .A1(net1485),
    .B1(net6355),
    .X(_09256_));
 sg13g2_nand2_1 _15121_ (.Y(_09257_),
    .A(_09255_),
    .B(_09256_));
 sg13g2_nor2_1 _15122_ (.A(net4947),
    .B(_09257_),
    .Y(_00044_));
 sg13g2_nor2_1 _15123_ (.A(_06652_),
    .B(_09255_),
    .Y(_09258_));
 sg13g2_and2_1 _15124_ (.A(_06652_),
    .B(_09255_),
    .X(_09259_));
 sg13g2_nor3_1 _15125_ (.A(net4947),
    .B(_09258_),
    .C(_09259_),
    .Y(_00045_));
 sg13g2_and2_1 _15126_ (.A(net3776),
    .B(_09258_),
    .X(_09260_));
 sg13g2_nor2_1 _15127_ (.A(net3776),
    .B(_09258_),
    .Y(_09261_));
 sg13g2_nor3_1 _15128_ (.A(net4948),
    .B(_09260_),
    .C(net3777),
    .Y(_00046_));
 sg13g2_xnor2_1 _15129_ (.Y(_09262_),
    .A(net4000),
    .B(_09260_));
 sg13g2_nor2_1 _15130_ (.A(net4947),
    .B(_09262_),
    .Y(_00047_));
 sg13g2_a21oi_1 _15131_ (.A1(\fpga_top.qspi_if.sck_cntr[5] ),
    .A2(_09260_),
    .Y(_09263_),
    .B1(net2003));
 sg13g2_and3_1 _15132_ (.X(_09264_),
    .A(net6603),
    .B(net2003),
    .C(_09260_));
 sg13g2_nor3_1 _15133_ (.A(net4948),
    .B(net2004),
    .C(_09264_),
    .Y(_00048_));
 sg13g2_nor2_1 _15134_ (.A(net3859),
    .B(_09264_),
    .Y(_09265_));
 sg13g2_and2_1 _15135_ (.A(net3859),
    .B(_09264_),
    .X(_09266_));
 sg13g2_nor3_1 _15136_ (.A(net4947),
    .B(net3860),
    .C(_09266_),
    .Y(_00049_));
 sg13g2_nor2_1 _15137_ (.A(net3956),
    .B(_09266_),
    .Y(_09267_));
 sg13g2_and2_1 _15138_ (.A(net3956),
    .B(_09266_),
    .X(_09268_));
 sg13g2_nor3_1 _15139_ (.A(net4947),
    .B(net3957),
    .C(_09268_),
    .Y(_00050_));
 sg13g2_a21oi_1 _15140_ (.A1(net6205),
    .A2(_09268_),
    .Y(_09269_),
    .B1(net4947));
 sg13g2_o21ai_1 _15141_ (.B1(_09269_),
    .Y(_09270_),
    .A1(net6205),
    .A2(_09268_));
 sg13g2_inv_1 _15142_ (.Y(_00051_),
    .A(_09270_));
 sg13g2_nor3_1 _15143_ (.A(net3932),
    .B(net3783),
    .C(net6266),
    .Y(_09271_));
 sg13g2_nor2b_1 _15144_ (.A(\fpga_top.uart_top.uart_if.sample_cntr[3] ),
    .B_N(_09271_),
    .Y(_09272_));
 sg13g2_nor2b_1 _15145_ (.A(net4026),
    .B_N(_09272_),
    .Y(_09273_));
 sg13g2_nor2b_1 _15146_ (.A(\fpga_top.uart_top.uart_if.sample_cntr[5] ),
    .B_N(_09273_),
    .Y(_09274_));
 sg13g2_nor2b_2 _15147_ (.A(net6122),
    .B_N(_09274_),
    .Y(_09275_));
 sg13g2_nand2b_2 _15148_ (.Y(_09276_),
    .B(_09275_),
    .A_N(\fpga_top.uart_top.uart_if.sample_cntr[7] ));
 sg13g2_nor4_2 _15149_ (.A(\fpga_top.uart_top.uart_if.sample_cntr[11] ),
    .B(\fpga_top.uart_top.uart_if.sample_cntr[10] ),
    .C(\fpga_top.uart_top.uart_if.sample_cntr[9] ),
    .Y(_09277_),
    .D(\fpga_top.uart_top.uart_if.sample_cntr[8] ));
 sg13g2_nor3_1 _15150_ (.A(\fpga_top.uart_top.uart_if.sample_cntr[9] ),
    .B(net3994),
    .C(_09276_),
    .Y(_09278_));
 sg13g2_nand2b_1 _15151_ (.Y(_09279_),
    .B(_09278_),
    .A_N(\fpga_top.uart_top.uart_if.sample_cntr[10] ));
 sg13g2_nand2b_2 _15152_ (.Y(_09280_),
    .B(_09277_),
    .A_N(_09276_));
 sg13g2_nor3_1 _15153_ (.A(net6171),
    .B(\fpga_top.uart_top.uart_if.sample_cntr[12] ),
    .C(_09280_),
    .Y(_09281_));
 sg13g2_nand2b_1 _15154_ (.Y(_09282_),
    .B(_09281_),
    .A_N(\fpga_top.uart_top.uart_if.sample_cntr[14] ));
 sg13g2_nor2_1 _15155_ (.A(\fpga_top.uart_top.uart_if.sample_cntr[15] ),
    .B(_09282_),
    .Y(_09283_));
 sg13g2_nor2_1 _15156_ (.A(_06672_),
    .B(\fpga_top.uart_top.uart_if.rx_state[2] ),
    .Y(_09284_));
 sg13g2_inv_1 _15157_ (.Y(_09285_),
    .A(_09284_));
 sg13g2_nor2b_1 _15158_ (.A(net6188),
    .B_N(net1602),
    .Y(_09286_));
 sg13g2_and2_1 _15159_ (.A(_09284_),
    .B(_09286_),
    .X(_09287_));
 sg13g2_or4_1 _15160_ (.A(\fpga_top.uart_top.uart_if.sample_cntr[3] ),
    .B(\fpga_top.uart_top.uart_if.sample_cntr[2] ),
    .C(\fpga_top.uart_top.uart_if.sample_cntr[7] ),
    .D(\fpga_top.uart_top.uart_if.sample_cntr[6] ),
    .X(_09288_));
 sg13g2_nand2b_1 _15161_ (.Y(_09289_),
    .B(\fpga_top.uart_top.uart_if.sample_cntr[0] ),
    .A_N(\fpga_top.uart_top.uart_if.sample_cntr[1] ));
 sg13g2_nor4_1 _15162_ (.A(\fpga_top.uart_top.uart_if.sample_cntr[14] ),
    .B(\fpga_top.uart_top.uart_if.sample_cntr[13] ),
    .C(_09288_),
    .D(_09289_),
    .Y(_09290_));
 sg13g2_nor4_1 _15163_ (.A(\fpga_top.uart_top.uart_if.sample_cntr[5] ),
    .B(net6599),
    .C(\fpga_top.uart_top.uart_if.sample_cntr[15] ),
    .D(\fpga_top.uart_top.uart_if.sample_cntr[12] ),
    .Y(_09291_));
 sg13g2_nand3_1 _15164_ (.B(_09290_),
    .C(_09291_),
    .A(_09277_),
    .Y(_09292_));
 sg13g2_nor2_2 _15165_ (.A(_09287_),
    .B(_09292_),
    .Y(_09293_));
 sg13g2_or2_1 _15166_ (.X(_09294_),
    .B(_09292_),
    .A(_09287_));
 sg13g2_nor2_1 _15167_ (.A(_09283_),
    .B(net5072),
    .Y(_09295_));
 sg13g2_nand2b_1 _15168_ (.Y(_09296_),
    .B(net4690),
    .A_N(net3932));
 sg13g2_nor2_1 _15169_ (.A(net6350),
    .B(net3928),
    .Y(_09297_));
 sg13g2_nor2_1 _15170_ (.A(\fpga_top.uart_top.uart_if.rx_state[1] ),
    .B(\fpga_top.uart_top.uart_if.rx_state[0] ),
    .Y(_09298_));
 sg13g2_nand2_1 _15171_ (.Y(_09299_),
    .A(net1383),
    .B(_09298_));
 sg13g2_nor4_1 _15172_ (.A(\fpga_top.uart_top.uart_if.rx_state[3] ),
    .B(net3928),
    .C(net1394),
    .D(_09299_),
    .Y(_09300_));
 sg13g2_a21oi_1 _15173_ (.A1(net3838),
    .A2(net5070),
    .Y(_09301_),
    .B1(net5170));
 sg13g2_a22oi_1 _15174_ (.Y(_00052_),
    .B1(_09301_),
    .B2(_09296_),
    .A2(net5169),
    .A1(_06832_));
 sg13g2_xnor2_1 _15175_ (.Y(_09302_),
    .A(\fpga_top.uart_top.uart_if.sample_cntr[0] ),
    .B(net3783));
 sg13g2_a221oi_1 _15176_ (.B2(net3784),
    .C1(net5169),
    .B1(net4690),
    .A1(net1973),
    .Y(_09303_),
    .A2(net5071));
 sg13g2_a21oi_1 _15177_ (.A1(_06833_),
    .A2(net5169),
    .Y(_00059_),
    .B1(_09303_));
 sg13g2_o21ai_1 _15178_ (.B1(net6266),
    .Y(_09304_),
    .A1(net3932),
    .A2(net3783));
 sg13g2_nand2b_1 _15179_ (.Y(_09305_),
    .B(_09304_),
    .A_N(_09271_));
 sg13g2_a221oi_1 _15180_ (.B2(_09305_),
    .C1(net5171),
    .B1(net4690),
    .A1(net2123),
    .Y(_09306_),
    .A2(net5071));
 sg13g2_a21oi_1 _15181_ (.A1(_06834_),
    .A2(net5169),
    .Y(_00060_),
    .B1(_09306_));
 sg13g2_xor2_1 _15182_ (.B(_09271_),
    .A(\fpga_top.uart_top.uart_if.sample_cntr[3] ),
    .X(_09307_));
 sg13g2_a221oi_1 _15183_ (.B2(_09307_),
    .C1(net5171),
    .B1(net4690),
    .A1(net2113),
    .Y(_09308_),
    .A2(net5071));
 sg13g2_a21oi_1 _15184_ (.A1(_06835_),
    .A2(net5169),
    .Y(_00061_),
    .B1(_09308_));
 sg13g2_xor2_1 _15185_ (.B(_09272_),
    .A(net4026),
    .X(_09309_));
 sg13g2_a221oi_1 _15186_ (.B2(net4027),
    .C1(net5172),
    .B1(net4691),
    .A1(net3973),
    .Y(_09310_),
    .A2(net5072));
 sg13g2_a21oi_1 _15187_ (.A1(_06836_),
    .A2(net5169),
    .Y(_00062_),
    .B1(_09310_));
 sg13g2_xor2_1 _15188_ (.B(_09273_),
    .A(net6216),
    .X(_09311_));
 sg13g2_a221oi_1 _15189_ (.B2(_09311_),
    .C1(net5169),
    .B1(net4690),
    .A1(net2373),
    .Y(_09312_),
    .A2(net5072));
 sg13g2_a21oi_1 _15190_ (.A1(_06837_),
    .A2(net5169),
    .Y(_00063_),
    .B1(_09312_));
 sg13g2_xor2_1 _15191_ (.B(_09274_),
    .A(net6122),
    .X(_09313_));
 sg13g2_a221oi_1 _15192_ (.B2(net6123),
    .C1(net5170),
    .B1(net4690),
    .A1(net3142),
    .Y(_09314_),
    .A2(net5072));
 sg13g2_a21oi_1 _15193_ (.A1(_06838_),
    .A2(net5172),
    .Y(_00064_),
    .B1(_09314_));
 sg13g2_xor2_1 _15194_ (.B(_09275_),
    .A(net6241),
    .X(_09315_));
 sg13g2_a221oi_1 _15195_ (.B2(_09315_),
    .C1(net5170),
    .B1(net4690),
    .A1(net3606),
    .Y(_09316_),
    .A2(net5071));
 sg13g2_a21oi_1 _15196_ (.A1(_06839_),
    .A2(net5170),
    .Y(_00065_),
    .B1(_09316_));
 sg13g2_xnor2_1 _15197_ (.Y(_09317_),
    .A(net3994),
    .B(_09276_));
 sg13g2_a221oi_1 _15198_ (.B2(net3995),
    .C1(net5173),
    .B1(net4691),
    .A1(net3965),
    .Y(_09318_),
    .A2(net5073));
 sg13g2_a21oi_1 _15199_ (.A1(_06840_),
    .A2(net5173),
    .Y(_00066_),
    .B1(net3996));
 sg13g2_o21ai_1 _15200_ (.B1(net6299),
    .Y(_09319_),
    .A1(net3994),
    .A2(_09276_));
 sg13g2_nand2b_1 _15201_ (.Y(_09320_),
    .B(_09319_),
    .A_N(_09278_));
 sg13g2_a221oi_1 _15202_ (.B2(net6300),
    .C1(net5171),
    .B1(net4691),
    .A1(net3305),
    .Y(_09321_),
    .A2(net5073));
 sg13g2_a21oi_1 _15203_ (.A1(_06841_),
    .A2(net5171),
    .Y(_00067_),
    .B1(_09321_));
 sg13g2_xor2_1 _15204_ (.B(_09278_),
    .A(net6206),
    .X(_09322_));
 sg13g2_a221oi_1 _15205_ (.B2(net6207),
    .C1(net5173),
    .B1(net4691),
    .A1(net3988),
    .Y(_09323_),
    .A2(net5073));
 sg13g2_a21oi_1 _15206_ (.A1(_06842_),
    .A2(net5173),
    .Y(_00053_),
    .B1(net6208));
 sg13g2_xnor2_1 _15207_ (.Y(_09324_),
    .A(\fpga_top.uart_top.uart_if.sample_cntr[11] ),
    .B(_09279_));
 sg13g2_a221oi_1 _15208_ (.B2(_09324_),
    .C1(net5173),
    .B1(net4691),
    .A1(net6174),
    .Y(_09325_),
    .A2(net5073));
 sg13g2_a21oi_1 _15209_ (.A1(_06843_),
    .A2(net5173),
    .Y(_00054_),
    .B1(net6175));
 sg13g2_xnor2_1 _15210_ (.Y(_09326_),
    .A(net6357),
    .B(_09280_));
 sg13g2_a221oi_1 _15211_ (.B2(net6358),
    .C1(net5171),
    .B1(net4691),
    .A1(net4022),
    .Y(_09327_),
    .A2(net5072));
 sg13g2_a21oi_1 _15212_ (.A1(_06844_),
    .A2(net5171),
    .Y(_00055_),
    .B1(_09327_));
 sg13g2_o21ai_1 _15213_ (.B1(net6171),
    .Y(_09328_),
    .A1(\fpga_top.uart_top.uart_if.sample_cntr[12] ),
    .A2(_09280_));
 sg13g2_nand2b_1 _15214_ (.Y(_09329_),
    .B(net6172),
    .A_N(_09281_));
 sg13g2_a221oi_1 _15215_ (.B2(net6173),
    .C1(net5171),
    .B1(net4691),
    .A1(net4043),
    .Y(_09330_),
    .A2(net5072));
 sg13g2_a21oi_1 _15216_ (.A1(_06845_),
    .A2(net5172),
    .Y(_00056_),
    .B1(_09330_));
 sg13g2_xor2_1 _15217_ (.B(_09281_),
    .A(\fpga_top.uart_top.uart_if.sample_cntr[14] ),
    .X(_09331_));
 sg13g2_a221oi_1 _15218_ (.B2(_09331_),
    .C1(net5170),
    .B1(net4690),
    .A1(net6111),
    .Y(_09332_),
    .A2(net5072));
 sg13g2_a21oi_1 _15219_ (.A1(_06846_),
    .A2(net5170),
    .Y(_00057_),
    .B1(_09332_));
 sg13g2_a22oi_1 _15220_ (.Y(_09333_),
    .B1(net5072),
    .B2(\fpga_top.io_uart_out.uart_term[15] ),
    .A2(_09282_),
    .A1(net3867));
 sg13g2_nor2_1 _15221_ (.A(net5170),
    .B(net3868),
    .Y(_00058_));
 sg13g2_nor4_1 _15222_ (.A(net3855),
    .B(net1536),
    .C(net3386),
    .D(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[3] ),
    .Y(_09334_));
 sg13g2_nor3_1 _15223_ (.A(net3730),
    .B(net3664),
    .C(_09334_),
    .Y(_09335_));
 sg13g2_or3_1 _15224_ (.A(net3730),
    .B(net3664),
    .C(_09334_),
    .X(_09336_));
 sg13g2_nor4_1 _15225_ (.A(\fpga_top.uart_top.uart_if.tx_out_cntr[0] ),
    .B(\fpga_top.uart_top.uart_if.tx_out_cntr[1] ),
    .C(\fpga_top.uart_top.uart_if.tx_out_cntr[3] ),
    .D(\fpga_top.uart_top.uart_if.tx_out_cntr[2] ),
    .Y(_09337_));
 sg13g2_nor4_1 _15226_ (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[3] ),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[2] ),
    .C(\fpga_top.uart_top.uart_if.tx_cycle_cntr[7] ),
    .D(net4010),
    .Y(_09338_));
 sg13g2_nor2_1 _15227_ (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[6] ),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[5] ),
    .Y(_09339_));
 sg13g2_nand4_1 _15228_ (.B(_06673_),
    .C(_09338_),
    .A(net1902),
    .Y(_09340_),
    .D(_09339_));
 sg13g2_nor4_1 _15229_ (.A(net6166),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[10] ),
    .C(\fpga_top.uart_top.uart_if.tx_cycle_cntr[9] ),
    .D(\fpga_top.uart_top.uart_if.tx_cycle_cntr[8] ),
    .Y(_09341_));
 sg13g2_nor4_1 _15230_ (.A(net1934),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[14] ),
    .C(\fpga_top.uart_top.uart_if.tx_cycle_cntr[13] ),
    .D(\fpga_top.uart_top.uart_if.tx_cycle_cntr[12] ),
    .Y(_09342_));
 sg13g2_nand2_1 _15231_ (.Y(_09343_),
    .A(_09341_),
    .B(_09342_));
 sg13g2_nor4_1 _15232_ (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[7] ),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[6] ),
    .C(\fpga_top.uart_top.uart_if.tx_cycle_cntr[5] ),
    .D(net4010),
    .Y(_09344_));
 sg13g2_nand3b_1 _15233_ (.B(_09341_),
    .C(_09342_),
    .Y(_09345_),
    .A_N(_09340_));
 sg13g2_or2_1 _15234_ (.X(_09346_),
    .B(_09345_),
    .A(_09337_));
 sg13g2_and2_1 _15235_ (.A(net5282),
    .B(_09346_),
    .X(_09347_));
 sg13g2_nand2_1 _15236_ (.Y(_09348_),
    .A(net5282),
    .B(_09346_));
 sg13g2_nor3_1 _15237_ (.A(net1902),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[1] ),
    .C(\fpga_top.uart_top.uart_if.tx_cycle_cntr[2] ),
    .Y(_09349_));
 sg13g2_nor2b_2 _15238_ (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[3] ),
    .B_N(_09349_),
    .Y(_09350_));
 sg13g2_nand2b_2 _15239_ (.Y(_09351_),
    .B(_09350_),
    .A_N(\fpga_top.uart_top.uart_if.tx_cycle_cntr[4] ));
 sg13g2_nor3_1 _15240_ (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[6] ),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[5] ),
    .C(_09351_),
    .Y(_09352_));
 sg13g2_nand2_2 _15241_ (.Y(_09353_),
    .A(_09344_),
    .B(_09350_));
 sg13g2_nor3_1 _15242_ (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[9] ),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[8] ),
    .C(_09353_),
    .Y(_09354_));
 sg13g2_nor2b_1 _15243_ (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[10] ),
    .B_N(_09354_),
    .Y(_09355_));
 sg13g2_nand3_1 _15244_ (.B(_09344_),
    .C(_09350_),
    .A(_09341_),
    .Y(_09356_));
 sg13g2_o21ai_1 _15245_ (.B1(_09347_),
    .Y(_09357_),
    .A1(_09343_),
    .A2(_09353_));
 sg13g2_nand2_1 _15246_ (.Y(_09358_),
    .A(\fpga_top.io_uart_out.uart_term[0] ),
    .B(net4944));
 sg13g2_o21ai_1 _15247_ (.B1(_09358_),
    .Y(_00068_),
    .A1(net1902),
    .A2(net4847));
 sg13g2_nand2_1 _15248_ (.Y(_09359_),
    .A(net1973),
    .B(net4942));
 sg13g2_xor2_1 _15249_ (.B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[1] ),
    .A(net1902),
    .X(_09360_));
 sg13g2_o21ai_1 _15250_ (.B1(_09359_),
    .Y(_00075_),
    .A1(net4847),
    .A2(_09360_));
 sg13g2_o21ai_1 _15251_ (.B1(\fpga_top.uart_top.uart_if.tx_cycle_cntr[2] ),
    .Y(_09361_),
    .A1(net1902),
    .A2(\fpga_top.uart_top.uart_if.tx_cycle_cntr[1] ));
 sg13g2_nor2b_1 _15252_ (.A(_09349_),
    .B_N(_09361_),
    .Y(_09362_));
 sg13g2_nand2_1 _15253_ (.Y(_09363_),
    .A(net2123),
    .B(net4942));
 sg13g2_o21ai_1 _15254_ (.B1(_09363_),
    .Y(_00076_),
    .A1(net4847),
    .A2(_09362_));
 sg13g2_xnor2_1 _15255_ (.Y(_09364_),
    .A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[3] ),
    .B(_09349_));
 sg13g2_nand2_1 _15256_ (.Y(_09365_),
    .A(net2113),
    .B(net4943));
 sg13g2_o21ai_1 _15257_ (.B1(_09365_),
    .Y(_00077_),
    .A1(net4847),
    .A2(_09364_));
 sg13g2_xnor2_1 _15258_ (.Y(_09366_),
    .A(net4010),
    .B(_09350_));
 sg13g2_nand2_1 _15259_ (.Y(_09367_),
    .A(net3973),
    .B(net4943));
 sg13g2_o21ai_1 _15260_ (.B1(_09367_),
    .Y(_00078_),
    .A1(net4848),
    .A2(net4011));
 sg13g2_xor2_1 _15261_ (.B(_09351_),
    .A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[5] ),
    .X(_09368_));
 sg13g2_nand2_1 _15262_ (.Y(_09369_),
    .A(net2373),
    .B(net4943));
 sg13g2_o21ai_1 _15263_ (.B1(_09369_),
    .Y(_00079_),
    .A1(net4848),
    .A2(_09368_));
 sg13g2_o21ai_1 _15264_ (.B1(\fpga_top.uart_top.uart_if.tx_cycle_cntr[6] ),
    .Y(_09370_),
    .A1(\fpga_top.uart_top.uart_if.tx_cycle_cntr[5] ),
    .A2(_09351_));
 sg13g2_nor2b_1 _15265_ (.A(_09352_),
    .B_N(_09370_),
    .Y(_09371_));
 sg13g2_nand2_1 _15266_ (.Y(_09372_),
    .A(net3142),
    .B(net4943));
 sg13g2_o21ai_1 _15267_ (.B1(_09372_),
    .Y(_00080_),
    .A1(net4848),
    .A2(_09371_));
 sg13g2_xnor2_1 _15268_ (.Y(_09373_),
    .A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[7] ),
    .B(_09352_));
 sg13g2_nand2_1 _15269_ (.Y(_09374_),
    .A(net3606),
    .B(net4943));
 sg13g2_o21ai_1 _15270_ (.B1(_09374_),
    .Y(_00081_),
    .A1(net4848),
    .A2(_09373_));
 sg13g2_xor2_1 _15271_ (.B(_09353_),
    .A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[8] ),
    .X(_09375_));
 sg13g2_nand2_1 _15272_ (.Y(_09376_),
    .A(net3965),
    .B(net4942));
 sg13g2_o21ai_1 _15273_ (.B1(_09376_),
    .Y(_00082_),
    .A1(net4847),
    .A2(_09375_));
 sg13g2_o21ai_1 _15274_ (.B1(\fpga_top.uart_top.uart_if.tx_cycle_cntr[9] ),
    .Y(_09377_),
    .A1(\fpga_top.uart_top.uart_if.tx_cycle_cntr[8] ),
    .A2(_09353_));
 sg13g2_nor2b_1 _15275_ (.A(_09354_),
    .B_N(_09377_),
    .Y(_09378_));
 sg13g2_nand2_1 _15276_ (.Y(_09379_),
    .A(net3305),
    .B(net4944));
 sg13g2_o21ai_1 _15277_ (.B1(_09379_),
    .Y(_00083_),
    .A1(net4847),
    .A2(_09378_));
 sg13g2_xnor2_1 _15278_ (.Y(_09380_),
    .A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[10] ),
    .B(_09354_));
 sg13g2_nand2_1 _15279_ (.Y(_09381_),
    .A(net3988),
    .B(net4944));
 sg13g2_o21ai_1 _15280_ (.B1(_09381_),
    .Y(_00069_),
    .A1(net4847),
    .A2(_09380_));
 sg13g2_xnor2_1 _15281_ (.Y(_09382_),
    .A(net6166),
    .B(_09355_));
 sg13g2_nand2_1 _15282_ (.Y(_09383_),
    .A(\fpga_top.io_uart_out.uart_term[11] ),
    .B(net4944));
 sg13g2_o21ai_1 _15283_ (.B1(_09383_),
    .Y(_00070_),
    .A1(net4847),
    .A2(net6167));
 sg13g2_xor2_1 _15284_ (.B(_09356_),
    .A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[12] ),
    .X(_09384_));
 sg13g2_nand2_1 _15285_ (.Y(_09385_),
    .A(net4022),
    .B(net4942));
 sg13g2_o21ai_1 _15286_ (.B1(_09385_),
    .Y(_00071_),
    .A1(net4848),
    .A2(_09384_));
 sg13g2_nor3_1 _15287_ (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[13] ),
    .B(\fpga_top.uart_top.uart_if.tx_cycle_cntr[12] ),
    .C(_09356_),
    .Y(_09386_));
 sg13g2_o21ai_1 _15288_ (.B1(\fpga_top.uart_top.uart_if.tx_cycle_cntr[13] ),
    .Y(_09387_),
    .A1(\fpga_top.uart_top.uart_if.tx_cycle_cntr[12] ),
    .A2(_09356_));
 sg13g2_nor2b_1 _15289_ (.A(_09386_),
    .B_N(_09387_),
    .Y(_09388_));
 sg13g2_nand2_1 _15290_ (.Y(_09389_),
    .A(net4043),
    .B(net4942));
 sg13g2_o21ai_1 _15291_ (.B1(_09389_),
    .Y(_00072_),
    .A1(net4848),
    .A2(_09388_));
 sg13g2_nand2b_1 _15292_ (.Y(_09390_),
    .B(_09386_),
    .A_N(\fpga_top.uart_top.uart_if.tx_cycle_cntr[14] ));
 sg13g2_xnor2_1 _15293_ (.Y(_09391_),
    .A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[14] ),
    .B(_09386_));
 sg13g2_nand2_1 _15294_ (.Y(_09392_),
    .A(net6111),
    .B(net4942));
 sg13g2_o21ai_1 _15295_ (.B1(_09392_),
    .Y(_00073_),
    .A1(net4848),
    .A2(_09391_));
 sg13g2_a21oi_1 _15296_ (.A1(net1934),
    .A2(_09390_),
    .Y(_09393_),
    .B1(net4942));
 sg13g2_a21oi_1 _15297_ (.A1(_06846_),
    .A2(net4942),
    .Y(_00074_),
    .B1(net1935));
 sg13g2_nor3_1 _15298_ (.A(net6219),
    .B(net6346),
    .C(_06680_),
    .Y(_09394_));
 sg13g2_nand2b_1 _15299_ (.Y(_09395_),
    .B(net5572),
    .A_N(net5280));
 sg13g2_nor2_2 _15300_ (.A(\fpga_top.bus_gather.u_read_adr[31] ),
    .B(net6608),
    .Y(_09396_));
 sg13g2_and2_1 _15301_ (.A(net5285),
    .B(_09396_),
    .X(_09397_));
 sg13g2_a21oi_1 _15302_ (.A1(\fpga_top.cpu_top.csr_uimm[0] ),
    .A2(net5280),
    .Y(_09398_),
    .B1(_09397_));
 sg13g2_a22oi_1 _15303_ (.Y(\fpga_top.cpu_top.register_file.inst_rs[8] ),
    .B1(_09398_),
    .B2(_09395_),
    .A2(_09397_),
    .A1(_06504_));
 sg13g2_nor2_1 _15304_ (.A(_06559_),
    .B(net5281),
    .Y(_09399_));
 sg13g2_a221oi_1 _15305_ (.B2(net5285),
    .C1(_09399_),
    .B1(_09396_),
    .A1(net6093),
    .Y(_09400_),
    .A2(net5280));
 sg13g2_a21oi_1 _15306_ (.A1(_06505_),
    .A2(_09397_),
    .Y(\fpga_top.cpu_top.register_file.inst_rs[7] ),
    .B1(_09400_));
 sg13g2_nor2_1 _15307_ (.A(_06548_),
    .B(net5280),
    .Y(_09401_));
 sg13g2_a221oi_1 _15308_ (.B2(net5285),
    .C1(_09401_),
    .B1(_09396_),
    .A1(net6211),
    .Y(_09402_),
    .A2(net5280));
 sg13g2_a21oi_2 _15309_ (.B1(_09402_),
    .Y(\fpga_top.cpu_top.register_file.inst_rs[6] ),
    .A2(_09397_),
    .A1(_06508_));
 sg13g2_nor2_1 _15310_ (.A(_06568_),
    .B(net5280),
    .Y(_09403_));
 sg13g2_a221oi_1 _15311_ (.B2(net5285),
    .C1(_09403_),
    .B1(_09396_),
    .A1(net6455),
    .Y(_09404_),
    .A2(net5281));
 sg13g2_a21oi_2 _15312_ (.B1(_09404_),
    .Y(\fpga_top.cpu_top.register_file.inst_rs[5] ),
    .A2(_09397_),
    .A1(_06507_));
 sg13g2_nor2_1 _15313_ (.A(_06575_),
    .B(net5280),
    .Y(_09405_));
 sg13g2_a221oi_1 _15314_ (.B2(\fpga_top.uart_top.uart_logics.radr_enable ),
    .C1(_09405_),
    .B1(_09396_),
    .A1(net6375),
    .Y(_09406_),
    .A2(net5280));
 sg13g2_a21oi_2 _15315_ (.B1(_09406_),
    .Y(\fpga_top.cpu_top.register_file.inst_rs[4] ),
    .A2(_09397_),
    .A1(_06514_));
 sg13g2_nand2_1 _15316_ (.Y(_09407_),
    .A(net6192),
    .B(net3827));
 sg13g2_nand2_1 _15317_ (.Y(_09408_),
    .A(\fpga_top.io_spi_lite.cs_all_status ),
    .B(_09407_));
 sg13g2_nor2b_2 _15318_ (.A(net6192),
    .B_N(net3827),
    .Y(_09409_));
 sg13g2_nand2b_2 _15319_ (.Y(_09410_),
    .B(net3827),
    .A_N(\fpga_top.io_spi_lite.spi_state[0] ));
 sg13g2_or3_1 _15320_ (.A(net1756),
    .B(net1681),
    .C(net1580),
    .X(_09411_));
 sg13g2_nand4_1 _15321_ (.B(net1975),
    .C(net1703),
    .A(net3201),
    .Y(_09412_),
    .D(net1915));
 sg13g2_or4_1 _15322_ (.A(_08972_),
    .B(_09410_),
    .C(_09411_),
    .D(_09412_),
    .X(_09413_));
 sg13g2_nand2b_1 _15323_ (.Y(_09414_),
    .B(_09413_),
    .A_N(_09408_));
 sg13g2_nor2_1 _15324_ (.A(net3827),
    .B(_06648_),
    .Y(_09415_));
 sg13g2_mux2_1 _15325_ (.A0(net1369),
    .A1(_09415_),
    .S(_09414_),
    .X(\fpga_top.io_spi_lite.org_spi_sck ));
 sg13g2_a21oi_1 _15326_ (.A1(net5826),
    .A2(_06926_),
    .Y(_09416_),
    .B1(\fpga_top.io_spi_lite.spi_mode[8] ));
 sg13g2_o21ai_1 _15327_ (.B1(_09416_),
    .Y(_09417_),
    .A1(net5826),
    .A2(\fpga_top.io_spi_lite.org_spi_sck ));
 sg13g2_o21ai_1 _15328_ (.B1(\fpga_top.io_spi_lite.spi_mode[8] ),
    .Y(_09418_),
    .A1(net5826),
    .A2(\fpga_top.io_spi_lite.sel_sck[2] ));
 sg13g2_a21oi_1 _15329_ (.A1(net5826),
    .A2(_06927_),
    .Y(_09419_),
    .B1(_09418_));
 sg13g2_nor2_1 _15330_ (.A(\fpga_top.io_spi_lite.spi_mode[9] ),
    .B(_09419_),
    .Y(_09420_));
 sg13g2_nor2b_1 _15331_ (.A(\fpga_top.io_spi_lite.sel_sck[5] ),
    .B_N(net5826),
    .Y(_09421_));
 sg13g2_nor2_1 _15332_ (.A(net5826),
    .B(\fpga_top.io_spi_lite.sel_sck[4] ),
    .Y(_09422_));
 sg13g2_nor3_1 _15333_ (.A(\fpga_top.io_spi_lite.spi_mode[8] ),
    .B(_09421_),
    .C(_09422_),
    .Y(_09423_));
 sg13g2_nor2b_1 _15334_ (.A(\fpga_top.io_spi_lite.sel_sck[7] ),
    .B_N(net5826),
    .Y(_09424_));
 sg13g2_o21ai_1 _15335_ (.B1(\fpga_top.io_spi_lite.spi_mode[8] ),
    .Y(_09425_),
    .A1(\fpga_top.io_spi_lite.spi_mode[7] ),
    .A2(\fpga_top.io_spi_lite.sel_sck[6] ));
 sg13g2_o21ai_1 _15336_ (.B1(\fpga_top.io_spi_lite.spi_mode[9] ),
    .Y(_09426_),
    .A1(_09424_),
    .A2(_09425_));
 sg13g2_o21ai_1 _15337_ (.B1(\fpga_top.io_spi_lite.spi_mode[0] ),
    .Y(_09427_),
    .A1(_09423_),
    .A2(_09426_));
 sg13g2_a21oi_2 _15338_ (.B1(_09427_),
    .Y(_09428_),
    .A2(_09420_),
    .A1(_09417_));
 sg13g2_a21o_2 _15339_ (.A2(_06875_),
    .A1(\fpga_top.io_led.led_value[0] ),
    .B1(_09428_),
    .X(uo_out[5]));
 sg13g2_mux4_1 _15340_ (.S0(\fpga_top.io_spi_lite.spi_mode[5] ),
    .A0(\fpga_top.io_spi_lite.cs_all_status ),
    .A1(\fpga_top.io_spi_lite.sel_cs[2] ),
    .A2(\fpga_top.io_spi_lite.sel_cs[1] ),
    .A3(\fpga_top.io_spi_lite.sel_cs[3] ),
    .S1(\fpga_top.io_spi_lite.spi_mode[4] ),
    .X(_09429_));
 sg13g2_nand2_1 _15341_ (.Y(_09430_),
    .A(_06913_),
    .B(_09429_));
 sg13g2_mux4_1 _15342_ (.S0(\fpga_top.io_spi_lite.spi_mode[4] ),
    .A0(\fpga_top.io_spi_lite.sel_cs[4] ),
    .A1(\fpga_top.io_spi_lite.sel_cs[5] ),
    .A2(\fpga_top.io_spi_lite.sel_cs[6] ),
    .A3(\fpga_top.io_spi_lite.sel_cs[7] ),
    .S1(\fpga_top.io_spi_lite.spi_mode[5] ),
    .X(_09431_));
 sg13g2_a21oi_1 _15343_ (.A1(\fpga_top.io_spi_lite.spi_mode[6] ),
    .A2(_09431_),
    .Y(_09432_),
    .B1(_06875_));
 sg13g2_nor2b_1 _15344_ (.A(\fpga_top.io_spi_lite.spi_mode[0] ),
    .B_N(\fpga_top.io_led.led_value[1] ),
    .Y(_09433_));
 sg13g2_a21o_2 _15345_ (.A2(_09432_),
    .A1(_09430_),
    .B1(_09433_),
    .X(uo_out[6]));
 sg13g2_nor3_1 _15346_ (.A(\fpga_top.dbg_bpoint_en[2] ),
    .B(\fpga_top.dbg_bpoint_en[1] ),
    .C(\fpga_top.dbg_bpoint_en[0] ),
    .Y(_09434_));
 sg13g2_mux2_1 _15347_ (.A0(\fpga_top.io_led.dbg_smpl_trgsig ),
    .A1(\fpga_top.io_led.led_value[2] ),
    .S(_09434_),
    .X(_09435_));
 sg13g2_mux2_1 _15348_ (.A0(\fpga_top.io_spi_lite.spi_mosi ),
    .A1(_09435_),
    .S(_06875_),
    .X(uo_out[7]));
 sg13g2_nor2b_2 _15349_ (.A(net6343),
    .B_N(\fpga_top.cpu_top.register_file.rfr_state[1] ),
    .Y(_09436_));
 sg13g2_and2_1 _15350_ (.A(_06680_),
    .B(_09436_),
    .X(_09437_));
 sg13g2_nor2b_1 _15351_ (.A(net6307),
    .B_N(net6496),
    .Y(_09438_));
 sg13g2_nand2b_2 _15352_ (.Y(_09439_),
    .B(net6496),
    .A_N(net6533));
 sg13g2_nand3_1 _15353_ (.B(net6514),
    .C(_09438_),
    .A(net5426),
    .Y(_09440_));
 sg13g2_nor2_1 _15354_ (.A(net6346),
    .B(net3894),
    .Y(_09441_));
 sg13g2_nor4_1 _15355_ (.A(net6219),
    .B(\fpga_top.cpu_top.register_file.rfr_state[1] ),
    .C(net3894),
    .D(_09440_),
    .Y(_09442_));
 sg13g2_a21o_1 _15356_ (.A2(_09437_),
    .A1(net5426),
    .B1(net6220),
    .X(\fpga_top.cpu_top.register_file.next_rfr_state[0] ));
 sg13g2_nor2_1 _15357_ (.A(net5281),
    .B(_09437_),
    .Y(_09443_));
 sg13g2_nor2b_1 _15358_ (.A(_09443_),
    .B_N(net5427),
    .Y(\fpga_top.cpu_top.register_file.next_rfr_state[1] ));
 sg13g2_nand2_1 _15359_ (.Y(_09444_),
    .A(net3894),
    .B(_09436_));
 sg13g2_o21ai_1 _15360_ (.B1(net3895),
    .Y(\fpga_top.cpu_top.register_file.next_rfr_state[2] ),
    .A1(net5427),
    .A2(_09443_));
 sg13g2_nor2_2 _15361_ (.A(net6496),
    .B(net6514),
    .Y(_09445_));
 sg13g2_nor3_2 _15362_ (.A(\fpga_top.cpu_top.cpu_state_machine.cpu_state[0] ),
    .B(net6400),
    .C(_09439_),
    .Y(_09446_));
 sg13g2_nor4_1 _15363_ (.A(net6514),
    .B(net1380),
    .C(_09439_),
    .D(_09446_),
    .Y(_09447_));
 sg13g2_o21ai_1 _15364_ (.B1(net5427),
    .Y(_09448_),
    .A1(_09445_),
    .A2(net6515));
 sg13g2_a21oi_1 _15365_ (.A1(net6219),
    .A2(_09441_),
    .Y(_09449_),
    .B1(_09440_));
 sg13g2_nor2b_2 _15366_ (.A(net6496),
    .B_N(\fpga_top.cpu_top.cpu_state_machine.cpu_state[0] ),
    .Y(_09450_));
 sg13g2_and2_1 _15367_ (.A(net6307),
    .B(_09450_),
    .X(_09451_));
 sg13g2_nor2_1 _15368_ (.A(_09449_),
    .B(_09451_),
    .Y(_09452_));
 sg13g2_nand2_1 _15369_ (.Y(\fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[0] ),
    .A(_09448_),
    .B(_09452_));
 sg13g2_nor2b_2 _15370_ (.A(net6307),
    .B_N(_09450_),
    .Y(_09453_));
 sg13g2_nand2b_2 _15371_ (.Y(_09454_),
    .B(_09450_),
    .A_N(net6533));
 sg13g2_nand3_1 _15372_ (.B(net6219),
    .C(_09441_),
    .A(net6514),
    .Y(_09455_));
 sg13g2_a21oi_1 _15373_ (.A1(_09438_),
    .A2(_09455_),
    .Y(_09456_),
    .B1(_09453_));
 sg13g2_nor2b_1 _15374_ (.A(net6497),
    .B_N(net5427),
    .Y(\fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[1] ));
 sg13g2_and3_1 _15375_ (.X(_09457_),
    .A(_08840_),
    .B(_08843_),
    .C(_08859_));
 sg13g2_nand3_1 _15376_ (.B(_08843_),
    .C(_08859_),
    .A(_08840_),
    .Y(_09458_));
 sg13g2_nand2_2 _15377_ (.Y(_09459_),
    .A(net6307),
    .B(_09445_));
 sg13g2_o21ai_1 _15378_ (.B1(net6308),
    .Y(_09460_),
    .A1(_09439_),
    .A2(_09455_));
 sg13g2_a22oi_1 _15379_ (.Y(_09461_),
    .B1(_09460_),
    .B2(net5427),
    .A2(net4480),
    .A1(_09451_));
 sg13g2_inv_1 _15380_ (.Y(\fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[2] ),
    .A(net6534));
 sg13g2_mux4_1 _15381_ (.S0(net5404),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][0] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][0] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][0] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][0] ),
    .S1(net5402),
    .X(_09462_));
 sg13g2_nor2b_1 _15382_ (.A(_09462_),
    .B_N(net5400),
    .Y(_09463_));
 sg13g2_xor2_1 _15383_ (.B(\fpga_top.io_spi_lite.bit_sel_org[0] ),
    .A(net5829),
    .X(_09464_));
 sg13g2_mux4_1 _15384_ (.S0(net5404),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][0] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][0] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][0] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][0] ),
    .S1(net5402),
    .X(_09465_));
 sg13g2_o21ai_1 _15385_ (.B1(_09464_),
    .Y(_09466_),
    .A1(net5399),
    .A2(_09465_));
 sg13g2_xnor2_1 _15386_ (.Y(_09467_),
    .A(net5830),
    .B(\fpga_top.io_spi_lite.bit_sel_org[1] ));
 sg13g2_mux4_1 _15387_ (.S0(net5405),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][1] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][1] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][1] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][1] ),
    .S1(net5403),
    .X(_09468_));
 sg13g2_nor2b_1 _15388_ (.A(_09468_),
    .B_N(net5401),
    .Y(_09469_));
 sg13g2_mux4_1 _15389_ (.S0(_00008_),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][1] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][1] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][1] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][1] ),
    .S1(_00009_),
    .X(_09470_));
 sg13g2_nor2_1 _15390_ (.A(net5399),
    .B(_09470_),
    .Y(_09471_));
 sg13g2_nor3_1 _15391_ (.A(_09464_),
    .B(_09469_),
    .C(_09471_),
    .Y(_09472_));
 sg13g2_nor2_1 _15392_ (.A(_09467_),
    .B(_09472_),
    .Y(_09473_));
 sg13g2_o21ai_1 _15393_ (.B1(_09473_),
    .Y(_09474_),
    .A1(_09463_),
    .A2(_09466_));
 sg13g2_xnor2_1 _15394_ (.Y(_09475_),
    .A(net5829),
    .B(\fpga_top.io_spi_lite.bit_sel_org[2] ));
 sg13g2_mux4_1 _15395_ (.S0(net5405),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][2] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][2] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][2] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][2] ),
    .S1(net5403),
    .X(_09476_));
 sg13g2_nor2b_1 _15396_ (.A(_09476_),
    .B_N(net5400),
    .Y(_09477_));
 sg13g2_mux4_1 _15397_ (.S0(net5404),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][2] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][2] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][2] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][2] ),
    .S1(net5402),
    .X(_09478_));
 sg13g2_o21ai_1 _15398_ (.B1(_09464_),
    .Y(_09479_),
    .A1(net5399),
    .A2(_09478_));
 sg13g2_mux4_1 _15399_ (.S0(net5404),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][3] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][3] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][3] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][3] ),
    .S1(net5402),
    .X(_09480_));
 sg13g2_nor2b_1 _15400_ (.A(_09480_),
    .B_N(net5400),
    .Y(_09481_));
 sg13g2_mux4_1 _15401_ (.S0(net5405),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][3] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][3] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][3] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][3] ),
    .S1(net5403),
    .X(_09482_));
 sg13g2_nor2_1 _15402_ (.A(net5399),
    .B(_09482_),
    .Y(_09483_));
 sg13g2_nor3_1 _15403_ (.A(_09464_),
    .B(_09481_),
    .C(_09483_),
    .Y(_09484_));
 sg13g2_o21ai_1 _15404_ (.B1(_09467_),
    .Y(_09485_),
    .A1(_09477_),
    .A2(_09479_));
 sg13g2_o21ai_1 _15405_ (.B1(_09474_),
    .Y(_09486_),
    .A1(_09484_),
    .A2(_09485_));
 sg13g2_mux4_1 _15406_ (.S0(net5405),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][7] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][7] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][7] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][7] ),
    .S1(net5403),
    .X(_09487_));
 sg13g2_nor2b_1 _15407_ (.A(_09487_),
    .B_N(net5399),
    .Y(_09488_));
 sg13g2_mux4_1 _15408_ (.S0(net5404),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][7] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][7] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][7] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][7] ),
    .S1(net5402),
    .X(_09489_));
 sg13g2_nor2_1 _15409_ (.A(net5399),
    .B(_09489_),
    .Y(_09490_));
 sg13g2_nor3_1 _15410_ (.A(_09464_),
    .B(_09488_),
    .C(_09490_),
    .Y(_09491_));
 sg13g2_mux4_1 _15411_ (.S0(net5404),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][6] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][6] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][6] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][6] ),
    .S1(net5402),
    .X(_09492_));
 sg13g2_nor2b_1 _15412_ (.A(_09492_),
    .B_N(net5400),
    .Y(_09493_));
 sg13g2_mux4_1 _15413_ (.S0(net5404),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][6] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][6] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][6] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][6] ),
    .S1(net5402),
    .X(_09494_));
 sg13g2_o21ai_1 _15414_ (.B1(_09464_),
    .Y(_09495_),
    .A1(net5399),
    .A2(_09494_));
 sg13g2_o21ai_1 _15415_ (.B1(_09467_),
    .Y(_09496_),
    .A1(_09493_),
    .A2(_09495_));
 sg13g2_mux4_1 _15416_ (.S0(net5405),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][4] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][4] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][4] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][4] ),
    .S1(net5403),
    .X(_09497_));
 sg13g2_nor2b_1 _15417_ (.A(_09497_),
    .B_N(net5401),
    .Y(_09498_));
 sg13g2_mux4_1 _15418_ (.S0(net5404),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][4] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][4] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][4] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][4] ),
    .S1(net5402),
    .X(_09499_));
 sg13g2_o21ai_1 _15419_ (.B1(_09464_),
    .Y(_09500_),
    .A1(net5399),
    .A2(_09499_));
 sg13g2_mux4_1 _15420_ (.S0(net5405),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][5] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][5] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][5] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][5] ),
    .S1(net5403),
    .X(_09501_));
 sg13g2_nor2b_1 _15421_ (.A(_09501_),
    .B_N(net5401),
    .Y(_09502_));
 sg13g2_mux4_1 _15422_ (.S0(net5405),
    .A0(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][5] ),
    .A1(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][5] ),
    .A2(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][5] ),
    .A3(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][5] ),
    .S1(net5403),
    .X(_09503_));
 sg13g2_nor2_1 _15423_ (.A(net5401),
    .B(_09503_),
    .Y(_09504_));
 sg13g2_nor3_1 _15424_ (.A(_09464_),
    .B(_09502_),
    .C(_09504_),
    .Y(_09505_));
 sg13g2_nor2_1 _15425_ (.A(_09467_),
    .B(_09505_),
    .Y(_09506_));
 sg13g2_o21ai_1 _15426_ (.B1(_09506_),
    .Y(_09507_),
    .A1(_09498_),
    .A2(_09500_));
 sg13g2_o21ai_1 _15427_ (.B1(_09507_),
    .Y(_09508_),
    .A1(_09491_),
    .A2(_09496_));
 sg13g2_mux2_1 _15428_ (.A0(_09486_),
    .A1(_09508_),
    .S(_09475_),
    .X(_09509_));
 sg13g2_nor2_2 _15429_ (.A(_09408_),
    .B(_09509_),
    .Y(\fpga_top.io_spi_lite.org_mosi ));
 sg13g2_mux4_1 _15430_ (.S0(\fpga_top.io_spi_lite.spi_mode[5] ),
    .A0(\fpga_top.io_spi_lite.org_mosi ),
    .A1(net1324),
    .A2(net1348),
    .A3(net1363),
    .S1(net6359),
    .X(_09510_));
 sg13g2_mux2_1 _15431_ (.A0(net1342),
    .A1(net1350),
    .S(\fpga_top.io_spi_lite.spi_mode[4] ),
    .X(_09511_));
 sg13g2_nor2b_1 _15432_ (.A(net6359),
    .B_N(net1343),
    .Y(_09512_));
 sg13g2_a21oi_1 _15433_ (.A1(net6359),
    .A2(net6430),
    .Y(_09513_),
    .B1(_09512_));
 sg13g2_o21ai_1 _15434_ (.B1(net3829),
    .Y(_09514_),
    .A1(net6332),
    .A2(_09511_));
 sg13g2_a21oi_1 _15435_ (.A1(net6332),
    .A2(_09513_),
    .Y(_09515_),
    .B1(_09514_));
 sg13g2_a21o_1 _15436_ (.A2(_09510_),
    .A1(_06913_),
    .B1(_09515_),
    .X(\fpga_top.io_spi_lite.spi_mosi_pre ));
 sg13g2_nand2b_1 _15437_ (.Y(_09516_),
    .B(net3664),
    .A_N(\fpga_top.uart_top.uart_if.tx_state[1] ));
 sg13g2_nand2_1 _15438_ (.Y(\fpga_top.uart_top.uart_if.next_tx_state[0] ),
    .A(net5284),
    .B(net3665));
 sg13g2_nor3_1 _15439_ (.A(net6283),
    .B(_09340_),
    .C(_09343_),
    .Y(_09517_));
 sg13g2_inv_1 _15440_ (.Y(_09518_),
    .A(_09517_));
 sg13g2_nor4_2 _15441_ (.A(net6447),
    .B(net1392),
    .C(net3946),
    .Y(_09519_),
    .D(_09518_));
 sg13g2_inv_1 _15442_ (.Y(_09520_),
    .A(net1393));
 sg13g2_nor2_1 _15443_ (.A(net3665),
    .B(_09520_),
    .Y(\fpga_top.uart_top.uart_if.next_tx_state[1] ));
 sg13g2_nand2b_1 _15444_ (.Y(_09521_),
    .B(net6188),
    .A_N(net1602));
 sg13g2_nor3_1 _15445_ (.A(\fpga_top.uart_top.uart_if.rx_state[3] ),
    .B(net3928),
    .C(_09521_),
    .Y(_09522_));
 sg13g2_nand2_1 _15446_ (.Y(_09523_),
    .A(net1602),
    .B(net6188));
 sg13g2_nand4_1 _15447_ (.B(net6188),
    .C(_06672_),
    .A(net1602),
    .Y(_09524_),
    .D(_09292_));
 sg13g2_a21oi_1 _15448_ (.A1(_09292_),
    .A2(net3929),
    .Y(_09525_),
    .B1(net5173));
 sg13g2_nor2b_2 _15449_ (.A(net6350),
    .B_N(net3928),
    .Y(_09526_));
 sg13g2_nor2_1 _15450_ (.A(_09284_),
    .B(_09526_),
    .Y(_09527_));
 sg13g2_nor2_1 _15451_ (.A(_09521_),
    .B(_09527_),
    .Y(_09528_));
 sg13g2_nand2_1 _15452_ (.Y(_09529_),
    .A(_06672_),
    .B(_09286_));
 sg13g2_o21ai_1 _15453_ (.B1(_09298_),
    .Y(_09530_),
    .A1(_09284_),
    .A2(_09526_));
 sg13g2_nand3_1 _15454_ (.B(_09529_),
    .C(_09530_),
    .A(net5073),
    .Y(_09531_));
 sg13g2_o21ai_1 _15455_ (.B1(_09531_),
    .Y(_09532_),
    .A1(net5073),
    .A2(_09528_));
 sg13g2_nand3_1 _15456_ (.B(_09525_),
    .C(_09532_),
    .A(net6189),
    .Y(\fpga_top.uart_top.uart_if.next_rx_state[0] ));
 sg13g2_nand2_1 _15457_ (.Y(_09533_),
    .A(_09287_),
    .B(_09292_));
 sg13g2_or2_1 _15458_ (.X(_09534_),
    .B(_00124_),
    .A(_00120_));
 sg13g2_and2_1 _15459_ (.A(_00120_),
    .B(_00124_),
    .X(_09535_));
 sg13g2_a21oi_1 _15460_ (.A1(_00122_),
    .A2(_09534_),
    .Y(_09536_),
    .B1(_09535_));
 sg13g2_o21ai_1 _15461_ (.B1(_00118_),
    .Y(_09537_),
    .A1(_00122_),
    .A2(_09534_));
 sg13g2_a21oi_1 _15462_ (.A1(_00122_),
    .A2(_09535_),
    .Y(_09538_),
    .B1(_00118_));
 sg13g2_nor2_1 _15463_ (.A(_09536_),
    .B(_09538_),
    .Y(_09539_));
 sg13g2_nor2_1 _15464_ (.A(net1394),
    .B(_09539_),
    .Y(_09540_));
 sg13g2_a21oi_2 _15465_ (.B1(_09540_),
    .Y(_09541_),
    .A2(_09537_),
    .A1(_09536_));
 sg13g2_nor2b_1 _15466_ (.A(_09292_),
    .B_N(_09541_),
    .Y(_09542_));
 sg13g2_and2_1 _15467_ (.A(_09522_),
    .B(_09542_),
    .X(_09543_));
 sg13g2_a21oi_1 _15468_ (.A1(net5073),
    .A2(_09528_),
    .Y(_09544_),
    .B1(_09543_));
 sg13g2_nand4_1 _15469_ (.B(_09529_),
    .C(_09533_),
    .A(net6189),
    .Y(\fpga_top.uart_top.uart_if.next_rx_state[1] ),
    .D(_09544_));
 sg13g2_nor2_1 _15470_ (.A(_09292_),
    .B(_09523_),
    .Y(_09545_));
 sg13g2_mux2_1 _15471_ (.A0(_09526_),
    .A1(_09297_),
    .S(_09545_),
    .X(\fpga_top.uart_top.uart_if.next_rx_state[2] ));
 sg13g2_a22oi_1 _15472_ (.Y(_09546_),
    .B1(_09526_),
    .B2(_09545_),
    .A2(_09292_),
    .A1(_09287_));
 sg13g2_o21ai_1 _15473_ (.B1(_09546_),
    .Y(\fpga_top.uart_top.uart_if.next_rx_state[3] ),
    .A1(net1602),
    .A2(_09285_));
 sg13g2_a21o_1 _15474_ (.A2(\fpga_top.uart_top.uart_logics.next_status_dump[1] ),
    .A1(_06997_),
    .B1(_08733_),
    .X(_09547_));
 sg13g2_inv_4 _15475_ (.A(net4569),
    .Y(_09548_));
 sg13g2_nor2b_1 _15476_ (.A(\fpga_top.cpu_top.inst_mem_read.imr_stat ),
    .B_N(_09446_),
    .Y(_09549_));
 sg13g2_nand2b_1 _15477_ (.Y(_09550_),
    .B(_09446_),
    .A_N(\fpga_top.cpu_top.inst_mem_read.imr_stat ));
 sg13g2_nand2_1 _15478_ (.Y(_09551_),
    .A(_09548_),
    .B(net5163));
 sg13g2_nand3_1 _15479_ (.B(_09548_),
    .C(net5163),
    .A(net4570),
    .Y(_09552_));
 sg13g2_nor2_1 _15480_ (.A(net1807),
    .B(net6306),
    .Y(_09553_));
 sg13g2_a22oi_1 _15481_ (.Y(_09554_),
    .B1(_09552_),
    .B2(_09553_),
    .A2(_08728_),
    .A1(_06933_));
 sg13g2_inv_1 _15482_ (.Y(\fpga_top.qspi_if.inner_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/qspi_if.v:768$329.$result[0] ),
    .A(_09554_));
 sg13g2_nor4_2 _15483_ (.A(net5632),
    .B(net5631),
    .C(_06546_),
    .Y(_09555_),
    .D(_06986_));
 sg13g2_nor2b_2 _15484_ (.A(net3315),
    .B_N(_00084_),
    .Y(_09556_));
 sg13g2_nor2_1 _15485_ (.A(_09555_),
    .B(_09556_),
    .Y(_09557_));
 sg13g2_nor2_1 _15486_ (.A(net1378),
    .B(_09557_),
    .Y(_09558_));
 sg13g2_o21ai_1 _15487_ (.B1(_06663_),
    .Y(_09559_),
    .A1(_09555_),
    .A2(_09556_));
 sg13g2_and2_1 _15488_ (.A(_08845_),
    .B(_09559_),
    .X(_09560_));
 sg13g2_nor4_1 _15489_ (.A(net1807),
    .B(\fpga_top.qspi_if.inner_state[1] ),
    .C(_09552_),
    .D(net4550),
    .Y(_09561_));
 sg13g2_a21oi_1 _15490_ (.A1(\fpga_top.qspi_if.inner_state[1] ),
    .A2(_08856_),
    .Y(_09562_),
    .B1(_09561_));
 sg13g2_a21oi_1 _15491_ (.A1(net1807),
    .A2(\fpga_top.qspi_if.inner_state[1] ),
    .Y(\fpga_top.qspi_if.inner_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/qspi_if.v:768$329.$result[1] ),
    .B1(_09562_));
 sg13g2_nand2_1 _15492_ (.Y(_09563_),
    .A(\fpga_top.bus_gather.u_read_adr[31] ),
    .B(net5285));
 sg13g2_and3_1 _15493_ (.X(_09564_),
    .A(\fpga_top.bus_gather.u_read_adr[31] ),
    .B(net5613),
    .C(net5285));
 sg13g2_nand2_1 _15494_ (.Y(_09565_),
    .A(\fpga_top.bus_gather.u_read_adr[13] ),
    .B(\fpga_top.bus_gather.u_read_adr[12] ));
 sg13g2_mux2_1 _15495_ (.A0(_08883_),
    .A1(_09565_),
    .S(net5158),
    .X(_09566_));
 sg13g2_nand2_1 _15496_ (.Y(_09567_),
    .A(\fpga_top.bus_gather.u_read_adr[10] ),
    .B(net5158));
 sg13g2_o21ai_1 _15497_ (.B1(_09567_),
    .Y(_09568_),
    .A1(_08012_),
    .A2(net5158));
 sg13g2_or2_1 _15498_ (.X(_09569_),
    .B(_09568_),
    .A(_09566_));
 sg13g2_nand3_1 _15499_ (.B(\fpga_top.bus_gather.u_read_adr[15] ),
    .C(net5159),
    .A(\fpga_top.bus_gather.u_read_adr[14] ),
    .Y(_09570_));
 sg13g2_o21ai_1 _15500_ (.B1(_09570_),
    .Y(_09571_),
    .A1(_08878_),
    .A2(net5159));
 sg13g2_nor2_1 _15501_ (.A(_08278_),
    .B(net5159),
    .Y(_09572_));
 sg13g2_a21oi_1 _15502_ (.A1(_06522_),
    .A2(net5159),
    .Y(_09573_),
    .B1(_09572_));
 sg13g2_nand2_1 _15503_ (.Y(_09574_),
    .A(_09571_),
    .B(_09573_));
 sg13g2_or2_1 _15504_ (.X(_09575_),
    .B(_09574_),
    .A(_09569_));
 sg13g2_nand3_1 _15505_ (.B(_06513_),
    .C(_06514_),
    .A(_06511_),
    .Y(_09576_));
 sg13g2_mux2_1 _15506_ (.A0(_08905_),
    .A1(_09576_),
    .S(net5158),
    .X(_09577_));
 sg13g2_nor2_1 _15507_ (.A(_08313_),
    .B(net5158),
    .Y(_09578_));
 sg13g2_a21oi_2 _15508_ (.B1(_09578_),
    .Y(_09579_),
    .A2(net5158),
    .A1(\fpga_top.bus_gather.u_read_adr[9] ));
 sg13g2_nand2_1 _15509_ (.Y(_09580_),
    .A(_06508_),
    .B(net5159));
 sg13g2_o21ai_1 _15510_ (.B1(_09580_),
    .Y(_09581_),
    .A1(_08222_),
    .A2(net5160));
 sg13g2_inv_1 _15511_ (.Y(_09582_),
    .A(_09581_));
 sg13g2_nor2_1 _15512_ (.A(_08101_),
    .B(net5158),
    .Y(_09583_));
 sg13g2_a21oi_2 _15513_ (.B1(_09583_),
    .Y(_09584_),
    .A2(net5159),
    .A1(\fpga_top.bus_gather.u_read_adr[5] ));
 sg13g2_and2_1 _15514_ (.A(_09581_),
    .B(_09584_),
    .X(_09585_));
 sg13g2_nand2_1 _15515_ (.Y(_09586_),
    .A(_09581_),
    .B(_09584_));
 sg13g2_nor3_1 _15516_ (.A(_09577_),
    .B(_09579_),
    .C(_09586_),
    .Y(_09587_));
 sg13g2_nand2_1 _15517_ (.Y(_09588_),
    .A(net5616),
    .B(net5159));
 sg13g2_o21ai_1 _15518_ (.B1(_09588_),
    .Y(_09589_),
    .A1(_08158_),
    .A2(net5160));
 sg13g2_nor2_2 _15519_ (.A(\fpga_top.cpu_top.data_rw_mem.dma_io_radr_en ),
    .B(net5158),
    .Y(_09590_));
 sg13g2_nor2_1 _15520_ (.A(_08191_),
    .B(net5159),
    .Y(_09591_));
 sg13g2_a21oi_2 _15521_ (.B1(_09591_),
    .Y(_09592_),
    .A2(net5160),
    .A1(net5615));
 sg13g2_nand2b_1 _15522_ (.Y(_09593_),
    .B(_09592_),
    .A_N(_09589_));
 sg13g2_nor2_2 _15523_ (.A(_09590_),
    .B(_09593_),
    .Y(_09594_));
 sg13g2_nand2_1 _15524_ (.Y(_09595_),
    .A(_09587_),
    .B(_09594_));
 sg13g2_nor2_1 _15525_ (.A(_09575_),
    .B(_09595_),
    .Y(\fpga_top.interrupter.re_int_enable ));
 sg13g2_nand2_1 _15526_ (.Y(_09596_),
    .A(_09589_),
    .B(_09592_));
 sg13g2_nor2_2 _15527_ (.A(_09590_),
    .B(_09596_),
    .Y(_09597_));
 sg13g2_nand2_2 _15528_ (.Y(_09598_),
    .A(_09587_),
    .B(_09597_));
 sg13g2_nor2_1 _15529_ (.A(_09575_),
    .B(_09598_),
    .Y(\fpga_top.interrupter.re_int_status ));
 sg13g2_nand2b_1 _15530_ (.Y(_09599_),
    .B(_09579_),
    .A_N(_09577_));
 sg13g2_nor2_1 _15531_ (.A(_09586_),
    .B(_09599_),
    .Y(_09600_));
 sg13g2_nand2_2 _15532_ (.Y(_09601_),
    .A(_09594_),
    .B(_09600_));
 sg13g2_nor2_1 _15533_ (.A(_09575_),
    .B(_09601_),
    .Y(\fpga_top.io_frc.re_frc_vallo ));
 sg13g2_nand2_1 _15534_ (.Y(_09602_),
    .A(_09597_),
    .B(_09600_));
 sg13g2_nor2_1 _15535_ (.A(_09575_),
    .B(_09602_),
    .Y(\fpga_top.io_frc.re_frc_valhi ));
 sg13g2_or2_1 _15536_ (.X(_09603_),
    .B(_09599_),
    .A(_09575_));
 sg13g2_nor2_1 _15537_ (.A(_09590_),
    .B(_09592_),
    .Y(_09604_));
 sg13g2_nor3_1 _15538_ (.A(_09589_),
    .B(_09590_),
    .C(_09592_),
    .Y(_09605_));
 sg13g2_nand2_2 _15539_ (.Y(_09606_),
    .A(_09585_),
    .B(_09605_));
 sg13g2_nor2_1 _15540_ (.A(_09603_),
    .B(_09606_),
    .Y(\fpga_top.io_frc.re_frc_cmplo ));
 sg13g2_nand3_1 _15541_ (.B(_09589_),
    .C(_09604_),
    .A(_09585_),
    .Y(_09607_));
 sg13g2_nor2_1 _15542_ (.A(_09603_),
    .B(_09607_),
    .Y(\fpga_top.io_frc.re_frc_cmphi ));
 sg13g2_nor2b_1 _15543_ (.A(_09581_),
    .B_N(_09584_),
    .Y(_09608_));
 sg13g2_inv_1 _15544_ (.Y(_09609_),
    .A(_09608_));
 sg13g2_nand2_1 _15545_ (.Y(_09610_),
    .A(_09594_),
    .B(_09608_));
 sg13g2_nor2_1 _15546_ (.A(_09603_),
    .B(_09610_),
    .Y(\fpga_top.io_frc.re_frc_cntrl ));
 sg13g2_nand2b_1 _15547_ (.Y(_09611_),
    .B(_09568_),
    .A_N(_09566_));
 sg13g2_or2_1 _15548_ (.X(_09612_),
    .B(_09611_),
    .A(_09574_));
 sg13g2_nor2_1 _15549_ (.A(_09601_),
    .B(_09612_),
    .Y(\fpga_top.io_uart_out.re_uart_char ));
 sg13g2_nor2_1 _15550_ (.A(_09602_),
    .B(_09612_),
    .Y(\fpga_top.io_uart_out.re_uart_full ));
 sg13g2_or2_1 _15551_ (.X(_09613_),
    .B(_09612_),
    .A(_09599_));
 sg13g2_nor2_1 _15552_ (.A(_09606_),
    .B(_09613_),
    .Y(\fpga_top.io_uart_out.re_uart_term ));
 sg13g2_nor2_1 _15553_ (.A(_09607_),
    .B(_09613_),
    .Y(\fpga_top.io_uart_out.re_uart_rxch ));
 sg13g2_nor2_1 _15554_ (.A(_09610_),
    .B(_09613_),
    .Y(\fpga_top.io_uart_out.re_uart_rxec ));
 sg13g2_nor2_1 _15555_ (.A(_08898_),
    .B(_08982_),
    .Y(_09614_));
 sg13g2_nand2_2 _15556_ (.Y(_09615_),
    .A(_08909_),
    .B(_09614_));
 sg13g2_and2_1 _15557_ (.A(_08886_),
    .B(_08888_),
    .X(_09616_));
 sg13g2_nand2_2 _15558_ (.Y(_09617_),
    .A(_08892_),
    .B(_09616_));
 sg13g2_nor2_1 _15559_ (.A(_09615_),
    .B(_09617_),
    .Y(_09618_));
 sg13g2_nor3_1 _15560_ (.A(net6117),
    .B(_09615_),
    .C(_09617_),
    .Y(_00041_));
 sg13g2_nor2_1 _15561_ (.A(_09595_),
    .B(_09612_),
    .Y(\fpga_top.io_led.re_led_value ));
 sg13g2_nor2_1 _15562_ (.A(_09598_),
    .B(_09612_),
    .Y(\fpga_top.io_led.re_gpi_value ));
 sg13g2_nor4_1 _15563_ (.A(_09577_),
    .B(_09579_),
    .C(_09609_),
    .D(_09612_),
    .Y(_09619_));
 sg13g2_and2_1 _15564_ (.A(_09594_),
    .B(_09619_),
    .X(\fpga_top.io_led.re_gpio_out_value ));
 sg13g2_and2_1 _15565_ (.A(_09597_),
    .B(_09619_),
    .X(\fpga_top.io_led.re_gpio_in_value ));
 sg13g2_and2_1 _15566_ (.A(_09605_),
    .B(_09619_),
    .X(\fpga_top.io_led.re_gpio_en_value ));
 sg13g2_o21ai_1 _15567_ (.B1(_09100_),
    .Y(_09620_),
    .A1(_09088_),
    .A2(net6571));
 sg13g2_nand2_1 _15568_ (.Y(\fpga_top.qspi_if.sio_out_enbl_pre ),
    .A(net5378),
    .B(net6572));
 sg13g2_nand2b_1 _15569_ (.Y(_09621_),
    .B(_09571_),
    .A_N(_09573_));
 sg13g2_or2_1 _15570_ (.X(_09622_),
    .B(_09621_),
    .A(_09611_));
 sg13g2_nor2_1 _15571_ (.A(_09601_),
    .B(_09622_),
    .Y(\fpga_top.qspi_if.re_qspi_latency0 ));
 sg13g2_nor2_1 _15572_ (.A(_09602_),
    .B(_09622_),
    .Y(\fpga_top.qspi_if.re_qspi_latency1 ));
 sg13g2_or2_1 _15573_ (.X(_09623_),
    .B(_09622_),
    .A(_09599_));
 sg13g2_nor2_1 _15574_ (.A(_09606_),
    .B(_09623_),
    .Y(\fpga_top.qspi_if.re_qspi_latency2 ));
 sg13g2_nor2_1 _15575_ (.A(_09607_),
    .B(_09623_),
    .Y(\fpga_top.qspi_if.re_qspi_sckdiv ));
 sg13g2_nor2_1 _15576_ (.A(_09609_),
    .B(_09623_),
    .Y(_09624_));
 sg13g2_and2_1 _15577_ (.A(_09594_),
    .B(_09624_),
    .X(\fpga_top.qspi_if.re_qspi_rdcmd0 ));
 sg13g2_and2_1 _15578_ (.A(_09597_),
    .B(_09624_),
    .X(\fpga_top.qspi_if.re_qspi_rdcmd1 ));
 sg13g2_and2_1 _15579_ (.A(_09605_),
    .B(_09624_),
    .X(\fpga_top.qspi_if.re_qspi_wrcmd0 ));
 sg13g2_and3_1 _15580_ (.X(\fpga_top.qspi_if.re_qspi_wrcmd1 ),
    .A(_09589_),
    .B(_09604_),
    .C(_09624_));
 sg13g2_nor3_1 _15581_ (.A(_09582_),
    .B(_09584_),
    .C(_09623_),
    .Y(_09625_));
 sg13g2_and2_1 _15582_ (.A(_09594_),
    .B(_09625_),
    .X(\fpga_top.qspi_if.re_qspi_rdwrch ));
 sg13g2_and2_1 _15583_ (.A(_09597_),
    .B(_09625_),
    .X(\fpga_top.qspi_if.re_qspi_rdedge ));
 sg13g2_o21ai_1 _15584_ (.B1(_00121_),
    .Y(\fpga_top.tx ),
    .A1(\fpga_top.uart_top.uart_if.tx_state[1] ),
    .A2(\fpga_top.uart_top.uart_if.tx_state[0] ));
 sg13g2_nor4_1 _15585_ (.A(_07007_),
    .B(_07009_),
    .C(_08688_),
    .D(_08703_),
    .Y(_09626_));
 sg13g2_nor2_1 _15586_ (.A(_07009_),
    .B(_07018_),
    .Y(_09627_));
 sg13g2_nand3_1 _15587_ (.B(_08694_),
    .C(_09626_),
    .A(_07019_),
    .Y(_09628_));
 sg13g2_nand3b_1 _15588_ (.B(_06956_),
    .C(\fpga_top.uart_top.uart_rec_char.pdata[4] ),
    .Y(_09629_),
    .A_N(\fpga_top.uart_top.uart_rec_char.pdata[6] ));
 sg13g2_nor2_2 _15589_ (.A(net5626),
    .B(_09629_),
    .Y(_09630_));
 sg13g2_nor3_1 _15590_ (.A(net5628),
    .B(_06960_),
    .C(_09629_),
    .Y(_09631_));
 sg13g2_o21ai_1 _15591_ (.B1(_06966_),
    .Y(_09632_),
    .A1(net5625),
    .A2(_06978_));
 sg13g2_nor2b_2 _15592_ (.A(_06957_),
    .B_N(_09632_),
    .Y(_09633_));
 sg13g2_nor4_2 _15593_ (.A(net5626),
    .B(_06957_),
    .C(_06964_),
    .Y(_09634_),
    .D(_06977_));
 sg13g2_nor3_2 _15594_ (.A(_09631_),
    .B(_09633_),
    .C(_09634_),
    .Y(_09635_));
 sg13g2_nand2b_1 _15595_ (.Y(_09636_),
    .B(_09635_),
    .A_N(_09630_));
 sg13g2_and3_2 _15596_ (.X(_09637_),
    .A(\fpga_top.uart_top.uart_rec_char.data_en ),
    .B(_09628_),
    .C(_09636_));
 sg13g2_inv_1 _15597_ (.Y(_09638_),
    .A(_09637_));
 sg13g2_nand2_1 _15598_ (.Y(_09639_),
    .A(net2790),
    .B(\fpga_top.uart_top.uart_rec_char.data_cntr[0] ));
 sg13g2_nand3_1 _15599_ (.B(net3513),
    .C(net2141),
    .A(net2790),
    .Y(_09640_));
 sg13g2_nor3_2 _15600_ (.A(net1396),
    .B(_09638_),
    .C(_09640_),
    .Y(\fpga_top.uart_top.uart_rec_char.word_valid_pre ));
 sg13g2_nor2_1 _15601_ (.A(_06771_),
    .B(_06773_),
    .Y(_00027_));
 sg13g2_nand4_1 _15602_ (.B(\fpga_top.cpu_top.decoder.illegal_ops_inst[1] ),
    .C(\fpga_top.cpu_top.cpu_state_machine.cpu_state[2] ),
    .A(net3864),
    .Y(_09641_),
    .D(_09445_));
 sg13g2_a21oi_1 _15603_ (.A1(\fpga_top.cpu_top.decoder.illegal_ops_inst[5] ),
    .A2(_07297_),
    .Y(_00026_),
    .B1(net3865));
 sg13g2_nor2_1 _15604_ (.A(_07377_),
    .B(net6308),
    .Y(_00025_));
 sg13g2_nor2_1 _15605_ (.A(_07371_),
    .B(net6308),
    .Y(_00024_));
 sg13g2_or2_1 _15606_ (.X(_09642_),
    .B(_09621_),
    .A(_09569_));
 sg13g2_nor2_1 _15607_ (.A(_09595_),
    .B(_09642_),
    .Y(\fpga_top.io_spi_lite.re_spi_mode ));
 sg13g2_nor2_1 _15608_ (.A(_09598_),
    .B(_09642_),
    .Y(\fpga_top.io_spi_lite.re_spi_sdiv ));
 sg13g2_or3_1 _15609_ (.A(_09577_),
    .B(_09579_),
    .C(_09642_),
    .X(_09643_));
 sg13g2_nor2_2 _15610_ (.A(_09606_),
    .B(_09643_),
    .Y(\fpga_top.io_spi_lite.re_spi_mosi ));
 sg13g2_nor2_1 _15611_ (.A(_09607_),
    .B(_09643_),
    .Y(\fpga_top.io_spi_lite.re_spi_miso ));
 sg13g2_and2_1 _15612_ (.A(_06649_),
    .B(_08970_),
    .X(_09644_));
 sg13g2_nand2b_1 _15613_ (.Y(_09645_),
    .B(net1777),
    .A_N(_08969_));
 sg13g2_nor2b_2 _15614_ (.A(_09644_),
    .B_N(_09645_),
    .Y(_09646_));
 sg13g2_nand2b_1 _15615_ (.Y(_09647_),
    .B(_09645_),
    .A_N(_09644_));
 sg13g2_and2_1 _15616_ (.A(net1655),
    .B(net1427),
    .X(_09648_));
 sg13g2_and3_1 _15617_ (.X(\fpga_top.io_spi_lite.miso_read_next_byte ),
    .A(net1407),
    .B(net1778),
    .C(_09648_));
 sg13g2_nand4_1 _15618_ (.B(_08843_),
    .C(_08859_),
    .A(\fpga_top.cpu_top.data_rw_mem.wbk_rd_reg_ma ),
    .Y(_09649_),
    .D(_09451_));
 sg13g2_a21oi_1 _15619_ (.A1(net5096),
    .A2(net4480),
    .Y(_09650_),
    .B1(net5436));
 sg13g2_and2_1 _15620_ (.A(_06664_),
    .B(_08874_),
    .X(_09651_));
 sg13g2_nor2b_2 _15621_ (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[31] ),
    .B_N(_09651_),
    .Y(_09652_));
 sg13g2_nor2_1 _15622_ (.A(_06564_),
    .B(net4937),
    .Y(_09653_));
 sg13g2_a21oi_1 _15623_ (.A1(net5665),
    .A2(net4936),
    .Y(_09654_),
    .B1(_09653_));
 sg13g2_a21oi_2 _15624_ (.B1(_09654_),
    .Y(_09655_),
    .A2(_09650_),
    .A1(_09649_));
 sg13g2_nand2_1 _15625_ (.Y(_09656_),
    .A(\fpga_top.cpu_top.csr_wadr_mon[1] ),
    .B(net4932));
 sg13g2_o21ai_1 _15626_ (.B1(_09656_),
    .Y(_09657_),
    .A1(_06560_),
    .A2(net4936));
 sg13g2_inv_2 _15627_ (.Y(_09658_),
    .A(_09657_));
 sg13g2_nand2_2 _15628_ (.Y(_09659_),
    .A(_09655_),
    .B(_09658_));
 sg13g2_nand2_1 _15629_ (.Y(_09660_),
    .A(\fpga_top.cpu_top.csr_wadr_mon[3] ),
    .B(net4937));
 sg13g2_o21ai_1 _15630_ (.B1(_09660_),
    .Y(_09661_),
    .A1(_06569_),
    .A2(net4937));
 sg13g2_nand2_1 _15631_ (.Y(_09662_),
    .A(\fpga_top.cpu_top.csr_wadr_mon[4] ),
    .B(net4936));
 sg13g2_o21ai_1 _15632_ (.B1(_09662_),
    .Y(_09663_),
    .A1(_06576_),
    .A2(net4936));
 sg13g2_inv_1 _15633_ (.Y(_09664_),
    .A(_09663_));
 sg13g2_nor2b_1 _15634_ (.A(net4937),
    .B_N(\fpga_top.cpu_top.br_ofs[2] ),
    .Y(_09665_));
 sg13g2_a21oi_2 _15635_ (.B1(_09665_),
    .Y(_09666_),
    .A2(net4937),
    .A1(\fpga_top.cpu_top.csr_wadr_mon[2] ));
 sg13g2_a21o_2 _15636_ (.A2(net4937),
    .A1(\fpga_top.cpu_top.csr_wadr_mon[2] ),
    .B1(_09665_),
    .X(_09667_));
 sg13g2_or3_1 _15637_ (.A(_09661_),
    .B(_09663_),
    .C(_09667_),
    .X(_09668_));
 sg13g2_or2_1 _15638_ (.X(_09669_),
    .B(_09668_),
    .A(_09659_));
 sg13g2_and2_1 _15639_ (.A(net5708),
    .B(net1402),
    .X(_09670_));
 sg13g2_a221oi_1 _15640_ (.B2(net3790),
    .C1(_09670_),
    .B1(net5330),
    .A1(net1910),
    .Y(_09671_),
    .A2(net5334));
 sg13g2_inv_1 _15641_ (.Y(_09672_),
    .A(_09671_));
 sg13g2_nor2_1 _15642_ (.A(\fpga_top.cpu_top.data_rw_mem.unsigned_bit_dly ),
    .B(net5439),
    .Y(_09673_));
 sg13g2_nand3b_1 _15643_ (.B(_09672_),
    .C(_09673_),
    .Y(_09674_),
    .A_N(\fpga_top.cpu_top.data_rw_mem.req_hw_dly ));
 sg13g2_a22oi_1 _15644_ (.Y(_09675_),
    .B1(net5333),
    .B2(\fpga_top.qspi_if.word_data[7] ),
    .A2(\fpga_top.qspi_if.word_data[23] ),
    .A1(net5704));
 sg13g2_nand2_1 _15645_ (.Y(_09676_),
    .A(\fpga_top.cpu_top.data_rw_mem.req_hw_dly ),
    .B(_09673_));
 sg13g2_o21ai_1 _15646_ (.B1(_09674_),
    .Y(_09677_),
    .A1(_09675_),
    .A2(_09676_));
 sg13g2_and2_1 _15647_ (.A(net5701),
    .B(\fpga_top.qspi_if.word_data[0] ),
    .X(_09678_));
 sg13g2_a21oi_1 _15648_ (.A1(net5440),
    .A2(_09678_),
    .Y(_09679_),
    .B1(net4925));
 sg13g2_a21oi_1 _15649_ (.A1(net4476),
    .A2(_09679_),
    .Y(_09680_),
    .B1(net5429));
 sg13g2_o21ai_1 _15650_ (.B1(_09680_),
    .Y(_09681_),
    .A1(_07907_),
    .A2(net4476));
 sg13g2_nand2_1 _15651_ (.Y(_09682_),
    .A(\fpga_top.io_spi_lite.spi_mode[10] ),
    .B(net5838));
 sg13g2_a21oi_1 _15652_ (.A1(\fpga_top.io_frc.frc_cmp_val[56] ),
    .A2(net5721),
    .Y(_09683_),
    .B1(net5729));
 sg13g2_a21o_1 _15653_ (.A2(net5729),
    .A1(_06722_),
    .B1(_09683_),
    .X(_09684_));
 sg13g2_a21oi_1 _15654_ (.A1(\fpga_top.io_frc.frc_cntr_val[56] ),
    .A2(net5738),
    .Y(_09685_),
    .B1(net5749));
 sg13g2_o21ai_1 _15655_ (.B1(_09685_),
    .Y(_09686_),
    .A1(net5741),
    .A2(_09684_));
 sg13g2_nor2_1 _15656_ (.A(\fpga_top.qspi_if.re_qspi_latency_dly[7] ),
    .B(net5691),
    .Y(_09687_));
 sg13g2_or2_1 _15657_ (.X(_09688_),
    .B(\fpga_top.qspi_if.re_qspi_latency_dly[6] ),
    .A(\fpga_top.qspi_if.re_qspi_latency_dly[7] ));
 sg13g2_nor2_2 _15658_ (.A(\fpga_top.qspi_if.re_qspi_latency_dly[9] ),
    .B(net5690),
    .Y(_09689_));
 sg13g2_or2_1 _15659_ (.X(_09690_),
    .B(net5690),
    .A(\fpga_top.qspi_if.re_qspi_latency_dly[9] ));
 sg13g2_nor2_2 _15660_ (.A(_09688_),
    .B(_09690_),
    .Y(_09691_));
 sg13g2_nor2_2 _15661_ (.A(\fpga_top.qspi_if.re_qspi_latency_dly[5] ),
    .B(net5693),
    .Y(_09692_));
 sg13g2_or2_1 _15662_ (.X(_09693_),
    .B(net5692),
    .A(\fpga_top.qspi_if.re_qspi_latency_dly[5] ));
 sg13g2_nand2_2 _15663_ (.Y(_09694_),
    .A(_09691_),
    .B(_09692_));
 sg13g2_nor2_2 _15664_ (.A(net5694),
    .B(_09693_),
    .Y(_09695_));
 sg13g2_nor2_2 _15665_ (.A(net5696),
    .B(_09694_),
    .Y(_09696_));
 sg13g2_nand2_2 _15666_ (.Y(_09697_),
    .A(_09691_),
    .B(_09695_));
 sg13g2_nor2_2 _15667_ (.A(\fpga_top.io_spi_lite.re_spi_value_dly[2] ),
    .B(net5834),
    .Y(_09698_));
 sg13g2_or2_1 _15668_ (.X(_09699_),
    .B(net5835),
    .A(\fpga_top.io_spi_lite.re_spi_value_dly[2] ));
 sg13g2_nor2_2 _15669_ (.A(net5837),
    .B(_09699_),
    .Y(_09700_));
 sg13g2_or2_1 _15670_ (.X(_09701_),
    .B(\fpga_top.interrupter.re_int_dly[0] ),
    .A(\fpga_top.interrupter.re_int_dly[1] ));
 sg13g2_or2_1 _15671_ (.X(_09702_),
    .B(\fpga_top.qspi_if.re_qspi_latency_dly[0] ),
    .A(\fpga_top.qspi_if.re_qspi_latency_dly[1] ));
 sg13g2_or3_1 _15672_ (.A(net5698),
    .B(_09701_),
    .C(net5329),
    .X(_09703_));
 sg13g2_nor2_2 _15673_ (.A(net5831),
    .B(_09703_),
    .Y(_09704_));
 sg13g2_nand2_2 _15674_ (.Y(_09705_),
    .A(_09700_),
    .B(_09704_));
 sg13g2_or2_1 _15675_ (.X(_09706_),
    .B(_09705_),
    .A(_09697_));
 sg13g2_o21ai_1 _15676_ (.B1(_09686_),
    .Y(_09707_),
    .A1(\fpga_top.io_frc.frc_cntr_val[24] ),
    .A2(_06871_));
 sg13g2_o21ai_1 _15677_ (.B1(_09682_),
    .Y(_09708_),
    .A1(net4922),
    .A2(_09707_));
 sg13g2_a21oi_1 _15678_ (.A1(net5430),
    .A2(_09708_),
    .Y(_09709_),
    .B1(net4930));
 sg13g2_a22oi_1 _15679_ (.Y(_09710_),
    .B1(_09681_),
    .B2(_09709_),
    .A2(net4930),
    .A1(_06805_));
 sg13g2_mux2_1 _15680_ (.A0(net4403),
    .A1(net2657),
    .S(net4208),
    .X(_00148_));
 sg13g2_and2_1 _15681_ (.A(net5707),
    .B(\fpga_top.qspi_if.word_data[1] ),
    .X(_09711_));
 sg13g2_nand2_1 _15682_ (.Y(_09712_),
    .A(net5702),
    .B(\fpga_top.qspi_if.word_data[1] ));
 sg13g2_a21oi_1 _15683_ (.A1(net5438),
    .A2(_09711_),
    .Y(_09713_),
    .B1(net4924));
 sg13g2_a21oi_1 _15684_ (.A1(net4474),
    .A2(_09713_),
    .Y(_09714_),
    .B1(net5431));
 sg13g2_o21ai_1 _15685_ (.B1(_09714_),
    .Y(_09715_),
    .A1(_08500_),
    .A2(net4475));
 sg13g2_nand2_1 _15686_ (.Y(_09716_),
    .A(\fpga_top.io_spi_lite.spi_mode[11] ),
    .B(net5838));
 sg13g2_nor2_1 _15687_ (.A(\fpga_top.io_uart_out.re_uart_rdflg_dly[3] ),
    .B(net5715),
    .Y(_09717_));
 sg13g2_nor2_1 _15688_ (.A(\fpga_top.io_uart_out.re_uart_rdflg_dly[1] ),
    .B(net5717),
    .Y(_09718_));
 sg13g2_nor4_1 _15689_ (.A(\fpga_top.io_uart_out.re_uart_rdflg_dly[1] ),
    .B(net5717),
    .C(\fpga_top.io_led.re_led_value_dly ),
    .D(\fpga_top.io_frc.re_frc_dly[4] ),
    .Y(_09719_));
 sg13g2_or2_1 _15690_ (.X(_09720_),
    .B(\fpga_top.io_led.re_gpio_value_dly[2] ),
    .A(\fpga_top.io_led.re_gpio_value_dly[3] ));
 sg13g2_nor3_1 _15691_ (.A(\fpga_top.io_led.re_gpio_value_dly[1] ),
    .B(net5710),
    .C(_09720_),
    .Y(_09721_));
 sg13g2_nand4_1 _15692_ (.B(_09717_),
    .C(_09719_),
    .A(_06867_),
    .Y(_09722_),
    .D(_09721_));
 sg13g2_a21oi_2 _15693_ (.B1(net5728),
    .Y(_09723_),
    .A2(_09722_),
    .A1(net5357));
 sg13g2_o21ai_1 _15694_ (.B1(net5068),
    .Y(_09724_),
    .A1(\fpga_top.io_frc.frc_cmp_val[57] ),
    .A2(net5356));
 sg13g2_a21oi_1 _15695_ (.A1(\fpga_top.io_frc.frc_cmp_val[25] ),
    .A2(net5728),
    .Y(_09725_),
    .B1(net5738));
 sg13g2_a22oi_1 _15696_ (.Y(_09726_),
    .B1(_09724_),
    .B2(_09725_),
    .A2(net5738),
    .A1(_06739_));
 sg13g2_a21oi_1 _15697_ (.A1(_06719_),
    .A2(net5752),
    .Y(_09727_),
    .B1(net4922));
 sg13g2_o21ai_1 _15698_ (.B1(_09727_),
    .Y(_09728_),
    .A1(net5750),
    .A2(_09726_));
 sg13g2_nand2_2 _15699_ (.Y(_09729_),
    .A(_09716_),
    .B(_09728_));
 sg13g2_a21oi_1 _15700_ (.A1(net5431),
    .A2(_09729_),
    .Y(_09730_),
    .B1(net4928));
 sg13g2_a22oi_1 _15701_ (.Y(_09731_),
    .B1(_09715_),
    .B2(_09730_),
    .A2(net4928),
    .A1(_06806_));
 sg13g2_mux2_1 _15702_ (.A0(net4400),
    .A1(net2433),
    .S(net4207),
    .X(_00149_));
 sg13g2_and2_1 _15703_ (.A(net5701),
    .B(\fpga_top.qspi_if.word_data[2] ),
    .X(_09732_));
 sg13g2_a21oi_1 _15704_ (.A1(net5439),
    .A2(_09732_),
    .Y(_09733_),
    .B1(net4925));
 sg13g2_o21ai_1 _15705_ (.B1(_06925_),
    .Y(_09734_),
    .A1(_08598_),
    .A2(net4474));
 sg13g2_a21o_1 _15706_ (.A2(_09733_),
    .A1(net4477),
    .B1(_09734_),
    .X(_09735_));
 sg13g2_nand2_1 _15707_ (.Y(_09736_),
    .A(\fpga_top.io_spi_lite.spi_mode[12] ),
    .B(net5838));
 sg13g2_o21ai_1 _15708_ (.B1(net5068),
    .Y(_09737_),
    .A1(\fpga_top.io_frc.frc_cmp_val[58] ),
    .A2(net5357));
 sg13g2_a21oi_1 _15709_ (.A1(\fpga_top.io_frc.frc_cmp_val[26] ),
    .A2(net5729),
    .Y(_09738_),
    .B1(net5741));
 sg13g2_a22oi_1 _15710_ (.Y(_09739_),
    .B1(_09737_),
    .B2(_09738_),
    .A2(net5738),
    .A1(_06738_));
 sg13g2_a21oi_1 _15711_ (.A1(_06718_),
    .A2(net5752),
    .Y(_09740_),
    .B1(net4922));
 sg13g2_o21ai_1 _15712_ (.B1(_09740_),
    .Y(_09741_),
    .A1(net5752),
    .A2(_09739_));
 sg13g2_nand2_2 _15713_ (.Y(_09742_),
    .A(_09736_),
    .B(_09741_));
 sg13g2_a21oi_1 _15714_ (.A1(net5432),
    .A2(_09742_),
    .Y(_09743_),
    .B1(net4931));
 sg13g2_a22oi_1 _15715_ (.Y(_09744_),
    .B1(_09735_),
    .B2(_09743_),
    .A2(net4931),
    .A1(_06807_));
 sg13g2_mux2_1 _15716_ (.A0(net4397),
    .A1(net2942),
    .S(net4206),
    .X(_00150_));
 sg13g2_nand2_1 _15717_ (.Y(_09745_),
    .A(_08452_),
    .B(net4483));
 sg13g2_and2_1 _15718_ (.A(net5705),
    .B(\fpga_top.qspi_if.word_data[3] ),
    .X(_09746_));
 sg13g2_a21o_1 _15719_ (.A2(_09746_),
    .A1(net5438),
    .B1(net4924),
    .X(_09747_));
 sg13g2_a21oi_1 _15720_ (.A1(net4478),
    .A2(_09747_),
    .Y(_09748_),
    .B1(net5435));
 sg13g2_nand2b_1 _15721_ (.Y(_09749_),
    .B(net5720),
    .A_N(\fpga_top.io_frc.frc_cmp_val[59] ));
 sg13g2_a22oi_1 _15722_ (.Y(_09750_),
    .B1(net5068),
    .B2(_09749_),
    .A2(net5728),
    .A1(\fpga_top.io_frc.frc_cmp_val[27] ));
 sg13g2_a21oi_1 _15723_ (.A1(\fpga_top.io_frc.frc_cntr_val[59] ),
    .A2(net5739),
    .Y(_09751_),
    .B1(net5750));
 sg13g2_o21ai_1 _15724_ (.B1(_09751_),
    .Y(_09752_),
    .A1(net5739),
    .A2(_09750_));
 sg13g2_a21oi_1 _15725_ (.A1(_06717_),
    .A2(net5749),
    .Y(_09753_),
    .B1(net4922));
 sg13g2_nand2_2 _15726_ (.Y(_09754_),
    .A(_09752_),
    .B(_09753_));
 sg13g2_a221oi_1 _15727_ (.B2(net5435),
    .C1(net4933),
    .B1(_09754_),
    .A1(_09745_),
    .Y(_09755_),
    .A2(_09748_));
 sg13g2_a21o_2 _15728_ (.A2(net4936),
    .A1(net5640),
    .B1(_09755_),
    .X(_09756_));
 sg13g2_mux2_1 _15729_ (.A0(net4388),
    .A1(net2757),
    .S(net4205),
    .X(_00151_));
 sg13g2_and2_1 _15730_ (.A(net5706),
    .B(net3288),
    .X(_09757_));
 sg13g2_a21oi_1 _15731_ (.A1(net5438),
    .A2(_09757_),
    .Y(_09758_),
    .B1(net4924));
 sg13g2_o21ai_1 _15732_ (.B1(_06925_),
    .Y(_09759_),
    .A1(_08574_),
    .A2(net4474));
 sg13g2_a21o_1 _15733_ (.A2(_09758_),
    .A1(net4474),
    .B1(_09759_),
    .X(_09760_));
 sg13g2_o21ai_1 _15734_ (.B1(_09723_),
    .Y(_09761_),
    .A1(\fpga_top.io_frc.frc_cmp_val[60] ),
    .A2(net5357));
 sg13g2_a21oi_1 _15735_ (.A1(\fpga_top.io_frc.frc_cmp_val[28] ),
    .A2(net5729),
    .Y(_09762_),
    .B1(net5741));
 sg13g2_a221oi_1 _15736_ (.B2(_09762_),
    .C1(net5749),
    .B1(_09761_),
    .A1(_06737_),
    .Y(_09763_),
    .A2(net5738));
 sg13g2_a21oi_1 _15737_ (.A1(\fpga_top.io_frc.frc_cntr_val[28] ),
    .A2(net5749),
    .Y(_09764_),
    .B1(_09763_));
 sg13g2_nor2_2 _15738_ (.A(net4922),
    .B(_09764_),
    .Y(_09765_));
 sg13g2_a21oi_1 _15739_ (.A1(net5431),
    .A2(_09765_),
    .Y(_09766_),
    .B1(net4931));
 sg13g2_a22oi_1 _15740_ (.Y(_09767_),
    .B1(_09760_),
    .B2(_09766_),
    .A2(net4931),
    .A1(_06808_));
 sg13g2_mux2_1 _15741_ (.A0(net4384),
    .A1(net3244),
    .S(net4206),
    .X(_00152_));
 sg13g2_nand2_1 _15742_ (.Y(_09768_),
    .A(_07798_),
    .B(net4483));
 sg13g2_and2_1 _15743_ (.A(net5703),
    .B(net2095),
    .X(_09769_));
 sg13g2_a21oi_1 _15744_ (.A1(net5438),
    .A2(_09769_),
    .Y(_09770_),
    .B1(_09677_));
 sg13g2_a21oi_1 _15745_ (.A1(net4480),
    .A2(_09770_),
    .Y(_09771_),
    .B1(net5436));
 sg13g2_nor2b_1 _15746_ (.A(\fpga_top.io_frc.frc_cmp_val[29] ),
    .B_N(net5729),
    .Y(_09772_));
 sg13g2_a21oi_1 _15747_ (.A1(\fpga_top.io_frc.frc_cmp_val[61] ),
    .A2(net5720),
    .Y(_09773_),
    .B1(net5728));
 sg13g2_or3_1 _15748_ (.A(net5738),
    .B(_09772_),
    .C(_09773_),
    .X(_09774_));
 sg13g2_a21oi_1 _15749_ (.A1(\fpga_top.io_frc.frc_cntr_val[61] ),
    .A2(net5738),
    .Y(_09775_),
    .B1(net5749));
 sg13g2_a221oi_1 _15750_ (.B2(_09775_),
    .C1(net4922),
    .B1(_09774_),
    .A1(_06714_),
    .Y(_09776_),
    .A2(net5749));
 sg13g2_a221oi_1 _15751_ (.B2(net5436),
    .C1(net4934),
    .B1(_09776_),
    .A1(_09768_),
    .Y(_09777_),
    .A2(_09771_));
 sg13g2_a21oi_2 _15752_ (.B1(_09777_),
    .Y(_09778_),
    .A2(net4934),
    .A1(_06809_));
 sg13g2_mux2_1 _15753_ (.A0(net4378),
    .A1(net3185),
    .S(net4208),
    .X(_00153_));
 sg13g2_nand2_1 _15754_ (.Y(_09779_),
    .A(net5707),
    .B(net3879));
 sg13g2_nand3_1 _15755_ (.B(\fpga_top.qspi_if.word_data[6] ),
    .C(net5438),
    .A(net5707),
    .Y(_09780_));
 sg13g2_nand3b_1 _15756_ (.B(_09780_),
    .C(net4480),
    .Y(_09781_),
    .A_N(_09677_));
 sg13g2_a21oi_1 _15757_ (.A1(_07750_),
    .A2(net4483),
    .Y(_09782_),
    .B1(net5435));
 sg13g2_o21ai_1 _15758_ (.B1(_09723_),
    .Y(_09783_),
    .A1(\fpga_top.io_frc.frc_cmp_val[62] ),
    .A2(net5357));
 sg13g2_a21oi_1 _15759_ (.A1(\fpga_top.io_frc.frc_cmp_val[30] ),
    .A2(net5727),
    .Y(_09784_),
    .B1(net5739));
 sg13g2_a221oi_1 _15760_ (.B2(_09784_),
    .C1(net5750),
    .B1(_09783_),
    .A1(_06734_),
    .Y(_09785_),
    .A2(net5739));
 sg13g2_a21oi_1 _15761_ (.A1(\fpga_top.io_frc.frc_cntr_val[30] ),
    .A2(net5750),
    .Y(_09786_),
    .B1(_09785_));
 sg13g2_nor2_2 _15762_ (.A(net4922),
    .B(_09786_),
    .Y(_09787_));
 sg13g2_a221oi_1 _15763_ (.B2(net5435),
    .C1(net4932),
    .B1(_09787_),
    .A1(_09781_),
    .Y(_09788_),
    .A2(_09782_));
 sg13g2_a21oi_2 _15764_ (.B1(_09788_),
    .Y(_09789_),
    .A2(net4936),
    .A1(_06810_));
 sg13g2_mux2_1 _15765_ (.A0(net4372),
    .A1(net2227),
    .S(net4207),
    .X(_00154_));
 sg13g2_nand2_1 _15766_ (.Y(_09790_),
    .A(net5707),
    .B(net3790));
 sg13g2_nand3_1 _15767_ (.B(\fpga_top.qspi_if.word_data[7] ),
    .C(net5439),
    .A(net5707),
    .Y(_09791_));
 sg13g2_nand3b_1 _15768_ (.B(_09791_),
    .C(net4476),
    .Y(_09792_),
    .A_N(net4924));
 sg13g2_o21ai_1 _15769_ (.B1(_06925_),
    .Y(_09793_),
    .A1(_07675_),
    .A2(net4474));
 sg13g2_nand2b_1 _15770_ (.Y(_09794_),
    .B(_09792_),
    .A_N(_09793_));
 sg13g2_o21ai_1 _15771_ (.B1(_09723_),
    .Y(_09795_),
    .A1(\fpga_top.io_frc.frc_cmp_val[63] ),
    .A2(net5357));
 sg13g2_a21oi_1 _15772_ (.A1(\fpga_top.io_frc.frc_cmp_val[31] ),
    .A2(net5729),
    .Y(_09796_),
    .B1(net5741));
 sg13g2_a221oi_1 _15773_ (.B2(_09796_),
    .C1(net5749),
    .B1(_09795_),
    .A1(_06733_),
    .Y(_09797_),
    .A2(net5738));
 sg13g2_a21oi_1 _15774_ (.A1(\fpga_top.io_frc.frc_cntr_val[31] ),
    .A2(net5749),
    .Y(_09798_),
    .B1(_09797_));
 sg13g2_nor2_2 _15775_ (.A(net4922),
    .B(_09798_),
    .Y(_09799_));
 sg13g2_a21oi_1 _15776_ (.A1(net5431),
    .A2(_09799_),
    .Y(_09800_),
    .B1(net4928));
 sg13g2_a22oi_1 _15777_ (.Y(_09801_),
    .B1(_09794_),
    .B2(_09800_),
    .A2(net4933),
    .A1(_06811_));
 sg13g2_mux2_1 _15778_ (.A0(net4368),
    .A1(net2865),
    .S(net4208),
    .X(_00155_));
 sg13g2_nor2_1 _15779_ (.A(_09661_),
    .B(_09664_),
    .Y(_09802_));
 sg13g2_nand2_1 _15780_ (.Y(_09803_),
    .A(_09666_),
    .B(_09802_));
 sg13g2_a221oi_1 _15781_ (.B2(\fpga_top.cpu_top.csr_wadr_mon[0] ),
    .C1(_09653_),
    .B1(net4936),
    .A1(_09649_),
    .Y(_09804_),
    .A2(_09650_));
 sg13g2_nand2_2 _15782_ (.Y(_09805_),
    .A(_09657_),
    .B(_09804_));
 sg13g2_or2_1 _15783_ (.X(_09806_),
    .B(_09805_),
    .A(_09803_));
 sg13g2_and2_1 _15784_ (.A(net5708),
    .B(\fpga_top.qspi_if.word_data[24] ),
    .X(_09807_));
 sg13g2_a221oi_1 _15785_ (.B2(\fpga_top.qspi_if.word_data[0] ),
    .C1(_09807_),
    .B1(net5330),
    .A1(\fpga_top.qspi_if.word_data[8] ),
    .Y(_09808_),
    .A2(net5335));
 sg13g2_inv_1 _15786_ (.Y(_09809_),
    .A(_09808_));
 sg13g2_nand2_1 _15787_ (.Y(_09810_),
    .A(net4476),
    .B(_09808_));
 sg13g2_mux4_1 _15788_ (.S0(net4995),
    .A0(net5820),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[0] ),
    .A2(net5816),
    .A3(net5823),
    .S1(net4976),
    .X(_09811_));
 sg13g2_nand2_1 _15789_ (.Y(_09812_),
    .A(net5003),
    .B(_09811_));
 sg13g2_a21oi_1 _15790_ (.A1(net5013),
    .A2(_08201_),
    .Y(_09813_),
    .B1(net4974));
 sg13g2_nand2_1 _15791_ (.Y(_09814_),
    .A(_09812_),
    .B(_09813_));
 sg13g2_o21ai_1 _15792_ (.B1(_09814_),
    .Y(_09815_),
    .A1(net4955),
    .A2(_08108_));
 sg13g2_o21ai_1 _15793_ (.B1(_07603_),
    .Y(_09816_),
    .A1(net4856),
    .A2(_08019_));
 sg13g2_a21oi_1 _15794_ (.A1(net4856),
    .A2(_09815_),
    .Y(_09817_),
    .B1(_09816_));
 sg13g2_nor3_1 _15795_ (.A(net4965),
    .B(net4784),
    .C(_07888_),
    .Y(_09818_));
 sg13g2_nand3_1 _15796_ (.B(net4977),
    .C(net5187),
    .A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[0] ),
    .Y(_09819_));
 sg13g2_o21ai_1 _15797_ (.B1(net5100),
    .Y(_09820_),
    .A1(\fpga_top.cpu_top.execution.csr_array.rs1_sel[0] ),
    .A2(net4977));
 sg13g2_o21ai_1 _15798_ (.B1(net5183),
    .Y(_09821_),
    .A1(_07395_),
    .A2(_07705_));
 sg13g2_nand4_1 _15799_ (.B(_09819_),
    .C(_09820_),
    .A(net5199),
    .Y(_09822_),
    .D(_09821_));
 sg13g2_or2_1 _15800_ (.X(_09823_),
    .B(_07718_),
    .A(_07570_));
 sg13g2_or2_1 _15801_ (.X(_09824_),
    .B(_07549_),
    .A(_06580_));
 sg13g2_nor2b_1 _15802_ (.A(_08484_),
    .B_N(net5770),
    .Y(_09825_));
 sg13g2_a22oi_1 _15803_ (.Y(_09826_),
    .B1(_07538_),
    .B2(_09825_),
    .A2(_07527_),
    .A1(net5767));
 sg13g2_nor2_1 _15804_ (.A(_08583_),
    .B(_09826_),
    .Y(_09827_));
 sg13g2_a21oi_1 _15805_ (.A1(net5765),
    .A2(_07533_),
    .Y(_09828_),
    .B1(_09827_));
 sg13g2_nor2_1 _15806_ (.A(_08440_),
    .B(_09828_),
    .Y(_09829_));
 sg13g2_a21oi_1 _15807_ (.A1(net5761),
    .A2(_07555_),
    .Y(_09830_),
    .B1(_09829_));
 sg13g2_or2_1 _15808_ (.X(_09831_),
    .B(_09830_),
    .A(_08563_));
 sg13g2_a21oi_1 _15809_ (.A1(_09824_),
    .A2(_09831_),
    .Y(_09832_),
    .B1(_07776_));
 sg13g2_a21oi_1 _15810_ (.A1(net5757),
    .A2(_07318_),
    .Y(_09833_),
    .B1(_09832_));
 sg13g2_nor3_1 _15811_ (.A(_08484_),
    .B(_08563_),
    .C(_08583_),
    .Y(_09834_));
 sg13g2_nor3_1 _15812_ (.A(_07776_),
    .B(_08440_),
    .C(_09823_),
    .Y(_09835_));
 sg13g2_nand3_1 _15813_ (.B(_09834_),
    .C(_09835_),
    .A(_07894_),
    .Y(_09836_));
 sg13g2_or2_1 _15814_ (.X(_09837_),
    .B(_08461_),
    .A(_07819_));
 sg13g2_nor2_1 _15815_ (.A(_07852_),
    .B(_08411_),
    .Y(_09838_));
 sg13g2_nand2_1 _15816_ (.Y(_09839_),
    .A(net5778),
    .B(_07331_));
 sg13g2_nand2_1 _15817_ (.Y(_09840_),
    .A(net5783),
    .B(_07494_));
 sg13g2_nand3_1 _15818_ (.B(_07505_),
    .C(_08359_),
    .A(net5786),
    .Y(_09841_));
 sg13g2_a21oi_1 _15819_ (.A1(_09840_),
    .A2(_09841_),
    .Y(_09842_),
    .B1(_08513_));
 sg13g2_a21oi_1 _15820_ (.A1(net5781),
    .A2(_07499_),
    .Y(_09843_),
    .B1(_09842_));
 sg13g2_o21ai_1 _15821_ (.B1(_09839_),
    .Y(_09844_),
    .A1(_08391_),
    .A2(_09843_));
 sg13g2_nor3_1 _15822_ (.A(_06578_),
    .B(_07335_),
    .C(_07852_),
    .Y(_09845_));
 sg13g2_a221oi_1 _15823_ (.B2(_09844_),
    .C1(_09845_),
    .B1(_09838_),
    .A1(net5775),
    .Y(_09846_),
    .A2(_07322_));
 sg13g2_nor3_1 _15824_ (.A(_06579_),
    .B(_07326_),
    .C(_08461_),
    .Y(_09847_));
 sg13g2_a21oi_1 _15825_ (.A1(net5771),
    .A2(_07520_),
    .Y(_09848_),
    .B1(_09847_));
 sg13g2_o21ai_1 _15826_ (.B1(_09848_),
    .Y(_09849_),
    .A1(_09837_),
    .A2(_09846_));
 sg13g2_nor2b_1 _15827_ (.A(_09836_),
    .B_N(_09849_),
    .Y(_09850_));
 sg13g2_nand2b_1 _15828_ (.Y(_09851_),
    .B(_08359_),
    .A_N(_08024_));
 sg13g2_or4_1 _15829_ (.A(_08391_),
    .B(_08513_),
    .C(_09837_),
    .D(_09851_),
    .X(_09852_));
 sg13g2_nor4_2 _15830_ (.A(_07852_),
    .B(_08411_),
    .C(_09836_),
    .Y(_09853_),
    .D(_09852_));
 sg13g2_or2_1 _15831_ (.X(_09854_),
    .B(_08538_),
    .A(_07929_));
 sg13g2_or3_1 _15832_ (.A(_07956_),
    .B(_08334_),
    .C(_09854_),
    .X(_09855_));
 sg13g2_or2_1 _15833_ (.X(_09856_),
    .B(_08265_),
    .A(_07988_));
 sg13g2_nor4_1 _15834_ (.A(_08114_),
    .B(_08300_),
    .C(_09855_),
    .D(_09856_),
    .Y(_09857_));
 sg13g2_nor2_1 _15835_ (.A(_08059_),
    .B(_08234_),
    .Y(_09858_));
 sg13g2_or2_1 _15836_ (.X(_09859_),
    .B(_08234_),
    .A(_08059_));
 sg13g2_and2_1 _15837_ (.A(_08148_),
    .B(_08176_),
    .X(_09860_));
 sg13g2_and3_1 _15838_ (.X(_09861_),
    .A(net5819),
    .B(net5004),
    .C(_08176_));
 sg13g2_nand3b_1 _15839_ (.B(net4860),
    .C(net5814),
    .Y(_09862_),
    .A_N(_08090_));
 sg13g2_o21ai_1 _15840_ (.B1(_09862_),
    .Y(_09863_),
    .A1(_06565_),
    .A2(_07423_));
 sg13g2_nand2_1 _15841_ (.Y(_09864_),
    .A(net5807),
    .B(_07417_));
 sg13g2_a22oi_1 _15842_ (.Y(_09865_),
    .B1(_09858_),
    .B2(_09863_),
    .A2(_07469_),
    .A1(net5806));
 sg13g2_o21ai_1 _15843_ (.B1(_09865_),
    .Y(_09866_),
    .A1(_08059_),
    .A2(_09864_));
 sg13g2_xnor2_1 _15844_ (.Y(_09867_),
    .A(net5822),
    .B(net4997));
 sg13g2_nor2_1 _15845_ (.A(_07395_),
    .B(_09867_),
    .Y(_09868_));
 sg13g2_nand2_1 _15846_ (.Y(_09869_),
    .A(_09860_),
    .B(_09868_));
 sg13g2_nor4_1 _15847_ (.A(_08090_),
    .B(_08209_),
    .C(_09859_),
    .D(_09869_),
    .Y(_09870_));
 sg13g2_a21o_1 _15848_ (.A2(net4997),
    .A1(net5822),
    .B1(_09868_),
    .X(_09871_));
 sg13g2_a221oi_1 _15849_ (.B2(_09871_),
    .C1(_09861_),
    .B1(_09860_),
    .A1(net5817),
    .Y(_09872_),
    .A2(net4963));
 sg13g2_nor4_1 _15850_ (.A(_08090_),
    .B(_08209_),
    .C(_09859_),
    .D(_09872_),
    .Y(_09873_));
 sg13g2_o21ai_1 _15851_ (.B1(_09857_),
    .Y(_09874_),
    .A1(_09866_),
    .A2(_09873_));
 sg13g2_nor2b_1 _15852_ (.A(_07956_),
    .B_N(net5795),
    .Y(_09875_));
 sg13g2_a22oi_1 _15853_ (.Y(_09876_),
    .B1(_07363_),
    .B2(_09875_),
    .A2(_07347_),
    .A1(net5791));
 sg13g2_nor3_1 _15854_ (.A(_06573_),
    .B(_07353_),
    .C(_08538_),
    .Y(_09877_));
 sg13g2_a21oi_1 _15855_ (.A1(net5787),
    .A2(_07488_),
    .Y(_09878_),
    .B1(_09877_));
 sg13g2_o21ai_1 _15856_ (.B1(_09878_),
    .Y(_09879_),
    .A1(_09854_),
    .A2(_09876_));
 sg13g2_nand3_1 _15857_ (.B(_07436_),
    .C(_07437_),
    .A(net5800),
    .Y(_09880_));
 sg13g2_nand3b_1 _15858_ (.B(_07461_),
    .C(net5803),
    .Y(_09881_),
    .A_N(_08300_));
 sg13g2_a21oi_1 _15859_ (.A1(_09880_),
    .A2(_09881_),
    .Y(_09882_),
    .B1(_09856_));
 sg13g2_nor3_1 _15860_ (.A(_06571_),
    .B(_07449_),
    .C(_08265_),
    .Y(_09883_));
 sg13g2_nor2_1 _15861_ (.A(_06572_),
    .B(_07359_),
    .Y(_09884_));
 sg13g2_nor3_1 _15862_ (.A(_09882_),
    .B(_09883_),
    .C(_09884_),
    .Y(_09885_));
 sg13g2_o21ai_1 _15863_ (.B1(_09874_),
    .Y(_09886_),
    .A1(_09855_),
    .A2(_09885_));
 sg13g2_o21ai_1 _15864_ (.B1(_09853_),
    .Y(_09887_),
    .A1(_09879_),
    .A2(_09886_));
 sg13g2_nor3_1 _15865_ (.A(_06581_),
    .B(_07311_),
    .C(_07570_),
    .Y(_09888_));
 sg13g2_nor2_1 _15866_ (.A(_09850_),
    .B(_09888_),
    .Y(_09889_));
 sg13g2_o21ai_1 _15867_ (.B1(_09889_),
    .Y(_09890_),
    .A1(_09823_),
    .A2(_09833_));
 sg13g2_nand2b_1 _15868_ (.Y(_09891_),
    .B(_09887_),
    .A_N(_09890_));
 sg13g2_a21oi_1 _15869_ (.A1(_06582_),
    .A2(_07569_),
    .Y(_09892_),
    .B1(_09891_));
 sg13g2_a21o_1 _15870_ (.A2(_07568_),
    .A1(net5754),
    .B1(_09891_),
    .X(_09893_));
 sg13g2_nor3_1 _15871_ (.A(net5382),
    .B(_06552_),
    .C(_09893_),
    .Y(_09894_));
 sg13g2_a21oi_1 _15872_ (.A1(_07606_),
    .A2(_09892_),
    .Y(_09895_),
    .B1(_09894_));
 sg13g2_nor2b_1 _15873_ (.A(_09895_),
    .B_N(_07579_),
    .Y(_09896_));
 sg13g2_nor4_1 _15874_ (.A(_09817_),
    .B(_09818_),
    .C(_09822_),
    .D(_09896_),
    .Y(_09897_));
 sg13g2_nor3_1 _15875_ (.A(_07395_),
    .B(net5198),
    .C(_07705_),
    .Y(_09898_));
 sg13g2_o21ai_1 _15876_ (.B1(net5193),
    .Y(_09899_),
    .A1(_09897_),
    .A2(_09898_));
 sg13g2_nor2_1 _15877_ (.A(net5308),
    .B(_08276_),
    .Y(_09900_));
 sg13g2_o21ai_1 _15878_ (.B1(_09900_),
    .Y(_09901_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[0] ),
    .A2(net5193));
 sg13g2_nand2b_2 _15879_ (.Y(_09902_),
    .B(_09899_),
    .A_N(_09901_));
 sg13g2_a21oi_1 _15880_ (.A1(net4484),
    .A2(_09902_),
    .Y(_09903_),
    .B1(net5429));
 sg13g2_nand2_1 _15881_ (.Y(_09904_),
    .A(\fpga_top.io_uart_out.re_uart_rdflg_dly[4] ),
    .B(_09717_));
 sg13g2_nand2_2 _15882_ (.Y(_09905_),
    .A(net5426),
    .B(\fpga_top.io_uart_out.rx_disable_echoback_value ));
 sg13g2_nand3_1 _15883_ (.B(_09717_),
    .C(_09905_),
    .A(\fpga_top.io_uart_out.re_uart_rdflg_dly[4] ),
    .Y(_09906_));
 sg13g2_nor2b_2 _15884_ (.A(net5715),
    .B_N(\fpga_top.io_uart_out.re_uart_rdflg_dly[3] ),
    .Y(_09907_));
 sg13g2_nand2b_2 _15885_ (.Y(_09908_),
    .B(\fpga_top.io_uart_out.re_uart_rdflg_dly[3] ),
    .A_N(net5715));
 sg13g2_a221oi_1 _15886_ (.B2(_06866_),
    .C1(\fpga_top.io_uart_out.re_uart_rdflg_dly[1] ),
    .B1(_09907_),
    .A1(_06831_),
    .Y(_09909_),
    .A2(net5715));
 sg13g2_a221oi_1 _15887_ (.B2(_09909_),
    .C1(net5717),
    .B1(_09906_),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[3] ),
    .Y(_09910_),
    .A2(\fpga_top.io_uart_out.re_uart_rdflg_dly[1] ));
 sg13g2_nor2b_1 _15888_ (.A(\fpga_top.io_uart_out.uart_io_char[0] ),
    .B_N(\fpga_top.io_uart_out.re_uart_rdflg_dly[0] ),
    .Y(_09911_));
 sg13g2_nor3_1 _15889_ (.A(_09720_),
    .B(_09910_),
    .C(_09911_),
    .Y(_09912_));
 sg13g2_nand2b_2 _15890_ (.Y(_09913_),
    .B(\fpga_top.io_led.re_gpio_value_dly[3] ),
    .A_N(\fpga_top.io_led.re_gpio_value_dly[2] ));
 sg13g2_nand2_1 _15891_ (.Y(_09914_),
    .A(\fpga_top.io_led.gpio_in_lat2[0] ),
    .B(\fpga_top.io_led.re_gpio_value_dly[2] ));
 sg13g2_o21ai_1 _15892_ (.B1(_09914_),
    .Y(_09915_),
    .A1(_06865_),
    .A2(_09913_));
 sg13g2_nor4_1 _15893_ (.A(\fpga_top.io_led.re_gpio_value_dly[1] ),
    .B(net5710),
    .C(_09912_),
    .D(_09915_),
    .Y(_09916_));
 sg13g2_nor2_1 _15894_ (.A(\fpga_top.io_led.gpi_init_lat2[0] ),
    .B(_06869_),
    .Y(_09917_));
 sg13g2_a21oi_1 _15895_ (.A1(\fpga_top.io_frc.frc_cntrl_val ),
    .A2(\fpga_top.io_frc.re_frc_dly[4] ),
    .Y(_09918_),
    .B1(net5719));
 sg13g2_nor3_1 _15896_ (.A(uio_out[4]),
    .B(_06868_),
    .C(net5710),
    .Y(_09919_));
 sg13g2_nor4_1 _15897_ (.A(\fpga_top.io_led.re_led_value_dly ),
    .B(_09916_),
    .C(_09917_),
    .D(_09919_),
    .Y(_09920_));
 sg13g2_a21oi_1 _15898_ (.A1(\fpga_top.io_led.led_value[0] ),
    .A2(\fpga_top.io_led.re_led_value_dly ),
    .Y(_09921_),
    .B1(_09920_));
 sg13g2_o21ai_1 _15899_ (.B1(_09918_),
    .Y(_09922_),
    .A1(\fpga_top.io_frc.re_frc_dly[4] ),
    .A2(_09921_));
 sg13g2_a21oi_1 _15900_ (.A1(_06768_),
    .A2(net5719),
    .Y(_09923_),
    .B1(net5723));
 sg13g2_a221oi_1 _15901_ (.B2(_09923_),
    .C1(net5732),
    .B1(_09922_),
    .A1(\fpga_top.io_frc.frc_cmp_val[0] ),
    .Y(_09924_),
    .A2(net5723));
 sg13g2_a21o_1 _15902_ (.A2(net5734),
    .A1(_06767_),
    .B1(net5745),
    .X(_09925_));
 sg13g2_a21oi_1 _15903_ (.A1(\fpga_top.io_frc.frc_cntr_val[0] ),
    .A2(net5743),
    .Y(_09926_),
    .B1(\fpga_top.qspi_if.re_qspi_latency_dly[9] ));
 sg13g2_o21ai_1 _15904_ (.B1(_09926_),
    .Y(_09927_),
    .A1(_09924_),
    .A2(_09925_));
 sg13g2_a21oi_1 _15905_ (.A1(_06677_),
    .A2(\fpga_top.qspi_if.re_qspi_latency_dly[9] ),
    .Y(_09928_),
    .B1(net5689));
 sg13g2_a221oi_1 _15906_ (.B2(_09928_),
    .C1(_09688_),
    .B1(_09927_),
    .A1(\fpga_top.qspi_if.rdwrch[0] ),
    .Y(_09929_),
    .A2(net5689));
 sg13g2_nor2b_2 _15907_ (.A(net5691),
    .B_N(\fpga_top.qspi_if.re_qspi_latency_dly[7] ),
    .Y(_09930_));
 sg13g2_nand2b_1 _15908_ (.Y(_09931_),
    .B(_09930_),
    .A_N(\fpga_top.qspi_if.wrcmd1[0] ));
 sg13g2_nand2b_1 _15909_ (.Y(_09932_),
    .B(net5691),
    .A_N(\fpga_top.qspi_if.wrcmd0[0] ));
 sg13g2_nand3_1 _15910_ (.B(_09931_),
    .C(_09932_),
    .A(_09695_),
    .Y(_09933_));
 sg13g2_nor2_2 _15911_ (.A(net5694),
    .B(_09692_),
    .Y(_09934_));
 sg13g2_nor2b_1 _15912_ (.A(net5692),
    .B_N(_00102_),
    .Y(_09935_));
 sg13g2_a21oi_1 _15913_ (.A1(_00108_),
    .A2(net5692),
    .Y(_09936_),
    .B1(_09935_));
 sg13g2_a221oi_1 _15914_ (.B2(_09936_),
    .C1(net5698),
    .B1(_09934_),
    .A1(_06497_),
    .Y(_09937_),
    .A2(net5694));
 sg13g2_o21ai_1 _15915_ (.B1(_09937_),
    .Y(_09938_),
    .A1(_09929_),
    .A2(_09933_));
 sg13g2_a21oi_1 _15916_ (.A1(_06830_),
    .A2(net5698),
    .Y(_09939_),
    .B1(net5329));
 sg13g2_mux2_1 _15917_ (.A0(\fpga_top.qspi_if.read_latency_1[0] ),
    .A1(\fpga_top.qspi_if.read_latency_0[0] ),
    .S(\fpga_top.qspi_if.re_qspi_latency_dly[0] ),
    .X(_09940_));
 sg13g2_a221oi_1 _15918_ (.B2(net5329),
    .C1(_09701_),
    .B1(_09940_),
    .A1(_09938_),
    .Y(_09941_),
    .A2(_09939_));
 sg13g2_nand2b_1 _15919_ (.Y(_09942_),
    .B(\fpga_top.interrupter.re_int_dly[0] ),
    .A_N(\fpga_top.interrupter.int_enable_rx ));
 sg13g2_o21ai_1 _15920_ (.B1(_09942_),
    .Y(_09943_),
    .A1(\fpga_top.interrupter.int_status_rx ),
    .A2(\fpga_top.interrupter.re_int_dly[0] ));
 sg13g2_a21oi_1 _15921_ (.A1(_09701_),
    .A2(_09943_),
    .Y(_09944_),
    .B1(_09941_));
 sg13g2_mux2_1 _15922_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][0] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][0] ),
    .S(net5395),
    .X(_09945_));
 sg13g2_nand2b_1 _15923_ (.Y(_09946_),
    .B(net5395),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][0] ));
 sg13g2_o21ai_1 _15924_ (.B1(_09946_),
    .Y(_09947_),
    .A1(net5395),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][0] ));
 sg13g2_o21ai_1 _15925_ (.B1(_06874_),
    .Y(_09948_),
    .A1(net5388),
    .A2(_09945_));
 sg13g2_a21oi_1 _15926_ (.A1(net5390),
    .A2(_09947_),
    .Y(_09949_),
    .B1(_09948_));
 sg13g2_nand2b_1 _15927_ (.Y(_09950_),
    .B(net5395),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][0] ));
 sg13g2_o21ai_1 _15928_ (.B1(_09950_),
    .Y(_09951_),
    .A1(net5395),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][0] ));
 sg13g2_mux2_1 _15929_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][0] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][0] ),
    .S(net5395),
    .X(_09952_));
 sg13g2_o21ai_1 _15930_ (.B1(net5387),
    .Y(_09953_),
    .A1(net5388),
    .A2(_09952_));
 sg13g2_a21oi_1 _15931_ (.A1(net5390),
    .A2(_09951_),
    .Y(_09954_),
    .B1(_09953_));
 sg13g2_nor3_1 _15932_ (.A(_06788_),
    .B(_09949_),
    .C(_09954_),
    .Y(_09955_));
 sg13g2_nor2_1 _15933_ (.A(_09699_),
    .B(_09955_),
    .Y(_09956_));
 sg13g2_o21ai_1 _15934_ (.B1(_09956_),
    .Y(_09957_),
    .A1(net5831),
    .A2(_09944_));
 sg13g2_a21oi_2 _15935_ (.B1(net5837),
    .Y(_09958_),
    .A2(net5835),
    .A1(\fpga_top.io_spi_lite.spi_sck_div[0] ));
 sg13g2_a22oi_1 _15936_ (.Y(_09959_),
    .B1(_09957_),
    .B2(_09958_),
    .A2(net5838),
    .A1(_06875_));
 sg13g2_a221oi_1 _15937_ (.B2(net5430),
    .C1(net4930),
    .B1(_09959_),
    .A1(_09810_),
    .Y(_09960_),
    .A2(_09903_));
 sg13g2_a21oi_2 _15938_ (.B1(_09960_),
    .Y(_09961_),
    .A2(net4929),
    .A1(_06683_));
 sg13g2_mux2_1 _15939_ (.A0(net4364),
    .A1(net3339),
    .S(net4200),
    .X(_00156_));
 sg13g2_and2_1 _15940_ (.A(net5704),
    .B(net1858),
    .X(_09962_));
 sg13g2_a221oi_1 _15941_ (.B2(\fpga_top.qspi_if.word_data[1] ),
    .C1(_09962_),
    .B1(net5330),
    .A1(\fpga_top.qspi_if.word_data[9] ),
    .Y(_09963_),
    .A2(net5333));
 sg13g2_nand2_1 _15942_ (.Y(_09964_),
    .A(net4477),
    .B(_09963_));
 sg13g2_and2_1 _15943_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[1] ),
    .B(net5293),
    .X(_09965_));
 sg13g2_mux4_1 _15944_ (.S0(net4991),
    .A0(net5823),
    .A1(net5817),
    .A2(net5820),
    .A3(net5813),
    .S1(net4980),
    .X(_09966_));
 sg13g2_a21oi_1 _15945_ (.A1(net5014),
    .A2(_08080_),
    .Y(_09967_),
    .B1(net4974));
 sg13g2_o21ai_1 _15946_ (.B1(_09967_),
    .Y(_09968_),
    .A1(net5013),
    .A2(_09966_));
 sg13g2_a21oi_1 _15947_ (.A1(net4968),
    .A2(_08284_),
    .Y(_09969_),
    .B1(net4950));
 sg13g2_a21oi_1 _15948_ (.A1(_09968_),
    .A2(_09969_),
    .Y(_09970_),
    .B1(_07604_));
 sg13g2_o21ai_1 _15949_ (.B1(_09970_),
    .Y(_09971_),
    .A1(net4856),
    .A2(_08353_));
 sg13g2_nand3_1 _15950_ (.B(net4990),
    .C(net5288),
    .A(net5822),
    .Y(_09972_));
 sg13g2_o21ai_1 _15951_ (.B1(net5099),
    .Y(_09973_),
    .A1(net5822),
    .A2(net4990));
 sg13g2_nand3_1 _15952_ (.B(_09972_),
    .C(_09973_),
    .A(net5199),
    .Y(_09974_));
 sg13g2_a221oi_1 _15953_ (.B2(net5184),
    .C1(_09974_),
    .B1(_09867_),
    .A1(net4855),
    .Y(_09975_),
    .A2(_08364_));
 sg13g2_xnor2_1 _15954_ (.Y(_09976_),
    .A(_07392_),
    .B(_07397_));
 sg13g2_a221oi_1 _15955_ (.B2(net5197),
    .C1(net5293),
    .B1(_09976_),
    .A1(_09971_),
    .Y(_09977_),
    .A2(_09975_));
 sg13g2_o21ai_1 _15956_ (.B1(_09900_),
    .Y(_09978_),
    .A1(_09965_),
    .A2(_09977_));
 sg13g2_a21oi_1 _15957_ (.A1(net4484),
    .A2(_09978_),
    .Y(_09979_),
    .B1(net5432));
 sg13g2_mux2_1 _15958_ (.A0(_06500_),
    .A1(\fpga_top.qspi_if.rdwrch[1] ),
    .S(net5689),
    .X(_09980_));
 sg13g2_o21ai_1 _15959_ (.B1(_09687_),
    .Y(_09981_),
    .A1(_09689_),
    .A2(_09980_));
 sg13g2_nand2_2 _15960_ (.Y(_09982_),
    .A(_09718_),
    .B(_09904_));
 sg13g2_a21oi_1 _15961_ (.A1(_06832_),
    .A2(net5716),
    .Y(_09983_),
    .B1(_09982_));
 sg13g2_o21ai_1 _15962_ (.B1(_09983_),
    .Y(_09984_),
    .A1(\fpga_top.io_uart_out.rx_data_latch[1] ),
    .A2(_09908_));
 sg13g2_a21oi_1 _15963_ (.A1(\fpga_top.io_uart_out.uart_io_char[1] ),
    .A2(net5717),
    .Y(_09985_),
    .B1(_09720_));
 sg13g2_a22oi_1 _15964_ (.Y(_09986_),
    .B1(_09984_),
    .B2(_09985_),
    .A2(_06880_),
    .A1(\fpga_top.io_led.re_gpio_value_dly[2] ));
 sg13g2_o21ai_1 _15965_ (.B1(_09986_),
    .Y(_09987_),
    .A1(uio_oe[5]),
    .A2(_09913_));
 sg13g2_nand2_1 _15966_ (.Y(_09988_),
    .A(_06868_),
    .B(_09987_));
 sg13g2_a21oi_1 _15967_ (.A1(\fpga_top.io_led.re_gpio_value_dly[1] ),
    .A2(_06879_),
    .Y(_09989_),
    .B1(net5710));
 sg13g2_a221oi_1 _15968_ (.B2(_09989_),
    .C1(\fpga_top.io_led.re_led_value_dly ),
    .B1(_09988_),
    .A1(net5710),
    .Y(_09990_),
    .A2(\fpga_top.io_led.gpi_init_lat2[1] ));
 sg13g2_nor2b_1 _15969_ (.A(\fpga_top.io_led.led_value[1] ),
    .B_N(\fpga_top.io_led.re_led_value_dly ),
    .Y(_09991_));
 sg13g2_nor4_1 _15970_ (.A(\fpga_top.io_frc.re_frc_dly[4] ),
    .B(net5718),
    .C(_09990_),
    .D(_09991_),
    .Y(_09992_));
 sg13g2_a21oi_1 _15971_ (.A1(\fpga_top.io_frc.frc_cmp_val[33] ),
    .A2(net5719),
    .Y(_09993_),
    .B1(_09992_));
 sg13g2_a21oi_1 _15972_ (.A1(\fpga_top.io_frc.frc_cmp_val[1] ),
    .A2(net5722),
    .Y(_09994_),
    .B1(net5733));
 sg13g2_o21ai_1 _15973_ (.B1(_09994_),
    .Y(_09995_),
    .A1(net5723),
    .A2(_09993_));
 sg13g2_a21oi_1 _15974_ (.A1(_06765_),
    .A2(net5732),
    .Y(_09996_),
    .B1(net5744));
 sg13g2_a221oi_1 _15975_ (.B2(_09996_),
    .C1(_09690_),
    .B1(_09995_),
    .A1(\fpga_top.io_frc.frc_cntr_val[1] ),
    .Y(_09997_),
    .A2(net5743));
 sg13g2_nor2_1 _15976_ (.A(_09981_),
    .B(_09997_),
    .Y(_09998_));
 sg13g2_a221oi_1 _15977_ (.B2(\fpga_top.qspi_if.wrcmd1[1] ),
    .C1(_09998_),
    .B1(_09930_),
    .A1(\fpga_top.qspi_if.wrcmd0[1] ),
    .Y(_09999_),
    .A2(net5691));
 sg13g2_nand2_1 _15978_ (.Y(_10000_),
    .A(_09695_),
    .B(_09999_));
 sg13g2_mux2_1 _15979_ (.A0(_00103_),
    .A1(_00109_),
    .S(net5692),
    .X(_10001_));
 sg13g2_a221oi_1 _15980_ (.B2(_10001_),
    .C1(net5698),
    .B1(_09934_),
    .A1(_06650_),
    .Y(_10002_),
    .A2(net5695));
 sg13g2_a221oi_1 _15981_ (.B2(_10002_),
    .C1(net5329),
    .B1(_10000_),
    .A1(\fpga_top.qspi_if.read_latency_2[1] ),
    .Y(_10003_),
    .A2(net5698));
 sg13g2_nand2b_1 _15982_ (.Y(_10004_),
    .B(\fpga_top.qspi_if.re_qspi_latency_dly[0] ),
    .A_N(\fpga_top.qspi_if.read_latency_0[1] ));
 sg13g2_o21ai_1 _15983_ (.B1(_10004_),
    .Y(_10005_),
    .A1(\fpga_top.qspi_if.read_latency_1[1] ),
    .A2(\fpga_top.qspi_if.re_qspi_latency_dly[0] ));
 sg13g2_a21o_1 _15984_ (.A2(_10005_),
    .A1(net5329),
    .B1(_09701_),
    .X(_10006_));
 sg13g2_nand2_1 _15985_ (.Y(_10007_),
    .A(\fpga_top.interrupter.int_enable_int0 ),
    .B(\fpga_top.interrupter.re_int_dly[0] ));
 sg13g2_o21ai_1 _15986_ (.B1(_10007_),
    .Y(_10008_),
    .A1(_06776_),
    .A2(\fpga_top.interrupter.re_int_dly[0] ));
 sg13g2_a21oi_1 _15987_ (.A1(_09701_),
    .A2(_10008_),
    .Y(_10009_),
    .B1(net5832));
 sg13g2_o21ai_1 _15988_ (.B1(_10009_),
    .Y(_10010_),
    .A1(_10003_),
    .A2(_10006_));
 sg13g2_nand2b_1 _15989_ (.Y(_10011_),
    .B(net5396),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][1] ));
 sg13g2_o21ai_1 _15990_ (.B1(_10011_),
    .Y(_10012_),
    .A1(net5397),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][1] ));
 sg13g2_mux2_1 _15991_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][1] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][1] ),
    .S(net5396),
    .X(_10013_));
 sg13g2_a21oi_1 _15992_ (.A1(net5391),
    .A2(_10012_),
    .Y(_10014_),
    .B1(_00007_));
 sg13g2_o21ai_1 _15993_ (.B1(_10014_),
    .Y(_10015_),
    .A1(net5391),
    .A2(_10013_));
 sg13g2_nand2b_1 _15994_ (.Y(_10016_),
    .B(net5396),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][1] ));
 sg13g2_o21ai_1 _15995_ (.B1(_10016_),
    .Y(_10017_),
    .A1(net5396),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][1] ));
 sg13g2_mux2_1 _15996_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][1] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][1] ),
    .S(net5396),
    .X(_10018_));
 sg13g2_o21ai_1 _15997_ (.B1(_00007_),
    .Y(_10019_),
    .A1(_00006_),
    .A2(_10018_));
 sg13g2_a21o_1 _15998_ (.A2(_10017_),
    .A1(net5391),
    .B1(_10019_),
    .X(_10020_));
 sg13g2_nand3_1 _15999_ (.B(_10015_),
    .C(_10020_),
    .A(net5831),
    .Y(_10021_));
 sg13g2_nand3_1 _16000_ (.B(_10010_),
    .C(_10021_),
    .A(_09698_),
    .Y(_10022_));
 sg13g2_a21oi_1 _16001_ (.A1(\fpga_top.io_spi_lite.spi_sck_div[1] ),
    .A2(net5834),
    .Y(_10023_),
    .B1(net5836));
 sg13g2_a22oi_1 _16002_ (.Y(_10024_),
    .B1(_10022_),
    .B2(_10023_),
    .A2(net5836),
    .A1(_06649_));
 sg13g2_a221oi_1 _16003_ (.B2(net5432),
    .C1(net4931),
    .B1(_10024_),
    .A1(_09964_),
    .Y(_10025_),
    .A2(_09979_));
 sg13g2_a21oi_2 _16004_ (.B1(_10025_),
    .Y(_10026_),
    .A2(net4931),
    .A1(_06681_));
 sg13g2_mux2_1 _16005_ (.A0(net4358),
    .A1(net2412),
    .S(net4202),
    .X(_00157_));
 sg13g2_and2_1 _16006_ (.A(net5703),
    .B(net1715),
    .X(_10027_));
 sg13g2_a221oi_1 _16007_ (.B2(\fpga_top.qspi_if.word_data[2] ),
    .C1(_10027_),
    .B1(net5330),
    .A1(net1863),
    .Y(_10028_),
    .A2(net5334));
 sg13g2_a21oi_1 _16008_ (.A1(net4476),
    .A2(_10028_),
    .Y(_10029_),
    .B1(net5429));
 sg13g2_o21ai_1 _16009_ (.B1(_10029_),
    .Y(_10030_),
    .A1(_08159_),
    .A2(net4476));
 sg13g2_nor3_2 _16010_ (.A(\fpga_top.io_led.re_led_value_dly ),
    .B(\fpga_top.io_frc.re_frc_dly[4] ),
    .C(net5718),
    .Y(_10031_));
 sg13g2_nand2b_1 _16011_ (.Y(_10032_),
    .B(\fpga_top.io_led.led_value[2] ),
    .A_N(\fpga_top.io_frc.re_frc_dly[4] ));
 sg13g2_a21oi_1 _16012_ (.A1(\fpga_top.cpu_top.execution.csr_array.frc_cntr_val_leq ),
    .A2(\fpga_top.io_frc.re_frc_dly[4] ),
    .Y(_10033_),
    .B1(net5721));
 sg13g2_a21oi_1 _16013_ (.A1(_10032_),
    .A2(_10033_),
    .Y(_10034_),
    .B1(_10031_));
 sg13g2_nand2_1 _16014_ (.Y(_10035_),
    .A(_06833_),
    .B(net5716));
 sg13g2_o21ai_1 _16015_ (.B1(_10035_),
    .Y(_10036_),
    .A1(\fpga_top.io_uart_out.rx_data_latch[2] ),
    .A2(_09908_));
 sg13g2_a21oi_1 _16016_ (.A1(\fpga_top.io_uart_out.uart_io_char[2] ),
    .A2(\fpga_top.io_uart_out.re_uart_rdflg_dly[0] ),
    .Y(_10037_),
    .B1(_09720_));
 sg13g2_o21ai_1 _16017_ (.B1(_10037_),
    .Y(_10038_),
    .A1(_09982_),
    .A2(_10036_));
 sg13g2_nand2b_1 _16018_ (.Y(_10039_),
    .B(\fpga_top.io_led.re_gpio_value_dly[2] ),
    .A_N(\fpga_top.io_led.gpio_in_lat2[2] ));
 sg13g2_o21ai_1 _16019_ (.B1(_10039_),
    .Y(_10040_),
    .A1(uio_oe[6]),
    .A2(_09913_));
 sg13g2_nor2_1 _16020_ (.A(\fpga_top.io_led.re_gpio_value_dly[1] ),
    .B(_10040_),
    .Y(_10041_));
 sg13g2_a221oi_1 _16021_ (.B2(_10041_),
    .C1(net5710),
    .B1(_10038_),
    .A1(\fpga_top.io_led.re_gpio_value_dly[1] ),
    .Y(_10042_),
    .A2(uio_out[6]));
 sg13g2_nor2_1 _16022_ (.A(_06869_),
    .B(\fpga_top.io_led.gpi_init_lat2[2] ),
    .Y(_10043_));
 sg13g2_nor4_1 _16023_ (.A(\fpga_top.io_led.re_led_value_dly ),
    .B(\fpga_top.io_frc.re_frc_dly[4] ),
    .C(_10042_),
    .D(_10043_),
    .Y(_10044_));
 sg13g2_nand2b_1 _16024_ (.Y(_10045_),
    .B(net5718),
    .A_N(\fpga_top.io_frc.frc_cmp_val[34] ));
 sg13g2_o21ai_1 _16025_ (.B1(_10045_),
    .Y(_10046_),
    .A1(_10034_),
    .A2(_10044_));
 sg13g2_a21oi_1 _16026_ (.A1(\fpga_top.io_frc.frc_cmp_val[2] ),
    .A2(net5722),
    .Y(_10047_),
    .B1(net5733));
 sg13g2_o21ai_1 _16027_ (.B1(_10047_),
    .Y(_10048_),
    .A1(net5723),
    .A2(_10046_));
 sg13g2_a21oi_1 _16028_ (.A1(_06764_),
    .A2(net5732),
    .Y(_10049_),
    .B1(net5743));
 sg13g2_a221oi_1 _16029_ (.B2(_10049_),
    .C1(_09690_),
    .B1(_10048_),
    .A1(\fpga_top.io_frc.frc_cntr_val[2] ),
    .Y(_10050_),
    .A2(net5743));
 sg13g2_nand2_1 _16030_ (.Y(_10051_),
    .A(\fpga_top.qspi_if.rdwrch[2] ),
    .B(net5689));
 sg13g2_o21ai_1 _16031_ (.B1(_10051_),
    .Y(_10052_),
    .A1(_06676_),
    .A2(net5689));
 sg13g2_o21ai_1 _16032_ (.B1(_09687_),
    .Y(_10053_),
    .A1(_09689_),
    .A2(_10052_));
 sg13g2_a221oi_1 _16033_ (.B2(\fpga_top.qspi_if.wrcmd1[2] ),
    .C1(\fpga_top.qspi_if.re_qspi_latency_dly[5] ),
    .B1(_09930_),
    .A1(\fpga_top.qspi_if.wrcmd0[2] ),
    .Y(_10054_),
    .A2(\fpga_top.qspi_if.re_qspi_latency_dly[6] ));
 sg13g2_o21ai_1 _16034_ (.B1(_10054_),
    .Y(_10055_),
    .A1(_10050_),
    .A2(_10053_));
 sg13g2_a21oi_1 _16035_ (.A1(_06818_),
    .A2(\fpga_top.qspi_if.re_qspi_latency_dly[5] ),
    .Y(_10056_),
    .B1(net5693));
 sg13g2_a221oi_1 _16036_ (.B2(_10056_),
    .C1(net5694),
    .B1(_10055_),
    .A1(\fpga_top.qspi_if.rdcmd0[2] ),
    .Y(_10057_),
    .A2(net5693));
 sg13g2_nor2_1 _16037_ (.A(\fpga_top.qspi_if.sck_div[2] ),
    .B(_06873_),
    .Y(_10058_));
 sg13g2_or3_1 _16038_ (.A(net5698),
    .B(_10057_),
    .C(_10058_),
    .X(_10059_));
 sg13g2_a21oi_1 _16039_ (.A1(\fpga_top.qspi_if.read_latency_2[2] ),
    .A2(net5698),
    .Y(_10060_),
    .B1(net5329));
 sg13g2_nand2b_1 _16040_ (.Y(_10061_),
    .B(\fpga_top.qspi_if.re_qspi_latency_dly[0] ),
    .A_N(\fpga_top.qspi_if.read_latency_0[2] ));
 sg13g2_o21ai_1 _16041_ (.B1(_10061_),
    .Y(_10062_),
    .A1(\fpga_top.qspi_if.read_latency_1[2] ),
    .A2(\fpga_top.qspi_if.re_qspi_latency_dly[0] ));
 sg13g2_a221oi_1 _16042_ (.B2(net5329),
    .C1(_09701_),
    .B1(_10062_),
    .A1(_10059_),
    .Y(_10063_),
    .A2(_10060_));
 sg13g2_mux2_1 _16043_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][2] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][2] ),
    .S(net5392),
    .X(_10064_));
 sg13g2_nand2b_1 _16044_ (.Y(_10065_),
    .B(net5392),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][2] ));
 sg13g2_o21ai_1 _16045_ (.B1(_10065_),
    .Y(_10066_),
    .A1(net5392),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][2] ));
 sg13g2_o21ai_1 _16046_ (.B1(_06874_),
    .Y(_10067_),
    .A1(net5388),
    .A2(_10064_));
 sg13g2_a21oi_1 _16047_ (.A1(net5388),
    .A2(_10066_),
    .Y(_10068_),
    .B1(_10067_));
 sg13g2_nand2b_1 _16048_ (.Y(_10069_),
    .B(net5393),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][2] ));
 sg13g2_o21ai_1 _16049_ (.B1(_10069_),
    .Y(_10070_),
    .A1(net5393),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][2] ));
 sg13g2_mux2_1 _16050_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][2] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][2] ),
    .S(net5392),
    .X(_10071_));
 sg13g2_o21ai_1 _16051_ (.B1(net5387),
    .Y(_10072_),
    .A1(net5389),
    .A2(_10071_));
 sg13g2_a21oi_1 _16052_ (.A1(net5388),
    .A2(_10070_),
    .Y(_10073_),
    .B1(_10072_));
 sg13g2_nor3_1 _16053_ (.A(_06788_),
    .B(_10068_),
    .C(_10073_),
    .Y(_10074_));
 sg13g2_nor2_1 _16054_ (.A(_09699_),
    .B(_10074_),
    .Y(_10075_));
 sg13g2_o21ai_1 _16055_ (.B1(_10075_),
    .Y(_10076_),
    .A1(net5831),
    .A2(_10063_));
 sg13g2_a21oi_1 _16056_ (.A1(\fpga_top.io_spi_lite.spi_sck_div[2] ),
    .A2(net5834),
    .Y(_10077_),
    .B1(net5836));
 sg13g2_a22oi_1 _16057_ (.Y(_10078_),
    .B1(_10076_),
    .B2(_10077_),
    .A2(net5836),
    .A1(_06648_));
 sg13g2_a21oi_1 _16058_ (.A1(net5430),
    .A2(_10078_),
    .Y(_10079_),
    .B1(net4930));
 sg13g2_a22oi_1 _16059_ (.Y(_10080_),
    .B1(_10030_),
    .B2(_10079_),
    .A2(net4930),
    .A1(_06684_));
 sg13g2_mux2_1 _16060_ (.A0(net4354),
    .A1(net3033),
    .S(net4201),
    .X(_00158_));
 sg13g2_and2_1 _16061_ (.A(net5706),
    .B(\fpga_top.qspi_if.word_data[27] ),
    .X(_10081_));
 sg13g2_a221oi_1 _16062_ (.B2(\fpga_top.qspi_if.word_data[3] ),
    .C1(_10081_),
    .B1(net5330),
    .A1(\fpga_top.qspi_if.word_data[11] ),
    .Y(_10082_),
    .A2(net5334));
 sg13g2_a21oi_1 _16063_ (.A1(net4474),
    .A2(_10082_),
    .Y(_10083_),
    .B1(net5431));
 sg13g2_o21ai_1 _16064_ (.B1(_10083_),
    .Y(_10084_),
    .A1(_08192_),
    .A2(net4474));
 sg13g2_nand2_1 _16065_ (.Y(_10085_),
    .A(_06834_),
    .B(net5716));
 sg13g2_o21ai_1 _16066_ (.B1(_10085_),
    .Y(_10086_),
    .A1(\fpga_top.io_uart_out.rx_data_latch[3] ),
    .A2(_09908_));
 sg13g2_a21oi_1 _16067_ (.A1(\fpga_top.io_uart_out.uart_io_char[3] ),
    .A2(\fpga_top.io_uart_out.re_uart_rdflg_dly[0] ),
    .Y(_10087_),
    .B1(_09720_));
 sg13g2_o21ai_1 _16068_ (.B1(_10087_),
    .Y(_10088_),
    .A1(_09982_),
    .A2(_10086_));
 sg13g2_nand2b_1 _16069_ (.Y(_10089_),
    .B(\fpga_top.io_led.re_gpio_value_dly[2] ),
    .A_N(\fpga_top.io_led.gpio_in_lat2[3] ));
 sg13g2_o21ai_1 _16070_ (.B1(_10089_),
    .Y(_10090_),
    .A1(uio_oe[7]),
    .A2(_09913_));
 sg13g2_nor2_1 _16071_ (.A(\fpga_top.io_led.re_gpio_value_dly[1] ),
    .B(_10090_),
    .Y(_10091_));
 sg13g2_a221oi_1 _16072_ (.B2(_10091_),
    .C1(net5710),
    .B1(_10088_),
    .A1(\fpga_top.io_led.re_gpio_value_dly[1] ),
    .Y(_10092_),
    .A2(uio_out[7]));
 sg13g2_o21ai_1 _16073_ (.B1(_10031_),
    .Y(_10093_),
    .A1(_06869_),
    .A2(\fpga_top.io_led.gpi_init_lat2[3] ));
 sg13g2_a21oi_1 _16074_ (.A1(\fpga_top.io_frc.frc_cmp_val[35] ),
    .A2(net5718),
    .Y(_10094_),
    .B1(net5731));
 sg13g2_o21ai_1 _16075_ (.B1(_10094_),
    .Y(_10095_),
    .A1(_10092_),
    .A2(_10093_));
 sg13g2_a21oi_1 _16076_ (.A1(_06688_),
    .A2(net5723),
    .Y(_10096_),
    .B1(net5732));
 sg13g2_a221oi_1 _16077_ (.B2(_10096_),
    .C1(net5743),
    .B1(_10095_),
    .A1(\fpga_top.io_frc.frc_cntr_val[35] ),
    .Y(_10097_),
    .A2(net5732));
 sg13g2_o21ai_1 _16078_ (.B1(_09689_),
    .Y(_10098_),
    .A1(\fpga_top.io_frc.frc_cntr_val[3] ),
    .A2(_06871_));
 sg13g2_a21oi_1 _16079_ (.A1(\fpga_top.qspi_if.rdwrch[3] ),
    .A2(net5690),
    .Y(_10099_),
    .B1(_09688_));
 sg13g2_o21ai_1 _16080_ (.B1(_10099_),
    .Y(_10100_),
    .A1(_10097_),
    .A2(_10098_));
 sg13g2_a221oi_1 _16081_ (.B2(_00096_),
    .C1(_09693_),
    .B1(_09930_),
    .A1(_00099_),
    .Y(_10101_),
    .A2(\fpga_top.qspi_if.re_qspi_latency_dly[6] ));
 sg13g2_nand2b_1 _16082_ (.Y(_10102_),
    .B(net5693),
    .A_N(_00110_));
 sg13g2_o21ai_1 _16083_ (.B1(_10102_),
    .Y(_10103_),
    .A1(_00104_),
    .A2(net5693));
 sg13g2_a221oi_1 _16084_ (.B2(_09693_),
    .C1(net5695),
    .B1(_10103_),
    .A1(_10100_),
    .Y(_10104_),
    .A2(_10101_));
 sg13g2_a21oi_1 _16085_ (.A1(_06653_),
    .A2(net5695),
    .Y(_10105_),
    .B1(net5698));
 sg13g2_nand2b_1 _16086_ (.Y(_10106_),
    .B(_10105_),
    .A_N(_10104_));
 sg13g2_a21oi_1 _16087_ (.A1(\fpga_top.qspi_if.read_latency_2[3] ),
    .A2(\fpga_top.qspi_if.re_qspi_latency_dly[2] ),
    .Y(_10107_),
    .B1(_09702_));
 sg13g2_nand2b_1 _16088_ (.Y(_10108_),
    .B(\fpga_top.qspi_if.re_qspi_latency_dly[0] ),
    .A_N(\fpga_top.qspi_if.read_latency_0[3] ));
 sg13g2_o21ai_1 _16089_ (.B1(_10108_),
    .Y(_10109_),
    .A1(\fpga_top.qspi_if.read_latency_1[3] ),
    .A2(\fpga_top.qspi_if.re_qspi_latency_dly[0] ));
 sg13g2_a221oi_1 _16090_ (.B2(net5329),
    .C1(_09701_),
    .B1(_10109_),
    .A1(_10106_),
    .Y(_10110_),
    .A2(_10107_));
 sg13g2_mux4_1 _16091_ (.S0(net5397),
    .A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][3] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][3] ),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][3] ),
    .A3(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][3] ),
    .S1(net5391),
    .X(_10111_));
 sg13g2_nand2b_1 _16092_ (.Y(_10112_),
    .B(net5396),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][3] ));
 sg13g2_o21ai_1 _16093_ (.B1(_10112_),
    .Y(_10113_),
    .A1(net5396),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][3] ));
 sg13g2_mux2_1 _16094_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][3] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][3] ),
    .S(net5396),
    .X(_10114_));
 sg13g2_a21oi_1 _16095_ (.A1(net5391),
    .A2(_10113_),
    .Y(_10115_),
    .B1(_06874_));
 sg13g2_o21ai_1 _16096_ (.B1(_10115_),
    .Y(_10116_),
    .A1(net5391),
    .A2(_10114_));
 sg13g2_a21oi_1 _16097_ (.A1(_06874_),
    .A2(_10111_),
    .Y(_10117_),
    .B1(_06788_));
 sg13g2_a21oi_1 _16098_ (.A1(_10116_),
    .A2(_10117_),
    .Y(_10118_),
    .B1(_09699_));
 sg13g2_o21ai_1 _16099_ (.B1(_10118_),
    .Y(_10119_),
    .A1(net5831),
    .A2(_10110_));
 sg13g2_a21oi_1 _16100_ (.A1(\fpga_top.io_spi_lite.spi_sck_div[3] ),
    .A2(net5834),
    .Y(_10120_),
    .B1(net5836));
 sg13g2_a22oi_1 _16101_ (.Y(_10121_),
    .B1(_10119_),
    .B2(_10120_),
    .A2(net5836),
    .A1(net5830));
 sg13g2_a21oi_1 _16102_ (.A1(net5428),
    .A2(_10121_),
    .Y(_10122_),
    .B1(net4928));
 sg13g2_a22oi_1 _16103_ (.Y(_10123_),
    .B1(_10084_),
    .B2(_10122_),
    .A2(net4928),
    .A1(_06789_));
 sg13g2_mux2_1 _16104_ (.A0(net4347),
    .A1(net3404),
    .S(net4200),
    .X(_00159_));
 sg13g2_nand2_1 _16105_ (.Y(_10124_),
    .A(_08222_),
    .B(net4482));
 sg13g2_a22oi_1 _16106_ (.Y(_10125_),
    .B1(net5331),
    .B2(\fpga_top.qspi_if.word_data[4] ),
    .A2(net5335),
    .A1(\fpga_top.qspi_if.word_data[12] ));
 sg13g2_o21ai_1 _16107_ (.B1(_10125_),
    .Y(_10126_),
    .A1(_06815_),
    .A2(_06828_));
 sg13g2_a21oi_1 _16108_ (.A1(net4474),
    .A2(_10126_),
    .Y(_10127_),
    .B1(net5431));
 sg13g2_nand2_1 _16109_ (.Y(_10128_),
    .A(\fpga_top.io_spi_lite.spi_sck_div[4] ),
    .B(net5835));
 sg13g2_a22oi_1 _16110_ (.Y(_10129_),
    .B1(\fpga_top.io_uart_out.rx_data_latch[4] ),
    .B2(_09907_),
    .A2(net5715),
    .A1(\fpga_top.io_uart_out.uart_term[4] ));
 sg13g2_inv_1 _16111_ (.Y(_10130_),
    .A(_10129_));
 sg13g2_and2_1 _16112_ (.A(_09721_),
    .B(_10031_),
    .X(_10131_));
 sg13g2_nand2_1 _16113_ (.Y(_10132_),
    .A(_09721_),
    .B(_10031_));
 sg13g2_and2_1 _16114_ (.A(_09718_),
    .B(_10131_),
    .X(_10133_));
 sg13g2_inv_1 _16115_ (.Y(_10134_),
    .A(_10133_));
 sg13g2_nand3_1 _16116_ (.B(\fpga_top.io_led.gpi_init_lat2[4] ),
    .C(_10031_),
    .A(\fpga_top.io_led.re_gpio_value_dly[0] ),
    .Y(_10135_));
 sg13g2_nand2_1 _16117_ (.Y(_10136_),
    .A(\fpga_top.io_uart_out.uart_io_char[4] ),
    .B(net5717));
 sg13g2_o21ai_1 _16118_ (.B1(_10135_),
    .Y(_10137_),
    .A1(_10132_),
    .A2(_10136_));
 sg13g2_a221oi_1 _16119_ (.B2(_10133_),
    .C1(_10137_),
    .B1(_10130_),
    .A1(\fpga_top.io_frc.frc_cmp_val[36] ),
    .Y(_10138_),
    .A2(net5718));
 sg13g2_a21oi_1 _16120_ (.A1(\fpga_top.io_frc.frc_cmp_val[4] ),
    .A2(net5722),
    .Y(_10139_),
    .B1(net5733));
 sg13g2_o21ai_1 _16121_ (.B1(_10139_),
    .Y(_10140_),
    .A1(net5722),
    .A2(_10138_));
 sg13g2_a21oi_1 _16122_ (.A1(_06761_),
    .A2(net5732),
    .Y(_10141_),
    .B1(net5743));
 sg13g2_a221oi_1 _16123_ (.B2(_10141_),
    .C1(\fpga_top.qspi_if.re_qspi_latency_dly[9] ),
    .B1(_10140_),
    .A1(\fpga_top.io_frc.frc_cntr_val[4] ),
    .Y(_10142_),
    .A2(net5743));
 sg13g2_a21oi_1 _16124_ (.A1(\fpga_top.qspi_if.wredge[0] ),
    .A2(_06872_),
    .Y(_10143_),
    .B1(_09689_));
 sg13g2_a21oi_1 _16125_ (.A1(net5687),
    .A2(net5690),
    .Y(_10144_),
    .B1(_09688_));
 sg13g2_o21ai_1 _16126_ (.B1(_10144_),
    .Y(_10145_),
    .A1(_10142_),
    .A2(_10143_));
 sg13g2_a221oi_1 _16127_ (.B2(_00097_),
    .C1(_09693_),
    .B1(_09930_),
    .A1(_00100_),
    .Y(_10146_),
    .A2(net5691));
 sg13g2_mux2_1 _16128_ (.A0(\fpga_top.qspi_if.rdcmd1[4] ),
    .A1(\fpga_top.qspi_if.rdcmd0[4] ),
    .S(net5692),
    .X(_10147_));
 sg13g2_a221oi_1 _16129_ (.B2(_09693_),
    .C1(net5694),
    .B1(_10147_),
    .A1(_10145_),
    .Y(_10148_),
    .A2(_10146_));
 sg13g2_nor2_1 _16130_ (.A(\fpga_top.qspi_if.sck_div[4] ),
    .B(_06873_),
    .Y(_10149_));
 sg13g2_nor3_1 _16131_ (.A(_09703_),
    .B(_10148_),
    .C(_10149_),
    .Y(_10150_));
 sg13g2_mux4_1 _16132_ (.S0(net5398),
    .A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][4] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][4] ),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][4] ),
    .A3(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][4] ),
    .S1(net5390),
    .X(_10151_));
 sg13g2_nand2b_1 _16133_ (.Y(_10152_),
    .B(net5397),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][4] ));
 sg13g2_o21ai_1 _16134_ (.B1(_10152_),
    .Y(_10153_),
    .A1(net5397),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][4] ));
 sg13g2_mux2_1 _16135_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][4] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][4] ),
    .S(net5395),
    .X(_10154_));
 sg13g2_a21oi_1 _16136_ (.A1(net5391),
    .A2(_10153_),
    .Y(_10155_),
    .B1(_06874_));
 sg13g2_o21ai_1 _16137_ (.B1(_10155_),
    .Y(_10156_),
    .A1(net5391),
    .A2(_10154_));
 sg13g2_a21oi_1 _16138_ (.A1(_06874_),
    .A2(_10151_),
    .Y(_10157_),
    .B1(_06788_));
 sg13g2_a21oi_1 _16139_ (.A1(_10156_),
    .A2(_10157_),
    .Y(_10158_),
    .B1(_09699_));
 sg13g2_o21ai_1 _16140_ (.B1(_10158_),
    .Y(_10159_),
    .A1(net5831),
    .A2(_10150_));
 sg13g2_a21o_2 _16141_ (.A2(_10159_),
    .A1(_10128_),
    .B1(net5836),
    .X(_10160_));
 sg13g2_a221oi_1 _16142_ (.B2(net5428),
    .C1(net4928),
    .B1(_10160_),
    .A1(_10124_),
    .Y(_10161_),
    .A2(_10127_));
 sg13g2_a21o_2 _16143_ (.A2(net4926),
    .A1(net5661),
    .B1(_10161_),
    .X(_10162_));
 sg13g2_mux2_1 _16144_ (.A0(net4341),
    .A1(net2569),
    .S(net4202),
    .X(_00160_));
 sg13g2_nor2_1 _16145_ (.A(_08101_),
    .B(net4478),
    .Y(_10163_));
 sg13g2_and2_1 _16146_ (.A(net5703),
    .B(net1615),
    .X(_10164_));
 sg13g2_a221oi_1 _16147_ (.B2(net6391),
    .C1(_10164_),
    .B1(net5330),
    .A1(\fpga_top.qspi_if.word_data[13] ),
    .Y(_10165_),
    .A2(net5333));
 sg13g2_or2_1 _16148_ (.X(_10166_),
    .B(_10165_),
    .A(net4484));
 sg13g2_nor2_1 _16149_ (.A(net5434),
    .B(_10163_),
    .Y(_10167_));
 sg13g2_nand2_1 _16150_ (.Y(_10168_),
    .A(\fpga_top.io_uart_out.uart_io_char[5] ),
    .B(net5717));
 sg13g2_nand2_1 _16151_ (.Y(_10169_),
    .A(_06836_),
    .B(net5716));
 sg13g2_o21ai_1 _16152_ (.B1(_10169_),
    .Y(_10170_),
    .A1(\fpga_top.io_uart_out.rx_data_latch[5] ),
    .A2(_09908_));
 sg13g2_o21ai_1 _16153_ (.B1(_10168_),
    .Y(_10171_),
    .A1(_09982_),
    .A2(_10170_));
 sg13g2_and3_1 _16154_ (.X(_10172_),
    .A(\fpga_top.io_led.re_gpio_value_dly[0] ),
    .B(\fpga_top.io_led.gpi_init_lat2[5] ),
    .C(_10031_));
 sg13g2_a221oi_1 _16155_ (.B2(_10171_),
    .C1(_10172_),
    .B1(_10131_),
    .A1(\fpga_top.io_frc.frc_cmp_val[37] ),
    .Y(_10173_),
    .A2(net5718));
 sg13g2_a21oi_1 _16156_ (.A1(\fpga_top.io_frc.frc_cmp_val[5] ),
    .A2(net5722),
    .Y(_10174_),
    .B1(net5733));
 sg13g2_o21ai_1 _16157_ (.B1(_10174_),
    .Y(_10175_),
    .A1(net5722),
    .A2(_10173_));
 sg13g2_a21oi_1 _16158_ (.A1(_06760_),
    .A2(net5732),
    .Y(_10176_),
    .B1(net5743));
 sg13g2_a221oi_1 _16159_ (.B2(_10176_),
    .C1(_09690_),
    .B1(_10175_),
    .A1(\fpga_top.io_frc.frc_cntr_val[5] ),
    .Y(_10177_),
    .A2(net5744));
 sg13g2_a21oi_1 _16160_ (.A1(net5685),
    .A2(net5690),
    .Y(_10178_),
    .B1(_09689_));
 sg13g2_o21ai_1 _16161_ (.B1(_10178_),
    .Y(_10179_),
    .A1(_00094_),
    .A2(net5689));
 sg13g2_nand3b_1 _16162_ (.B(_10179_),
    .C(_09687_),
    .Y(_10180_),
    .A_N(_10177_));
 sg13g2_nand2b_1 _16163_ (.Y(_10181_),
    .B(_09930_),
    .A_N(_00098_));
 sg13g2_nand2b_1 _16164_ (.Y(_10182_),
    .B(net5691),
    .A_N(_00101_));
 sg13g2_nand4_1 _16165_ (.B(_10180_),
    .C(_10181_),
    .A(_09695_),
    .Y(_10183_),
    .D(_10182_));
 sg13g2_nor2_1 _16166_ (.A(_00105_),
    .B(net5692),
    .Y(_10184_));
 sg13g2_a21oi_1 _16167_ (.A1(_06498_),
    .A2(net5692),
    .Y(_10185_),
    .B1(_10184_));
 sg13g2_a221oi_1 _16168_ (.B2(_10185_),
    .C1(_09703_),
    .B1(_09934_),
    .A1(_06655_),
    .Y(_10186_),
    .A2(net5694));
 sg13g2_a21oi_1 _16169_ (.A1(_10183_),
    .A2(_10186_),
    .Y(_10187_),
    .B1(net5831));
 sg13g2_o21ai_1 _16170_ (.B1(net5390),
    .Y(_10188_),
    .A1(net5393),
    .A2(_06891_));
 sg13g2_a21oi_1 _16171_ (.A1(net5395),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][5] ),
    .Y(_10189_),
    .B1(_10188_));
 sg13g2_mux2_1 _16172_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][5] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][5] ),
    .S(net5394),
    .X(_10190_));
 sg13g2_o21ai_1 _16173_ (.B1(net5387),
    .Y(_10191_),
    .A1(net5390),
    .A2(_10190_));
 sg13g2_mux4_1 _16174_ (.S0(net5394),
    .A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][5] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][5] ),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][5] ),
    .A3(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][5] ),
    .S1(net5389),
    .X(_10192_));
 sg13g2_o21ai_1 _16175_ (.B1(net5833),
    .Y(_10193_),
    .A1(_10189_),
    .A2(_10191_));
 sg13g2_a21oi_1 _16176_ (.A1(_06874_),
    .A2(_10192_),
    .Y(_10194_),
    .B1(_10193_));
 sg13g2_nor2_2 _16177_ (.A(_10187_),
    .B(_10194_),
    .Y(_10195_));
 sg13g2_a22oi_1 _16178_ (.Y(_10196_),
    .B1(_09698_),
    .B2(_10195_),
    .A2(net5835),
    .A1(\fpga_top.io_spi_lite.spi_sck_div[5] ));
 sg13g2_or2_1 _16179_ (.X(_10197_),
    .B(_10196_),
    .A(net5838));
 sg13g2_a221oi_1 _16180_ (.B2(net5434),
    .C1(net4927),
    .B1(_10197_),
    .A1(_10166_),
    .Y(_10198_),
    .A2(_10167_));
 sg13g2_a21o_2 _16181_ (.A2(net4926),
    .A1(net5658),
    .B1(_10198_),
    .X(_10199_));
 sg13g2_mux2_1 _16182_ (.A0(net4198),
    .A1(net3423),
    .S(net4202),
    .X(_00161_));
 sg13g2_nand2_1 _16183_ (.Y(_10200_),
    .A(_08247_),
    .B(net4483));
 sg13g2_and2_1 _16184_ (.A(net5703),
    .B(net1442),
    .X(_10201_));
 sg13g2_a221oi_1 _16185_ (.B2(\fpga_top.qspi_if.word_data[6] ),
    .C1(_10201_),
    .B1(net5330),
    .A1(\fpga_top.qspi_if.word_data[14] ),
    .Y(_10202_),
    .A2(net5333));
 sg13g2_a21oi_1 _16186_ (.A1(net4479),
    .A2(_10202_),
    .Y(_10203_),
    .B1(net5434));
 sg13g2_nand2_1 _16187_ (.Y(_10204_),
    .A(\fpga_top.io_uart_out.uart_io_char[6] ),
    .B(net5717));
 sg13g2_nand2_1 _16188_ (.Y(_10205_),
    .A(_06837_),
    .B(net5716));
 sg13g2_o21ai_1 _16189_ (.B1(_10205_),
    .Y(_10206_),
    .A1(\fpga_top.io_uart_out.rx_data_latch[6] ),
    .A2(_09908_));
 sg13g2_o21ai_1 _16190_ (.B1(_10204_),
    .Y(_10207_),
    .A1(_09982_),
    .A2(_10206_));
 sg13g2_a22oi_1 _16191_ (.Y(_10208_),
    .B1(_10131_),
    .B2(_10207_),
    .A2(net5718),
    .A1(\fpga_top.io_frc.frc_cmp_val[38] ));
 sg13g2_a21oi_1 _16192_ (.A1(\fpga_top.io_frc.frc_cmp_val[6] ),
    .A2(net5722),
    .Y(_10209_),
    .B1(net5733));
 sg13g2_o21ai_1 _16193_ (.B1(_10209_),
    .Y(_10210_),
    .A1(net5723),
    .A2(_10208_));
 sg13g2_a21oi_1 _16194_ (.A1(_06758_),
    .A2(net5732),
    .Y(_10211_),
    .B1(net5745));
 sg13g2_a221oi_1 _16195_ (.B2(_10211_),
    .C1(\fpga_top.qspi_if.re_qspi_latency_dly[9] ),
    .B1(_10210_),
    .A1(\fpga_top.io_frc.frc_cntr_val[6] ),
    .Y(_10212_),
    .A2(net5744));
 sg13g2_nor2b_1 _16196_ (.A(\fpga_top.qspi_if.wredge[2] ),
    .B_N(\fpga_top.qspi_if.re_qspi_latency_dly[9] ),
    .Y(_10213_));
 sg13g2_or4_1 _16197_ (.A(net5689),
    .B(_09688_),
    .C(_10212_),
    .D(_10213_),
    .X(_10214_));
 sg13g2_a22oi_1 _16198_ (.Y(_10215_),
    .B1(_09930_),
    .B2(\fpga_top.qspi_if.wrcmd1[6] ),
    .A2(net5691),
    .A1(\fpga_top.qspi_if.wrcmd0[6] ));
 sg13g2_nand3_1 _16199_ (.B(_10214_),
    .C(_10215_),
    .A(_09695_),
    .Y(_10216_));
 sg13g2_mux2_1 _16200_ (.A0(_00106_),
    .A1(_00112_),
    .S(net5692),
    .X(_10217_));
 sg13g2_a221oi_1 _16201_ (.B2(_10217_),
    .C1(_09703_),
    .B1(_09934_),
    .A1(_06657_),
    .Y(_10218_),
    .A2(net5694));
 sg13g2_nand2_1 _16202_ (.Y(_10219_),
    .A(_10216_),
    .B(_10218_));
 sg13g2_nand2b_1 _16203_ (.Y(_10220_),
    .B(net5392),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][6] ));
 sg13g2_o21ai_1 _16204_ (.B1(_10220_),
    .Y(_10221_),
    .A1(net5392),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][6] ));
 sg13g2_mux2_1 _16205_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][6] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][6] ),
    .S(net5392),
    .X(_10222_));
 sg13g2_a21oi_1 _16206_ (.A1(net5389),
    .A2(_10221_),
    .Y(_10223_),
    .B1(net5387));
 sg13g2_o21ai_1 _16207_ (.B1(_10223_),
    .Y(_10224_),
    .A1(net5389),
    .A2(_10222_));
 sg13g2_mux2_1 _16208_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][6] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][6] ),
    .S(net5392),
    .X(_10225_));
 sg13g2_nand2b_1 _16209_ (.Y(_10226_),
    .B(net5393),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][6] ));
 sg13g2_o21ai_1 _16210_ (.B1(_10226_),
    .Y(_10227_),
    .A1(net5393),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][6] ));
 sg13g2_o21ai_1 _16211_ (.B1(net5387),
    .Y(_10228_),
    .A1(net5389),
    .A2(_10225_));
 sg13g2_a21oi_1 _16212_ (.A1(net5388),
    .A2(_10227_),
    .Y(_10229_),
    .B1(_10228_));
 sg13g2_nor2_1 _16213_ (.A(_06788_),
    .B(_10229_),
    .Y(_10230_));
 sg13g2_a22oi_1 _16214_ (.Y(_10231_),
    .B1(_10224_),
    .B2(_10230_),
    .A2(_10219_),
    .A1(_06788_));
 sg13g2_a22oi_1 _16215_ (.Y(_10232_),
    .B1(_09698_),
    .B2(_10231_),
    .A2(net5835),
    .A1(\fpga_top.io_spi_lite.spi_sck_div[6] ));
 sg13g2_nor2_2 _16216_ (.A(net5838),
    .B(_10232_),
    .Y(_10233_));
 sg13g2_a221oi_1 _16217_ (.B2(net5437),
    .C1(net4926),
    .B1(_10233_),
    .A1(_10200_),
    .Y(_10234_),
    .A2(_10203_));
 sg13g2_a21oi_2 _16218_ (.B1(_10234_),
    .Y(_10235_),
    .A2(net4938),
    .A1(_06790_));
 sg13g2_mux2_1 _16219_ (.A0(net4336),
    .A1(net3038),
    .S(net4200),
    .X(_00162_));
 sg13g2_nand2_1 _16220_ (.Y(_10236_),
    .A(_08073_),
    .B(net4482));
 sg13g2_a21oi_1 _16221_ (.A1(net4477),
    .A2(_09671_),
    .Y(_10237_),
    .B1(net5432));
 sg13g2_a221oi_1 _16222_ (.B2(_09907_),
    .C1(_09982_),
    .B1(_06895_),
    .A1(_06838_),
    .Y(_10238_),
    .A2(net5714));
 sg13g2_a21oi_1 _16223_ (.A1(\fpga_top.io_uart_out.uart_io_char[7] ),
    .A2(net5717),
    .Y(_10239_),
    .B1(_10238_));
 sg13g2_a21oi_1 _16224_ (.A1(\fpga_top.io_frc.frc_cmp_val[39] ),
    .A2(net5718),
    .Y(_10240_),
    .B1(net5731));
 sg13g2_o21ai_1 _16225_ (.B1(_10240_),
    .Y(_10241_),
    .A1(_10132_),
    .A2(_10239_));
 sg13g2_a21oi_1 _16226_ (.A1(_06691_),
    .A2(net5722),
    .Y(_10242_),
    .B1(net5733));
 sg13g2_a221oi_1 _16227_ (.B2(_10242_),
    .C1(net5745),
    .B1(_10241_),
    .A1(\fpga_top.io_frc.frc_cntr_val[39] ),
    .Y(_10243_),
    .A2(net5733));
 sg13g2_o21ai_1 _16228_ (.B1(_09691_),
    .Y(_10244_),
    .A1(\fpga_top.io_frc.frc_cntr_val[7] ),
    .A2(_06871_));
 sg13g2_a22oi_1 _16229_ (.Y(_10245_),
    .B1(_09930_),
    .B2(\fpga_top.qspi_if.wrcmd1[7] ),
    .A2(net5691),
    .A1(\fpga_top.qspi_if.wrcmd0[7] ));
 sg13g2_and2_1 _16230_ (.A(_09695_),
    .B(_10245_),
    .X(_10246_));
 sg13g2_o21ai_1 _16231_ (.B1(_10246_),
    .Y(_10247_),
    .A1(_10243_),
    .A2(_10244_));
 sg13g2_nand2b_1 _16232_ (.Y(_10248_),
    .B(net5694),
    .A_N(\fpga_top.qspi_if.sck_div[7] ));
 sg13g2_nand2b_1 _16233_ (.Y(_10249_),
    .B(\fpga_top.qspi_if.rdcmd1[7] ),
    .A_N(net5693));
 sg13g2_nand2b_1 _16234_ (.Y(_10250_),
    .B(net5693),
    .A_N(_00113_));
 sg13g2_nand3_1 _16235_ (.B(_10249_),
    .C(_10250_),
    .A(_09934_),
    .Y(_10251_));
 sg13g2_nand4_1 _16236_ (.B(_10247_),
    .C(_10248_),
    .A(_09704_),
    .Y(_10252_),
    .D(_10251_));
 sg13g2_nand2b_1 _16237_ (.Y(_10253_),
    .B(net5394),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][7] ));
 sg13g2_o21ai_1 _16238_ (.B1(_10253_),
    .Y(_10254_),
    .A1(net5393),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][7] ));
 sg13g2_mux2_1 _16239_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][7] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][7] ),
    .S(net5394),
    .X(_10255_));
 sg13g2_o21ai_1 _16240_ (.B1(net5387),
    .Y(_10256_),
    .A1(net5388),
    .A2(_10254_));
 sg13g2_a21oi_1 _16241_ (.A1(net5388),
    .A2(_10255_),
    .Y(_10257_),
    .B1(_10256_));
 sg13g2_nand2b_1 _16242_ (.Y(_10258_),
    .B(net5393),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][7] ));
 sg13g2_o21ai_1 _16243_ (.B1(_10258_),
    .Y(_10259_),
    .A1(net5393),
    .A2(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][7] ));
 sg13g2_mux2_1 _16244_ (.A0(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][7] ),
    .A1(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][7] ),
    .S(net5394),
    .X(_10260_));
 sg13g2_a21oi_1 _16245_ (.A1(net5389),
    .A2(_10260_),
    .Y(_10261_),
    .B1(net5387));
 sg13g2_o21ai_1 _16246_ (.B1(_10261_),
    .Y(_10262_),
    .A1(net5389),
    .A2(_10259_));
 sg13g2_nand2_1 _16247_ (.Y(_10263_),
    .A(net5833),
    .B(_10262_));
 sg13g2_o21ai_1 _16248_ (.B1(_10252_),
    .Y(_10264_),
    .A1(_10257_),
    .A2(_10263_));
 sg13g2_nand2_1 _16249_ (.Y(_10265_),
    .A(_09700_),
    .B(_10264_));
 sg13g2_nand2_1 _16250_ (.Y(_10266_),
    .A(\fpga_top.io_spi_lite.spi_sck_div[7] ),
    .B(net5834));
 sg13g2_o21ai_1 _16251_ (.B1(_10265_),
    .Y(_10267_),
    .A1(net5837),
    .A2(_10266_));
 sg13g2_a221oi_1 _16252_ (.B2(net5431),
    .C1(net4928),
    .B1(_10267_),
    .A1(_10236_),
    .Y(_10268_),
    .A2(_10237_));
 sg13g2_a21oi_2 _16253_ (.B1(_10268_),
    .Y(_10269_),
    .A2(net4931),
    .A1(_06791_));
 sg13g2_mux2_1 _16254_ (.A0(net4332),
    .A1(net3215),
    .S(net4203),
    .X(_00163_));
 sg13g2_nand2_1 _16255_ (.Y(_10270_),
    .A(_08129_),
    .B(net4482));
 sg13g2_nor2_2 _16256_ (.A(\fpga_top.cpu_top.data_rw_mem.req_hw_dly ),
    .B(net5438),
    .Y(_10271_));
 sg13g2_a22oi_1 _16257_ (.Y(_10272_),
    .B1(net5334),
    .B2(\fpga_top.qspi_if.word_data[0] ),
    .A2(\fpga_top.qspi_if.word_data[16] ),
    .A1(net5706));
 sg13g2_o21ai_1 _16258_ (.B1(_09674_),
    .Y(_10273_),
    .A1(_10271_),
    .A2(_10272_));
 sg13g2_a21oi_1 _16259_ (.A1(net4475),
    .A2(_10273_),
    .Y(_10274_),
    .B1(net5431));
 sg13g2_xnor2_1 _16260_ (.Y(_10275_),
    .A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[2] ),
    .B(\fpga_top.io_spi_lite.miso_fifo.radr[2] ));
 sg13g2_nand2b_1 _16261_ (.Y(_10276_),
    .B(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[0] ),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.radr[0] ));
 sg13g2_nor3_1 _16262_ (.A(_06786_),
    .B(\fpga_top.io_spi_lite.miso_fifo.radr[1] ),
    .C(_10275_),
    .Y(_10277_));
 sg13g2_nor2b_1 _16263_ (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ),
    .B_N(\fpga_top.io_spi_lite.miso_fifo.radr[1] ),
    .Y(_10278_));
 sg13g2_a21oi_1 _16264_ (.A1(_10275_),
    .A2(_10278_),
    .Y(_10279_),
    .B1(_10277_));
 sg13g2_xnor2_1 _16265_ (.Y(_10280_),
    .A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ),
    .B(\fpga_top.io_spi_lite.miso_fifo.radr[1] ));
 sg13g2_nor2b_1 _16266_ (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[0] ),
    .B_N(\fpga_top.io_spi_lite.miso_fifo.radr[0] ),
    .Y(_10281_));
 sg13g2_nand3_1 _16267_ (.B(_10280_),
    .C(_10281_),
    .A(_10275_),
    .Y(_10282_));
 sg13g2_o21ai_1 _16268_ (.B1(_10282_),
    .Y(_10283_),
    .A1(_10276_),
    .A2(_10279_));
 sg13g2_nand2_1 _16269_ (.Y(_10284_),
    .A(\fpga_top.qspi_if.sck_div[8] ),
    .B(net5695));
 sg13g2_a22oi_1 _16270_ (.Y(_10285_),
    .B1(_09907_),
    .B2(\fpga_top.io_uart_out.rx_first_read ),
    .A2(net5715),
    .A1(\fpga_top.io_uart_out.uart_term[8] ));
 sg13g2_a21oi_1 _16271_ (.A1(\fpga_top.io_frc.frc_cmp_val[40] ),
    .A2(net5719),
    .Y(_10286_),
    .B1(net5724));
 sg13g2_o21ai_1 _16272_ (.B1(_10286_),
    .Y(_10287_),
    .A1(_10134_),
    .A2(_10285_));
 sg13g2_a21oi_1 _16273_ (.A1(_06711_),
    .A2(net5724),
    .Y(_10288_),
    .B1(net5734));
 sg13g2_a221oi_1 _16274_ (.B2(_10288_),
    .C1(net5753),
    .B1(_10287_),
    .A1(\fpga_top.io_frc.frc_cntr_val[40] ),
    .Y(_10289_),
    .A2(net5734));
 sg13g2_o21ai_1 _16275_ (.B1(_09696_),
    .Y(_10290_),
    .A1(\fpga_top.io_frc.frc_cntr_val[8] ),
    .A2(_06871_));
 sg13g2_o21ai_1 _16276_ (.B1(_10284_),
    .Y(_10291_),
    .A1(_10289_),
    .A2(_10290_));
 sg13g2_a22oi_1 _16277_ (.Y(_10292_),
    .B1(_10291_),
    .B2(_09704_),
    .A2(_10283_),
    .A1(net5832));
 sg13g2_nor3_1 _16278_ (.A(\fpga_top.io_spi_lite.mosi_pp_cntr[0] ),
    .B(\fpga_top.io_spi_lite.mosi_pp_cntr[1] ),
    .C(\fpga_top.io_spi_lite.mosi_pp_cntr[2] ),
    .Y(_10293_));
 sg13g2_and2_1 _16279_ (.A(\fpga_top.io_spi_lite.mosi_pp_cntr[3] ),
    .B(_10293_),
    .X(_10294_));
 sg13g2_a21oi_1 _16280_ (.A1(\fpga_top.io_spi_lite.re_spi_value_dly[2] ),
    .A2(_10294_),
    .Y(_10295_),
    .B1(net5834));
 sg13g2_o21ai_1 _16281_ (.B1(_10295_),
    .Y(_10296_),
    .A1(\fpga_top.io_spi_lite.re_spi_value_dly[2] ),
    .A2(_10292_));
 sg13g2_nand2b_1 _16282_ (.Y(_10297_),
    .B(net5834),
    .A_N(\fpga_top.io_spi_lite.spi_sck_div[8] ));
 sg13g2_nand3b_1 _16283_ (.B(_10296_),
    .C(_10297_),
    .Y(_10298_),
    .A_N(net5836));
 sg13g2_a221oi_1 _16284_ (.B2(net5433),
    .C1(net4928),
    .B1(_10298_),
    .A1(_10270_),
    .Y(_10299_),
    .A2(_10274_));
 sg13g2_a21o_2 _16285_ (.A2(net4926),
    .A1(net5655),
    .B1(_10299_),
    .X(_10300_));
 sg13g2_mux2_1 _16286_ (.A0(net4328),
    .A1(net2737),
    .S(net4202),
    .X(_00164_));
 sg13g2_a22oi_1 _16287_ (.Y(_10301_),
    .B1(net5333),
    .B2(\fpga_top.qspi_if.word_data[1] ),
    .A2(net1610),
    .A1(net5703));
 sg13g2_o21ai_1 _16288_ (.B1(_09674_),
    .Y(_10302_),
    .A1(_10271_),
    .A2(_10301_));
 sg13g2_a21oi_1 _16289_ (.A1(_08313_),
    .A2(net4484),
    .Y(_10303_),
    .B1(net5435));
 sg13g2_o21ai_1 _16290_ (.B1(_10303_),
    .Y(_10304_),
    .A1(net4484),
    .A2(_10302_));
 sg13g2_xnor2_1 _16291_ (.Y(_10305_),
    .A(_08990_),
    .B(_10275_));
 sg13g2_o21ai_1 _16292_ (.B1(net5832),
    .Y(_10306_),
    .A1(_10280_),
    .A2(_10281_));
 sg13g2_a21oi_1 _16293_ (.A1(_10276_),
    .A2(_10280_),
    .Y(_10307_),
    .B1(_10306_));
 sg13g2_nand2_1 _16294_ (.Y(_10308_),
    .A(\fpga_top.qspi_if.sck_div[9] ),
    .B(net5696));
 sg13g2_a22oi_1 _16295_ (.Y(_10309_),
    .B1(_06903_),
    .B2(_09907_),
    .A2(net5715),
    .A1(_06840_));
 sg13g2_nand2_2 _16296_ (.Y(_10310_),
    .A(_09904_),
    .B(_10309_));
 sg13g2_a21oi_1 _16297_ (.A1(\fpga_top.io_frc.frc_cmp_val[41] ),
    .A2(net5719),
    .Y(_10311_),
    .B1(net5724));
 sg13g2_o21ai_1 _16298_ (.B1(_10311_),
    .Y(_10312_),
    .A1(_10134_),
    .A2(_10310_));
 sg13g2_a21oi_1 _16299_ (.A1(_06709_),
    .A2(net5724),
    .Y(_10313_),
    .B1(net5734));
 sg13g2_a221oi_1 _16300_ (.B2(_10313_),
    .C1(net5753),
    .B1(_10312_),
    .A1(\fpga_top.io_frc.frc_cntr_val[41] ),
    .Y(_10314_),
    .A2(net5734));
 sg13g2_o21ai_1 _16301_ (.B1(_09696_),
    .Y(_10315_),
    .A1(\fpga_top.io_frc.frc_cntr_val[9] ),
    .A2(_06871_));
 sg13g2_o21ai_1 _16302_ (.B1(_10308_),
    .Y(_10316_),
    .A1(_10314_),
    .A2(_10315_));
 sg13g2_a22oi_1 _16303_ (.Y(_10317_),
    .B1(_10316_),
    .B2(_09704_),
    .A2(_10307_),
    .A1(_10305_));
 sg13g2_or2_1 _16304_ (.X(_10318_),
    .B(_10317_),
    .A(\fpga_top.io_spi_lite.re_spi_value_dly[2] ));
 sg13g2_nor2b_2 _16305_ (.A(net1681),
    .B_N(_10293_),
    .Y(_10319_));
 sg13g2_a21oi_1 _16306_ (.A1(\fpga_top.io_spi_lite.re_spi_value_dly[2] ),
    .A2(_10319_),
    .Y(_10320_),
    .B1(net5834));
 sg13g2_a221oi_1 _16307_ (.B2(_10320_),
    .C1(net5837),
    .B1(_10318_),
    .A1(_06785_),
    .Y(_10321_),
    .A2(net5835));
 sg13g2_a21oi_1 _16308_ (.A1(net5436),
    .A2(_10321_),
    .Y(_10322_),
    .B1(net4934));
 sg13g2_a22oi_1 _16309_ (.Y(_10323_),
    .B1(_10304_),
    .B2(_10322_),
    .A2(net4934),
    .A1(_06792_));
 sg13g2_mux2_1 _16310_ (.A0(net4318),
    .A1(net2848),
    .S(net4201),
    .X(_00165_));
 sg13g2_a22oi_1 _16311_ (.Y(_10324_),
    .B1(net5334),
    .B2(\fpga_top.qspi_if.word_data[2] ),
    .A2(net1784),
    .A1(net5703));
 sg13g2_o21ai_1 _16312_ (.B1(_09674_),
    .Y(_10325_),
    .A1(_10271_),
    .A2(_10324_));
 sg13g2_o21ai_1 _16313_ (.B1(_06925_),
    .Y(_10326_),
    .A1(_08012_),
    .A2(net4478));
 sg13g2_a21oi_1 _16314_ (.A1(net4478),
    .A2(_10325_),
    .Y(_10327_),
    .B1(_10326_));
 sg13g2_nand2b_1 _16315_ (.Y(_10328_),
    .B(\fpga_top.io_uart_out.re_uart_rdflg_dly[4] ),
    .A_N(net5714));
 sg13g2_nand3_1 _16316_ (.B(_10133_),
    .C(_10328_),
    .A(_09908_),
    .Y(_10329_));
 sg13g2_nor2b_2 _16317_ (.A(\fpga_top.io_uart_out.uart_term[10] ),
    .B_N(net5714),
    .Y(_10330_));
 sg13g2_a21oi_1 _16318_ (.A1(\fpga_top.io_frc.frc_cmp_val[42] ),
    .A2(net5719),
    .Y(_10331_),
    .B1(net5724));
 sg13g2_o21ai_1 _16319_ (.B1(_10331_),
    .Y(_10332_),
    .A1(_10329_),
    .A2(_10330_));
 sg13g2_a21oi_1 _16320_ (.A1(_06707_),
    .A2(net5730),
    .Y(_10333_),
    .B1(net5742));
 sg13g2_a221oi_1 _16321_ (.B2(_10333_),
    .C1(net5753),
    .B1(_10332_),
    .A1(\fpga_top.io_frc.frc_cntr_val[42] ),
    .Y(_10334_),
    .A2(net5742));
 sg13g2_nor2_1 _16322_ (.A(\fpga_top.io_frc.frc_cntr_val[10] ),
    .B(_06871_),
    .Y(_10335_));
 sg13g2_nor3_2 _16323_ (.A(net4923),
    .B(_10334_),
    .C(_10335_),
    .Y(_10336_));
 sg13g2_nor2_1 _16324_ (.A(_06925_),
    .B(_10336_),
    .Y(_10337_));
 sg13g2_nor3_1 _16325_ (.A(net4932),
    .B(_10327_),
    .C(_10337_),
    .Y(_10338_));
 sg13g2_a21o_2 _16326_ (.A2(net4932),
    .A1(net5652),
    .B1(_10338_),
    .X(_10339_));
 sg13g2_mux2_1 _16327_ (.A0(net4193),
    .A1(net2572),
    .S(net4203),
    .X(_00166_));
 sg13g2_a22oi_1 _16328_ (.Y(_10340_),
    .B1(net5333),
    .B2(\fpga_top.qspi_if.word_data[3] ),
    .A2(net1846),
    .A1(net5704));
 sg13g2_o21ai_1 _16329_ (.B1(_09674_),
    .Y(_10341_),
    .A1(_10271_),
    .A2(_10340_));
 sg13g2_o21ai_1 _16330_ (.B1(_06925_),
    .Y(_10342_),
    .A1(_08279_),
    .A2(net4479));
 sg13g2_a21oi_1 _16331_ (.A1(net4478),
    .A2(_10341_),
    .Y(_10343_),
    .B1(_10342_));
 sg13g2_nor2b_1 _16332_ (.A(\fpga_top.io_uart_out.uart_term[11] ),
    .B_N(net5714),
    .Y(_10344_));
 sg13g2_a21oi_1 _16333_ (.A1(\fpga_top.io_frc.frc_cmp_val[43] ),
    .A2(net5719),
    .Y(_10345_),
    .B1(net5724));
 sg13g2_o21ai_1 _16334_ (.B1(_10345_),
    .Y(_10346_),
    .A1(_10329_),
    .A2(_10344_));
 sg13g2_a21oi_1 _16335_ (.A1(_06705_),
    .A2(net5726),
    .Y(_10347_),
    .B1(net5737));
 sg13g2_a221oi_1 _16336_ (.B2(_10347_),
    .C1(net5748),
    .B1(_10346_),
    .A1(\fpga_top.io_frc.frc_cntr_val[43] ),
    .Y(_10348_),
    .A2(net5737));
 sg13g2_nor2_1 _16337_ (.A(\fpga_top.io_frc.frc_cntr_val[11] ),
    .B(_06871_),
    .Y(_10349_));
 sg13g2_nor3_2 _16338_ (.A(net4923),
    .B(_10348_),
    .C(_10349_),
    .Y(_10350_));
 sg13g2_nor2_1 _16339_ (.A(_06925_),
    .B(_10350_),
    .Y(_10351_));
 sg13g2_nor3_1 _16340_ (.A(net4934),
    .B(_10343_),
    .C(_10351_),
    .Y(_10352_));
 sg13g2_a21o_2 _16341_ (.A2(net4934),
    .A1(net5651),
    .B1(_10352_),
    .X(_10353_));
 sg13g2_mux2_1 _16342_ (.A0(net4189),
    .A1(net3346),
    .S(net4201),
    .X(_00167_));
 sg13g2_a22oi_1 _16343_ (.Y(_10354_),
    .B1(net5334),
    .B2(\fpga_top.qspi_if.word_data[4] ),
    .A2(\fpga_top.qspi_if.word_data[20] ),
    .A1(net5706));
 sg13g2_o21ai_1 _16344_ (.B1(_09674_),
    .Y(_10355_),
    .A1(_10271_),
    .A2(_10354_));
 sg13g2_inv_1 _16345_ (.Y(_10356_),
    .A(_10355_));
 sg13g2_a21oi_1 _16346_ (.A1(net4479),
    .A2(_10356_),
    .Y(_10357_),
    .B1(net5435));
 sg13g2_o21ai_1 _16347_ (.B1(_10357_),
    .Y(_10358_),
    .A1(_08345_),
    .A2(net4479));
 sg13g2_a21oi_2 _16348_ (.B1(_10329_),
    .Y(_10359_),
    .A2(net5714),
    .A1(_06843_));
 sg13g2_a21o_1 _16349_ (.A2(net5720),
    .A1(\fpga_top.io_frc.frc_cmp_val[44] ),
    .B1(net5727),
    .X(_10360_));
 sg13g2_a21oi_1 _16350_ (.A1(_06704_),
    .A2(net5727),
    .Y(_10361_),
    .B1(net5740));
 sg13g2_o21ai_1 _16351_ (.B1(_10361_),
    .Y(_10362_),
    .A1(_10359_),
    .A2(_10360_));
 sg13g2_a21oi_1 _16352_ (.A1(\fpga_top.io_frc.frc_cntr_val[44] ),
    .A2(net5740),
    .Y(_10363_),
    .B1(net5751));
 sg13g2_a221oi_1 _16353_ (.B2(_10363_),
    .C1(net4923),
    .B1(_10362_),
    .A1(_06703_),
    .Y(_10364_),
    .A2(net5751));
 sg13g2_a21oi_1 _16354_ (.A1(net5434),
    .A2(_10364_),
    .Y(_10365_),
    .B1(net4932));
 sg13g2_a22oi_1 _16355_ (.Y(_10366_),
    .B1(_10358_),
    .B2(_10365_),
    .A2(net4932),
    .A1(net5376));
 sg13g2_mux2_1 _16356_ (.A0(net4317),
    .A1(net3451),
    .S(net4203),
    .X(_00168_));
 sg13g2_a22oi_1 _16357_ (.Y(_10367_),
    .B1(net5333),
    .B2(net2095),
    .A2(net1660),
    .A1(net5703));
 sg13g2_o21ai_1 _16358_ (.B1(_09674_),
    .Y(_10368_),
    .A1(_10271_),
    .A2(_10367_));
 sg13g2_inv_1 _16359_ (.Y(_10369_),
    .A(_10368_));
 sg13g2_a21oi_1 _16360_ (.A1(net4479),
    .A2(_10369_),
    .Y(_10370_),
    .B1(net5435));
 sg13g2_o21ai_1 _16361_ (.B1(_10370_),
    .Y(_10371_),
    .A1(_07970_),
    .A2(net4480));
 sg13g2_a21oi_2 _16362_ (.B1(_10329_),
    .Y(_10372_),
    .A2(net5714),
    .A1(_06844_));
 sg13g2_a21o_1 _16363_ (.A2(net5720),
    .A1(\fpga_top.io_frc.frc_cmp_val[45] ),
    .B1(net5727),
    .X(_10373_));
 sg13g2_a21oi_1 _16364_ (.A1(_06702_),
    .A2(net5727),
    .Y(_10374_),
    .B1(net5740));
 sg13g2_o21ai_1 _16365_ (.B1(_10374_),
    .Y(_10375_),
    .A1(_10372_),
    .A2(_10373_));
 sg13g2_a21oi_1 _16366_ (.A1(\fpga_top.io_frc.frc_cntr_val[45] ),
    .A2(net5740),
    .Y(_10376_),
    .B1(net5751));
 sg13g2_a221oi_1 _16367_ (.B2(_10376_),
    .C1(net4923),
    .B1(_10375_),
    .A1(_06701_),
    .Y(_10377_),
    .A2(net5750));
 sg13g2_a21oi_1 _16368_ (.A1(net5435),
    .A2(_10377_),
    .Y(_10378_),
    .B1(net4932));
 sg13g2_a22oi_1 _16369_ (.Y(_10379_),
    .B1(_10371_),
    .B2(_10378_),
    .A2(net4936),
    .A1(net5374));
 sg13g2_mux2_1 _16370_ (.A0(net4311),
    .A1(net3100),
    .S(net4201),
    .X(_00169_));
 sg13g2_nand2_1 _16371_ (.Y(_10380_),
    .A(_07944_),
    .B(net4483));
 sg13g2_a22oi_1 _16372_ (.Y(_10381_),
    .B1(net5333),
    .B2(\fpga_top.qspi_if.word_data[6] ),
    .A2(net1669),
    .A1(net5703));
 sg13g2_o21ai_1 _16373_ (.B1(_09674_),
    .Y(_10382_),
    .A1(_10271_),
    .A2(_10381_));
 sg13g2_a21oi_1 _16374_ (.A1(net4479),
    .A2(_10382_),
    .Y(_10383_),
    .B1(net5436));
 sg13g2_nand3_1 _16375_ (.B(net5714),
    .C(_10133_),
    .A(\fpga_top.io_uart_out.uart_term[14] ),
    .Y(_10384_));
 sg13g2_a21oi_1 _16376_ (.A1(\fpga_top.io_frc.frc_cmp_val[46] ),
    .A2(net5720),
    .Y(_10385_),
    .B1(net5727));
 sg13g2_a22oi_1 _16377_ (.Y(_10386_),
    .B1(_10384_),
    .B2(_10385_),
    .A2(net5727),
    .A1(_06700_));
 sg13g2_nand2b_1 _16378_ (.Y(_10387_),
    .B(_10386_),
    .A_N(net5740));
 sg13g2_a21oi_1 _16379_ (.A1(\fpga_top.io_frc.frc_cntr_val[46] ),
    .A2(net5740),
    .Y(_10388_),
    .B1(net5751));
 sg13g2_a21oi_1 _16380_ (.A1(_10387_),
    .A2(_10388_),
    .Y(_10389_),
    .B1(net4923));
 sg13g2_o21ai_1 _16381_ (.B1(_10389_),
    .Y(_10390_),
    .A1(\fpga_top.io_frc.frc_cntr_val[14] ),
    .A2(_06871_));
 sg13g2_a221oi_1 _16382_ (.B2(net5434),
    .C1(net4927),
    .B1(_10390_),
    .A1(_10380_),
    .Y(_10391_),
    .A2(_10383_));
 sg13g2_a21o_2 _16383_ (.A2(net4926),
    .A1(net5650),
    .B1(_10391_),
    .X(_10392_));
 sg13g2_mux2_1 _16384_ (.A0(net4303),
    .A1(net2418),
    .S(net4200),
    .X(_00170_));
 sg13g2_nor3_1 _16385_ (.A(_09673_),
    .B(_09675_),
    .C(_10271_),
    .Y(_10393_));
 sg13g2_nor2_1 _16386_ (.A(net4924),
    .B(_10393_),
    .Y(_10394_));
 sg13g2_a21oi_1 _16387_ (.A1(net4479),
    .A2(_10394_),
    .Y(_10395_),
    .B1(net5436));
 sg13g2_o21ai_1 _16388_ (.B1(_10395_),
    .Y(_10396_),
    .A1(_08548_),
    .A2(net4478));
 sg13g2_a21oi_2 _16389_ (.B1(_10329_),
    .Y(_10397_),
    .A2(net5714),
    .A1(_06846_));
 sg13g2_a21o_1 _16390_ (.A2(net5720),
    .A1(\fpga_top.io_frc.frc_cmp_val[47] ),
    .B1(net5727),
    .X(_10398_));
 sg13g2_a21oi_1 _16391_ (.A1(_06698_),
    .A2(net5728),
    .Y(_10399_),
    .B1(net5739));
 sg13g2_o21ai_1 _16392_ (.B1(_10399_),
    .Y(_10400_),
    .A1(_10397_),
    .A2(_10398_));
 sg13g2_a21oi_1 _16393_ (.A1(\fpga_top.io_frc.frc_cntr_val[47] ),
    .A2(net5739),
    .Y(_10401_),
    .B1(net5750));
 sg13g2_a221oi_1 _16394_ (.B2(_10401_),
    .C1(net4923),
    .B1(_10400_),
    .A1(_06697_),
    .Y(_10402_),
    .A2(net5750));
 sg13g2_a21oi_1 _16395_ (.A1(net5434),
    .A2(_10402_),
    .Y(_10403_),
    .B1(net4933));
 sg13g2_a22oi_1 _16396_ (.Y(_10404_),
    .B1(_10396_),
    .B2(_10403_),
    .A2(net4932),
    .A1(net5373));
 sg13g2_mux2_1 _16397_ (.A0(net4299),
    .A1(net2426),
    .S(net4203),
    .X(_00171_));
 sg13g2_nand2_2 _16398_ (.Y(_10405_),
    .A(net5702),
    .B(net3837));
 sg13g2_nand3_1 _16399_ (.B(\fpga_top.qspi_if.word_data[8] ),
    .C(net5440),
    .A(net5702),
    .Y(_10406_));
 sg13g2_nor2b_1 _16400_ (.A(net4925),
    .B_N(_10406_),
    .Y(_10407_));
 sg13g2_a21oi_1 _16401_ (.A1(net4475),
    .A2(_10407_),
    .Y(_10408_),
    .B1(net5429));
 sg13g2_o21ai_1 _16402_ (.B1(_10408_),
    .Y(_10409_),
    .A1(_08038_),
    .A2(net4475));
 sg13g2_o21ai_1 _16403_ (.B1(net5068),
    .Y(_10410_),
    .A1(\fpga_top.io_frc.frc_cmp_val[48] ),
    .A2(net5356));
 sg13g2_a21oi_1 _16404_ (.A1(\fpga_top.io_frc.frc_cmp_val[16] ),
    .A2(net5725),
    .Y(_10411_),
    .B1(net5735));
 sg13g2_a22oi_1 _16405_ (.Y(_10412_),
    .B1(_10410_),
    .B2(_10411_),
    .A2(net5736),
    .A1(_06742_));
 sg13g2_a21oi_1 _16406_ (.A1(_06730_),
    .A2(net5747),
    .Y(_10413_),
    .B1(_09694_));
 sg13g2_o21ai_1 _16407_ (.B1(_10413_),
    .Y(_10414_),
    .A1(net5746),
    .A2(_10412_));
 sg13g2_nand2b_1 _16408_ (.Y(_10415_),
    .B(net5696),
    .A_N(\fpga_top.qspi_if.dbg_2div_wirte_half_end ));
 sg13g2_nand3_1 _16409_ (.B(_09704_),
    .C(_10415_),
    .A(_09700_),
    .Y(_10416_));
 sg13g2_a21oi_2 _16410_ (.B1(_10416_),
    .Y(_10417_),
    .A2(_10414_),
    .A1(_06873_));
 sg13g2_a21o_2 _16411_ (.A2(\fpga_top.io_spi_lite.spi_mode[4] ),
    .A1(net5838),
    .B1(_10417_),
    .X(_10418_));
 sg13g2_a21oi_1 _16412_ (.A1(net5429),
    .A2(_10418_),
    .Y(_10419_),
    .B1(net4929));
 sg13g2_a22oi_1 _16413_ (.Y(_10420_),
    .B1(_10409_),
    .B2(_10419_),
    .A2(net4929),
    .A1(_06798_));
 sg13g2_mux2_1 _16414_ (.A0(net4293),
    .A1(net3397),
    .S(net4203),
    .X(_00172_));
 sg13g2_nand2_2 _16415_ (.Y(_10421_),
    .A(net5707),
    .B(net2241));
 sg13g2_and3_1 _16416_ (.X(_10422_),
    .A(net5707),
    .B(\fpga_top.qspi_if.word_data[9] ),
    .C(net5438));
 sg13g2_o21ai_1 _16417_ (.B1(net4477),
    .Y(_10423_),
    .A1(net4924),
    .A2(_10422_));
 sg13g2_a21oi_1 _16418_ (.A1(_08377_),
    .A2(net4482),
    .Y(_10424_),
    .B1(net5428));
 sg13g2_nor3_1 _16419_ (.A(_06741_),
    .B(net5356),
    .C(net5725),
    .Y(_10425_));
 sg13g2_a21oi_1 _16420_ (.A1(\fpga_top.io_frc.frc_cmp_val[17] ),
    .A2(net5725),
    .Y(_10426_),
    .B1(_10425_));
 sg13g2_a21oi_1 _16421_ (.A1(\fpga_top.io_frc.frc_cntr_val[49] ),
    .A2(net5735),
    .Y(_10427_),
    .B1(net5747));
 sg13g2_o21ai_1 _16422_ (.B1(_10427_),
    .Y(_10428_),
    .A1(net5735),
    .A2(_10426_));
 sg13g2_a21oi_1 _16423_ (.A1(_06729_),
    .A2(net5747),
    .Y(_10429_),
    .B1(_09697_));
 sg13g2_a22oi_1 _16424_ (.Y(_10430_),
    .B1(_10428_),
    .B2(_10429_),
    .A2(net5696),
    .A1(\fpga_top.qspi_if.dbg_2div_read_half_end ));
 sg13g2_nor2_2 _16425_ (.A(_09705_),
    .B(_10430_),
    .Y(_10431_));
 sg13g2_a21oi_2 _16426_ (.B1(_10431_),
    .Y(_10432_),
    .A2(\fpga_top.io_spi_lite.spi_mode[5] ),
    .A1(net5838));
 sg13g2_a221oi_1 _16427_ (.B2(net5432),
    .C1(net4929),
    .B1(_10432_),
    .A1(_10423_),
    .Y(_10433_),
    .A2(_10424_));
 sg13g2_a21o_2 _16428_ (.A2(net4933),
    .A1(net5648),
    .B1(_10433_),
    .X(_10434_));
 sg13g2_mux2_1 _16429_ (.A0(net4287),
    .A1(net2662),
    .S(net4200),
    .X(_00173_));
 sg13g2_nand2_1 _16430_ (.Y(_10435_),
    .A(_08526_),
    .B(net4482));
 sg13g2_and2_1 _16431_ (.A(net5705),
    .B(net1863),
    .X(_10436_));
 sg13g2_a21oi_1 _16432_ (.A1(net5439),
    .A2(_10436_),
    .Y(_10437_),
    .B1(net4925));
 sg13g2_a21oi_1 _16433_ (.A1(net4475),
    .A2(_10437_),
    .Y(_10438_),
    .B1(net5430));
 sg13g2_nand2_1 _16434_ (.Y(_10439_),
    .A(\fpga_top.io_spi_lite.re_spi_value_dly[0] ),
    .B(\fpga_top.io_spi_lite.spi_mode[6] ));
 sg13g2_o21ai_1 _16435_ (.B1(net5068),
    .Y(_10440_),
    .A1(\fpga_top.io_frc.frc_cmp_val[50] ),
    .A2(net5356));
 sg13g2_a21oi_1 _16436_ (.A1(\fpga_top.io_frc.frc_cmp_val[18] ),
    .A2(net5725),
    .Y(_10441_),
    .B1(net5735));
 sg13g2_a22oi_1 _16437_ (.Y(_10442_),
    .B1(_10440_),
    .B2(_10441_),
    .A2(net5735),
    .A1(_06746_));
 sg13g2_a21oi_1 _16438_ (.A1(_06732_),
    .A2(net5746),
    .Y(_10443_),
    .B1(_09694_));
 sg13g2_o21ai_1 _16439_ (.B1(_10443_),
    .Y(_10444_),
    .A1(net5746),
    .A2(_10442_));
 sg13g2_nand2_1 _16440_ (.Y(_10445_),
    .A(_06873_),
    .B(_10444_));
 sg13g2_o21ai_1 _16441_ (.B1(_10445_),
    .Y(_10446_),
    .A1(\fpga_top.qspi_if.dbg_reg_2div_cec_write ),
    .A2(_06873_));
 sg13g2_o21ai_1 _16442_ (.B1(_10439_),
    .Y(_10447_),
    .A1(_09705_),
    .A2(_10446_));
 sg13g2_a221oi_1 _16443_ (.B2(net5429),
    .C1(net4930),
    .B1(_10447_),
    .A1(_10435_),
    .Y(_10448_),
    .A2(_10438_));
 sg13g2_a21oi_2 _16444_ (.B1(_10448_),
    .Y(_10449_),
    .A2(net4931),
    .A1(_06800_));
 sg13g2_mux2_1 _16445_ (.A0(net4282),
    .A1(net2723),
    .S(net4203),
    .X(_00174_));
 sg13g2_and2_1 _16446_ (.A(net5705),
    .B(net1999),
    .X(_10450_));
 sg13g2_a21oi_1 _16447_ (.A1(net5438),
    .A2(_10450_),
    .Y(_10451_),
    .B1(net4924));
 sg13g2_a21oi_1 _16448_ (.A1(net4478),
    .A2(_10451_),
    .Y(_10452_),
    .B1(net5434));
 sg13g2_o21ai_1 _16449_ (.B1(_10452_),
    .Y(_10453_),
    .A1(_08405_),
    .A2(net4478));
 sg13g2_o21ai_1 _16450_ (.B1(net5068),
    .Y(_10454_),
    .A1(\fpga_top.io_frc.frc_cmp_val[51] ),
    .A2(net5356));
 sg13g2_a21oi_1 _16451_ (.A1(\fpga_top.io_frc.frc_cmp_val[19] ),
    .A2(net5725),
    .Y(_10455_),
    .B1(net5736));
 sg13g2_a22oi_1 _16452_ (.Y(_10456_),
    .B1(_10454_),
    .B2(_10455_),
    .A2(net5736),
    .A1(_06744_));
 sg13g2_nor2_1 _16453_ (.A(net5746),
    .B(_10456_),
    .Y(_10457_));
 sg13g2_a21oi_1 _16454_ (.A1(_06731_),
    .A2(net5746),
    .Y(_10458_),
    .B1(_10457_));
 sg13g2_a22oi_1 _16455_ (.Y(_10459_),
    .B1(_09696_),
    .B2(_10458_),
    .A2(net5696),
    .A1(\fpga_top.qspi_if.dbg_reg_2div_cec_read ));
 sg13g2_nor2_2 _16456_ (.A(_09705_),
    .B(_10459_),
    .Y(_10460_));
 sg13g2_a21oi_1 _16457_ (.A1(net5434),
    .A2(_10460_),
    .Y(_10461_),
    .B1(net4926));
 sg13g2_a22oi_1 _16458_ (.Y(_10462_),
    .B1(_10453_),
    .B2(_10461_),
    .A2(net4926),
    .A1(_06801_));
 sg13g2_mux2_1 _16459_ (.A0(net4278),
    .A1(net3030),
    .S(net4200),
    .X(_00175_));
 sg13g2_nand2_1 _16460_ (.Y(_10463_),
    .A(net5702),
    .B(net3728));
 sg13g2_and3_1 _16461_ (.X(_10464_),
    .A(net5702),
    .B(\fpga_top.qspi_if.word_data[12] ),
    .C(net5440));
 sg13g2_o21ai_1 _16462_ (.B1(net4476),
    .Y(_10465_),
    .A1(net4925),
    .A2(_10464_));
 sg13g2_a21oi_1 _16463_ (.A1(_08428_),
    .A2(net4482),
    .Y(_10466_),
    .B1(net5428));
 sg13g2_nor3_1 _16464_ (.A(_06753_),
    .B(net5356),
    .C(net5725),
    .Y(_10467_));
 sg13g2_a21oi_1 _16465_ (.A1(\fpga_top.io_frc.frc_cmp_val[20] ),
    .A2(net5725),
    .Y(_10468_),
    .B1(_10467_));
 sg13g2_a21oi_1 _16466_ (.A1(\fpga_top.io_frc.frc_cntr_val[52] ),
    .A2(net5735),
    .Y(_10469_),
    .B1(net5746));
 sg13g2_o21ai_1 _16467_ (.B1(_10469_),
    .Y(_10470_),
    .A1(net5736),
    .A2(_10468_));
 sg13g2_a21oi_1 _16468_ (.A1(_06728_),
    .A2(net5747),
    .Y(_10471_),
    .B1(_09697_));
 sg13g2_a22oi_1 _16469_ (.Y(_10472_),
    .B1(_10470_),
    .B2(_10471_),
    .A2(net5696),
    .A1(\fpga_top.qspi_if.dbg_2div_trt ));
 sg13g2_nor2_1 _16470_ (.A(_09705_),
    .B(_10472_),
    .Y(_10473_));
 sg13g2_a21oi_2 _16471_ (.B1(_10473_),
    .Y(_10474_),
    .A2(\fpga_top.io_spi_lite.spi_mode[7] ),
    .A1(net5837));
 sg13g2_a221oi_1 _16472_ (.B2(net5428),
    .C1(net4927),
    .B1(_10474_),
    .A1(_10465_),
    .Y(_10475_),
    .A2(_10466_));
 sg13g2_a21o_2 _16473_ (.A2(net4927),
    .A1(net5646),
    .B1(_10475_),
    .X(_10476_));
 sg13g2_mux2_1 _16474_ (.A0(net4271),
    .A1(net2956),
    .S(net4202),
    .X(_00176_));
 sg13g2_and2_1 _16475_ (.A(net5704),
    .B(net1718),
    .X(_10477_));
 sg13g2_a21oi_1 _16476_ (.A1(net5439),
    .A2(_10477_),
    .Y(_10478_),
    .B1(net4924));
 sg13g2_or2_1 _16477_ (.X(_10479_),
    .B(_10478_),
    .A(net4484));
 sg13g2_a21oi_1 _16478_ (.A1(_07867_),
    .A2(net4482),
    .Y(_10480_),
    .B1(net5428));
 sg13g2_o21ai_1 _16479_ (.B1(net5068),
    .Y(_10481_),
    .A1(\fpga_top.io_frc.frc_cmp_val[53] ),
    .A2(net5356));
 sg13g2_a21oi_1 _16480_ (.A1(\fpga_top.io_frc.frc_cmp_val[21] ),
    .A2(net5725),
    .Y(_10482_),
    .B1(net5735));
 sg13g2_a22oi_1 _16481_ (.Y(_10483_),
    .B1(_10481_),
    .B2(_10482_),
    .A2(net5735),
    .A1(_06751_));
 sg13g2_a21oi_1 _16482_ (.A1(_06726_),
    .A2(net5746),
    .Y(_10484_),
    .B1(_09694_));
 sg13g2_o21ai_1 _16483_ (.B1(_10484_),
    .Y(_10485_),
    .A1(net5746),
    .A2(_10483_));
 sg13g2_nand2_1 _16484_ (.Y(_10486_),
    .A(_06873_),
    .B(_10485_));
 sg13g2_a21oi_1 _16485_ (.A1(_06770_),
    .A2(net5696),
    .Y(_10487_),
    .B1(_09705_));
 sg13g2_a22oi_1 _16486_ (.Y(_10488_),
    .B1(_10486_),
    .B2(_10487_),
    .A2(\fpga_top.io_spi_lite.spi_mode[8] ),
    .A1(net5837));
 sg13g2_a221oi_1 _16487_ (.B2(net5428),
    .C1(net4927),
    .B1(_10488_),
    .A1(_10479_),
    .Y(_10489_),
    .A2(_10480_));
 sg13g2_a21o_2 _16488_ (.A2(net4926),
    .A1(net5644),
    .B1(_10489_),
    .X(_10490_));
 sg13g2_mux2_1 _16489_ (.A0(net4264),
    .A1(net3043),
    .S(net4200),
    .X(_00177_));
 sg13g2_nand2_1 _16490_ (.Y(_10491_),
    .A(net5702),
    .B(net3207));
 sg13g2_nand3_1 _16491_ (.B(\fpga_top.qspi_if.word_data[14] ),
    .C(net5440),
    .A(net5702),
    .Y(_10492_));
 sg13g2_nand3b_1 _16492_ (.B(_10492_),
    .C(net4475),
    .Y(_10493_),
    .A_N(net4925));
 sg13g2_a21oi_1 _16493_ (.A1(_07837_),
    .A2(net4482),
    .Y(_10494_),
    .B1(net5433));
 sg13g2_a21oi_1 _16494_ (.A1(\fpga_top.io_frc.frc_cmp_val[54] ),
    .A2(net5720),
    .Y(_10495_),
    .B1(net5726));
 sg13g2_a21o_1 _16495_ (.A2(net5726),
    .A1(_06725_),
    .B1(_10495_),
    .X(_10496_));
 sg13g2_a21oi_1 _16496_ (.A1(\fpga_top.io_frc.frc_cntr_val[54] ),
    .A2(net5737),
    .Y(_10497_),
    .B1(net5748));
 sg13g2_o21ai_1 _16497_ (.B1(_10497_),
    .Y(_10498_),
    .A1(net5737),
    .A2(_10496_));
 sg13g2_a21oi_1 _16498_ (.A1(_06724_),
    .A2(net5748),
    .Y(_10499_),
    .B1(_09697_));
 sg13g2_a22oi_1 _16499_ (.Y(_10500_),
    .B1(_10498_),
    .B2(_10499_),
    .A2(net5697),
    .A1(\fpga_top.dbg_bpoint_en[1] ));
 sg13g2_nand2_1 _16500_ (.Y(_10501_),
    .A(net5837),
    .B(\fpga_top.io_spi_lite.spi_mode[9] ));
 sg13g2_o21ai_1 _16501_ (.B1(_10501_),
    .Y(_10502_),
    .A1(_09705_),
    .A2(_10500_));
 sg13g2_a221oi_1 _16502_ (.B2(net5428),
    .C1(net4927),
    .B1(_10502_),
    .A1(_10493_),
    .Y(_10503_),
    .A2(_10494_));
 sg13g2_a21oi_2 _16503_ (.B1(_10503_),
    .Y(_10504_),
    .A2(net4927),
    .A1(_06803_));
 sg13g2_mux2_1 _16504_ (.A0(net4262),
    .A1(net3752),
    .S(net4204),
    .X(_00178_));
 sg13g2_and2_1 _16505_ (.A(net5702),
    .B(net1910),
    .X(_10505_));
 sg13g2_a21oi_1 _16506_ (.A1(net5440),
    .A2(_10505_),
    .Y(_10506_),
    .B1(net4925));
 sg13g2_a21oi_1 _16507_ (.A1(net4476),
    .A2(_10506_),
    .Y(_10507_),
    .B1(net5429));
 sg13g2_o21ai_1 _16508_ (.B1(_10507_),
    .Y(_10508_),
    .A1(_08475_),
    .A2(net4475));
 sg13g2_o21ai_1 _16509_ (.B1(net5068),
    .Y(_10509_),
    .A1(\fpga_top.io_frc.frc_cmp_val[55] ),
    .A2(net5356));
 sg13g2_a21oi_1 _16510_ (.A1(\fpga_top.io_frc.frc_cmp_val[23] ),
    .A2(net5726),
    .Y(_10510_),
    .B1(net5737));
 sg13g2_a22oi_1 _16511_ (.Y(_10511_),
    .B1(_10509_),
    .B2(_10510_),
    .A2(net5737),
    .A1(_06748_));
 sg13g2_nor2_1 _16512_ (.A(net5748),
    .B(_10511_),
    .Y(_10512_));
 sg13g2_a21oi_1 _16513_ (.A1(_06723_),
    .A2(net5748),
    .Y(_10513_),
    .B1(_10512_));
 sg13g2_a22oi_1 _16514_ (.Y(_10514_),
    .B1(_09696_),
    .B2(_10513_),
    .A2(net5697),
    .A1(\fpga_top.dbg_bpoint_en[2] ));
 sg13g2_nor2_2 _16515_ (.A(_09705_),
    .B(_10514_),
    .Y(_10515_));
 sg13g2_a21oi_1 _16516_ (.A1(net5429),
    .A2(_10515_),
    .Y(_10516_),
    .B1(net4930));
 sg13g2_a22oi_1 _16517_ (.Y(_10517_),
    .B1(_10508_),
    .B2(_10516_),
    .A2(net4930),
    .A1(_06804_));
 sg13g2_mux2_1 _16518_ (.A0(net4258),
    .A1(net3238),
    .S(net4203),
    .X(_00179_));
 sg13g2_mux2_1 _16519_ (.A0(net4406),
    .A1(net3452),
    .S(net4204),
    .X(_00180_));
 sg13g2_mux2_1 _16520_ (.A0(net4401),
    .A1(net2798),
    .S(net4202),
    .X(_00181_));
 sg13g2_mux2_1 _16521_ (.A0(net4396),
    .A1(net3465),
    .S(net4201),
    .X(_00182_));
 sg13g2_mux2_1 _16522_ (.A0(net4390),
    .A1(net2384),
    .S(net4201),
    .X(_00183_));
 sg13g2_mux2_1 _16523_ (.A0(net4382),
    .A1(net2650),
    .S(net4200),
    .X(_00184_));
 sg13g2_mux2_1 _16524_ (.A0(net4380),
    .A1(net2615),
    .S(net4203),
    .X(_00185_));
 sg13g2_mux2_1 _16525_ (.A0(net4374),
    .A1(net2244),
    .S(net4202),
    .X(_00186_));
 sg13g2_mux2_1 _16526_ (.A0(net4371),
    .A1(net2799),
    .S(net4202),
    .X(_00187_));
 sg13g2_nand2b_1 _16527_ (.Y(_10518_),
    .B(_08978_),
    .A_N(_08898_));
 sg13g2_or2_1 _16528_ (.X(_10519_),
    .B(_10518_),
    .A(_08982_));
 sg13g2_nor2_2 _16529_ (.A(_09617_),
    .B(_10519_),
    .Y(_10520_));
 sg13g2_and2_1 _16530_ (.A(_08888_),
    .B(_08988_),
    .X(_10521_));
 sg13g2_nand2_2 _16531_ (.Y(_10522_),
    .A(_08892_),
    .B(_10521_));
 sg13g2_nor2_1 _16532_ (.A(net3153),
    .B(_10520_),
    .Y(_10523_));
 sg13g2_nand2_1 _16533_ (.Y(_10524_),
    .A(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .B(net5085));
 sg13g2_mux2_1 _16534_ (.A0(_06562_),
    .A1(_06683_),
    .S(net5086),
    .X(_10525_));
 sg13g2_o21ai_1 _16535_ (.B1(_10524_),
    .Y(_10526_),
    .A1(_06562_),
    .A2(net5085));
 sg13g2_a21oi_1 _16536_ (.A1(_10520_),
    .A2(net4920),
    .Y(_00188_),
    .B1(_10523_));
 sg13g2_nor2_1 _16537_ (.A(net2119),
    .B(_10520_),
    .Y(_10527_));
 sg13g2_nand2_1 _16538_ (.Y(_10528_),
    .A(\fpga_top.cpu_top.csr_wdata_mon[1] ),
    .B(net5087));
 sg13g2_mux2_1 _16539_ (.A0(_06561_),
    .A1(_06681_),
    .S(net5088),
    .X(_10529_));
 sg13g2_o21ai_1 _16540_ (.B1(_10528_),
    .Y(_10530_),
    .A1(_06561_),
    .A2(net5087));
 sg13g2_a21oi_1 _16541_ (.A1(_10520_),
    .A2(net4918),
    .Y(_00189_),
    .B1(_10527_));
 sg13g2_nor2_1 _16542_ (.A(net3831),
    .B(_10520_),
    .Y(_10531_));
 sg13g2_a21oi_1 _16543_ (.A1(net4852),
    .A2(_10520_),
    .Y(_00190_),
    .B1(_10531_));
 sg13g2_nand3_1 _16544_ (.B(net1777),
    .C(_08835_),
    .A(net3181),
    .Y(_10532_));
 sg13g2_or3_1 _16545_ (.A(_08972_),
    .B(_10319_),
    .C(_10532_),
    .X(_10533_));
 sg13g2_nand2_1 _16546_ (.Y(_10534_),
    .A(net6192),
    .B(_08972_));
 sg13g2_nand3_1 _16547_ (.B(_10533_),
    .C(_10534_),
    .A(_09413_),
    .Y(_00191_));
 sg13g2_nand2_1 _16548_ (.Y(_10535_),
    .A(_08835_),
    .B(_10319_));
 sg13g2_nand3_1 _16549_ (.B(_10532_),
    .C(_10535_),
    .A(_09407_),
    .Y(_10536_));
 sg13g2_nand2_1 _16550_ (.Y(_10537_),
    .A(net3827),
    .B(_08972_));
 sg13g2_o21ai_1 _16551_ (.B1(_10537_),
    .Y(_00192_),
    .A1(_08972_),
    .A2(_10536_));
 sg13g2_nor2_2 _16552_ (.A(_09410_),
    .B(_09646_),
    .Y(_10538_));
 sg13g2_nand2_1 _16553_ (.Y(_10539_),
    .A(_09409_),
    .B(_09647_));
 sg13g2_mux4_1 _16554_ (.S0(\fpga_top.io_spi_lite.spi_mode[10] ),
    .A0(\fpga_top.io_spi_lite.miso_lat[4] ),
    .A1(\fpga_top.io_spi_lite.miso_lat[5] ),
    .A2(\fpga_top.io_spi_lite.miso_lat[6] ),
    .A3(\fpga_top.io_spi_lite.miso_lat[7] ),
    .S1(\fpga_top.io_spi_lite.spi_mode[11] ),
    .X(_10540_));
 sg13g2_nor2_1 _16555_ (.A(_09410_),
    .B(_09647_),
    .Y(_10541_));
 sg13g2_mux4_1 _16556_ (.S0(\fpga_top.io_spi_lite.spi_mode[10] ),
    .A0(\fpga_top.io_led.gpi_init_lat1[0] ),
    .A1(\fpga_top.io_led.gpi_init_lat2[0] ),
    .A2(\fpga_top.io_spi_lite.miso_lat[2] ),
    .A3(\fpga_top.io_spi_lite.miso_lat[3] ),
    .S1(\fpga_top.io_spi_lite.spi_mode[11] ),
    .X(_10542_));
 sg13g2_mux2_1 _16557_ (.A0(_10542_),
    .A1(_10540_),
    .S(\fpga_top.io_spi_lite.spi_mode[12] ),
    .X(_10543_));
 sg13g2_a22oi_1 _16558_ (.Y(_10544_),
    .B1(net5067),
    .B2(_10543_),
    .A2(_10538_),
    .A1(net3733));
 sg13g2_inv_1 _16559_ (.Y(_00193_),
    .A(_10544_));
 sg13g2_a22oi_1 _16560_ (.Y(_10545_),
    .B1(net5067),
    .B2(net3733),
    .A2(_10538_),
    .A1(net3713));
 sg13g2_inv_1 _16561_ (.Y(_00194_),
    .A(net3734));
 sg13g2_a22oi_1 _16562_ (.Y(_10546_),
    .B1(net5067),
    .B2(net3713),
    .A2(_10538_),
    .A1(net3651));
 sg13g2_inv_1 _16563_ (.Y(_00195_),
    .A(net3714));
 sg13g2_a22oi_1 _16564_ (.Y(_10547_),
    .B1(net5067),
    .B2(net3651),
    .A2(_10538_),
    .A1(net3574));
 sg13g2_inv_1 _16565_ (.Y(_00196_),
    .A(net3652));
 sg13g2_a22oi_1 _16566_ (.Y(_10548_),
    .B1(net5067),
    .B2(net3574),
    .A2(_10538_),
    .A1(net3509));
 sg13g2_inv_1 _16567_ (.Y(_00197_),
    .A(net3575));
 sg13g2_a22oi_1 _16568_ (.Y(_10549_),
    .B1(net5067),
    .B2(net3509),
    .A2(_10538_),
    .A1(\fpga_top.io_spi_lite.miso_byte_org[5] ));
 sg13g2_inv_1 _16569_ (.Y(_00198_),
    .A(net3510));
 sg13g2_a22oi_1 _16570_ (.Y(_10550_),
    .B1(net5067),
    .B2(net3692),
    .A2(_10538_),
    .A1(\fpga_top.io_spi_lite.miso_byte_org[6] ));
 sg13g2_inv_1 _16571_ (.Y(_00199_),
    .A(net3693));
 sg13g2_a22oi_1 _16572_ (.Y(_10551_),
    .B1(net5067),
    .B2(net3841),
    .A2(_10538_),
    .A1(\fpga_top.io_spi_lite.miso_byte_org[7] ));
 sg13g2_inv_1 _16573_ (.Y(_00200_),
    .A(net3842));
 sg13g2_nor2b_1 _16574_ (.A(_08895_),
    .B_N(_08897_),
    .Y(_10552_));
 sg13g2_nor2b_2 _16575_ (.A(_08982_),
    .B_N(_10552_),
    .Y(_10553_));
 sg13g2_inv_1 _16576_ (.Y(_10554_),
    .A(_10553_));
 sg13g2_nand3b_1 _16577_ (.B(_10553_),
    .C(_08978_),
    .Y(_10555_),
    .A_N(_10294_));
 sg13g2_nor4_2 _16578_ (.A(_08979_),
    .B(_08985_),
    .C(_10294_),
    .Y(_10556_),
    .D(_10554_));
 sg13g2_nor2_2 _16579_ (.A(_08989_),
    .B(_10555_),
    .Y(_10557_));
 sg13g2_nor2_1 _16580_ (.A(_08975_),
    .B(_10557_),
    .Y(_10558_));
 sg13g2_nand2_1 _16581_ (.Y(_10559_),
    .A(_08975_),
    .B(_10556_));
 sg13g2_nor2b_1 _16582_ (.A(_10558_),
    .B_N(_10559_),
    .Y(_10560_));
 sg13g2_xnor2_1 _16583_ (.Y(_00201_),
    .A(net3201),
    .B(_10560_));
 sg13g2_or4_1 _16584_ (.A(\fpga_top.io_spi_lite.mosi_pp_cntr[0] ),
    .B(\fpga_top.io_spi_lite.mosi_pp_cntr[1] ),
    .C(_08975_),
    .D(_10557_),
    .X(_10561_));
 sg13g2_nand2_1 _16585_ (.Y(_10562_),
    .A(\fpga_top.io_spi_lite.mosi_pp_cntr[0] ),
    .B(_10559_));
 sg13g2_o21ai_1 _16586_ (.B1(_10562_),
    .Y(_10563_),
    .A1(\fpga_top.io_spi_lite.mosi_pp_cntr[0] ),
    .A2(_10558_));
 sg13g2_xnor2_1 _16587_ (.Y(_00202_),
    .A(net1756),
    .B(_10563_));
 sg13g2_nand4_1 _16588_ (.B(\fpga_top.io_spi_lite.mosi_pp_cntr[1] ),
    .C(_08975_),
    .A(\fpga_top.io_spi_lite.mosi_pp_cntr[0] ),
    .Y(_10564_),
    .D(_10556_));
 sg13g2_nand2_1 _16589_ (.Y(_10565_),
    .A(_10561_),
    .B(_10564_));
 sg13g2_xor2_1 _16590_ (.B(_10565_),
    .A(net1580),
    .X(_00203_));
 sg13g2_mux2_1 _16591_ (.A0(_10561_),
    .A1(_10564_),
    .S(net1580),
    .X(_10566_));
 sg13g2_xnor2_1 _16592_ (.Y(_00204_),
    .A(net1681),
    .B(_10566_));
 sg13g2_nor2_1 _16593_ (.A(net1655),
    .B(_10541_),
    .Y(_10567_));
 sg13g2_a21oi_1 _16594_ (.A1(net1655),
    .A2(_10539_),
    .Y(_00205_),
    .B1(_10567_));
 sg13g2_a21oi_1 _16595_ (.A1(\fpga_top.io_spi_lite.miso_bit_cntr[0] ),
    .A2(_10539_),
    .Y(_10568_),
    .B1(net1427));
 sg13g2_a21oi_1 _16596_ (.A1(_09646_),
    .A2(_09648_),
    .Y(_10569_),
    .B1(_09410_));
 sg13g2_nor2b_1 _16597_ (.A(net1428),
    .B_N(_10569_),
    .Y(_00206_));
 sg13g2_a21oi_1 _16598_ (.A1(_09648_),
    .A2(_10539_),
    .Y(_10570_),
    .B1(net1407));
 sg13g2_nor3_1 _16599_ (.A(_09410_),
    .B(\fpga_top.io_spi_lite.miso_read_next_byte ),
    .C(net1408),
    .Y(_00207_));
 sg13g2_nand2_1 _16600_ (.Y(_10571_),
    .A(_08972_),
    .B(_09409_));
 sg13g2_nor2_1 _16601_ (.A(_08972_),
    .B(_09410_),
    .Y(_10572_));
 sg13g2_nor2_1 _16602_ (.A(net1703),
    .B(_10572_),
    .Y(_10573_));
 sg13g2_a21oi_1 _16603_ (.A1(net1703),
    .A2(_10571_),
    .Y(_00208_),
    .B1(_10573_));
 sg13g2_a21oi_1 _16604_ (.A1(net1703),
    .A2(_10571_),
    .Y(_10574_),
    .B1(net1975));
 sg13g2_nor3_1 _16605_ (.A(_08973_),
    .B(_09410_),
    .C(net1976),
    .Y(_00209_));
 sg13g2_o21ai_1 _16606_ (.B1(_09409_),
    .Y(_10575_),
    .A1(net1915),
    .A2(_08973_));
 sg13g2_nor2_1 _16607_ (.A(_08974_),
    .B(_10575_),
    .Y(_00210_));
 sg13g2_nand2_2 _16608_ (.Y(_10576_),
    .A(net6414),
    .B(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[0] ));
 sg13g2_or2_1 _16609_ (.X(_10577_),
    .B(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[0] ),
    .A(net6414));
 sg13g2_nand2b_2 _16610_ (.Y(_10578_),
    .B(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wen ),
    .A_N(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[0] ));
 sg13g2_and3_1 _16611_ (.X(_00211_),
    .A(_08987_),
    .B(net6415),
    .C(_10577_));
 sg13g2_nand3_1 _16612_ (.B(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[0] ),
    .C(net6491),
    .A(net6414),
    .Y(_10579_));
 sg13g2_nand2_1 _16613_ (.Y(_10580_),
    .A(_06786_),
    .B(net6415));
 sg13g2_and3_1 _16614_ (.X(_00212_),
    .A(_08987_),
    .B(_10579_),
    .C(_10580_));
 sg13g2_or2_1 _16615_ (.X(_10581_),
    .B(_10579_),
    .A(_06787_));
 sg13g2_nand2_1 _16616_ (.Y(_10582_),
    .A(_06787_),
    .B(_10579_));
 sg13g2_and3_1 _16617_ (.X(_00213_),
    .A(_08987_),
    .B(net5270),
    .C(net6537));
 sg13g2_or2_1 _16618_ (.X(_10583_),
    .B(_09803_),
    .A(_09659_));
 sg13g2_mux2_1 _16619_ (.A0(net4364),
    .A1(net2849),
    .S(net4180),
    .X(_00214_));
 sg13g2_mux2_1 _16620_ (.A0(net4358),
    .A1(net3576),
    .S(net4182),
    .X(_00215_));
 sg13g2_mux2_1 _16621_ (.A0(net4354),
    .A1(net2320),
    .S(net4181),
    .X(_00216_));
 sg13g2_mux2_1 _16622_ (.A0(net4347),
    .A1(net2969),
    .S(net4180),
    .X(_00217_));
 sg13g2_mux2_1 _16623_ (.A0(net4341),
    .A1(net2254),
    .S(net4182),
    .X(_00218_));
 sg13g2_mux2_1 _16624_ (.A0(net4199),
    .A1(net3403),
    .S(net4182),
    .X(_00219_));
 sg13g2_mux2_1 _16625_ (.A0(net4336),
    .A1(net2681),
    .S(net4180),
    .X(_00220_));
 sg13g2_mux2_1 _16626_ (.A0(net4332),
    .A1(net2267),
    .S(net4183),
    .X(_00221_));
 sg13g2_mux2_1 _16627_ (.A0(net4328),
    .A1(net2460),
    .S(net4182),
    .X(_00222_));
 sg13g2_mux2_1 _16628_ (.A0(net4318),
    .A1(net2953),
    .S(net4181),
    .X(_00223_));
 sg13g2_mux2_1 _16629_ (.A0(net4193),
    .A1(net2225),
    .S(net4183),
    .X(_00224_));
 sg13g2_mux2_1 _16630_ (.A0(net4187),
    .A1(net2389),
    .S(net4181),
    .X(_00225_));
 sg13g2_mux2_1 _16631_ (.A0(net4317),
    .A1(net2903),
    .S(net4183),
    .X(_00226_));
 sg13g2_mux2_1 _16632_ (.A0(net4311),
    .A1(net2510),
    .S(net4181),
    .X(_00227_));
 sg13g2_mux2_1 _16633_ (.A0(net4303),
    .A1(net2172),
    .S(net4180),
    .X(_00228_));
 sg13g2_mux2_1 _16634_ (.A0(net4299),
    .A1(net3216),
    .S(net4183),
    .X(_00229_));
 sg13g2_mux2_1 _16635_ (.A0(net4293),
    .A1(net2366),
    .S(net4183),
    .X(_00230_));
 sg13g2_mux2_1 _16636_ (.A0(net4288),
    .A1(net3241),
    .S(net4180),
    .X(_00231_));
 sg13g2_mux2_1 _16637_ (.A0(net4282),
    .A1(net2322),
    .S(net4183),
    .X(_00232_));
 sg13g2_mux2_1 _16638_ (.A0(net4278),
    .A1(net3416),
    .S(net4180),
    .X(_00233_));
 sg13g2_mux2_1 _16639_ (.A0(net4271),
    .A1(net2512),
    .S(net4182),
    .X(_00234_));
 sg13g2_mux2_1 _16640_ (.A0(net4264),
    .A1(net2739),
    .S(net4180),
    .X(_00235_));
 sg13g2_mux2_1 _16641_ (.A0(net4262),
    .A1(net3099),
    .S(net4184),
    .X(_00236_));
 sg13g2_mux2_1 _16642_ (.A0(net4258),
    .A1(net3014),
    .S(net4183),
    .X(_00237_));
 sg13g2_mux2_1 _16643_ (.A0(net4406),
    .A1(net3420),
    .S(net4184),
    .X(_00238_));
 sg13g2_mux2_1 _16644_ (.A0(net4401),
    .A1(net2447),
    .S(net4182),
    .X(_00239_));
 sg13g2_mux2_1 _16645_ (.A0(net4396),
    .A1(net2438),
    .S(net4181),
    .X(_00240_));
 sg13g2_mux2_1 _16646_ (.A0(net4390),
    .A1(net2715),
    .S(net4181),
    .X(_00241_));
 sg13g2_mux2_1 _16647_ (.A0(net4382),
    .A1(net3485),
    .S(net4180),
    .X(_00242_));
 sg13g2_mux2_1 _16648_ (.A0(net4380),
    .A1(net3271),
    .S(net4183),
    .X(_00243_));
 sg13g2_mux2_1 _16649_ (.A0(net4374),
    .A1(net3247),
    .S(net4182),
    .X(_00244_));
 sg13g2_mux2_1 _16650_ (.A0(net4371),
    .A1(net3062),
    .S(net4182),
    .X(_00245_));
 sg13g2_nor2_2 _16651_ (.A(_08985_),
    .B(_10519_),
    .Y(_10584_));
 sg13g2_nor2_1 _16652_ (.A(net6089),
    .B(net4471),
    .Y(_10585_));
 sg13g2_a21oi_1 _16653_ (.A1(net4920),
    .A2(net4471),
    .Y(_00246_),
    .B1(_10585_));
 sg13g2_nor2_1 _16654_ (.A(net1777),
    .B(net4469),
    .Y(_10586_));
 sg13g2_a21oi_1 _16655_ (.A1(net4917),
    .A2(net4469),
    .Y(_00247_),
    .B1(_10586_));
 sg13g2_nor2_1 _16656_ (.A(net3181),
    .B(net4469),
    .Y(_10587_));
 sg13g2_a21oi_1 _16657_ (.A1(net4852),
    .A2(net4469),
    .Y(_00248_),
    .B1(_10587_));
 sg13g2_nor2_1 _16658_ (.A(net5830),
    .B(net4469),
    .Y(_10588_));
 sg13g2_nand2_1 _16659_ (.Y(_10589_),
    .A(net5662),
    .B(net5087));
 sg13g2_o21ai_1 _16660_ (.B1(_10589_),
    .Y(_10590_),
    .A1(_06570_),
    .A2(net5087));
 sg13g2_a21oi_1 _16661_ (.A1(net4469),
    .A2(net4844),
    .Y(_00249_),
    .B1(_10588_));
 sg13g2_nor2_1 _16662_ (.A(net6359),
    .B(net4471),
    .Y(_10591_));
 sg13g2_nor2_2 _16663_ (.A(\fpga_top.bus_gather.d_write_data[16] ),
    .B(net5078),
    .Y(_10592_));
 sg13g2_nand2_1 _16664_ (.Y(_10593_),
    .A(_06798_),
    .B(net5080));
 sg13g2_nor2b_2 _16665_ (.A(_10592_),
    .B_N(_10593_),
    .Y(_10594_));
 sg13g2_nand2b_2 _16666_ (.Y(_10595_),
    .B(_10593_),
    .A_N(_10592_));
 sg13g2_a21oi_1 _16667_ (.A1(net4471),
    .A2(_10595_),
    .Y(_00250_),
    .B1(_10591_));
 sg13g2_nor2_1 _16668_ (.A(net6332),
    .B(net4471),
    .Y(_10596_));
 sg13g2_nor2_1 _16669_ (.A(\fpga_top.bus_gather.d_write_data[17] ),
    .B(net5080),
    .Y(_10597_));
 sg13g2_nand2_1 _16670_ (.Y(_10598_),
    .A(_06799_),
    .B(net5080));
 sg13g2_nor2b_2 _16671_ (.A(_10597_),
    .B_N(_10598_),
    .Y(_10599_));
 sg13g2_nand2b_2 _16672_ (.Y(_10600_),
    .B(_10598_),
    .A_N(_10597_));
 sg13g2_a21oi_1 _16673_ (.A1(net4471),
    .A2(_10600_),
    .Y(_00251_),
    .B1(_10596_));
 sg13g2_nor2_1 _16674_ (.A(net3829),
    .B(net4471),
    .Y(_10601_));
 sg13g2_nand2_1 _16675_ (.Y(_10602_),
    .A(_06800_),
    .B(net5090));
 sg13g2_o21ai_1 _16676_ (.B1(_10602_),
    .Y(_10603_),
    .A1(\fpga_top.bus_gather.d_write_data[18] ),
    .A2(net5090));
 sg13g2_a21oi_1 _16677_ (.A1(net4471),
    .A2(_10603_),
    .Y(_00252_),
    .B1(_10601_));
 sg13g2_nor2_1 _16678_ (.A(net5826),
    .B(net4470),
    .Y(_10604_));
 sg13g2_mux2_1 _16679_ (.A0(_06619_),
    .A1(_06802_),
    .S(net5083),
    .X(_10605_));
 sg13g2_inv_1 _16680_ (.Y(_10606_),
    .A(_10605_));
 sg13g2_a21oi_1 _16681_ (.A1(net4470),
    .A2(_10605_),
    .Y(_00253_),
    .B1(_10604_));
 sg13g2_nor2_1 _16682_ (.A(net3892),
    .B(net4470),
    .Y(_10607_));
 sg13g2_nand2b_1 _16683_ (.Y(_10608_),
    .B(net5086),
    .A_N(net5644));
 sg13g2_o21ai_1 _16684_ (.B1(_10608_),
    .Y(_10609_),
    .A1(\fpga_top.bus_gather.d_write_data[21] ),
    .A2(net5086));
 sg13g2_a21oi_1 _16685_ (.A1(net4469),
    .A2(_10609_),
    .Y(_00254_),
    .B1(_10607_));
 sg13g2_nor2_1 _16686_ (.A(net3502),
    .B(net4469),
    .Y(_10610_));
 sg13g2_mux2_1 _16687_ (.A0(_06624_),
    .A1(_06803_),
    .S(net5084),
    .X(_10611_));
 sg13g2_inv_1 _16688_ (.Y(_10612_),
    .A(_10611_));
 sg13g2_a21oi_1 _16689_ (.A1(net4470),
    .A2(_10611_),
    .Y(_00255_),
    .B1(_10610_));
 sg13g2_nor2_1 _16690_ (.A(net6312),
    .B(net4472),
    .Y(_10613_));
 sg13g2_nand2_1 _16691_ (.Y(_10614_),
    .A(_06805_),
    .B(net5089));
 sg13g2_o21ai_1 _16692_ (.B1(_10614_),
    .Y(_10615_),
    .A1(\fpga_top.bus_gather.d_write_data[24] ),
    .A2(net5090));
 sg13g2_a21oi_1 _16693_ (.A1(net4472),
    .A2(_10615_),
    .Y(_00256_),
    .B1(_10613_));
 sg13g2_nor2_1 _16694_ (.A(net6288),
    .B(net4472),
    .Y(_10616_));
 sg13g2_nand2_1 _16695_ (.Y(_10617_),
    .A(_06806_),
    .B(net5089));
 sg13g2_o21ai_1 _16696_ (.B1(_10617_),
    .Y(_10618_),
    .A1(\fpga_top.bus_gather.d_write_data[25] ),
    .A2(net5089));
 sg13g2_inv_2 _16697_ (.Y(_10619_),
    .A(_10618_));
 sg13g2_a21oi_1 _16698_ (.A1(net4472),
    .A2(_10618_),
    .Y(_00257_),
    .B1(_10616_));
 sg13g2_nor2_1 _16699_ (.A(net6085),
    .B(net4473),
    .Y(_10620_));
 sg13g2_nand2_1 _16700_ (.Y(_10621_),
    .A(_06807_),
    .B(net5090));
 sg13g2_o21ai_1 _16701_ (.B1(_10621_),
    .Y(_10622_),
    .A1(\fpga_top.bus_gather.d_write_data[26] ),
    .A2(net5090));
 sg13g2_a21oi_1 _16702_ (.A1(net4473),
    .A2(_10622_),
    .Y(_00258_),
    .B1(_10620_));
 sg13g2_nor3_1 _16703_ (.A(\fpga_top.cpu_top.csr_uimm[0] ),
    .B(\fpga_top.cpu_top.csr_uimm[1] ),
    .C(\fpga_top.cpu_top.csr_uimm[3] ),
    .Y(_10623_));
 sg13g2_nand3b_1 _16704_ (.B(_06618_),
    .C(_10623_),
    .Y(_10624_),
    .A_N(\fpga_top.cpu_top.csr_uimm[2] ));
 sg13g2_nor2b_1 _16705_ (.A(_09437_),
    .B_N(_10624_),
    .Y(_10625_));
 sg13g2_nand2_1 _16706_ (.Y(_10626_),
    .A(net5825),
    .B(net5157));
 sg13g2_nand2_1 _16707_ (.Y(_10627_),
    .A(_09437_),
    .B(_10624_));
 sg13g2_mux4_1 _16708_ (.S0(net5535),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][0] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][0] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][0] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][0] ),
    .S1(net5490),
    .X(_10628_));
 sg13g2_mux4_1 _16709_ (.S0(net5538),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][0] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][0] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][0] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][0] ),
    .S1(net5493),
    .X(_10629_));
 sg13g2_mux2_1 _16710_ (.A0(_10628_),
    .A1(_10629_),
    .S(net5362),
    .X(_10630_));
 sg13g2_mux4_1 _16711_ (.S0(net5526),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][0] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][0] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][0] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][0] ),
    .S1(net5481),
    .X(_10631_));
 sg13g2_nor2_1 _16712_ (.A(net5464),
    .B(_10631_),
    .Y(_10632_));
 sg13g2_mux4_1 _16713_ (.S0(net5535),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][0] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][0] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][0] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][0] ),
    .S1(net5490),
    .X(_10633_));
 sg13g2_o21ai_1 _16714_ (.B1(net5453),
    .Y(_10634_),
    .A1(net5362),
    .A2(_10633_));
 sg13g2_o21ai_1 _16715_ (.B1(net5442),
    .Y(_10635_),
    .A1(_10632_),
    .A2(_10634_));
 sg13g2_a21o_1 _16716_ (.A2(_10630_),
    .A1(net5359),
    .B1(_10635_),
    .X(_10636_));
 sg13g2_mux4_1 _16717_ (.S0(net5524),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][0] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][0] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][0] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][0] ),
    .S1(net5479),
    .X(_10637_));
 sg13g2_mux4_1 _16718_ (.S0(net5524),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][0] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][0] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][0] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][0] ),
    .S1(net5479),
    .X(_10638_));
 sg13g2_mux4_1 _16719_ (.S0(net5524),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][0] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][0] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][0] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][0] ),
    .S1(net5479),
    .X(_10639_));
 sg13g2_mux4_1 _16720_ (.S0(net5527),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][0] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][0] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][0] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][0] ),
    .S1(net5482),
    .X(_10640_));
 sg13g2_mux4_1 _16721_ (.S0(net5362),
    .A0(_10637_),
    .A1(_10638_),
    .A2(_10639_),
    .A3(_10640_),
    .S1(net5453),
    .X(_10641_));
 sg13g2_o21ai_1 _16722_ (.B1(_10636_),
    .Y(_10642_),
    .A1(net5442),
    .A2(_10641_));
 sg13g2_o21ai_1 _16723_ (.B1(_10626_),
    .Y(_00259_),
    .A1(net5151),
    .A2(_10642_));
 sg13g2_nand2_1 _16724_ (.Y(_10643_),
    .A(net5824),
    .B(net5157));
 sg13g2_mux4_1 _16725_ (.S0(net5559),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][1] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][1] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][1] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][1] ),
    .S1(net5514),
    .X(_10644_));
 sg13g2_inv_1 _16726_ (.Y(_10645_),
    .A(_10644_));
 sg13g2_mux4_1 _16727_ (.S0(net5559),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][1] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][1] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][1] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][1] ),
    .S1(net5514),
    .X(_10646_));
 sg13g2_a21oi_1 _16728_ (.A1(net5470),
    .A2(_10645_),
    .Y(_10647_),
    .B1(net5458));
 sg13g2_o21ai_1 _16729_ (.B1(_10647_),
    .Y(_10648_),
    .A1(net5470),
    .A2(_10646_));
 sg13g2_mux4_1 _16730_ (.S0(net5559),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][1] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][1] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][1] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][1] ),
    .S1(net5514),
    .X(_10649_));
 sg13g2_mux4_1 _16731_ (.S0(net5559),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][1] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][1] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][1] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][1] ),
    .S1(net5514),
    .X(_10650_));
 sg13g2_nor2_1 _16732_ (.A(net5369),
    .B(_10650_),
    .Y(_10651_));
 sg13g2_o21ai_1 _16733_ (.B1(net5458),
    .Y(_10652_),
    .A1(net5470),
    .A2(_10649_));
 sg13g2_o21ai_1 _16734_ (.B1(net5449),
    .Y(_10653_),
    .A1(_10651_),
    .A2(_10652_));
 sg13g2_nand2b_2 _16735_ (.Y(_10654_),
    .B(_10648_),
    .A_N(_10653_));
 sg13g2_mux4_1 _16736_ (.S0(net5548),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][1] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][1] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][1] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][1] ),
    .S1(net5503),
    .X(_10655_));
 sg13g2_mux4_1 _16737_ (.S0(net5547),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][1] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][1] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][1] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][1] ),
    .S1(net5502),
    .X(_10656_));
 sg13g2_mux4_1 _16738_ (.S0(net5549),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][1] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][1] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][1] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][1] ),
    .S1(net5504),
    .X(_10657_));
 sg13g2_mux4_1 _16739_ (.S0(net5548),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][1] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][1] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][1] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][1] ),
    .S1(net5503),
    .X(_10658_));
 sg13g2_mux4_1 _16740_ (.S0(net5368),
    .A0(_10655_),
    .A1(_10656_),
    .A2(_10657_),
    .A3(_10658_),
    .S1(net5457),
    .X(_10659_));
 sg13g2_o21ai_1 _16741_ (.B1(_10654_),
    .Y(_10660_),
    .A1(net5446),
    .A2(_10659_));
 sg13g2_o21ai_1 _16742_ (.B1(_10643_),
    .Y(_00260_),
    .A1(net5151),
    .A2(_10660_));
 sg13g2_nand2_1 _16743_ (.Y(_10661_),
    .A(net5819),
    .B(net5157));
 sg13g2_mux4_1 _16744_ (.S0(net5543),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][2] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][2] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][2] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][2] ),
    .S1(net5498),
    .X(_10662_));
 sg13g2_nor2_1 _16745_ (.A(net5366),
    .B(_10662_),
    .Y(_10663_));
 sg13g2_mux4_1 _16746_ (.S0(net5543),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][2] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][2] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][2] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][2] ),
    .S1(net5498),
    .X(_10664_));
 sg13g2_o21ai_1 _16747_ (.B1(net5455),
    .Y(_10665_),
    .A1(net5467),
    .A2(_10664_));
 sg13g2_nor2_1 _16748_ (.A(_10663_),
    .B(_10665_),
    .Y(_10666_));
 sg13g2_mux4_1 _16749_ (.S0(net5543),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][2] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][2] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][2] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][2] ),
    .S1(net5498),
    .X(_10667_));
 sg13g2_mux4_1 _16750_ (.S0(net5543),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][2] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][2] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][2] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][2] ),
    .S1(net5498),
    .X(_10668_));
 sg13g2_nor2_1 _16751_ (.A(net5467),
    .B(_10668_),
    .Y(_10669_));
 sg13g2_o21ai_1 _16752_ (.B1(net5358),
    .Y(_10670_),
    .A1(net5366),
    .A2(_10667_));
 sg13g2_o21ai_1 _16753_ (.B1(net5444),
    .Y(_10671_),
    .A1(_10669_),
    .A2(_10670_));
 sg13g2_mux4_1 _16754_ (.S0(net5532),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][2] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][2] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][2] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][2] ),
    .S1(net5487),
    .X(_10672_));
 sg13g2_mux4_1 _16755_ (.S0(net5532),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][2] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][2] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][2] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][2] ),
    .S1(net5487),
    .X(_10673_));
 sg13g2_mux4_1 _16756_ (.S0(net5539),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][2] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][2] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][2] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][2] ),
    .S1(net5494),
    .X(_10674_));
 sg13g2_mux4_1 _16757_ (.S0(net5539),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][2] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][2] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][2] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][2] ),
    .S1(net5494),
    .X(_10675_));
 sg13g2_mux4_1 _16758_ (.S0(net5468),
    .A0(_10672_),
    .A1(_10673_),
    .A2(_10675_),
    .A3(_10674_),
    .S1(net5358),
    .X(_10676_));
 sg13g2_or2_1 _16759_ (.X(_10677_),
    .B(_10676_),
    .A(net5444));
 sg13g2_o21ai_1 _16760_ (.B1(_10677_),
    .Y(_10678_),
    .A1(_10666_),
    .A2(_10671_));
 sg13g2_o21ai_1 _16761_ (.B1(_10661_),
    .Y(_00261_),
    .A1(net5151),
    .A2(_10678_));
 sg13g2_nand2_1 _16762_ (.Y(_10679_),
    .A(net5818),
    .B(net5157));
 sg13g2_mux4_1 _16763_ (.S0(net5534),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][3] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][3] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][3] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][3] ),
    .S1(net5489),
    .X(_10680_));
 sg13g2_nor2_1 _16764_ (.A(net5365),
    .B(_10680_),
    .Y(_10681_));
 sg13g2_mux4_1 _16765_ (.S0(net5535),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][3] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][3] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][3] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][3] ),
    .S1(net5490),
    .X(_10682_));
 sg13g2_o21ai_1 _16766_ (.B1(net5359),
    .Y(_10683_),
    .A1(net5465),
    .A2(_10682_));
 sg13g2_nor2_1 _16767_ (.A(_10681_),
    .B(_10683_),
    .Y(_10684_));
 sg13g2_mux4_1 _16768_ (.S0(net5538),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][3] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][3] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][3] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][3] ),
    .S1(net5493),
    .X(_10685_));
 sg13g2_nor2_1 _16769_ (.A(net5465),
    .B(_10685_),
    .Y(_10686_));
 sg13g2_mux4_1 _16770_ (.S0(net5534),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][3] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][3] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][3] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][3] ),
    .S1(net5489),
    .X(_10687_));
 sg13g2_o21ai_1 _16771_ (.B1(net5454),
    .Y(_10688_),
    .A1(net5365),
    .A2(_10687_));
 sg13g2_o21ai_1 _16772_ (.B1(net5443),
    .Y(_10689_),
    .A1(_10686_),
    .A2(_10688_));
 sg13g2_mux4_1 _16773_ (.S0(net5535),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][3] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][3] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][3] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][3] ),
    .S1(net5490),
    .X(_10690_));
 sg13g2_mux4_1 _16774_ (.S0(net5534),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][3] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][3] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][3] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][3] ),
    .S1(net5489),
    .X(_10691_));
 sg13g2_mux4_1 _16775_ (.S0(net5534),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][3] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][3] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][3] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][3] ),
    .S1(net5489),
    .X(_10692_));
 sg13g2_mux4_1 _16776_ (.S0(net5534),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][3] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][3] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][3] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][3] ),
    .S1(net5489),
    .X(_10693_));
 sg13g2_mux4_1 _16777_ (.S0(net5365),
    .A0(_10690_),
    .A1(_10691_),
    .A2(_10692_),
    .A3(_10693_),
    .S1(net5454),
    .X(_10694_));
 sg13g2_or2_1 _16778_ (.X(_10695_),
    .B(_10694_),
    .A(net5443));
 sg13g2_o21ai_1 _16779_ (.B1(_10695_),
    .Y(_10696_),
    .A1(_10684_),
    .A2(_10689_));
 sg13g2_o21ai_1 _16780_ (.B1(_10679_),
    .Y(_00262_),
    .A1(net5151),
    .A2(_10696_));
 sg13g2_nand2_1 _16781_ (.Y(_10697_),
    .A(net5815),
    .B(net5157));
 sg13g2_mux4_1 _16782_ (.S0(net5560),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][4] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][4] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][4] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][4] ),
    .S1(net5515),
    .X(_10698_));
 sg13g2_nor2_1 _16783_ (.A(net5369),
    .B(_10698_),
    .Y(_10699_));
 sg13g2_mux4_1 _16784_ (.S0(net5559),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][4] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][4] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][4] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][4] ),
    .S1(net5514),
    .X(_10700_));
 sg13g2_o21ai_1 _16785_ (.B1(net5461),
    .Y(_10701_),
    .A1(net5470),
    .A2(_10700_));
 sg13g2_nor2_1 _16786_ (.A(_10699_),
    .B(_10701_),
    .Y(_10702_));
 sg13g2_mux4_1 _16787_ (.S0(net5560),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][4] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][4] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][4] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][4] ),
    .S1(net5515),
    .X(_10703_));
 sg13g2_mux4_1 _16788_ (.S0(net5560),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][4] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][4] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][4] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][4] ),
    .S1(net5515),
    .X(_10704_));
 sg13g2_nor2_1 _16789_ (.A(net5470),
    .B(_10704_),
    .Y(_10705_));
 sg13g2_o21ai_1 _16790_ (.B1(net5360),
    .Y(_10706_),
    .A1(net5371),
    .A2(_10703_));
 sg13g2_o21ai_1 _16791_ (.B1(net5449),
    .Y(_10707_),
    .A1(_10705_),
    .A2(_10706_));
 sg13g2_mux4_1 _16792_ (.S0(net5547),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][4] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][4] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][4] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][4] ),
    .S1(net5502),
    .X(_10708_));
 sg13g2_mux4_1 _16793_ (.S0(net5547),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][4] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][4] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][4] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][4] ),
    .S1(net5502),
    .X(_10709_));
 sg13g2_mux4_1 _16794_ (.S0(net5547),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][4] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][4] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][4] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][4] ),
    .S1(net5502),
    .X(_10710_));
 sg13g2_mux4_1 _16795_ (.S0(net5547),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][4] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][4] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][4] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][4] ),
    .S1(net5502),
    .X(_10711_));
 sg13g2_mux4_1 _16796_ (.S0(net5368),
    .A0(_10708_),
    .A1(_10709_),
    .A2(_10710_),
    .A3(_10711_),
    .S1(net5457),
    .X(_10712_));
 sg13g2_or2_1 _16797_ (.X(_10713_),
    .B(_10712_),
    .A(net5449));
 sg13g2_o21ai_1 _16798_ (.B1(_10713_),
    .Y(_10714_),
    .A1(_10702_),
    .A2(_10707_));
 sg13g2_o21ai_1 _16799_ (.B1(_10697_),
    .Y(_00263_),
    .A1(net5151),
    .A2(_10714_));
 sg13g2_nand2_1 _16800_ (.Y(_10715_),
    .A(net5812),
    .B(net5157));
 sg13g2_mux4_1 _16801_ (.S0(net5549),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][5] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][5] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][5] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][5] ),
    .S1(net5504),
    .X(_10716_));
 sg13g2_nor2_1 _16802_ (.A(net5369),
    .B(_10716_),
    .Y(_10717_));
 sg13g2_mux4_1 _16803_ (.S0(net5548),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][5] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][5] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][5] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][5] ),
    .S1(net5503),
    .X(_10718_));
 sg13g2_o21ai_1 _16804_ (.B1(net5457),
    .Y(_10719_),
    .A1(net5471),
    .A2(_10718_));
 sg13g2_nor2_1 _16805_ (.A(_10717_),
    .B(_10719_),
    .Y(_10720_));
 sg13g2_mux4_1 _16806_ (.S0(net5548),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][5] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][5] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][5] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][5] ),
    .S1(net5503),
    .X(_10721_));
 sg13g2_mux4_1 _16807_ (.S0(net5548),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][5] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][5] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][5] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][5] ),
    .S1(net5503),
    .X(_10722_));
 sg13g2_nor2_1 _16808_ (.A(net5469),
    .B(_10722_),
    .Y(_10723_));
 sg13g2_o21ai_1 _16809_ (.B1(net5360),
    .Y(_10724_),
    .A1(net5368),
    .A2(_10721_));
 sg13g2_o21ai_1 _16810_ (.B1(net5446),
    .Y(_10725_),
    .A1(_10723_),
    .A2(_10724_));
 sg13g2_mux4_1 _16811_ (.S0(net5546),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][5] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][5] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][5] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][5] ),
    .S1(net5501),
    .X(_10726_));
 sg13g2_mux4_1 _16812_ (.S0(net5546),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][5] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][5] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][5] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][5] ),
    .S1(net5501),
    .X(_10727_));
 sg13g2_mux4_1 _16813_ (.S0(net5546),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][5] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][5] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][5] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][5] ),
    .S1(net5501),
    .X(_10728_));
 sg13g2_mux4_1 _16814_ (.S0(net5546),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][5] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][5] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][5] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][5] ),
    .S1(net5501),
    .X(_10729_));
 sg13g2_mux4_1 _16815_ (.S0(net5368),
    .A0(_10726_),
    .A1(_10727_),
    .A2(_10728_),
    .A3(_10729_),
    .S1(net5457),
    .X(_10730_));
 sg13g2_or2_1 _16816_ (.X(_10731_),
    .B(_10730_),
    .A(net5446));
 sg13g2_o21ai_1 _16817_ (.B1(_10731_),
    .Y(_10732_),
    .A1(_10720_),
    .A2(_10725_));
 sg13g2_o21ai_1 _16818_ (.B1(_10715_),
    .Y(_00264_),
    .A1(net5151),
    .A2(_10732_));
 sg13g2_nand2_1 _16819_ (.Y(_10733_),
    .A(net5809),
    .B(net5157));
 sg13g2_mux4_1 _16820_ (.S0(net5537),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][6] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][6] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][6] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][6] ),
    .S1(net5492),
    .X(_10734_));
 sg13g2_inv_1 _16821_ (.Y(_10735_),
    .A(_10734_));
 sg13g2_mux4_1 _16822_ (.S0(net5546),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][6] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][6] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][6] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][6] ),
    .S1(net5501),
    .X(_10736_));
 sg13g2_a21oi_1 _16823_ (.A1(net5466),
    .A2(_10735_),
    .Y(_10737_),
    .B1(net5454));
 sg13g2_o21ai_1 _16824_ (.B1(_10737_),
    .Y(_10738_),
    .A1(net5466),
    .A2(_10736_));
 sg13g2_mux4_1 _16825_ (.S0(net5546),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][6] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][6] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][6] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][6] ),
    .S1(net5501),
    .X(_10739_));
 sg13g2_mux4_1 _16826_ (.S0(net5546),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][6] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][6] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][6] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][6] ),
    .S1(net5501),
    .X(_10740_));
 sg13g2_nor2_1 _16827_ (.A(net5368),
    .B(_10740_),
    .Y(_10741_));
 sg13g2_o21ai_1 _16828_ (.B1(net5457),
    .Y(_10742_),
    .A1(net5469),
    .A2(_10739_));
 sg13g2_o21ai_1 _16829_ (.B1(net5446),
    .Y(_10743_),
    .A1(_10741_),
    .A2(_10742_));
 sg13g2_nand2b_2 _16830_ (.Y(_10744_),
    .B(_10738_),
    .A_N(_10743_));
 sg13g2_mux4_1 _16831_ (.S0(net5530),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][6] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][6] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][6] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][6] ),
    .S1(net5485),
    .X(_10745_));
 sg13g2_mux4_1 _16832_ (.S0(net5530),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][6] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][6] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][6] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][6] ),
    .S1(net5485),
    .X(_10746_));
 sg13g2_mux4_1 _16833_ (.S0(net5530),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][6] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][6] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][6] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][6] ),
    .S1(net5485),
    .X(_10747_));
 sg13g2_mux4_1 _16834_ (.S0(net5530),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][6] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][6] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][6] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][6] ),
    .S1(net5485),
    .X(_10748_));
 sg13g2_mux4_1 _16835_ (.S0(net5363),
    .A0(_10745_),
    .A1(_10746_),
    .A2(_10747_),
    .A3(_10748_),
    .S1(net5452),
    .X(_10749_));
 sg13g2_o21ai_1 _16836_ (.B1(_10744_),
    .Y(_10750_),
    .A1(net5441),
    .A2(_10749_));
 sg13g2_o21ai_1 _16837_ (.B1(_10733_),
    .Y(_00265_),
    .A1(net5151),
    .A2(_10750_));
 sg13g2_nand2_1 _16838_ (.Y(_10751_),
    .A(net5806),
    .B(net5152));
 sg13g2_mux4_1 _16839_ (.S0(net5566),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][7] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][7] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][7] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][7] ),
    .S1(net5521),
    .X(_10752_));
 sg13g2_inv_1 _16840_ (.Y(_10753_),
    .A(_10752_));
 sg13g2_mux4_1 _16841_ (.S0(net5566),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][7] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][7] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][7] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][7] ),
    .S1(net5521),
    .X(_10754_));
 sg13g2_a21oi_1 _16842_ (.A1(net5474),
    .A2(_10753_),
    .Y(_10755_),
    .B1(net5459));
 sg13g2_o21ai_1 _16843_ (.B1(_10755_),
    .Y(_10756_),
    .A1(net5474),
    .A2(_10754_));
 sg13g2_mux4_1 _16844_ (.S0(net5566),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][7] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][7] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][7] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][7] ),
    .S1(net5521),
    .X(_10757_));
 sg13g2_mux4_1 _16845_ (.S0(net5566),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][7] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][7] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][7] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][7] ),
    .S1(net5521),
    .X(_10758_));
 sg13g2_nor2_1 _16846_ (.A(net5370),
    .B(_10758_),
    .Y(_10759_));
 sg13g2_o21ai_1 _16847_ (.B1(net5459),
    .Y(_10760_),
    .A1(net5474),
    .A2(_10757_));
 sg13g2_o21ai_1 _16848_ (.B1(net5448),
    .Y(_10761_),
    .A1(_10759_),
    .A2(_10760_));
 sg13g2_nand2b_2 _16849_ (.Y(_10762_),
    .B(_10756_),
    .A_N(_10761_));
 sg13g2_mux4_1 _16850_ (.S0(net5550),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][7] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][7] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][7] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][7] ),
    .S1(net5505),
    .X(_10763_));
 sg13g2_mux4_1 _16851_ (.S0(net5551),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][7] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][7] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][7] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][7] ),
    .S1(net5506),
    .X(_10764_));
 sg13g2_mux4_1 _16852_ (.S0(net5552),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][7] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][7] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][7] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][7] ),
    .S1(net5507),
    .X(_10765_));
 sg13g2_mux4_1 _16853_ (.S0(net5551),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][7] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][7] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][7] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][7] ),
    .S1(net5506),
    .X(_10766_));
 sg13g2_mux4_1 _16854_ (.S0(net5469),
    .A0(_10763_),
    .A1(_10764_),
    .A2(_10766_),
    .A3(_10765_),
    .S1(net5361),
    .X(_10767_));
 sg13g2_o21ai_1 _16855_ (.B1(_10762_),
    .Y(_10768_),
    .A1(net5447),
    .A2(_10767_));
 sg13g2_o21ai_1 _16856_ (.B1(_10751_),
    .Y(_00266_),
    .A1(net5149),
    .A2(_10768_));
 sg13g2_nand2_1 _16857_ (.Y(_10769_),
    .A(net5804),
    .B(net5155));
 sg13g2_mux4_1 _16858_ (.S0(net5558),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][8] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][8] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][8] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][8] ),
    .S1(net5513),
    .X(_10770_));
 sg13g2_mux4_1 _16859_ (.S0(net5557),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][8] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][8] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][8] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][8] ),
    .S1(net5512),
    .X(_10771_));
 sg13g2_mux2_1 _16860_ (.A0(_10770_),
    .A1(_10771_),
    .S(net5369),
    .X(_10772_));
 sg13g2_mux4_1 _16861_ (.S0(net5558),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][8] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][8] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][8] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][8] ),
    .S1(net5513),
    .X(_10773_));
 sg13g2_nor2_1 _16862_ (.A(net5471),
    .B(_10773_),
    .Y(_10774_));
 sg13g2_mux4_1 _16863_ (.S0(net5558),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][8] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][8] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][8] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][8] ),
    .S1(net5513),
    .X(_10775_));
 sg13g2_o21ai_1 _16864_ (.B1(net5458),
    .Y(_10776_),
    .A1(net5369),
    .A2(_10775_));
 sg13g2_o21ai_1 _16865_ (.B1(net5449),
    .Y(_10777_),
    .A1(_10774_),
    .A2(_10776_));
 sg13g2_a21o_2 _16866_ (.A2(_10772_),
    .A1(net5360),
    .B1(_10777_),
    .X(_10778_));
 sg13g2_mux4_1 _16867_ (.S0(net5537),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][8] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][8] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][8] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][8] ),
    .S1(net5492),
    .X(_10779_));
 sg13g2_mux4_1 _16868_ (.S0(net5537),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][8] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][8] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][8] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][8] ),
    .S1(net5492),
    .X(_10780_));
 sg13g2_mux4_1 _16869_ (.S0(net5537),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][8] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][8] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][8] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][8] ),
    .S1(net5492),
    .X(_10781_));
 sg13g2_mux4_1 _16870_ (.S0(net5537),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][8] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][8] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][8] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][8] ),
    .S1(net5492),
    .X(_10782_));
 sg13g2_mux4_1 _16871_ (.S0(net5366),
    .A0(_10779_),
    .A1(_10780_),
    .A2(_10781_),
    .A3(_10782_),
    .S1(net5454),
    .X(_10783_));
 sg13g2_o21ai_1 _16872_ (.B1(_10778_),
    .Y(_10784_),
    .A1(net5443),
    .A2(_10783_));
 sg13g2_o21ai_1 _16873_ (.B1(_10769_),
    .Y(_00267_),
    .A1(net5150),
    .A2(_10784_));
 sg13g2_nand2_1 _16874_ (.Y(_10785_),
    .A(net5802),
    .B(net5155));
 sg13g2_mux4_1 _16875_ (.S0(net5529),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][9] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][9] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][9] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][9] ),
    .S1(net5484),
    .X(_10786_));
 sg13g2_inv_1 _16876_ (.Y(_10787_),
    .A(_10786_));
 sg13g2_mux4_1 _16877_ (.S0(net5531),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][9] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][9] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][9] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][9] ),
    .S1(net5486),
    .X(_10788_));
 sg13g2_a21oi_1 _16878_ (.A1(net5463),
    .A2(_10787_),
    .Y(_10789_),
    .B1(net5452));
 sg13g2_o21ai_1 _16879_ (.B1(_10789_),
    .Y(_10790_),
    .A1(net5463),
    .A2(_10788_));
 sg13g2_mux4_1 _16880_ (.S0(net5531),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][9] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][9] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][9] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][9] ),
    .S1(net5486),
    .X(_10791_));
 sg13g2_mux4_1 _16881_ (.S0(net5531),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][9] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][9] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][9] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][9] ),
    .S1(net5486),
    .X(_10792_));
 sg13g2_nor2_1 _16882_ (.A(net5363),
    .B(_10792_),
    .Y(_10793_));
 sg13g2_o21ai_1 _16883_ (.B1(net5452),
    .Y(_10794_),
    .A1(net5463),
    .A2(_10791_));
 sg13g2_o21ai_1 _16884_ (.B1(net5441),
    .Y(_10795_),
    .A1(_10793_),
    .A2(_10794_));
 sg13g2_nand2b_1 _16885_ (.Y(_10796_),
    .B(_10790_),
    .A_N(_10795_));
 sg13g2_mux4_1 _16886_ (.S0(net5532),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][9] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][9] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][9] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][9] ),
    .S1(net5487),
    .X(_10797_));
 sg13g2_mux4_1 _16887_ (.S0(net5541),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][9] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][9] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][9] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][9] ),
    .S1(net5496),
    .X(_10798_));
 sg13g2_mux4_1 _16888_ (.S0(net5539),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][9] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][9] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][9] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][9] ),
    .S1(net5494),
    .X(_10799_));
 sg13g2_mux4_1 _16889_ (.S0(net5539),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][9] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][9] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][9] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][9] ),
    .S1(net5494),
    .X(_10800_));
 sg13g2_mux4_1 _16890_ (.S0(net5466),
    .A0(_10797_),
    .A1(_10798_),
    .A2(_10800_),
    .A3(_10799_),
    .S1(net5359),
    .X(_10801_));
 sg13g2_o21ai_1 _16891_ (.B1(_10796_),
    .Y(_10802_),
    .A1(net5441),
    .A2(_10801_));
 sg13g2_o21ai_1 _16892_ (.B1(_10785_),
    .Y(_00268_),
    .A1(net5150),
    .A2(_10802_));
 sg13g2_nand2_1 _16893_ (.Y(_10803_),
    .A(net5799),
    .B(net5154));
 sg13g2_mux4_1 _16894_ (.S0(net5562),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][10] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][10] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][10] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][10] ),
    .S1(net5517),
    .X(_10804_));
 sg13g2_nor2_1 _16895_ (.A(net5370),
    .B(_10804_),
    .Y(_10805_));
 sg13g2_mux4_1 _16896_ (.S0(net5562),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][10] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][10] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][10] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][10] ),
    .S1(net5517),
    .X(_10806_));
 sg13g2_o21ai_1 _16897_ (.B1(net5360),
    .Y(_10807_),
    .A1(net5472),
    .A2(_10806_));
 sg13g2_nor2_1 _16898_ (.A(_10805_),
    .B(_10807_),
    .Y(_10808_));
 sg13g2_mux4_1 _16899_ (.S0(net5564),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][10] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][10] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][10] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][10] ),
    .S1(net5519),
    .X(_10809_));
 sg13g2_nor2_1 _16900_ (.A(net5472),
    .B(_10809_),
    .Y(_10810_));
 sg13g2_mux4_1 _16901_ (.S0(net5564),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][10] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][10] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][10] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][10] ),
    .S1(net5519),
    .X(_10811_));
 sg13g2_o21ai_1 _16902_ (.B1(net5460),
    .Y(_10812_),
    .A1(net5370),
    .A2(_10811_));
 sg13g2_o21ai_1 _16903_ (.B1(net5448),
    .Y(_10813_),
    .A1(_10810_),
    .A2(_10812_));
 sg13g2_mux4_1 _16904_ (.S0(net5553),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][10] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][10] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][10] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][10] ),
    .S1(net5508),
    .X(_10814_));
 sg13g2_mux4_1 _16905_ (.S0(net5553),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][10] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][10] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][10] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][10] ),
    .S1(net5508),
    .X(_10815_));
 sg13g2_mux4_1 _16906_ (.S0(net5553),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][10] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][10] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][10] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][10] ),
    .S1(net5508),
    .X(_10816_));
 sg13g2_mux4_1 _16907_ (.S0(net5553),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][10] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][10] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][10] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][10] ),
    .S1(net5508),
    .X(_10817_));
 sg13g2_mux4_1 _16908_ (.S0(net5469),
    .A0(_10814_),
    .A1(_10815_),
    .A2(_10817_),
    .A3(_10816_),
    .S1(net5360),
    .X(_10818_));
 sg13g2_or2_1 _16909_ (.X(_10819_),
    .B(_10818_),
    .A(net5448));
 sg13g2_o21ai_1 _16910_ (.B1(_10819_),
    .Y(_10820_),
    .A1(_10808_),
    .A2(_10813_));
 sg13g2_o21ai_1 _16911_ (.B1(_10803_),
    .Y(_00269_),
    .A1(net5147),
    .A2(_10820_));
 sg13g2_nand2_1 _16912_ (.Y(_10821_),
    .A(net1919),
    .B(net5155));
 sg13g2_mux4_1 _16913_ (.S0(net5532),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][11] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][11] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][11] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][11] ),
    .S1(net5487),
    .X(_10822_));
 sg13g2_nor2_1 _16914_ (.A(net5363),
    .B(_10822_),
    .Y(_10823_));
 sg13g2_mux4_1 _16915_ (.S0(net5532),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][11] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][11] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][11] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][11] ),
    .S1(net5487),
    .X(_10824_));
 sg13g2_o21ai_1 _16916_ (.B1(net5452),
    .Y(_10825_),
    .A1(net5463),
    .A2(_10824_));
 sg13g2_nor2_1 _16917_ (.A(_10823_),
    .B(_10825_),
    .Y(_10826_));
 sg13g2_mux4_1 _16918_ (.S0(net5529),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][11] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][11] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][11] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][11] ),
    .S1(net5484),
    .X(_10827_));
 sg13g2_nor2_1 _16919_ (.A(net5363),
    .B(_10827_),
    .Y(_10828_));
 sg13g2_mux4_1 _16920_ (.S0(net5529),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][11] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][11] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][11] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][11] ),
    .S1(net5484),
    .X(_10829_));
 sg13g2_o21ai_1 _16921_ (.B1(net5358),
    .Y(_10830_),
    .A1(net5463),
    .A2(_10829_));
 sg13g2_o21ai_1 _16922_ (.B1(net5441),
    .Y(_10831_),
    .A1(_10828_),
    .A2(_10830_));
 sg13g2_mux4_1 _16923_ (.S0(net5528),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][11] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][11] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][11] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][11] ),
    .S1(net5483),
    .X(_10832_));
 sg13g2_mux4_1 _16924_ (.S0(net5529),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][11] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][11] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][11] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][11] ),
    .S1(net5484),
    .X(_10833_));
 sg13g2_mux4_1 _16925_ (.S0(net5528),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][11] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][11] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][11] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][11] ),
    .S1(net5483),
    .X(_10834_));
 sg13g2_mux4_1 _16926_ (.S0(net5528),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][11] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][11] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][11] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][11] ),
    .S1(net5483),
    .X(_10835_));
 sg13g2_mux4_1 _16927_ (.S0(net5363),
    .A0(_10832_),
    .A1(_10833_),
    .A2(_10834_),
    .A3(_10835_),
    .S1(net5452),
    .X(_10836_));
 sg13g2_or2_1 _16928_ (.X(_10837_),
    .B(_10836_),
    .A(net5441));
 sg13g2_o21ai_1 _16929_ (.B1(_10837_),
    .Y(_10838_),
    .A1(_10826_),
    .A2(_10831_));
 sg13g2_o21ai_1 _16930_ (.B1(_10821_),
    .Y(_00270_),
    .A1(net5149),
    .A2(_10838_));
 sg13g2_nand2_1 _16931_ (.Y(_10839_),
    .A(net5796),
    .B(net5155));
 sg13g2_mux4_1 _16932_ (.S0(net5565),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][12] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][12] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][12] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][12] ),
    .S1(net5520),
    .X(_10840_));
 sg13g2_inv_1 _16933_ (.Y(_10841_),
    .A(_10840_));
 sg13g2_mux4_1 _16934_ (.S0(net5565),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][12] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][12] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][12] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][12] ),
    .S1(net5520),
    .X(_10842_));
 sg13g2_a21oi_1 _16935_ (.A1(net5475),
    .A2(_10841_),
    .Y(_10843_),
    .B1(net5459));
 sg13g2_o21ai_1 _16936_ (.B1(_10843_),
    .Y(_10844_),
    .A1(net5475),
    .A2(_10842_));
 sg13g2_mux4_1 _16937_ (.S0(net5565),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][12] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][12] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][12] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][12] ),
    .S1(net5520),
    .X(_10845_));
 sg13g2_mux4_1 _16938_ (.S0(net5565),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][12] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][12] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][12] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][12] ),
    .S1(net5520),
    .X(_10846_));
 sg13g2_nor2_1 _16939_ (.A(net5370),
    .B(_10846_),
    .Y(_10847_));
 sg13g2_o21ai_1 _16940_ (.B1(net5459),
    .Y(_10848_),
    .A1(net5475),
    .A2(_10845_));
 sg13g2_o21ai_1 _16941_ (.B1(net5448),
    .Y(_10849_),
    .A1(_10847_),
    .A2(_10848_));
 sg13g2_nand2b_2 _16942_ (.Y(_10850_),
    .B(_10844_),
    .A_N(_10849_));
 sg13g2_mux4_1 _16943_ (.S0(net5550),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][12] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][12] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][12] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][12] ),
    .S1(net5505),
    .X(_10851_));
 sg13g2_mux4_1 _16944_ (.S0(net5550),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][12] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][12] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][12] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][12] ),
    .S1(net5505),
    .X(_10852_));
 sg13g2_mux4_1 _16945_ (.S0(net5550),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][12] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][12] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][12] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][12] ),
    .S1(net5505),
    .X(_10853_));
 sg13g2_mux4_1 _16946_ (.S0(net5550),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][12] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][12] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][12] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][12] ),
    .S1(net5505),
    .X(_10854_));
 sg13g2_mux4_1 _16947_ (.S0(net5372),
    .A0(_10851_),
    .A1(_10852_),
    .A2(_10853_),
    .A3(_10854_),
    .S1(net5462),
    .X(_10855_));
 sg13g2_o21ai_1 _16948_ (.B1(_10850_),
    .Y(_10856_),
    .A1(net5447),
    .A2(_10855_));
 sg13g2_o21ai_1 _16949_ (.B1(_10839_),
    .Y(_00271_),
    .A1(net5149),
    .A2(_10856_));
 sg13g2_nand2_1 _16950_ (.Y(_10857_),
    .A(net5793),
    .B(net5154));
 sg13g2_mux4_1 _16951_ (.S0(net5540),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][13] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][13] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][13] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][13] ),
    .S1(net5495),
    .X(_10858_));
 sg13g2_nor2_1 _16952_ (.A(net5363),
    .B(_10858_),
    .Y(_10859_));
 sg13g2_mux4_1 _16953_ (.S0(net5539),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][13] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][13] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][13] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][13] ),
    .S1(net5494),
    .X(_10860_));
 sg13g2_o21ai_1 _16954_ (.B1(net5452),
    .Y(_10861_),
    .A1(net5463),
    .A2(_10860_));
 sg13g2_nor2_1 _16955_ (.A(_10859_),
    .B(_10861_),
    .Y(_10862_));
 sg13g2_mux4_1 _16956_ (.S0(net5541),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][13] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][13] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][13] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][13] ),
    .S1(net5496),
    .X(_10863_));
 sg13g2_mux4_1 _16957_ (.S0(net5531),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][13] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][13] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][13] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][13] ),
    .S1(net5486),
    .X(_10864_));
 sg13g2_nor2_1 _16958_ (.A(net5463),
    .B(_10864_),
    .Y(_10865_));
 sg13g2_o21ai_1 _16959_ (.B1(net5358),
    .Y(_10866_),
    .A1(net5363),
    .A2(_10863_));
 sg13g2_o21ai_1 _16960_ (.B1(net5441),
    .Y(_10867_),
    .A1(_10865_),
    .A2(_10866_));
 sg13g2_mux4_1 _16961_ (.S0(net5528),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][13] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][13] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][13] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][13] ),
    .S1(net5483),
    .X(_10868_));
 sg13g2_mux4_1 _16962_ (.S0(net5530),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][13] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][13] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][13] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][13] ),
    .S1(net5485),
    .X(_10869_));
 sg13g2_mux4_1 _16963_ (.S0(net5528),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][13] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][13] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][13] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][13] ),
    .S1(net5483),
    .X(_10870_));
 sg13g2_mux4_1 _16964_ (.S0(net5530),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][13] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][13] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][13] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][13] ),
    .S1(net5485),
    .X(_10871_));
 sg13g2_mux4_1 _16965_ (.S0(net5363),
    .A0(_10868_),
    .A1(_10869_),
    .A2(_10870_),
    .A3(_10871_),
    .S1(net5452),
    .X(_10872_));
 sg13g2_or2_1 _16966_ (.X(_10873_),
    .B(_10872_),
    .A(net5441));
 sg13g2_o21ai_1 _16967_ (.B1(_10873_),
    .Y(_10874_),
    .A1(_10862_),
    .A2(_10867_));
 sg13g2_o21ai_1 _16968_ (.B1(_10857_),
    .Y(_00272_),
    .A1(net5147),
    .A2(_10874_));
 sg13g2_nand2_1 _16969_ (.Y(_10875_),
    .A(net5790),
    .B(net5154));
 sg13g2_mux4_1 _16970_ (.S0(net5525),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][14] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][14] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][14] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][14] ),
    .S1(net5480),
    .X(_10876_));
 sg13g2_inv_1 _16971_ (.Y(_10877_),
    .A(_10876_));
 sg13g2_mux4_1 _16972_ (.S0(net5525),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][14] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][14] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][14] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][14] ),
    .S1(net5480),
    .X(_10878_));
 sg13g2_a21oi_1 _16973_ (.A1(net5464),
    .A2(_10877_),
    .Y(_10879_),
    .B1(net5453));
 sg13g2_o21ai_1 _16974_ (.B1(_10879_),
    .Y(_10880_),
    .A1(net5464),
    .A2(_10878_));
 sg13g2_mux4_1 _16975_ (.S0(net5525),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][14] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][14] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][14] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][14] ),
    .S1(net5480),
    .X(_10881_));
 sg13g2_mux4_1 _16976_ (.S0(net5525),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][14] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][14] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][14] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][14] ),
    .S1(net5480),
    .X(_10882_));
 sg13g2_nor2_1 _16977_ (.A(net5362),
    .B(_10882_),
    .Y(_10883_));
 sg13g2_o21ai_1 _16978_ (.B1(net5453),
    .Y(_10884_),
    .A1(net5464),
    .A2(_10881_));
 sg13g2_o21ai_1 _16979_ (.B1(net5442),
    .Y(_10885_),
    .A1(_10883_),
    .A2(_10884_));
 sg13g2_nand2b_1 _16980_ (.Y(_10886_),
    .B(_10880_),
    .A_N(_10885_));
 sg13g2_mux4_1 _16981_ (.S0(net5534),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][14] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][14] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][14] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][14] ),
    .S1(net5489),
    .X(_10887_));
 sg13g2_mux4_1 _16982_ (.S0(net5526),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][14] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][14] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][14] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][14] ),
    .S1(net5481),
    .X(_10888_));
 sg13g2_mux4_1 _16983_ (.S0(net5525),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][14] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][14] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][14] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][14] ),
    .S1(net5480),
    .X(_10889_));
 sg13g2_mux4_1 _16984_ (.S0(net5524),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][14] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][14] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][14] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][14] ),
    .S1(net5479),
    .X(_10890_));
 sg13g2_mux4_1 _16985_ (.S0(net5362),
    .A0(_10887_),
    .A1(_10888_),
    .A2(_10889_),
    .A3(_10890_),
    .S1(net5453),
    .X(_10891_));
 sg13g2_o21ai_1 _16986_ (.B1(_10886_),
    .Y(_10892_),
    .A1(net5442),
    .A2(_10891_));
 sg13g2_o21ai_1 _16987_ (.B1(_10875_),
    .Y(_00273_),
    .A1(net5147),
    .A2(_10892_));
 sg13g2_nand2_1 _16988_ (.Y(_10893_),
    .A(net5789),
    .B(net5152));
 sg13g2_mux4_1 _16989_ (.S0(net5566),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][15] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][15] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][15] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][15] ),
    .S1(net5521),
    .X(_10894_));
 sg13g2_inv_1 _16990_ (.Y(_10895_),
    .A(_10894_));
 sg13g2_mux4_1 _16991_ (.S0(net5565),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][15] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][15] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][15] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][15] ),
    .S1(net5520),
    .X(_10896_));
 sg13g2_a21oi_1 _16992_ (.A1(net5475),
    .A2(_10895_),
    .Y(_10897_),
    .B1(net5459));
 sg13g2_o21ai_1 _16993_ (.B1(_10897_),
    .Y(_10898_),
    .A1(net5475),
    .A2(_10896_));
 sg13g2_mux4_1 _16994_ (.S0(net5565),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][15] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][15] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][15] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][15] ),
    .S1(net5520),
    .X(_10899_));
 sg13g2_mux4_1 _16995_ (.S0(net5559),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][15] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][15] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][15] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][15] ),
    .S1(net5514),
    .X(_10900_));
 sg13g2_nor2_1 _16996_ (.A(net5371),
    .B(_10900_),
    .Y(_10901_));
 sg13g2_o21ai_1 _16997_ (.B1(net5459),
    .Y(_10902_),
    .A1(net5475),
    .A2(_10899_));
 sg13g2_o21ai_1 _16998_ (.B1(net5450),
    .Y(_10903_),
    .A1(_10901_),
    .A2(_10902_));
 sg13g2_nand2b_2 _16999_ (.Y(_10904_),
    .B(_10898_),
    .A_N(_10903_));
 sg13g2_mux4_1 _17000_ (.S0(net5553),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][15] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][15] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][15] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][15] ),
    .S1(net5508),
    .X(_10905_));
 sg13g2_mux4_1 _17001_ (.S0(net5553),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][15] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][15] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][15] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][15] ),
    .S1(net5508),
    .X(_10906_));
 sg13g2_mux4_1 _17002_ (.S0(net5553),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][15] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][15] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][15] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][15] ),
    .S1(net5508),
    .X(_10907_));
 sg13g2_mux4_1 _17003_ (.S0(net5553),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][15] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][15] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][15] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][15] ),
    .S1(net5508),
    .X(_10908_));
 sg13g2_mux4_1 _17004_ (.S0(net5469),
    .A0(_10905_),
    .A1(_10906_),
    .A2(_10908_),
    .A3(_10907_),
    .S1(net5360),
    .X(_10909_));
 sg13g2_o21ai_1 _17005_ (.B1(_10904_),
    .Y(_10910_),
    .A1(net5447),
    .A2(_10909_));
 sg13g2_o21ai_1 _17006_ (.B1(_10893_),
    .Y(_00274_),
    .A1(net5147),
    .A2(_10910_));
 sg13g2_nand2_1 _17007_ (.Y(_10911_),
    .A(net3641),
    .B(net5154));
 sg13g2_mux4_1 _17008_ (.S0(net5562),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][16] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][16] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][16] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][16] ),
    .S1(net5517),
    .X(_10912_));
 sg13g2_inv_1 _17009_ (.Y(_10913_),
    .A(_10912_));
 sg13g2_mux4_1 _17010_ (.S0(net5562),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][16] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][16] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][16] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][16] ),
    .S1(net5517),
    .X(_10914_));
 sg13g2_a21oi_1 _17011_ (.A1(net5472),
    .A2(_10913_),
    .Y(_10915_),
    .B1(net5460));
 sg13g2_o21ai_1 _17012_ (.B1(_10915_),
    .Y(_10916_),
    .A1(net5472),
    .A2(_10914_));
 sg13g2_mux4_1 _17013_ (.S0(net5562),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][16] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][16] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][16] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][16] ),
    .S1(net5517),
    .X(_10917_));
 sg13g2_mux4_1 _17014_ (.S0(net5562),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][16] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][16] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][16] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][16] ),
    .S1(net5517),
    .X(_10918_));
 sg13g2_nor2_1 _17015_ (.A(net5370),
    .B(_10918_),
    .Y(_10919_));
 sg13g2_o21ai_1 _17016_ (.B1(net5460),
    .Y(_10920_),
    .A1(net5472),
    .A2(_10917_));
 sg13g2_o21ai_1 _17017_ (.B1(net5448),
    .Y(_10921_),
    .A1(_10919_),
    .A2(_10920_));
 sg13g2_nand2b_2 _17018_ (.Y(_10922_),
    .B(_10916_),
    .A_N(_10921_));
 sg13g2_mux4_1 _17019_ (.S0(net5542),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][16] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][16] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][16] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][16] ),
    .S1(net5497),
    .X(_10923_));
 sg13g2_mux4_1 _17020_ (.S0(net5542),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][16] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][16] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][16] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][16] ),
    .S1(net5497),
    .X(_10924_));
 sg13g2_mux4_1 _17021_ (.S0(net5542),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][16] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][16] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][16] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][16] ),
    .S1(net5497),
    .X(_10925_));
 sg13g2_mux4_1 _17022_ (.S0(net5542),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][16] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][16] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][16] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][16] ),
    .S1(net5497),
    .X(_10926_));
 sg13g2_mux4_1 _17023_ (.S0(net5366),
    .A0(_10923_),
    .A1(_10924_),
    .A2(_10925_),
    .A3(_10926_),
    .S1(net5455),
    .X(_10927_));
 sg13g2_o21ai_1 _17024_ (.B1(_10922_),
    .Y(_10928_),
    .A1(net5443),
    .A2(_10927_));
 sg13g2_o21ai_1 _17025_ (.B1(_10911_),
    .Y(_00275_),
    .A1(net5147),
    .A2(_10928_));
 sg13g2_nand2_1 _17026_ (.Y(_10929_),
    .A(net5785),
    .B(net5154));
 sg13g2_mux4_1 _17027_ (.S0(net5526),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][17] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][17] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][17] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][17] ),
    .S1(net5481),
    .X(_10930_));
 sg13g2_mux4_1 _17028_ (.S0(net5526),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][17] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][17] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][17] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][17] ),
    .S1(net5481),
    .X(_10931_));
 sg13g2_mux2_1 _17029_ (.A0(_10930_),
    .A1(_10931_),
    .S(net5362),
    .X(_10932_));
 sg13g2_mux4_1 _17030_ (.S0(net5526),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][17] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][17] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][17] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][17] ),
    .S1(net5481),
    .X(_10933_));
 sg13g2_nor2_1 _17031_ (.A(net5464),
    .B(_10933_),
    .Y(_10934_));
 sg13g2_mux4_1 _17032_ (.S0(net5526),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][17] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][17] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][17] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][17] ),
    .S1(net5481),
    .X(_10935_));
 sg13g2_o21ai_1 _17033_ (.B1(net5453),
    .Y(_10936_),
    .A1(net5362),
    .A2(_10935_));
 sg13g2_o21ai_1 _17034_ (.B1(net5442),
    .Y(_10937_),
    .A1(_10934_),
    .A2(_10936_));
 sg13g2_a21o_1 _17035_ (.A2(_10932_),
    .A1(net5358),
    .B1(_10937_),
    .X(_10938_));
 sg13g2_mux4_1 _17036_ (.S0(net5524),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][17] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][17] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][17] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][17] ),
    .S1(net5479),
    .X(_10939_));
 sg13g2_mux4_1 _17037_ (.S0(net5524),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][17] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][17] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][17] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][17] ),
    .S1(net5479),
    .X(_10940_));
 sg13g2_mux4_1 _17038_ (.S0(net5524),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][17] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][17] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][17] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][17] ),
    .S1(net5479),
    .X(_10941_));
 sg13g2_mux4_1 _17039_ (.S0(net5525),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][17] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][17] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][17] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][17] ),
    .S1(net5480),
    .X(_10942_));
 sg13g2_mux4_1 _17040_ (.S0(net5464),
    .A0(_10939_),
    .A1(_10940_),
    .A2(_10942_),
    .A3(_10941_),
    .S1(net5358),
    .X(_10943_));
 sg13g2_o21ai_1 _17041_ (.B1(_10938_),
    .Y(_10944_),
    .A1(net5442),
    .A2(_10943_));
 sg13g2_o21ai_1 _17042_ (.B1(_10929_),
    .Y(_00276_),
    .A1(net5147),
    .A2(_10944_));
 sg13g2_nand2_1 _17043_ (.Y(_10945_),
    .A(net5782),
    .B(net5153));
 sg13g2_mux4_1 _17044_ (.S0(net5567),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][18] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][18] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][18] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][18] ),
    .S1(net5522),
    .X(_10946_));
 sg13g2_inv_1 _17045_ (.Y(_10947_),
    .A(_10946_));
 sg13g2_mux4_1 _17046_ (.S0(net5566),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][18] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][18] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][18] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][18] ),
    .S1(net5521),
    .X(_10948_));
 sg13g2_a21oi_1 _17047_ (.A1(net5474),
    .A2(_10947_),
    .Y(_10949_),
    .B1(net5461));
 sg13g2_o21ai_1 _17048_ (.B1(_10949_),
    .Y(_10950_),
    .A1(net5476),
    .A2(_10948_));
 sg13g2_mux4_1 _17049_ (.S0(net5566),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][18] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][18] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][18] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][18] ),
    .S1(net5521),
    .X(_10951_));
 sg13g2_mux4_1 _17050_ (.S0(net5567),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][18] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][18] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][18] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][18] ),
    .S1(net5522),
    .X(_10952_));
 sg13g2_nor2_1 _17051_ (.A(net5371),
    .B(_10952_),
    .Y(_10953_));
 sg13g2_o21ai_1 _17052_ (.B1(net5461),
    .Y(_10954_),
    .A1(net5474),
    .A2(_10951_));
 sg13g2_o21ai_1 _17053_ (.B1(net5448),
    .Y(_10955_),
    .A1(_10953_),
    .A2(_10954_));
 sg13g2_nand2b_2 _17054_ (.Y(_10956_),
    .B(_10950_),
    .A_N(_10955_));
 sg13g2_mux4_1 _17055_ (.S0(net5552),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][18] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][18] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][18] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][18] ),
    .S1(net5507),
    .X(_10957_));
 sg13g2_mux4_1 _17056_ (.S0(net5554),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][18] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][18] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][18] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][18] ),
    .S1(net5509),
    .X(_10958_));
 sg13g2_mux4_1 _17057_ (.S0(net5552),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][18] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][18] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][18] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][18] ),
    .S1(net5507),
    .X(_10959_));
 sg13g2_mux4_1 _17058_ (.S0(net5552),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][18] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][18] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][18] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][18] ),
    .S1(net5507),
    .X(_10960_));
 sg13g2_mux4_1 _17059_ (.S0(net5469),
    .A0(_10957_),
    .A1(_10958_),
    .A2(_10960_),
    .A3(_10959_),
    .S1(net5361),
    .X(_10961_));
 sg13g2_o21ai_1 _17060_ (.B1(_10956_),
    .Y(_10962_),
    .A1(net5447),
    .A2(_10961_));
 sg13g2_o21ai_1 _17061_ (.B1(_10945_),
    .Y(_00277_),
    .A1(net5149),
    .A2(_10962_));
 sg13g2_nand2_1 _17062_ (.Y(_10963_),
    .A(net5780),
    .B(net5152));
 sg13g2_mux4_1 _17063_ (.S0(net5536),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][19] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][19] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][19] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][19] ),
    .S1(net5491),
    .X(_10964_));
 sg13g2_nor2_1 _17064_ (.A(net5365),
    .B(_10964_),
    .Y(_10965_));
 sg13g2_mux4_1 _17065_ (.S0(net5536),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][19] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][19] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][19] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][19] ),
    .S1(net5491),
    .X(_10966_));
 sg13g2_o21ai_1 _17066_ (.B1(net5454),
    .Y(_10967_),
    .A1(net5465),
    .A2(_10966_));
 sg13g2_nor2_1 _17067_ (.A(_10965_),
    .B(_10967_),
    .Y(_10968_));
 sg13g2_mux4_1 _17068_ (.S0(net5536),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][19] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][19] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][19] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][19] ),
    .S1(net5491),
    .X(_10969_));
 sg13g2_nor2_1 _17069_ (.A(net5365),
    .B(_10969_),
    .Y(_10970_));
 sg13g2_mux4_1 _17070_ (.S0(net5536),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][19] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][19] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][19] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][19] ),
    .S1(net5491),
    .X(_10971_));
 sg13g2_o21ai_1 _17071_ (.B1(net5359),
    .Y(_10972_),
    .A1(net5466),
    .A2(_10971_));
 sg13g2_o21ai_1 _17072_ (.B1(net5443),
    .Y(_10973_),
    .A1(_10970_),
    .A2(_10972_));
 sg13g2_mux4_1 _17073_ (.S0(net5536),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][19] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][19] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][19] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][19] ),
    .S1(net5491),
    .X(_10974_));
 sg13g2_mux4_1 _17074_ (.S0(net5536),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][19] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][19] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][19] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][19] ),
    .S1(net5491),
    .X(_10975_));
 sg13g2_mux4_1 _17075_ (.S0(net5536),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][19] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][19] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][19] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][19] ),
    .S1(net5491),
    .X(_10976_));
 sg13g2_mux4_1 _17076_ (.S0(net5536),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][19] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][19] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][19] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][19] ),
    .S1(net5491),
    .X(_10977_));
 sg13g2_mux4_1 _17077_ (.S0(net5365),
    .A0(_10974_),
    .A1(_10975_),
    .A2(_10976_),
    .A3(_10977_),
    .S1(net5454),
    .X(_10978_));
 sg13g2_or2_1 _17078_ (.X(_10979_),
    .B(_10978_),
    .A(net5443));
 sg13g2_o21ai_1 _17079_ (.B1(_10979_),
    .Y(_10980_),
    .A1(_10968_),
    .A2(_10973_));
 sg13g2_o21ai_1 _17080_ (.B1(_10963_),
    .Y(_00278_),
    .A1(net5148),
    .A2(_10980_));
 sg13g2_nand2_1 _17081_ (.Y(_10981_),
    .A(net5777),
    .B(net5154));
 sg13g2_mux4_1 _17082_ (.S0(net5560),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][20] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][20] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][20] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][20] ),
    .S1(net5515),
    .X(_10982_));
 sg13g2_inv_1 _17083_ (.Y(_10983_),
    .A(_10982_));
 sg13g2_mux4_1 _17084_ (.S0(net5560),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][20] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][20] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][20] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][20] ),
    .S1(net5515),
    .X(_10984_));
 sg13g2_a21oi_1 _17085_ (.A1(net5470),
    .A2(_10983_),
    .Y(_10985_),
    .B1(net5461));
 sg13g2_o21ai_1 _17086_ (.B1(_10985_),
    .Y(_10986_),
    .A1(net5470),
    .A2(_10984_));
 sg13g2_mux4_1 _17087_ (.S0(net5560),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][20] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][20] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][20] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][20] ),
    .S1(net5515),
    .X(_10987_));
 sg13g2_nor2_1 _17088_ (.A(net5470),
    .B(_10987_),
    .Y(_10988_));
 sg13g2_mux4_1 _17089_ (.S0(net5560),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][20] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][20] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][20] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][20] ),
    .S1(net5515),
    .X(_10989_));
 sg13g2_o21ai_1 _17090_ (.B1(net5461),
    .Y(_10990_),
    .A1(net5371),
    .A2(_10989_));
 sg13g2_o21ai_1 _17091_ (.B1(net5449),
    .Y(_10991_),
    .A1(_10988_),
    .A2(_10990_));
 sg13g2_nand2b_2 _17092_ (.Y(_10992_),
    .B(_10986_),
    .A_N(_10991_));
 sg13g2_mux4_1 _17093_ (.S0(net5545),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][20] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][20] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][20] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][20] ),
    .S1(net5500),
    .X(_10993_));
 sg13g2_mux4_1 _17094_ (.S0(net5545),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][20] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][20] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][20] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][20] ),
    .S1(net5500),
    .X(_10994_));
 sg13g2_mux4_1 _17095_ (.S0(net5545),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][20] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][20] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][20] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][20] ),
    .S1(net5500),
    .X(_10995_));
 sg13g2_mux4_1 _17096_ (.S0(net5545),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][20] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][20] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][20] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][20] ),
    .S1(net5500),
    .X(_10996_));
 sg13g2_mux4_1 _17097_ (.S0(net5368),
    .A0(_10993_),
    .A1(_10994_),
    .A2(_10995_),
    .A3(_10996_),
    .S1(net5457),
    .X(_10997_));
 sg13g2_o21ai_1 _17098_ (.B1(_10992_),
    .Y(_10998_),
    .A1(net5446),
    .A2(_10997_));
 sg13g2_o21ai_1 _17099_ (.B1(_10981_),
    .Y(_00279_),
    .A1(net5147),
    .A2(_10998_));
 sg13g2_nand2_1 _17100_ (.Y(_02536_),
    .A(net5776),
    .B(net5152));
 sg13g2_mux4_1 _17101_ (.S0(net5534),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][21] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][21] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][21] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][21] ),
    .S1(net5489),
    .X(_02537_));
 sg13g2_nor2_1 _17102_ (.A(net5365),
    .B(_02537_),
    .Y(_02538_));
 sg13g2_mux4_1 _17103_ (.S0(net5538),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][21] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][21] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][21] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][21] ),
    .S1(net5493),
    .X(_02539_));
 sg13g2_o21ai_1 _17104_ (.B1(net5453),
    .Y(_02540_),
    .A1(net5465),
    .A2(_02539_));
 sg13g2_nor2_1 _17105_ (.A(_02538_),
    .B(_02540_),
    .Y(_02541_));
 sg13g2_mux4_1 _17106_ (.S0(net5526),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][21] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][21] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][21] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][21] ),
    .S1(net5481),
    .X(_02542_));
 sg13g2_mux4_1 _17107_ (.S0(net5525),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][21] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][21] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][21] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][21] ),
    .S1(net5480),
    .X(_02543_));
 sg13g2_nor2_1 _17108_ (.A(net5464),
    .B(_02543_),
    .Y(_02544_));
 sg13g2_o21ai_1 _17109_ (.B1(net5358),
    .Y(_02545_),
    .A1(net5362),
    .A2(_02542_));
 sg13g2_o21ai_1 _17110_ (.B1(net5442),
    .Y(_02546_),
    .A1(_02544_),
    .A2(_02545_));
 sg13g2_mux4_1 _17111_ (.S0(net5527),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][21] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][21] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][21] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][21] ),
    .S1(net5482),
    .X(_02547_));
 sg13g2_mux4_1 _17112_ (.S0(net5534),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][21] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][21] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][21] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][21] ),
    .S1(net5489),
    .X(_02548_));
 sg13g2_mux4_1 _17113_ (.S0(net5524),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][21] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][21] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][21] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][21] ),
    .S1(net5479),
    .X(_02549_));
 sg13g2_mux4_1 _17114_ (.S0(net5525),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][21] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][21] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][21] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][21] ),
    .S1(net5480),
    .X(_02550_));
 sg13g2_mux4_1 _17115_ (.S0(net5364),
    .A0(_02547_),
    .A1(_02548_),
    .A2(_02549_),
    .A3(_02550_),
    .S1(net5453),
    .X(_02551_));
 sg13g2_or2_1 _17116_ (.X(_02552_),
    .B(_02551_),
    .A(net5442));
 sg13g2_o21ai_1 _17117_ (.B1(_02552_),
    .Y(_02553_),
    .A1(_02541_),
    .A2(_02546_));
 sg13g2_o21ai_1 _17118_ (.B1(_02536_),
    .Y(_00280_),
    .A1(net5148),
    .A2(_02553_));
 sg13g2_nand2_1 _17119_ (.Y(_02554_),
    .A(net5774),
    .B(net5154));
 sg13g2_mux4_1 _17120_ (.S0(net5557),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][22] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][22] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][22] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][22] ),
    .S1(net5512),
    .X(_02555_));
 sg13g2_inv_1 _17121_ (.Y(_02556_),
    .A(_02555_));
 sg13g2_mux4_1 _17122_ (.S0(net5557),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][22] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][22] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][22] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][22] ),
    .S1(net5512),
    .X(_02557_));
 sg13g2_a21oi_1 _17123_ (.A1(net5471),
    .A2(_02556_),
    .Y(_02558_),
    .B1(net5458));
 sg13g2_o21ai_1 _17124_ (.B1(_02558_),
    .Y(_02559_),
    .A1(net5471),
    .A2(_02557_));
 sg13g2_mux4_1 _17125_ (.S0(net5558),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][22] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][22] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][22] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][22] ),
    .S1(net5513),
    .X(_02560_));
 sg13g2_mux4_1 _17126_ (.S0(net5557),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][22] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][22] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][22] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][22] ),
    .S1(net5512),
    .X(_02561_));
 sg13g2_nor2_1 _17127_ (.A(net5369),
    .B(_02561_),
    .Y(_02562_));
 sg13g2_o21ai_1 _17128_ (.B1(net5458),
    .Y(_02563_),
    .A1(net5471),
    .A2(_02560_));
 sg13g2_o21ai_1 _17129_ (.B1(net5449),
    .Y(_02564_),
    .A1(_02562_),
    .A2(_02563_));
 sg13g2_nand2b_2 _17130_ (.Y(_02565_),
    .B(_02559_),
    .A_N(_02564_));
 sg13g2_mux4_1 _17131_ (.S0(net5545),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][22] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][22] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][22] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][22] ),
    .S1(net5500),
    .X(_02566_));
 sg13g2_mux4_1 _17132_ (.S0(net5545),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][22] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][22] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][22] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][22] ),
    .S1(net5500),
    .X(_02567_));
 sg13g2_mux4_1 _17133_ (.S0(net5545),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][22] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][22] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][22] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][22] ),
    .S1(net5500),
    .X(_02568_));
 sg13g2_mux4_1 _17134_ (.S0(net5545),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][22] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][22] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][22] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][22] ),
    .S1(net5500),
    .X(_02569_));
 sg13g2_mux4_1 _17135_ (.S0(net5368),
    .A0(_02566_),
    .A1(_02567_),
    .A2(_02568_),
    .A3(_02569_),
    .S1(net5457),
    .X(_02570_));
 sg13g2_o21ai_1 _17136_ (.B1(_02565_),
    .Y(_02571_),
    .A1(net5446),
    .A2(_02570_));
 sg13g2_o21ai_1 _17137_ (.B1(_02554_),
    .Y(_00281_),
    .A1(net5148),
    .A2(_02571_));
 sg13g2_nand2_1 _17138_ (.Y(_02572_),
    .A(net5771),
    .B(net5153));
 sg13g2_mux4_1 _17139_ (.S0(net5563),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][23] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][23] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][23] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][23] ),
    .S1(net5518),
    .X(_02573_));
 sg13g2_inv_1 _17140_ (.Y(_02574_),
    .A(_02573_));
 sg13g2_mux4_1 _17141_ (.S0(net5552),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][23] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][23] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][23] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][23] ),
    .S1(net5507),
    .X(_02575_));
 sg13g2_a21oi_1 _17142_ (.A1(net5473),
    .A2(_02574_),
    .Y(_02576_),
    .B1(net5460));
 sg13g2_o21ai_1 _17143_ (.B1(_02576_),
    .Y(_02577_),
    .A1(net5472),
    .A2(_02575_));
 sg13g2_mux4_1 _17144_ (.S0(net5552),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][23] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][23] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][23] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][23] ),
    .S1(net5507),
    .X(_02578_));
 sg13g2_mux4_1 _17145_ (.S0(net5563),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][23] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][23] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][23] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][23] ),
    .S1(net5518),
    .X(_02579_));
 sg13g2_nor2_1 _17146_ (.A(net5370),
    .B(_02579_),
    .Y(_02580_));
 sg13g2_o21ai_1 _17147_ (.B1(net5462),
    .Y(_02581_),
    .A1(net5473),
    .A2(_02578_));
 sg13g2_o21ai_1 _17148_ (.B1(net5448),
    .Y(_02582_),
    .A1(_02580_),
    .A2(_02581_));
 sg13g2_nand2b_2 _17149_ (.Y(_02583_),
    .B(_02577_),
    .A_N(_02582_));
 sg13g2_mux4_1 _17150_ (.S0(net5551),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][23] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][23] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][23] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][23] ),
    .S1(net5506),
    .X(_02584_));
 sg13g2_mux4_1 _17151_ (.S0(net5551),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][23] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][23] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][23] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][23] ),
    .S1(net5506),
    .X(_02585_));
 sg13g2_mux4_1 _17152_ (.S0(net5551),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][23] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][23] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][23] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][23] ),
    .S1(net5506),
    .X(_02586_));
 sg13g2_mux4_1 _17153_ (.S0(net5551),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][23] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][23] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][23] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][23] ),
    .S1(net5506),
    .X(_02587_));
 sg13g2_mux4_1 _17154_ (.S0(net5469),
    .A0(_02584_),
    .A1(_02585_),
    .A2(_02587_),
    .A3(_02586_),
    .S1(net5361),
    .X(_02588_));
 sg13g2_o21ai_1 _17155_ (.B1(_02583_),
    .Y(_02589_),
    .A1(net5447),
    .A2(_02588_));
 sg13g2_o21ai_1 _17156_ (.B1(_02572_),
    .Y(_00282_),
    .A1(net5149),
    .A2(_02589_));
 sg13g2_nand2_1 _17157_ (.Y(_02590_),
    .A(net5769),
    .B(net5153));
 sg13g2_mux4_1 _17158_ (.S0(net5563),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][24] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][24] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][24] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][24] ),
    .S1(net5518),
    .X(_02591_));
 sg13g2_inv_1 _17159_ (.Y(_02592_),
    .A(_02591_));
 sg13g2_mux4_1 _17160_ (.S0(net5563),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][24] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][24] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][24] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][24] ),
    .S1(net5518),
    .X(_02593_));
 sg13g2_a21oi_1 _17161_ (.A1(net5473),
    .A2(_02592_),
    .Y(_02594_),
    .B1(net5460));
 sg13g2_o21ai_1 _17162_ (.B1(_02594_),
    .Y(_02595_),
    .A1(net5472),
    .A2(_02593_));
 sg13g2_mux4_1 _17163_ (.S0(net5563),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][24] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][24] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][24] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][24] ),
    .S1(net5518),
    .X(_02596_));
 sg13g2_mux4_1 _17164_ (.S0(net5563),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][24] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][24] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][24] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][24] ),
    .S1(net5518),
    .X(_02597_));
 sg13g2_nor2_1 _17165_ (.A(net5370),
    .B(_02597_),
    .Y(_02598_));
 sg13g2_o21ai_1 _17166_ (.B1(net5460),
    .Y(_02599_),
    .A1(net5473),
    .A2(_02596_));
 sg13g2_o21ai_1 _17167_ (.B1(net5448),
    .Y(_02600_),
    .A1(_02598_),
    .A2(_02599_));
 sg13g2_nand2b_2 _17168_ (.Y(_02601_),
    .B(_02595_),
    .A_N(_02600_));
 sg13g2_mux4_1 _17169_ (.S0(net5543),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][24] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][24] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][24] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][24] ),
    .S1(net5498),
    .X(_02602_));
 sg13g2_mux4_1 _17170_ (.S0(net5542),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][24] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][24] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][24] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][24] ),
    .S1(net5497),
    .X(_02603_));
 sg13g2_mux4_1 _17171_ (.S0(net5542),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][24] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][24] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][24] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][24] ),
    .S1(net5497),
    .X(_02604_));
 sg13g2_mux4_1 _17172_ (.S0(net5551),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][24] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][24] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][24] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][24] ),
    .S1(net5506),
    .X(_02605_));
 sg13g2_mux4_1 _17173_ (.S0(net5366),
    .A0(_02602_),
    .A1(_02603_),
    .A2(_02604_),
    .A3(_02605_),
    .S1(net5454),
    .X(_02606_));
 sg13g2_o21ai_1 _17174_ (.B1(_02601_),
    .Y(_02607_),
    .A1(net5447),
    .A2(_02606_));
 sg13g2_o21ai_1 _17175_ (.B1(_02590_),
    .Y(_00283_),
    .A1(net5149),
    .A2(_02607_));
 sg13g2_nand2_1 _17176_ (.Y(_02608_),
    .A(net5768),
    .B(net5152));
 sg13g2_mux4_1 _17177_ (.S0(net5557),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][25] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][25] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][25] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][25] ),
    .S1(net5512),
    .X(_02609_));
 sg13g2_mux4_1 _17178_ (.S0(net5557),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][25] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][25] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][25] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][25] ),
    .S1(net5512),
    .X(_02610_));
 sg13g2_mux2_1 _17179_ (.A0(_02609_),
    .A1(_02610_),
    .S(net5369),
    .X(_02611_));
 sg13g2_mux4_1 _17180_ (.S0(net5557),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][25] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][25] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][25] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][25] ),
    .S1(net5512),
    .X(_02612_));
 sg13g2_nor2_1 _17181_ (.A(net5471),
    .B(_02612_),
    .Y(_02613_));
 sg13g2_mux4_1 _17182_ (.S0(net5557),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][25] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][25] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][25] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][25] ),
    .S1(net5512),
    .X(_02614_));
 sg13g2_o21ai_1 _17183_ (.B1(net5458),
    .Y(_02615_),
    .A1(net5371),
    .A2(_02614_));
 sg13g2_o21ai_1 _17184_ (.B1(net5449),
    .Y(_02616_),
    .A1(_02613_),
    .A2(_02615_));
 sg13g2_a21o_1 _17185_ (.A2(_02611_),
    .A1(net5360),
    .B1(_02616_),
    .X(_02617_));
 sg13g2_mux4_1 _17186_ (.S0(net5547),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][25] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][25] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][25] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][25] ),
    .S1(net5502),
    .X(_02618_));
 sg13g2_mux4_1 _17187_ (.S0(net5547),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][25] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][25] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][25] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][25] ),
    .S1(net5502),
    .X(_02619_));
 sg13g2_mux4_1 _17188_ (.S0(net5547),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][25] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][25] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][25] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][25] ),
    .S1(net5502),
    .X(_02620_));
 sg13g2_mux4_1 _17189_ (.S0(net5549),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][25] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][25] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][25] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][25] ),
    .S1(net5504),
    .X(_02621_));
 sg13g2_mux4_1 _17190_ (.S0(net5469),
    .A0(_02618_),
    .A1(_02619_),
    .A2(_02621_),
    .A3(_02620_),
    .S1(net5360),
    .X(_02622_));
 sg13g2_o21ai_1 _17191_ (.B1(_02617_),
    .Y(_02623_),
    .A1(net5446),
    .A2(_02622_));
 sg13g2_o21ai_1 _17192_ (.B1(_02608_),
    .Y(_00284_),
    .A1(net5148),
    .A2(_02623_));
 sg13g2_nand2_1 _17193_ (.Y(_02624_),
    .A(net5765),
    .B(net5153));
 sg13g2_mux4_1 _17194_ (.S0(net5539),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][26] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][26] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][26] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][26] ),
    .S1(net5494),
    .X(_02625_));
 sg13g2_inv_1 _17195_ (.Y(_02626_),
    .A(_02625_));
 sg13g2_mux4_1 _17196_ (.S0(net5541),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][26] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][26] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][26] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][26] ),
    .S1(net5496),
    .X(_02627_));
 sg13g2_a21oi_1 _17197_ (.A1(net5466),
    .A2(_02626_),
    .Y(_02628_),
    .B1(net5455));
 sg13g2_o21ai_1 _17198_ (.B1(_02628_),
    .Y(_02629_),
    .A1(net5467),
    .A2(_02627_));
 sg13g2_mux4_1 _17199_ (.S0(net5539),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][26] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][26] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][26] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][26] ),
    .S1(net5494),
    .X(_02630_));
 sg13g2_nor2_1 _17200_ (.A(net5466),
    .B(_02630_),
    .Y(_02631_));
 sg13g2_mux4_1 _17201_ (.S0(net5539),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][26] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][26] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][26] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][26] ),
    .S1(net5494),
    .X(_02632_));
 sg13g2_o21ai_1 _17202_ (.B1(net5455),
    .Y(_02633_),
    .A1(net5366),
    .A2(_02632_));
 sg13g2_o21ai_1 _17203_ (.B1(net5443),
    .Y(_02634_),
    .A1(_02631_),
    .A2(_02633_));
 sg13g2_nand2b_2 _17204_ (.Y(_02635_),
    .B(_02629_),
    .A_N(_02634_));
 sg13g2_mux4_1 _17205_ (.S0(net5528),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][26] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][26] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][26] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][26] ),
    .S1(net5483),
    .X(_02636_));
 sg13g2_mux4_1 _17206_ (.S0(net5528),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][26] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][26] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][26] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][26] ),
    .S1(net5483),
    .X(_02637_));
 sg13g2_mux4_1 _17207_ (.S0(net5528),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][26] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][26] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][26] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][26] ),
    .S1(net5483),
    .X(_02638_));
 sg13g2_mux4_1 _17208_ (.S0(net5532),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][26] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][26] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][26] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][26] ),
    .S1(net5487),
    .X(_02639_));
 sg13g2_mux4_1 _17209_ (.S0(net5463),
    .A0(_02636_),
    .A1(_02637_),
    .A2(_02639_),
    .A3(_02638_),
    .S1(net5358),
    .X(_02640_));
 sg13g2_o21ai_1 _17210_ (.B1(_02635_),
    .Y(_02641_),
    .A1(net5441),
    .A2(_02640_));
 sg13g2_o21ai_1 _17211_ (.B1(_02624_),
    .Y(_00285_),
    .A1(net5149),
    .A2(_02641_));
 sg13g2_nand2_1 _17212_ (.Y(_02642_),
    .A(net5763),
    .B(net5152));
 sg13g2_mux4_1 _17213_ (.S0(net5542),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][27] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][27] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][27] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][27] ),
    .S1(net5497),
    .X(_02643_));
 sg13g2_mux4_1 _17214_ (.S0(net5540),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][27] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][27] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][27] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][27] ),
    .S1(net5495),
    .X(_02644_));
 sg13g2_nor2_1 _17215_ (.A(net5467),
    .B(_02644_),
    .Y(_02645_));
 sg13g2_o21ai_1 _17216_ (.B1(net5455),
    .Y(_02646_),
    .A1(net5367),
    .A2(_02643_));
 sg13g2_mux4_1 _17217_ (.S0(net5535),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][27] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][27] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][27] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][27] ),
    .S1(net5490),
    .X(_02647_));
 sg13g2_nor2_1 _17218_ (.A(net5365),
    .B(_02647_),
    .Y(_02648_));
 sg13g2_mux4_1 _17219_ (.S0(net5537),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][27] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][27] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][27] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][27] ),
    .S1(net5492),
    .X(_02649_));
 sg13g2_o21ai_1 _17220_ (.B1(net5359),
    .Y(_02650_),
    .A1(net5465),
    .A2(_02649_));
 sg13g2_nor2_1 _17221_ (.A(_02648_),
    .B(_02650_),
    .Y(_02651_));
 sg13g2_o21ai_1 _17222_ (.B1(net5444),
    .Y(_02652_),
    .A1(_02645_),
    .A2(_02646_));
 sg13g2_mux4_1 _17223_ (.S0(net5531),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][27] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][27] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][27] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][27] ),
    .S1(net5486),
    .X(_02653_));
 sg13g2_mux4_1 _17224_ (.S0(net5531),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][27] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][27] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][27] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][27] ),
    .S1(net5486),
    .X(_02654_));
 sg13g2_mux4_1 _17225_ (.S0(net5531),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][27] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][27] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][27] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][27] ),
    .S1(net5486),
    .X(_02655_));
 sg13g2_mux4_1 _17226_ (.S0(net5531),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][27] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][27] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][27] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][27] ),
    .S1(net5486),
    .X(_02656_));
 sg13g2_mux4_1 _17227_ (.S0(net5364),
    .A0(_02653_),
    .A1(_02654_),
    .A2(_02655_),
    .A3(_02656_),
    .S1(net5456),
    .X(_02657_));
 sg13g2_or2_1 _17228_ (.X(_02658_),
    .B(_02657_),
    .A(net5445));
 sg13g2_o21ai_1 _17229_ (.B1(_02658_),
    .Y(_02659_),
    .A1(_02651_),
    .A2(_02652_));
 sg13g2_o21ai_1 _17230_ (.B1(_02642_),
    .Y(_00286_),
    .A1(net5148),
    .A2(_02659_));
 sg13g2_nand2_1 _17231_ (.Y(_02660_),
    .A(net5760),
    .B(net5152));
 sg13g2_mux4_1 _17232_ (.S0(net5540),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][28] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][28] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][28] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][28] ),
    .S1(net5495),
    .X(_02661_));
 sg13g2_inv_1 _17233_ (.Y(_02662_),
    .A(_02661_));
 sg13g2_mux4_1 _17234_ (.S0(net5535),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][28] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][28] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][28] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][28] ),
    .S1(net5490),
    .X(_02663_));
 sg13g2_a21oi_1 _17235_ (.A1(net5465),
    .A2(_02662_),
    .Y(_02664_),
    .B1(net5455));
 sg13g2_o21ai_1 _17236_ (.B1(_02664_),
    .Y(_02665_),
    .A1(net5466),
    .A2(_02663_));
 sg13g2_mux4_1 _17237_ (.S0(net5535),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][28] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][28] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][28] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][28] ),
    .S1(net5490),
    .X(_02666_));
 sg13g2_mux4_1 _17238_ (.S0(net5540),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][28] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][28] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][28] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][28] ),
    .S1(net5495),
    .X(_02667_));
 sg13g2_nor2_1 _17239_ (.A(net5366),
    .B(_02667_),
    .Y(_02668_));
 sg13g2_o21ai_1 _17240_ (.B1(net5454),
    .Y(_02669_),
    .A1(net5465),
    .A2(_02666_));
 sg13g2_o21ai_1 _17241_ (.B1(net5443),
    .Y(_02670_),
    .A1(_02668_),
    .A2(_02669_));
 sg13g2_nand2b_1 _17242_ (.Y(_02671_),
    .B(_02665_),
    .A_N(_02670_));
 sg13g2_mux4_1 _17243_ (.S0(net5540),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][28] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][28] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][28] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][28] ),
    .S1(net5495),
    .X(_02672_));
 sg13g2_mux4_1 _17244_ (.S0(net5540),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][28] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][28] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][28] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][28] ),
    .S1(net5495),
    .X(_02673_));
 sg13g2_mux4_1 _17245_ (.S0(net5540),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][28] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][28] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][28] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][28] ),
    .S1(net5495),
    .X(_02674_));
 sg13g2_mux4_1 _17246_ (.S0(net5540),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][28] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][28] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][28] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][28] ),
    .S1(net5495),
    .X(_02675_));
 sg13g2_mux4_1 _17247_ (.S0(net5367),
    .A0(_02672_),
    .A1(_02673_),
    .A2(_02674_),
    .A3(_02675_),
    .S1(net5455),
    .X(_02676_));
 sg13g2_o21ai_1 _17248_ (.B1(_02671_),
    .Y(_02677_),
    .A1(net5444),
    .A2(_02676_));
 sg13g2_o21ai_1 _17249_ (.B1(_02660_),
    .Y(_00287_),
    .A1(net5148),
    .A2(_02677_));
 sg13g2_nand2_1 _17250_ (.Y(_02678_),
    .A(net5759),
    .B(net5155));
 sg13g2_mux4_1 _17251_ (.S0(net5562),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][29] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][29] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][29] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][29] ),
    .S1(net5517),
    .X(_02679_));
 sg13g2_mux4_1 _17252_ (.S0(net5563),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][29] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][29] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][29] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][29] ),
    .S1(net5518),
    .X(_02680_));
 sg13g2_nor2_1 _17253_ (.A(net5474),
    .B(_02680_),
    .Y(_02681_));
 sg13g2_nor2_1 _17254_ (.A(net5361),
    .B(_02681_),
    .Y(_02682_));
 sg13g2_o21ai_1 _17255_ (.B1(_02682_),
    .Y(_02683_),
    .A1(net5370),
    .A2(_02679_));
 sg13g2_mux4_1 _17256_ (.S0(net5564),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][29] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][29] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][29] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][29] ),
    .S1(net5519),
    .X(_02684_));
 sg13g2_inv_1 _17257_ (.Y(_02685_),
    .A(_02684_));
 sg13g2_mux4_1 _17258_ (.S0(net5563),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][29] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][29] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][29] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][29] ),
    .S1(net5518),
    .X(_02686_));
 sg13g2_a21oi_1 _17259_ (.A1(net5474),
    .A2(_02685_),
    .Y(_02687_),
    .B1(net5460));
 sg13g2_o21ai_1 _17260_ (.B1(_02687_),
    .Y(_02688_),
    .A1(net5474),
    .A2(_02686_));
 sg13g2_nand3_1 _17261_ (.B(_02683_),
    .C(_02688_),
    .A(net5450),
    .Y(_02689_));
 sg13g2_mux4_1 _17262_ (.S0(net5552),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][29] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][29] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][29] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][29] ),
    .S1(net5507),
    .X(_02690_));
 sg13g2_mux4_1 _17263_ (.S0(net5554),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][29] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][29] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][29] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][29] ),
    .S1(net5509),
    .X(_02691_));
 sg13g2_mux4_1 _17264_ (.S0(net5554),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][29] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][29] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][29] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][29] ),
    .S1(net5509),
    .X(_02692_));
 sg13g2_mux4_1 _17265_ (.S0(net5552),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][29] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][29] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][29] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][29] ),
    .S1(net5507),
    .X(_02693_));
 sg13g2_mux4_1 _17266_ (.S0(net5372),
    .A0(_02690_),
    .A1(_02691_),
    .A2(_02692_),
    .A3(_02693_),
    .S1(net5462),
    .X(_02694_));
 sg13g2_o21ai_1 _17267_ (.B1(_02689_),
    .Y(_02695_),
    .A1(net5447),
    .A2(_02694_));
 sg13g2_o21ai_1 _17268_ (.B1(_02678_),
    .Y(_00288_),
    .A1(net5149),
    .A2(_02695_));
 sg13g2_nand2_1 _17269_ (.Y(_02696_),
    .A(net5756),
    .B(net5152));
 sg13g2_mux4_1 _17270_ (.S0(net5561),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][30] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][30] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][30] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][30] ),
    .S1(net5516),
    .X(_02697_));
 sg13g2_inv_1 _17271_ (.Y(_02698_),
    .A(_02697_));
 sg13g2_mux4_1 _17272_ (.S0(net5559),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][30] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][30] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][30] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][30] ),
    .S1(net5514),
    .X(_02699_));
 sg13g2_a21oi_1 _17273_ (.A1(net5477),
    .A2(_02698_),
    .Y(_02700_),
    .B1(net5458));
 sg13g2_o21ai_1 _17274_ (.B1(_02700_),
    .Y(_02701_),
    .A1(net5477),
    .A2(_02699_));
 sg13g2_mux4_1 _17275_ (.S0(net5561),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][30] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][30] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][30] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][30] ),
    .S1(net5516),
    .X(_02702_));
 sg13g2_mux4_1 _17276_ (.S0(net5561),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][30] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][30] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][30] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][30] ),
    .S1(net5516),
    .X(_02703_));
 sg13g2_nor2_1 _17277_ (.A(net5369),
    .B(_02703_),
    .Y(_02704_));
 sg13g2_o21ai_1 _17278_ (.B1(net5458),
    .Y(_02705_),
    .A1(net5471),
    .A2(_02702_));
 sg13g2_o21ai_1 _17279_ (.B1(net5449),
    .Y(_02706_),
    .A1(_02704_),
    .A2(_02705_));
 sg13g2_nand2b_2 _17280_ (.Y(_02707_),
    .B(_02701_),
    .A_N(_02706_));
 sg13g2_mux4_1 _17281_ (.S0(net5548),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][30] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][30] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][30] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][30] ),
    .S1(net5503),
    .X(_02708_));
 sg13g2_mux4_1 _17282_ (.S0(net5548),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][30] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][30] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][30] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][30] ),
    .S1(net5503),
    .X(_02709_));
 sg13g2_mux4_1 _17283_ (.S0(net5549),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][30] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][30] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][30] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][30] ),
    .S1(net5504),
    .X(_02710_));
 sg13g2_mux4_1 _17284_ (.S0(net5548),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][30] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][30] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][30] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][30] ),
    .S1(net5503),
    .X(_02711_));
 sg13g2_mux4_1 _17285_ (.S0(net5368),
    .A0(_02708_),
    .A1(_02709_),
    .A2(_02710_),
    .A3(_02711_),
    .S1(net5457),
    .X(_02712_));
 sg13g2_o21ai_1 _17286_ (.B1(_02707_),
    .Y(_02713_),
    .A1(net5446),
    .A2(_02712_));
 sg13g2_o21ai_1 _17287_ (.B1(_02696_),
    .Y(_00289_),
    .A1(net5148),
    .A2(_02713_));
 sg13g2_nand2_1 _17288_ (.Y(_02714_),
    .A(net5755),
    .B(net5154));
 sg13g2_mux4_1 _17289_ (.S0(net5559),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][31] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][31] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][31] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][31] ),
    .S1(net5514),
    .X(_02715_));
 sg13g2_inv_1 _17290_ (.Y(_02716_),
    .A(_02715_));
 sg13g2_mux4_1 _17291_ (.S0(net5562),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][31] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][31] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][31] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][31] ),
    .S1(net5517),
    .X(_02717_));
 sg13g2_a21oi_1 _17292_ (.A1(net5475),
    .A2(_02716_),
    .Y(_02718_),
    .B1(net5459));
 sg13g2_o21ai_1 _17293_ (.B1(_02718_),
    .Y(_02719_),
    .A1(net5472),
    .A2(_02717_));
 sg13g2_mux4_1 _17294_ (.S0(net5565),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][31] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][31] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][31] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][31] ),
    .S1(net5520),
    .X(_02720_));
 sg13g2_nor2_1 _17295_ (.A(net5475),
    .B(_02720_),
    .Y(_02721_));
 sg13g2_mux4_1 _17296_ (.S0(net5565),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][31] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][31] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][31] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][31] ),
    .S1(net5520),
    .X(_02722_));
 sg13g2_o21ai_1 _17297_ (.B1(net5459),
    .Y(_02723_),
    .A1(net5371),
    .A2(_02722_));
 sg13g2_o21ai_1 _17298_ (.B1(net5450),
    .Y(_02724_),
    .A1(_02721_),
    .A2(_02723_));
 sg13g2_nand2b_2 _17299_ (.Y(_02725_),
    .B(_02719_),
    .A_N(_02724_));
 sg13g2_mux4_1 _17300_ (.S0(net5550),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][31] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][31] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][31] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][31] ),
    .S1(net5505),
    .X(_02726_));
 sg13g2_mux4_1 _17301_ (.S0(net5542),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][31] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][31] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][31] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][31] ),
    .S1(net5497),
    .X(_02727_));
 sg13g2_mux4_1 _17302_ (.S0(net5550),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][31] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][31] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][31] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][31] ),
    .S1(net5505),
    .X(_02728_));
 sg13g2_mux4_1 _17303_ (.S0(net5550),
    .A0(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][31] ),
    .A1(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][31] ),
    .A2(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][31] ),
    .A3(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][31] ),
    .S1(net5505),
    .X(_02729_));
 sg13g2_mux4_1 _17304_ (.S0(net5478),
    .A0(_02726_),
    .A1(_02727_),
    .A2(_02729_),
    .A3(_02728_),
    .S1(net5361),
    .X(_02730_));
 sg13g2_o21ai_1 _17305_ (.B1(_02725_),
    .Y(_02731_),
    .A1(net5447),
    .A2(_02730_));
 sg13g2_o21ai_1 _17306_ (.B1(_02714_),
    .Y(_00290_),
    .A1(net5147),
    .A2(_02731_));
 sg13g2_nand4_1 _17307_ (.B(net1781),
    .C(_06682_),
    .A(\fpga_top.cpu_top.csr_meie ),
    .Y(_02732_),
    .D(net1373));
 sg13g2_nand2b_2 _17308_ (.Y(_02733_),
    .B(_08895_),
    .A_N(_08897_));
 sg13g2_nor2_1 _17309_ (.A(_08982_),
    .B(_02733_),
    .Y(_02734_));
 sg13g2_nand2_1 _17310_ (.Y(_02735_),
    .A(_08978_),
    .B(_02734_));
 sg13g2_nor2_1 _17311_ (.A(net4560),
    .B(_02735_),
    .Y(_02736_));
 sg13g2_a22oi_1 _17312_ (.Y(_00291_),
    .B1(_02736_),
    .B2(net4917),
    .A2(net3969),
    .A1(_06776_));
 sg13g2_nand2_1 _17313_ (.Y(_02737_),
    .A(net5426),
    .B(net5666));
 sg13g2_inv_2 _17314_ (.Y(_02738_),
    .A(net5327));
 sg13g2_nand3_1 _17315_ (.B(net1834),
    .C(_02738_),
    .A(\fpga_top.cpu_top.csr_meie ),
    .Y(_02739_));
 sg13g2_a22oi_1 _17316_ (.Y(_00292_),
    .B1(_02739_),
    .B2(_06777_),
    .A2(_02736_),
    .A1(net4919));
 sg13g2_nand2_2 _17317_ (.Y(_02740_),
    .A(_08909_),
    .B(_08984_));
 sg13g2_nor2_2 _17318_ (.A(net4560),
    .B(_02740_),
    .Y(_02741_));
 sg13g2_nor2_1 _17319_ (.A(net2189),
    .B(net4517),
    .Y(_02742_));
 sg13g2_a21oi_1 _17320_ (.A1(net4919),
    .A2(net4517),
    .Y(_00293_),
    .B1(_02742_));
 sg13g2_nor2_1 _17321_ (.A(net3768),
    .B(net4518),
    .Y(_02743_));
 sg13g2_a21oi_1 _17322_ (.A1(net4917),
    .A2(net4518),
    .Y(_00294_),
    .B1(_02743_));
 sg13g2_nor2_1 _17323_ (.A(net3421),
    .B(net4518),
    .Y(_02744_));
 sg13g2_a21oi_1 _17324_ (.A1(net4852),
    .A2(net4518),
    .Y(_00295_),
    .B1(_02744_));
 sg13g2_nand2_1 _17325_ (.Y(_02745_),
    .A(net4844),
    .B(net4519));
 sg13g2_o21ai_1 _17326_ (.B1(_02745_),
    .Y(_00296_),
    .A1(_06763_),
    .A2(net4519));
 sg13g2_nand2_1 _17327_ (.Y(_02746_),
    .A(net5660),
    .B(net5088));
 sg13g2_o21ai_1 _17328_ (.B1(_02746_),
    .Y(_02747_),
    .A1(_06577_),
    .A2(net5088));
 sg13g2_nand2_1 _17329_ (.Y(_02748_),
    .A(net4518),
    .B(net4839));
 sg13g2_o21ai_1 _17330_ (.B1(_02748_),
    .Y(_00297_),
    .A1(_06762_),
    .A2(net4518));
 sg13g2_nor2_1 _17331_ (.A(net3826),
    .B(net4517),
    .Y(_02749_));
 sg13g2_nor2_1 _17332_ (.A(_06586_),
    .B(net5077),
    .Y(_02750_));
 sg13g2_a21oi_2 _17333_ (.B1(_02750_),
    .Y(_02751_),
    .A2(net5077),
    .A1(net5658));
 sg13g2_a21o_2 _17334_ (.A2(net5077),
    .A1(net5658),
    .B1(_02750_),
    .X(_02752_));
 sg13g2_a21oi_1 _17335_ (.A1(net4517),
    .A2(net4836),
    .Y(_00298_),
    .B1(_02749_));
 sg13g2_nor2_1 _17336_ (.A(net3755),
    .B(net4517),
    .Y(_02753_));
 sg13g2_nor2b_1 _17337_ (.A(net5077),
    .B_N(\fpga_top.bus_gather.d_write_data[6] ),
    .Y(_02754_));
 sg13g2_a21oi_2 _17338_ (.B1(_02754_),
    .Y(_02755_),
    .A2(net5077),
    .A1(\fpga_top.cpu_start_adr[6] ));
 sg13g2_a21o_2 _17339_ (.A2(net5079),
    .A1(\fpga_top.cpu_start_adr[6] ),
    .B1(_02754_),
    .X(_02756_));
 sg13g2_a21oi_1 _17340_ (.A1(net4517),
    .A2(net4833),
    .Y(_00299_),
    .B1(_02753_));
 sg13g2_nor2_1 _17341_ (.A(net3717),
    .B(net4517),
    .Y(_02757_));
 sg13g2_nor2b_1 _17342_ (.A(net5077),
    .B_N(\fpga_top.bus_gather.d_write_data[7] ),
    .Y(_02758_));
 sg13g2_a21oi_2 _17343_ (.B1(_02758_),
    .Y(_02759_),
    .A2(net5077),
    .A1(net5656));
 sg13g2_a21o_2 _17344_ (.A2(net5079),
    .A1(net5656),
    .B1(_02758_),
    .X(_02760_));
 sg13g2_a21oi_1 _17345_ (.A1(net4517),
    .A2(net4831),
    .Y(_00300_),
    .B1(_02757_));
 sg13g2_nor2_1 _17346_ (.A(net3667),
    .B(net4523),
    .Y(_02761_));
 sg13g2_nor2b_2 _17347_ (.A(net5078),
    .B_N(\fpga_top.bus_gather.d_write_data[8] ),
    .Y(_02762_));
 sg13g2_a21oi_2 _17348_ (.B1(_02762_),
    .Y(_02763_),
    .A2(net5080),
    .A1(net5654));
 sg13g2_a21o_2 _17349_ (.A2(net5080),
    .A1(net5654),
    .B1(_02762_),
    .X(_02764_));
 sg13g2_a21oi_1 _17350_ (.A1(net4523),
    .A2(_02763_),
    .Y(_00301_),
    .B1(_02761_));
 sg13g2_nor2_1 _17351_ (.A(net3699),
    .B(net4523),
    .Y(_02765_));
 sg13g2_nor2b_2 _17352_ (.A(net5079),
    .B_N(\fpga_top.bus_gather.d_write_data[9] ),
    .Y(_02766_));
 sg13g2_a21oi_2 _17353_ (.B1(_02766_),
    .Y(_02767_),
    .A2(net5080),
    .A1(net5653));
 sg13g2_a21o_2 _17354_ (.A2(net5077),
    .A1(net5653),
    .B1(_02766_),
    .X(_02768_));
 sg13g2_a21oi_1 _17355_ (.A1(net4523),
    .A2(_02767_),
    .Y(_00302_),
    .B1(_02765_));
 sg13g2_mux2_1 _17356_ (.A0(net6101),
    .A1(_08981_),
    .S(net4519),
    .X(_00303_));
 sg13g2_nor2_1 _17357_ (.A(net2957),
    .B(net4519),
    .Y(_02769_));
 sg13g2_nand2_1 _17358_ (.Y(_02770_),
    .A(_06793_),
    .B(net5084));
 sg13g2_o21ai_1 _17359_ (.B1(_02770_),
    .Y(_02771_),
    .A1(\fpga_top.bus_gather.d_write_data[11] ),
    .A2(net5082));
 sg13g2_a21oi_1 _17360_ (.A1(net4519),
    .A2(_02771_),
    .Y(_00304_),
    .B1(_02769_));
 sg13g2_nor2_1 _17361_ (.A(net2856),
    .B(net4526),
    .Y(_02772_));
 sg13g2_nor2_1 _17362_ (.A(\fpga_top.bus_gather.d_write_data[12] ),
    .B(net5086),
    .Y(_02773_));
 sg13g2_a21oi_2 _17363_ (.B1(_02773_),
    .Y(_02774_),
    .A2(net5081),
    .A1(net5375));
 sg13g2_a21o_2 _17364_ (.A2(net5085),
    .A1(net5375),
    .B1(_02773_),
    .X(_02775_));
 sg13g2_a21oi_1 _17365_ (.A1(net4526),
    .A2(_02775_),
    .Y(_00305_),
    .B1(_02772_));
 sg13g2_nor2_1 _17366_ (.A(net3704),
    .B(net4526),
    .Y(_02776_));
 sg13g2_nand2_1 _17367_ (.Y(_02777_),
    .A(net5374),
    .B(net5085));
 sg13g2_o21ai_1 _17368_ (.B1(_02777_),
    .Y(_02778_),
    .A1(\fpga_top.bus_gather.d_write_data[13] ),
    .A2(net5087));
 sg13g2_a21oi_1 _17369_ (.A1(net4526),
    .A2(_02778_),
    .Y(_00306_),
    .B1(_02776_));
 sg13g2_nor2_1 _17370_ (.A(net3658),
    .B(net4526),
    .Y(_02779_));
 sg13g2_nand2_1 _17371_ (.Y(_02780_),
    .A(_06796_),
    .B(net5084));
 sg13g2_o21ai_1 _17372_ (.B1(_02780_),
    .Y(_02781_),
    .A1(\fpga_top.bus_gather.d_write_data[14] ),
    .A2(net5084));
 sg13g2_inv_1 _17373_ (.Y(_02782_),
    .A(_02781_));
 sg13g2_a21oi_1 _17374_ (.A1(net4527),
    .A2(_02781_),
    .Y(_00307_),
    .B1(_02779_));
 sg13g2_nor2_1 _17375_ (.A(net3234),
    .B(net4527),
    .Y(_02783_));
 sg13g2_mux2_1 _17376_ (.A0(_06604_),
    .A1(net5373),
    .S(net5089),
    .X(_02784_));
 sg13g2_a21oi_1 _17377_ (.A1(net4527),
    .A2(_02784_),
    .Y(_00308_),
    .B1(_02783_));
 sg13g2_nor2_1 _17378_ (.A(net3580),
    .B(net4521),
    .Y(_02785_));
 sg13g2_a21oi_1 _17379_ (.A1(_10595_),
    .A2(net4520),
    .Y(_00309_),
    .B1(_02785_));
 sg13g2_nor2_1 _17380_ (.A(net3297),
    .B(net4521),
    .Y(_02786_));
 sg13g2_a21oi_1 _17381_ (.A1(_10600_),
    .A2(net4521),
    .Y(_00310_),
    .B1(_02786_));
 sg13g2_nor2_1 _17382_ (.A(net3808),
    .B(net4520),
    .Y(_02787_));
 sg13g2_a21oi_1 _17383_ (.A1(_10603_),
    .A2(net4520),
    .Y(_00311_),
    .B1(_02787_));
 sg13g2_nor2_1 _17384_ (.A(net3685),
    .B(net4520),
    .Y(_02788_));
 sg13g2_mux2_1 _17385_ (.A0(_06616_),
    .A1(_06801_),
    .S(net5084),
    .X(_02789_));
 sg13g2_a21oi_1 _17386_ (.A1(net4520),
    .A2(_02789_),
    .Y(_00312_),
    .B1(_02788_));
 sg13g2_nor2_1 _17387_ (.A(net2869),
    .B(net4520),
    .Y(_02790_));
 sg13g2_a21oi_1 _17388_ (.A1(_10605_),
    .A2(net4521),
    .Y(_00313_),
    .B1(_02790_));
 sg13g2_nor2_1 _17389_ (.A(net3390),
    .B(net4520),
    .Y(_02791_));
 sg13g2_a21oi_1 _17390_ (.A1(_10609_),
    .A2(net4520),
    .Y(_00314_),
    .B1(_02791_));
 sg13g2_nor2_1 _17391_ (.A(net3711),
    .B(net4522),
    .Y(_02792_));
 sg13g2_a21oi_1 _17392_ (.A1(_10611_),
    .A2(net4522),
    .Y(_00315_),
    .B1(_02792_));
 sg13g2_nor2_1 _17393_ (.A(net3528),
    .B(net4522),
    .Y(_02793_));
 sg13g2_nand2_1 _17394_ (.Y(_02794_),
    .A(_06804_),
    .B(net5089));
 sg13g2_o21ai_1 _17395_ (.B1(_02794_),
    .Y(_02795_),
    .A1(\fpga_top.bus_gather.d_write_data[23] ),
    .A2(net5089));
 sg13g2_a21oi_1 _17396_ (.A1(net4522),
    .A2(_02795_),
    .Y(_00316_),
    .B1(_02793_));
 sg13g2_nor2_1 _17397_ (.A(net3686),
    .B(net4524),
    .Y(_02796_));
 sg13g2_a21oi_1 _17398_ (.A1(_10615_),
    .A2(net4527),
    .Y(_00317_),
    .B1(_02796_));
 sg13g2_nor2_1 _17399_ (.A(net3741),
    .B(net4524),
    .Y(_02797_));
 sg13g2_a21oi_1 _17400_ (.A1(_10618_),
    .A2(net4525),
    .Y(_00318_),
    .B1(_02797_));
 sg13g2_nor2_1 _17401_ (.A(net3861),
    .B(net4524),
    .Y(_02798_));
 sg13g2_a21oi_1 _17402_ (.A1(_10622_),
    .A2(net4524),
    .Y(_00319_),
    .B1(_02798_));
 sg13g2_nor2_1 _17403_ (.A(net3157),
    .B(net4525),
    .Y(_02799_));
 sg13g2_nor2_1 _17404_ (.A(\fpga_top.bus_gather.d_write_data[27] ),
    .B(net5078),
    .Y(_02800_));
 sg13g2_nand2b_1 _17405_ (.Y(_02801_),
    .B(net5078),
    .A_N(net5640));
 sg13g2_nor2b_2 _17406_ (.A(_02800_),
    .B_N(_02801_),
    .Y(_02802_));
 sg13g2_nand2b_1 _17407_ (.Y(_02803_),
    .B(_02801_),
    .A_N(_02800_));
 sg13g2_a21oi_1 _17408_ (.A1(net4525),
    .A2(_02803_),
    .Y(_00320_),
    .B1(_02799_));
 sg13g2_nor2_1 _17409_ (.A(net3419),
    .B(net4525),
    .Y(_02804_));
 sg13g2_mux2_1 _17410_ (.A0(_06639_),
    .A1(_06808_),
    .S(net5085),
    .X(_02805_));
 sg13g2_a21oi_1 _17411_ (.A1(net4525),
    .A2(_02805_),
    .Y(_00321_),
    .B1(_02804_));
 sg13g2_nor2_1 _17412_ (.A(net3669),
    .B(net4524),
    .Y(_02806_));
 sg13g2_nor2_1 _17413_ (.A(\fpga_top.bus_gather.d_write_data[29] ),
    .B(net5078),
    .Y(_02807_));
 sg13g2_a21oi_2 _17414_ (.B1(_02807_),
    .Y(_02808_),
    .A2(net5078),
    .A1(_06809_));
 sg13g2_a21o_1 _17415_ (.A2(net5078),
    .A1(_06809_),
    .B1(_02807_),
    .X(_02809_));
 sg13g2_a21oi_1 _17416_ (.A1(net4524),
    .A2(_02809_),
    .Y(_00322_),
    .B1(_02806_));
 sg13g2_nor2_1 _17417_ (.A(net3587),
    .B(net4525),
    .Y(_02810_));
 sg13g2_nor2_1 _17418_ (.A(\fpga_top.bus_gather.d_write_data[30] ),
    .B(net5085),
    .Y(_02811_));
 sg13g2_nand2_1 _17419_ (.Y(_02812_),
    .A(_06810_),
    .B(net5078));
 sg13g2_nor2b_2 _17420_ (.A(_02811_),
    .B_N(_02812_),
    .Y(_02813_));
 sg13g2_nand2b_1 _17421_ (.Y(_02814_),
    .B(_02812_),
    .A_N(_02811_));
 sg13g2_a21oi_1 _17422_ (.A1(net4525),
    .A2(_02814_),
    .Y(_00323_),
    .B1(_02810_));
 sg13g2_nor2_1 _17423_ (.A(net3436),
    .B(net4524),
    .Y(_02815_));
 sg13g2_nand2_1 _17424_ (.Y(_02816_),
    .A(_06811_),
    .B(net5089));
 sg13g2_o21ai_1 _17425_ (.B1(_02816_),
    .Y(_02817_),
    .A1(\fpga_top.bus_gather.d_write_data[31] ),
    .A2(net5089));
 sg13g2_a21oi_1 _17426_ (.A1(net4524),
    .A2(_02817_),
    .Y(_00324_),
    .B1(_02815_));
 sg13g2_or2_1 _17427_ (.X(_02818_),
    .B(_10519_),
    .A(net4560));
 sg13g2_nand2_1 _17428_ (.Y(_02819_),
    .A(net1834),
    .B(_02818_));
 sg13g2_o21ai_1 _17429_ (.B1(_02819_),
    .Y(_00325_),
    .A1(net4919),
    .A2(_02818_));
 sg13g2_nand2_1 _17430_ (.Y(_02820_),
    .A(net1781),
    .B(_02818_));
 sg13g2_o21ai_1 _17431_ (.B1(_02820_),
    .Y(_00326_),
    .A1(net4917),
    .A2(_02818_));
 sg13g2_nor2_1 _17432_ (.A(net6203),
    .B(_08912_),
    .Y(_02821_));
 sg13g2_a21oi_1 _17433_ (.A1(_08912_),
    .A2(net4919),
    .Y(_00327_),
    .B1(_02821_));
 sg13g2_a22oi_1 _17434_ (.Y(_02822_),
    .B1(_06756_),
    .B2(\fpga_top.io_frc.frc_cmp_val[46] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[47] ),
    .A1(_06755_));
 sg13g2_nand2b_1 _17435_ (.Y(_02823_),
    .B(\fpga_top.io_frc.frc_cmp_val[44] ),
    .A_N(\fpga_top.io_frc.frc_cntr_val[44] ));
 sg13g2_nand2b_1 _17436_ (.Y(_02824_),
    .B(\fpga_top.io_frc.frc_cmp_val[45] ),
    .A_N(\fpga_top.io_frc.frc_cntr_val[45] ));
 sg13g2_nand3_1 _17437_ (.B(_02823_),
    .C(_02824_),
    .A(_02822_),
    .Y(_02825_));
 sg13g2_inv_1 _17438_ (.Y(_02826_),
    .A(_02825_));
 sg13g2_nand2b_1 _17439_ (.Y(_02827_),
    .B(\fpga_top.io_frc.frc_cntr_val[42] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[42] ));
 sg13g2_nand2b_1 _17440_ (.Y(_02828_),
    .B(\fpga_top.io_frc.frc_cmp_val[41] ),
    .A_N(\fpga_top.io_frc.frc_cntr_val[41] ));
 sg13g2_nand2b_1 _17441_ (.Y(_02829_),
    .B(\fpga_top.io_frc.frc_cmp_val[42] ),
    .A_N(\fpga_top.io_frc.frc_cntr_val[42] ));
 sg13g2_nand2b_1 _17442_ (.Y(_02830_),
    .B(\fpga_top.io_frc.frc_cntr_val[43] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[43] ));
 sg13g2_nand3_1 _17443_ (.B(_02829_),
    .C(_02830_),
    .A(_02828_),
    .Y(_02831_));
 sg13g2_nand2b_1 _17444_ (.Y(_02832_),
    .B(\fpga_top.io_frc.frc_cmp_val[43] ),
    .A_N(\fpga_top.io_frc.frc_cntr_val[43] ));
 sg13g2_nor2b_1 _17445_ (.A(\fpga_top.io_frc.frc_cmp_val[41] ),
    .B_N(\fpga_top.io_frc.frc_cntr_val[41] ),
    .Y(_02833_));
 sg13g2_o21ai_1 _17446_ (.B1(_02827_),
    .Y(_02834_),
    .A1(_06754_),
    .A2(\fpga_top.io_frc.frc_cmp_val[40] ));
 sg13g2_o21ai_1 _17447_ (.B1(_02832_),
    .Y(_02835_),
    .A1(_02833_),
    .A2(_02834_));
 sg13g2_a21oi_1 _17448_ (.A1(_02827_),
    .A2(_02831_),
    .Y(_02836_),
    .B1(_02835_));
 sg13g2_nand2b_1 _17449_ (.Y(_02837_),
    .B(\fpga_top.io_frc.frc_cntr_val[44] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[44] ));
 sg13g2_nand2_1 _17450_ (.Y(_02838_),
    .A(_02830_),
    .B(_02837_));
 sg13g2_o21ai_1 _17451_ (.B1(_02826_),
    .Y(_02839_),
    .A1(_02836_),
    .A2(_02838_));
 sg13g2_nor2_1 _17452_ (.A(_06755_),
    .B(\fpga_top.io_frc.frc_cmp_val[47] ),
    .Y(_02840_));
 sg13g2_nand2b_1 _17453_ (.Y(_02841_),
    .B(\fpga_top.io_frc.frc_cntr_val[45] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[45] ));
 sg13g2_o21ai_1 _17454_ (.B1(_02841_),
    .Y(_02842_),
    .A1(_06756_),
    .A2(\fpga_top.io_frc.frc_cmp_val[46] ));
 sg13g2_a21oi_1 _17455_ (.A1(_02822_),
    .A2(_02842_),
    .Y(_02843_),
    .B1(_02840_));
 sg13g2_a22oi_1 _17456_ (.Y(_02844_),
    .B1(\fpga_top.io_frc.frc_cntr_val[38] ),
    .B2(_06759_),
    .A2(_06757_),
    .A1(\fpga_top.io_frc.frc_cntr_val[39] ));
 sg13g2_nor2_1 _17457_ (.A(_06760_),
    .B(\fpga_top.io_frc.frc_cmp_val[37] ),
    .Y(_02845_));
 sg13g2_a22oi_1 _17458_ (.Y(_02846_),
    .B1(_06761_),
    .B2(\fpga_top.io_frc.frc_cmp_val[36] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[37] ),
    .A1(_06760_));
 sg13g2_a22oi_1 _17459_ (.Y(_02847_),
    .B1(\fpga_top.io_frc.frc_cntr_val[35] ),
    .B2(_06763_),
    .A2(_06762_),
    .A1(\fpga_top.io_frc.frc_cntr_val[36] ));
 sg13g2_nor2_1 _17460_ (.A(\fpga_top.io_frc.frc_cntr_val[35] ),
    .B(_06763_),
    .Y(_02848_));
 sg13g2_nor2_1 _17461_ (.A(_06764_),
    .B(\fpga_top.io_frc.frc_cmp_val[34] ),
    .Y(_02849_));
 sg13g2_a22oi_1 _17462_ (.Y(_02850_),
    .B1(\fpga_top.io_frc.frc_cntr_val[32] ),
    .B2(_06768_),
    .A2(_06766_),
    .A1(\fpga_top.io_frc.frc_cntr_val[33] ));
 sg13g2_a22oi_1 _17463_ (.Y(_02851_),
    .B1(_06765_),
    .B2(\fpga_top.io_frc.frc_cmp_val[33] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[34] ),
    .A1(_06764_));
 sg13g2_nor2b_1 _17464_ (.A(_02850_),
    .B_N(_02851_),
    .Y(_02852_));
 sg13g2_nor2_1 _17465_ (.A(_02849_),
    .B(_02852_),
    .Y(_02853_));
 sg13g2_o21ai_1 _17466_ (.B1(_02847_),
    .Y(_02854_),
    .A1(_02848_),
    .A2(_02853_));
 sg13g2_a21oi_1 _17467_ (.A1(_02846_),
    .A2(_02854_),
    .Y(_02855_),
    .B1(_02845_));
 sg13g2_a21oi_1 _17468_ (.A1(_06758_),
    .A2(\fpga_top.io_frc.frc_cmp_val[38] ),
    .Y(_02856_),
    .B1(_02855_));
 sg13g2_nor2b_1 _17469_ (.A(_02856_),
    .B_N(_02844_),
    .Y(_02857_));
 sg13g2_nor2_1 _17470_ (.A(_06712_),
    .B(\fpga_top.io_frc.frc_cmp_val[31] ),
    .Y(_02858_));
 sg13g2_a22oi_1 _17471_ (.Y(_02859_),
    .B1(_06713_),
    .B2(\fpga_top.io_frc.frc_cmp_val[30] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[31] ),
    .A1(_06712_));
 sg13g2_nand2_1 _17472_ (.Y(_02860_),
    .A(_06717_),
    .B(\fpga_top.io_frc.frc_cmp_val[27] ));
 sg13g2_nand2b_1 _17473_ (.Y(_02861_),
    .B(\fpga_top.io_frc.frc_cntr_val[26] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[26] ));
 sg13g2_nor2_1 _17474_ (.A(_06717_),
    .B(\fpga_top.io_frc.frc_cmp_val[27] ),
    .Y(_02862_));
 sg13g2_a21oi_1 _17475_ (.A1(_06718_),
    .A2(\fpga_top.io_frc.frc_cmp_val[26] ),
    .Y(_02863_),
    .B1(_02862_));
 sg13g2_o21ai_1 _17476_ (.B1(_02863_),
    .Y(_02864_),
    .A1(\fpga_top.io_frc.frc_cntr_val[25] ),
    .A2(_06720_));
 sg13g2_a22oi_1 _17477_ (.Y(_02865_),
    .B1(\fpga_top.io_frc.frc_cntr_val[24] ),
    .B2(_06722_),
    .A2(_06720_),
    .A1(\fpga_top.io_frc.frc_cntr_val[25] ));
 sg13g2_o21ai_1 _17478_ (.B1(_02861_),
    .Y(_02866_),
    .A1(_02864_),
    .A2(_02865_));
 sg13g2_a221oi_1 _17479_ (.B2(_02866_),
    .C1(_02862_),
    .B1(_02860_),
    .A1(\fpga_top.io_frc.frc_cntr_val[28] ),
    .Y(_02867_),
    .A2(_06716_));
 sg13g2_a221oi_1 _17480_ (.B2(\fpga_top.io_frc.frc_cmp_val[28] ),
    .C1(_02867_),
    .B1(_06715_),
    .A1(_06714_),
    .Y(_02868_),
    .A2(\fpga_top.io_frc.frc_cmp_val[29] ));
 sg13g2_nand2b_1 _17481_ (.Y(_02869_),
    .B(\fpga_top.io_frc.frc_cntr_val[29] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[29] ));
 sg13g2_o21ai_1 _17482_ (.B1(_02869_),
    .Y(_02870_),
    .A1(_06713_),
    .A2(\fpga_top.io_frc.frc_cmp_val[30] ));
 sg13g2_o21ai_1 _17483_ (.B1(_02859_),
    .Y(_02871_),
    .A1(_02868_),
    .A2(_02870_));
 sg13g2_nand2b_1 _17484_ (.Y(_02872_),
    .B(_02871_),
    .A_N(_02858_));
 sg13g2_nor2_1 _17485_ (.A(\fpga_top.io_frc.frc_cntr_val[15] ),
    .B(_06698_),
    .Y(_02873_));
 sg13g2_a22oi_1 _17486_ (.Y(_02874_),
    .B1(\fpga_top.io_frc.frc_cntr_val[14] ),
    .B2(_06700_),
    .A2(_06698_),
    .A1(\fpga_top.io_frc.frc_cntr_val[15] ));
 sg13g2_a22oi_1 _17487_ (.Y(_02875_),
    .B1(_06701_),
    .B2(\fpga_top.io_frc.frc_cmp_val[13] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[14] ),
    .A1(_06699_));
 sg13g2_nand2_1 _17488_ (.Y(_02876_),
    .A(\fpga_top.io_frc.frc_cntr_val[12] ),
    .B(_06704_));
 sg13g2_o21ai_1 _17489_ (.B1(_02876_),
    .Y(_02877_),
    .A1(_06701_),
    .A2(\fpga_top.io_frc.frc_cmp_val[13] ));
 sg13g2_nand2_1 _17490_ (.Y(_02878_),
    .A(_02875_),
    .B(_02877_));
 sg13g2_a21oi_1 _17491_ (.A1(_02874_),
    .A2(_02878_),
    .Y(_02879_),
    .B1(_02873_));
 sg13g2_nand2_1 _17492_ (.Y(_02880_),
    .A(\fpga_top.io_frc.frc_cntr_val[7] ),
    .B(_06691_));
 sg13g2_nor2_1 _17493_ (.A(\fpga_top.io_frc.frc_cntr_val[6] ),
    .B(_06692_),
    .Y(_02881_));
 sg13g2_nand2b_1 _17494_ (.Y(_02882_),
    .B(\fpga_top.io_frc.frc_cntr_val[1] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[1] ));
 sg13g2_a22oi_1 _17495_ (.Y(_02883_),
    .B1(_06686_),
    .B2(\fpga_top.io_frc.frc_cmp_val[1] ),
    .A2(_06685_),
    .A1(\fpga_top.io_frc.frc_cmp_val[0] ));
 sg13g2_o21ai_1 _17496_ (.B1(_02882_),
    .Y(_02884_),
    .A1(_06689_),
    .A2(\fpga_top.io_frc.frc_cmp_val[2] ));
 sg13g2_nor2_1 _17497_ (.A(_02883_),
    .B(_02884_),
    .Y(_02885_));
 sg13g2_a221oi_1 _17498_ (.B2(\fpga_top.io_frc.frc_cmp_val[2] ),
    .C1(_02885_),
    .B1(_06689_),
    .A1(_06687_),
    .Y(_02886_),
    .A2(\fpga_top.io_frc.frc_cmp_val[3] ));
 sg13g2_a221oi_1 _17499_ (.B2(_06696_),
    .C1(_02886_),
    .B1(\fpga_top.io_frc.frc_cntr_val[4] ),
    .A1(\fpga_top.io_frc.frc_cntr_val[3] ),
    .Y(_02887_),
    .A2(_06688_));
 sg13g2_a221oi_1 _17500_ (.B2(\fpga_top.io_frc.frc_cmp_val[4] ),
    .C1(_02887_),
    .B1(_06695_),
    .A1(_06693_),
    .Y(_02888_),
    .A2(\fpga_top.io_frc.frc_cmp_val[5] ));
 sg13g2_a221oi_1 _17501_ (.B2(_06694_),
    .C1(_02888_),
    .B1(\fpga_top.io_frc.frc_cntr_val[5] ),
    .A1(\fpga_top.io_frc.frc_cntr_val[6] ),
    .Y(_02889_),
    .A2(_06692_));
 sg13g2_o21ai_1 _17502_ (.B1(_02880_),
    .Y(_02890_),
    .A1(_02881_),
    .A2(_02889_));
 sg13g2_a22oi_1 _17503_ (.Y(_02891_),
    .B1(_06710_),
    .B2(\fpga_top.io_frc.frc_cmp_val[8] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[7] ),
    .A1(_06690_));
 sg13g2_nor2_1 _17504_ (.A(_06710_),
    .B(\fpga_top.io_frc.frc_cmp_val[8] ),
    .Y(_02892_));
 sg13g2_a221oi_1 _17505_ (.B2(_02891_),
    .C1(_02892_),
    .B1(_02890_),
    .A1(\fpga_top.io_frc.frc_cntr_val[9] ),
    .Y(_02893_),
    .A2(_06709_));
 sg13g2_a221oi_1 _17506_ (.B2(\fpga_top.io_frc.frc_cmp_val[9] ),
    .C1(_02893_),
    .B1(_06708_),
    .A1(_06706_),
    .Y(_02894_),
    .A2(\fpga_top.io_frc.frc_cmp_val[10] ));
 sg13g2_a221oi_1 _17507_ (.B2(_06707_),
    .C1(_02894_),
    .B1(\fpga_top.io_frc.frc_cntr_val[10] ),
    .A1(\fpga_top.io_frc.frc_cntr_val[11] ),
    .Y(_02895_),
    .A2(_06705_));
 sg13g2_nand2_1 _17508_ (.Y(_02896_),
    .A(_06703_),
    .B(\fpga_top.io_frc.frc_cmp_val[12] ));
 sg13g2_o21ai_1 _17509_ (.B1(_02896_),
    .Y(_02897_),
    .A1(\fpga_top.io_frc.frc_cntr_val[11] ),
    .A2(_06705_));
 sg13g2_and2_1 _17510_ (.A(_02874_),
    .B(_02875_),
    .X(_02898_));
 sg13g2_nor4_1 _17511_ (.A(_02873_),
    .B(_02877_),
    .C(_02895_),
    .D(_02897_),
    .Y(_02899_));
 sg13g2_a21oi_1 _17512_ (.A1(_02898_),
    .A2(_02899_),
    .Y(_02900_),
    .B1(_02879_));
 sg13g2_a22oi_1 _17513_ (.Y(_02901_),
    .B1(\fpga_top.io_frc.frc_cntr_val[21] ),
    .B2(_06727_),
    .A2(_06725_),
    .A1(\fpga_top.io_frc.frc_cntr_val[22] ));
 sg13g2_a22oi_1 _17514_ (.Y(_02902_),
    .B1(_06728_),
    .B2(\fpga_top.io_frc.frc_cmp_val[20] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[21] ),
    .A1(_06726_));
 sg13g2_nand2b_1 _17515_ (.Y(_02903_),
    .B(\fpga_top.io_frc.frc_cntr_val[16] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[16] ));
 sg13g2_o21ai_1 _17516_ (.B1(_02903_),
    .Y(_02904_),
    .A1(_06729_),
    .A2(\fpga_top.io_frc.frc_cmp_val[17] ));
 sg13g2_nor2_1 _17517_ (.A(_06731_),
    .B(\fpga_top.io_frc.frc_cmp_val[19] ),
    .Y(_02905_));
 sg13g2_a21oi_1 _17518_ (.A1(_06732_),
    .A2(\fpga_top.io_frc.frc_cmp_val[18] ),
    .Y(_02906_),
    .B1(_02905_));
 sg13g2_nand3_1 _17519_ (.B(_02902_),
    .C(_02906_),
    .A(_02901_),
    .Y(_02907_));
 sg13g2_nor2b_1 _17520_ (.A(\fpga_top.io_frc.frc_cntr_val[17] ),
    .B_N(\fpga_top.io_frc.frc_cmp_val[17] ),
    .Y(_02908_));
 sg13g2_nand2_1 _17521_ (.Y(_02909_),
    .A(_06729_),
    .B(\fpga_top.io_frc.frc_cmp_val[17] ));
 sg13g2_nor2_1 _17522_ (.A(_06728_),
    .B(\fpga_top.io_frc.frc_cmp_val[20] ),
    .Y(_02910_));
 sg13g2_nor2_1 _17523_ (.A(_06723_),
    .B(\fpga_top.io_frc.frc_cmp_val[23] ),
    .Y(_02911_));
 sg13g2_nor2b_1 _17524_ (.A(\fpga_top.io_frc.frc_cntr_val[16] ),
    .B_N(\fpga_top.io_frc.frc_cmp_val[16] ),
    .Y(_02912_));
 sg13g2_nor4_1 _17525_ (.A(_02908_),
    .B(_02910_),
    .C(_02911_),
    .D(_02912_),
    .Y(_02913_));
 sg13g2_a22oi_1 _17526_ (.Y(_02914_),
    .B1(_06724_),
    .B2(\fpga_top.io_frc.frc_cmp_val[22] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[23] ),
    .A1(_06723_));
 sg13g2_nand2_1 _17527_ (.Y(_02915_),
    .A(_06731_),
    .B(\fpga_top.io_frc.frc_cmp_val[19] ));
 sg13g2_nand2b_1 _17528_ (.Y(_02916_),
    .B(\fpga_top.io_frc.frc_cntr_val[18] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[18] ));
 sg13g2_nand4_1 _17529_ (.B(_02914_),
    .C(_02915_),
    .A(_02913_),
    .Y(_02917_),
    .D(_02916_));
 sg13g2_nor4_1 _17530_ (.A(_02900_),
    .B(_02904_),
    .C(_02907_),
    .D(_02917_),
    .Y(_02918_));
 sg13g2_nand3_1 _17531_ (.B(_02906_),
    .C(_02909_),
    .A(_02904_),
    .Y(_02919_));
 sg13g2_a22oi_1 _17532_ (.Y(_02920_),
    .B1(_02916_),
    .B2(_02919_),
    .A2(\fpga_top.io_frc.frc_cmp_val[19] ),
    .A1(_06731_));
 sg13g2_or2_1 _17533_ (.X(_02921_),
    .B(_02910_),
    .A(_02905_));
 sg13g2_o21ai_1 _17534_ (.B1(_02902_),
    .Y(_02922_),
    .A1(_02920_),
    .A2(_02921_));
 sg13g2_nand2_1 _17535_ (.Y(_02923_),
    .A(_02901_),
    .B(_02922_));
 sg13g2_a21oi_1 _17536_ (.A1(_02914_),
    .A2(_02923_),
    .Y(_02924_),
    .B1(_02911_));
 sg13g2_nor2b_2 _17537_ (.A(_02918_),
    .B_N(_02924_),
    .Y(_02925_));
 sg13g2_a221oi_1 _17538_ (.B2(\fpga_top.io_frc.frc_cmp_val[28] ),
    .C1(_02870_),
    .B1(_06715_),
    .A1(_06714_),
    .Y(_02926_),
    .A2(\fpga_top.io_frc.frc_cmp_val[29] ));
 sg13g2_nand2_1 _17539_ (.Y(_02927_),
    .A(_02865_),
    .B(_02926_));
 sg13g2_a221oi_1 _17540_ (.B2(\fpga_top.io_frc.frc_cmp_val[24] ),
    .C1(_02858_),
    .B1(_06721_),
    .A1(\fpga_top.io_frc.frc_cntr_val[28] ),
    .Y(_02928_),
    .A2(_06716_));
 sg13g2_nand4_1 _17541_ (.B(_02860_),
    .C(_02861_),
    .A(_02859_),
    .Y(_02929_),
    .D(_02928_));
 sg13g2_nor4_1 _17542_ (.A(_02864_),
    .B(_02925_),
    .C(_02927_),
    .D(_02929_),
    .Y(_02930_));
 sg13g2_nor2_1 _17543_ (.A(_02872_),
    .B(_02930_),
    .Y(_02931_));
 sg13g2_and4_1 _17544_ (.A(_02846_),
    .B(_02847_),
    .C(_02850_),
    .D(_02851_),
    .X(_02932_));
 sg13g2_a221oi_1 _17545_ (.B2(\fpga_top.io_frc.frc_cmp_val[32] ),
    .C1(_02845_),
    .B1(_06767_),
    .A1(_06758_),
    .Y(_02933_),
    .A2(\fpga_top.io_frc.frc_cmp_val[38] ));
 sg13g2_nor2_1 _17546_ (.A(_02848_),
    .B(_02849_),
    .Y(_02934_));
 sg13g2_nand4_1 _17547_ (.B(_02932_),
    .C(_02933_),
    .A(_02844_),
    .Y(_02935_),
    .D(_02934_));
 sg13g2_o21ai_1 _17548_ (.B1(_02857_),
    .Y(_02936_),
    .A1(_02931_),
    .A2(_02935_));
 sg13g2_nand2b_1 _17549_ (.Y(_02937_),
    .B(\fpga_top.io_frc.frc_cmp_val[39] ),
    .A_N(\fpga_top.io_frc.frc_cntr_val[39] ));
 sg13g2_nand3_1 _17550_ (.B(_02837_),
    .C(_02937_),
    .A(_02832_),
    .Y(_02938_));
 sg13g2_nor2b_1 _17551_ (.A(\fpga_top.io_frc.frc_cntr_val[40] ),
    .B_N(\fpga_top.io_frc.frc_cmp_val[40] ),
    .Y(_02939_));
 sg13g2_nor4_1 _17552_ (.A(_02840_),
    .B(_02842_),
    .C(_02938_),
    .D(_02939_),
    .Y(_02940_));
 sg13g2_nor4_1 _17553_ (.A(_02825_),
    .B(_02831_),
    .C(_02833_),
    .D(_02834_),
    .Y(_02941_));
 sg13g2_nand3_1 _17554_ (.B(_02940_),
    .C(_02941_),
    .A(_02936_),
    .Y(_02942_));
 sg13g2_nand3_1 _17555_ (.B(_02843_),
    .C(_02942_),
    .A(_02839_),
    .Y(_02943_));
 sg13g2_nand2b_1 _17556_ (.Y(_02944_),
    .B(\fpga_top.io_frc.frc_cmp_val[60] ),
    .A_N(\fpga_top.io_frc.frc_cntr_val[60] ));
 sg13g2_o21ai_1 _17557_ (.B1(_02944_),
    .Y(_02945_),
    .A1(\fpga_top.io_frc.frc_cntr_val[61] ),
    .A2(_06736_));
 sg13g2_nor2b_1 _17558_ (.A(\fpga_top.io_frc.frc_cmp_val[60] ),
    .B_N(\fpga_top.io_frc.frc_cntr_val[60] ),
    .Y(_02946_));
 sg13g2_nor2_1 _17559_ (.A(_06738_),
    .B(\fpga_top.io_frc.frc_cmp_val[58] ),
    .Y(_02947_));
 sg13g2_nand2b_1 _17560_ (.Y(_02948_),
    .B(\fpga_top.io_frc.frc_cntr_val[57] ),
    .A_N(\fpga_top.io_frc.frc_cmp_val[57] ));
 sg13g2_o21ai_1 _17561_ (.B1(_02948_),
    .Y(_02949_),
    .A1(_06740_),
    .A2(\fpga_top.io_frc.frc_cmp_val[56] ));
 sg13g2_a22oi_1 _17562_ (.Y(_02950_),
    .B1(_06734_),
    .B2(\fpga_top.io_frc.frc_cmp_val[62] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[63] ),
    .A1(_06733_));
 sg13g2_nor2_1 _17563_ (.A(_06733_),
    .B(\fpga_top.io_frc.frc_cmp_val[63] ),
    .Y(_02951_));
 sg13g2_nor2b_1 _17564_ (.A(\fpga_top.io_frc.frc_cntr_val[59] ),
    .B_N(\fpga_top.io_frc.frc_cmp_val[59] ),
    .Y(_02952_));
 sg13g2_nor2b_1 _17565_ (.A(\fpga_top.io_frc.frc_cntr_val[57] ),
    .B_N(\fpga_top.io_frc.frc_cmp_val[57] ),
    .Y(_02953_));
 sg13g2_nor2b_1 _17566_ (.A(\fpga_top.io_frc.frc_cntr_val[56] ),
    .B_N(\fpga_top.io_frc.frc_cmp_val[56] ),
    .Y(_02954_));
 sg13g2_a22oi_1 _17567_ (.Y(_02955_),
    .B1(\fpga_top.io_frc.frc_cntr_val[61] ),
    .B2(_06736_),
    .A2(_06735_),
    .A1(\fpga_top.io_frc.frc_cntr_val[62] ));
 sg13g2_nor2b_1 _17568_ (.A(\fpga_top.io_frc.frc_cmp_val[59] ),
    .B_N(\fpga_top.io_frc.frc_cntr_val[59] ),
    .Y(_02956_));
 sg13g2_nor2b_1 _17569_ (.A(\fpga_top.io_frc.frc_cntr_val[58] ),
    .B_N(\fpga_top.io_frc.frc_cmp_val[58] ),
    .Y(_02957_));
 sg13g2_nor4_1 _17570_ (.A(_02946_),
    .B(_02947_),
    .C(_02952_),
    .D(_02954_),
    .Y(_02958_));
 sg13g2_nor3_1 _17571_ (.A(_02945_),
    .B(_02956_),
    .C(_02957_),
    .Y(_02959_));
 sg13g2_nand4_1 _17572_ (.B(_02955_),
    .C(_02958_),
    .A(_02950_),
    .Y(_02960_),
    .D(_02959_));
 sg13g2_nor4_2 _17573_ (.A(_02949_),
    .B(_02951_),
    .C(_02953_),
    .Y(_02961_),
    .D(_02960_));
 sg13g2_a22oi_1 _17574_ (.Y(_02962_),
    .B1(\fpga_top.io_frc.frc_cntr_val[54] ),
    .B2(_06750_),
    .A2(_06749_),
    .A1(\fpga_top.io_frc.frc_cntr_val[55] ));
 sg13g2_a22oi_1 _17575_ (.Y(_02963_),
    .B1(\fpga_top.io_frc.frc_cntr_val[52] ),
    .B2(_06753_),
    .A2(_06745_),
    .A1(\fpga_top.io_frc.frc_cntr_val[51] ));
 sg13g2_a22oi_1 _17576_ (.Y(_02964_),
    .B1(_06746_),
    .B2(\fpga_top.io_frc.frc_cmp_val[50] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[51] ),
    .A1(_06744_));
 sg13g2_a22oi_1 _17577_ (.Y(_02965_),
    .B1(\fpga_top.io_frc.frc_cntr_val[50] ),
    .B2(_06747_),
    .A2(_06743_),
    .A1(\fpga_top.io_frc.frc_cntr_val[48] ));
 sg13g2_nand4_1 _17578_ (.B(_02963_),
    .C(_02964_),
    .A(_02962_),
    .Y(_02966_),
    .D(_02965_));
 sg13g2_nor2_1 _17579_ (.A(\fpga_top.io_frc.frc_cntr_val[49] ),
    .B(_06741_),
    .Y(_02967_));
 sg13g2_nor2_1 _17580_ (.A(\fpga_top.io_frc.frc_cntr_val[48] ),
    .B(_06743_),
    .Y(_02968_));
 sg13g2_nor2_1 _17581_ (.A(\fpga_top.io_frc.frc_cntr_val[54] ),
    .B(_06750_),
    .Y(_02969_));
 sg13g2_nor2b_1 _17582_ (.A(\fpga_top.io_frc.frc_cmp_val[49] ),
    .B_N(\fpga_top.io_frc.frc_cntr_val[49] ),
    .Y(_02970_));
 sg13g2_or4_1 _17583_ (.A(_02967_),
    .B(_02968_),
    .C(_02969_),
    .D(_02970_),
    .X(_02971_));
 sg13g2_a22oi_1 _17584_ (.Y(_02972_),
    .B1(_06752_),
    .B2(\fpga_top.io_frc.frc_cmp_val[52] ),
    .A2(\fpga_top.io_frc.frc_cmp_val[53] ),
    .A1(_06751_));
 sg13g2_nor2_1 _17585_ (.A(_06751_),
    .B(\fpga_top.io_frc.frc_cmp_val[53] ),
    .Y(_02973_));
 sg13g2_nand2_1 _17586_ (.Y(_02974_),
    .A(_06748_),
    .B(\fpga_top.io_frc.frc_cmp_val[55] ));
 sg13g2_nand3b_1 _17587_ (.B(_02974_),
    .C(_02972_),
    .Y(_02975_),
    .A_N(_02973_));
 sg13g2_nor3_1 _17588_ (.A(_02966_),
    .B(_02971_),
    .C(_02975_),
    .Y(_02976_));
 sg13g2_nand3_1 _17589_ (.B(_02961_),
    .C(_02976_),
    .A(_02943_),
    .Y(_02977_));
 sg13g2_nor2b_1 _17590_ (.A(_02970_),
    .B_N(_02965_),
    .Y(_02978_));
 sg13g2_o21ai_1 _17591_ (.B1(_02967_),
    .Y(_02979_),
    .A1(_06746_),
    .A2(\fpga_top.io_frc.frc_cmp_val[50] ));
 sg13g2_nand2_1 _17592_ (.Y(_02980_),
    .A(_02964_),
    .B(_02979_));
 sg13g2_o21ai_1 _17593_ (.B1(_02963_),
    .Y(_02981_),
    .A1(_02978_),
    .A2(_02980_));
 sg13g2_a21oi_1 _17594_ (.A1(_02972_),
    .A2(_02981_),
    .Y(_02982_),
    .B1(_02973_));
 sg13g2_o21ai_1 _17595_ (.B1(_02962_),
    .Y(_02983_),
    .A1(_02969_),
    .A2(_02982_));
 sg13g2_nand3_1 _17596_ (.B(_02974_),
    .C(_02983_),
    .A(_02961_),
    .Y(_02984_));
 sg13g2_nor3_1 _17597_ (.A(_02953_),
    .B(_02956_),
    .C(_02957_),
    .Y(_02985_));
 sg13g2_a21oi_1 _17598_ (.A1(_02949_),
    .A2(_02985_),
    .Y(_02986_),
    .B1(_02947_));
 sg13g2_nor2_1 _17599_ (.A(_02952_),
    .B(_02986_),
    .Y(_02987_));
 sg13g2_nor3_1 _17600_ (.A(_02946_),
    .B(_02956_),
    .C(_02987_),
    .Y(_02988_));
 sg13g2_o21ai_1 _17601_ (.B1(_02955_),
    .Y(_02989_),
    .A1(_02945_),
    .A2(_02988_));
 sg13g2_a21oi_1 _17602_ (.A1(_02950_),
    .A2(_02989_),
    .Y(_02990_),
    .B1(_02951_));
 sg13g2_nand3_1 _17603_ (.B(_02984_),
    .C(_02990_),
    .A(_02977_),
    .Y(_02991_));
 sg13g2_nand3_1 _17604_ (.B(\fpga_top.io_frc.frc_cntrl_val ),
    .C(_02991_),
    .A(\fpga_top.cpu_top.csr_mtie ),
    .Y(_02992_));
 sg13g2_a221oi_1 _17605_ (.B2(_06773_),
    .C1(net1381),
    .B1(_02992_),
    .A1(_08912_),
    .Y(_00328_),
    .A2(net4852));
 sg13g2_nand2_2 _17606_ (.Y(_02993_),
    .A(_09658_),
    .B(_09804_));
 sg13g2_or2_1 _17607_ (.X(_02994_),
    .B(_02993_),
    .A(_09803_));
 sg13g2_mux2_1 _17608_ (.A0(net4364),
    .A1(net2933),
    .S(net4175),
    .X(_00329_));
 sg13g2_mux2_1 _17609_ (.A0(net4360),
    .A1(net2843),
    .S(net4177),
    .X(_00330_));
 sg13g2_mux2_1 _17610_ (.A0(net4354),
    .A1(net2746),
    .S(net4176),
    .X(_00331_));
 sg13g2_mux2_1 _17611_ (.A0(net4348),
    .A1(net2617),
    .S(net4175),
    .X(_00332_));
 sg13g2_mux2_1 _17612_ (.A0(net4341),
    .A1(net2308),
    .S(net4177),
    .X(_00333_));
 sg13g2_mux2_1 _17613_ (.A0(net4199),
    .A1(net2350),
    .S(net4177),
    .X(_00334_));
 sg13g2_mux2_1 _17614_ (.A0(net4336),
    .A1(net2954),
    .S(net4175),
    .X(_00335_));
 sg13g2_mux2_1 _17615_ (.A0(net4332),
    .A1(net2575),
    .S(net4178),
    .X(_00336_));
 sg13g2_mux2_1 _17616_ (.A0(net4328),
    .A1(net3564),
    .S(net4177),
    .X(_00337_));
 sg13g2_mux2_1 _17617_ (.A0(net4318),
    .A1(net2409),
    .S(net4176),
    .X(_00338_));
 sg13g2_mux2_1 _17618_ (.A0(net4193),
    .A1(net2882),
    .S(net4178),
    .X(_00339_));
 sg13g2_mux2_1 _17619_ (.A0(net4189),
    .A1(net2346),
    .S(net4176),
    .X(_00340_));
 sg13g2_mux2_1 _17620_ (.A0(net4317),
    .A1(net3124),
    .S(net4178),
    .X(_00341_));
 sg13g2_mux2_1 _17621_ (.A0(net4311),
    .A1(net2735),
    .S(net4176),
    .X(_00342_));
 sg13g2_mux2_1 _17622_ (.A0(net4303),
    .A1(net2638),
    .S(net4175),
    .X(_00343_));
 sg13g2_mux2_1 _17623_ (.A0(net4299),
    .A1(net3640),
    .S(net4178),
    .X(_00344_));
 sg13g2_mux2_1 _17624_ (.A0(net4293),
    .A1(net2237),
    .S(net4178),
    .X(_00345_));
 sg13g2_mux2_1 _17625_ (.A0(net4287),
    .A1(net2778),
    .S(net4175),
    .X(_00346_));
 sg13g2_mux2_1 _17626_ (.A0(net4282),
    .A1(net2913),
    .S(net4178),
    .X(_00347_));
 sg13g2_mux2_1 _17627_ (.A0(net4278),
    .A1(net2161),
    .S(net4175),
    .X(_00348_));
 sg13g2_mux2_1 _17628_ (.A0(net4271),
    .A1(net2140),
    .S(net4177),
    .X(_00349_));
 sg13g2_mux2_1 _17629_ (.A0(net4264),
    .A1(net2326),
    .S(net4175),
    .X(_00350_));
 sg13g2_mux2_1 _17630_ (.A0(net4262),
    .A1(net2472),
    .S(net4179),
    .X(_00351_));
 sg13g2_mux2_1 _17631_ (.A0(net4258),
    .A1(net2256),
    .S(net4178),
    .X(_00352_));
 sg13g2_mux2_1 _17632_ (.A0(net4406),
    .A1(net2767),
    .S(net4179),
    .X(_00353_));
 sg13g2_mux2_1 _17633_ (.A0(net4401),
    .A1(net2770),
    .S(net4177),
    .X(_00354_));
 sg13g2_mux2_1 _17634_ (.A0(net4396),
    .A1(net3668),
    .S(net4176),
    .X(_00355_));
 sg13g2_mux2_1 _17635_ (.A0(net4390),
    .A1(net2644),
    .S(net4176),
    .X(_00356_));
 sg13g2_mux2_1 _17636_ (.A0(net4382),
    .A1(net2459),
    .S(net4175),
    .X(_00357_));
 sg13g2_mux2_1 _17637_ (.A0(net4380),
    .A1(net2483),
    .S(net4178),
    .X(_00358_));
 sg13g2_mux2_1 _17638_ (.A0(net4374),
    .A1(net2349),
    .S(net4177),
    .X(_00359_));
 sg13g2_mux2_1 _17639_ (.A0(net4371),
    .A1(net2503),
    .S(net4177),
    .X(_00360_));
 sg13g2_nand2_2 _17640_ (.Y(_02995_),
    .A(_08909_),
    .B(_10553_));
 sg13g2_nor2_2 _17641_ (.A(_09617_),
    .B(_02995_),
    .Y(_02996_));
 sg13g2_nor2b_2 _17642_ (.A(net4460),
    .B_N(net5601),
    .Y(_02997_));
 sg13g2_o21ai_1 _17643_ (.B1(net5603),
    .Y(_02998_),
    .A1(_09617_),
    .A2(_02995_));
 sg13g2_nand2_2 _17644_ (.Y(_02999_),
    .A(net5600),
    .B(_10526_));
 sg13g2_o21ai_1 _17645_ (.B1(_02999_),
    .Y(_03000_),
    .A1(net8),
    .A2(net5599));
 sg13g2_nor2_1 _17646_ (.A(_02997_),
    .B(_03000_),
    .Y(_03001_));
 sg13g2_a21oi_1 _17647_ (.A1(_06831_),
    .A2(_02997_),
    .Y(_00361_),
    .B1(_03001_));
 sg13g2_nand2_1 _17648_ (.Y(_03002_),
    .A(net5599),
    .B(net4845));
 sg13g2_nand3_1 _17649_ (.B(net4845),
    .C(net4460),
    .A(net5602),
    .Y(_03003_));
 sg13g2_o21ai_1 _17650_ (.B1(_03003_),
    .Y(_00362_),
    .A1(_06832_),
    .A2(net4458));
 sg13g2_nor2_1 _17651_ (.A(_06812_),
    .B(net5602),
    .Y(_03004_));
 sg13g2_nor3_1 _17652_ (.A(net8),
    .B(net7),
    .C(net5602),
    .Y(_03005_));
 sg13g2_a221oi_1 _17653_ (.B2(net7),
    .C1(_03005_),
    .B1(_03004_),
    .A1(net5602),
    .Y(_03006_),
    .A2(net4851));
 sg13g2_nand2_1 _17654_ (.Y(_03007_),
    .A(net4458),
    .B(_03006_));
 sg13g2_o21ai_1 _17655_ (.B1(_03007_),
    .Y(_00363_),
    .A1(_06833_),
    .A2(net4458));
 sg13g2_nand2_1 _17656_ (.Y(_03008_),
    .A(net5599),
    .B(net4842));
 sg13g2_nand3_1 _17657_ (.B(net4844),
    .C(net4460),
    .A(net5602),
    .Y(_03009_));
 sg13g2_a21oi_1 _17658_ (.A1(net2113),
    .A2(_02997_),
    .Y(_03010_),
    .B1(_03004_));
 sg13g2_nand2_1 _17659_ (.Y(_00364_),
    .A(_03009_),
    .B(_03010_));
 sg13g2_a21oi_1 _17660_ (.A1(_06812_),
    .A2(net7),
    .Y(_03011_),
    .B1(net5601));
 sg13g2_nand2_1 _17661_ (.Y(_03012_),
    .A(net5601),
    .B(net4838));
 sg13g2_a21oi_1 _17662_ (.A1(net5601),
    .A2(net4838),
    .Y(_03013_),
    .B1(_03011_));
 sg13g2_nor2_1 _17663_ (.A(net3973),
    .B(net4458),
    .Y(_03014_));
 sg13g2_a21oi_1 _17664_ (.A1(net4458),
    .A2(_03013_),
    .Y(_00365_),
    .B1(_03014_));
 sg13g2_nand2_1 _17665_ (.Y(_03015_),
    .A(net5601),
    .B(net4834));
 sg13g2_a221oi_1 _17666_ (.B2(net7),
    .C1(_02997_),
    .B1(_03004_),
    .A1(net5602),
    .Y(_03016_),
    .A2(net4834));
 sg13g2_a21oi_1 _17667_ (.A1(_06836_),
    .A2(_02997_),
    .Y(_00366_),
    .B1(_03016_));
 sg13g2_a21oi_1 _17668_ (.A1(net5602),
    .A2(_02756_),
    .Y(_03017_),
    .B1(_03005_));
 sg13g2_nor2_1 _17669_ (.A(net3142),
    .B(net4458),
    .Y(_03018_));
 sg13g2_a21oi_1 _17670_ (.A1(net4458),
    .A2(_03017_),
    .Y(_00367_),
    .B1(_03018_));
 sg13g2_nand3_1 _17671_ (.B(_02760_),
    .C(net4460),
    .A(net5601),
    .Y(_03019_));
 sg13g2_a21oi_1 _17672_ (.A1(net3606),
    .A2(_02997_),
    .Y(_03020_),
    .B1(_03011_));
 sg13g2_nand2_1 _17673_ (.Y(_00368_),
    .A(_03019_),
    .B(_03020_));
 sg13g2_and2_1 _17674_ (.A(net5603),
    .B(_02763_),
    .X(_03021_));
 sg13g2_a221oi_1 _17675_ (.B2(net4460),
    .C1(_03011_),
    .B1(_03021_),
    .A1(_06839_),
    .Y(_00369_),
    .A2(_02997_));
 sg13g2_nand3_1 _17676_ (.B(_02768_),
    .C(net4459),
    .A(net5604),
    .Y(_03022_));
 sg13g2_o21ai_1 _17677_ (.B1(_03022_),
    .Y(_00370_),
    .A1(_06840_),
    .A2(net4458));
 sg13g2_nand3_1 _17678_ (.B(_08981_),
    .C(net4460),
    .A(net5603),
    .Y(_03023_));
 sg13g2_o21ai_1 _17679_ (.B1(_03023_),
    .Y(_00371_),
    .A1(_06841_),
    .A2(_02998_));
 sg13g2_o21ai_1 _17680_ (.B1(net5603),
    .Y(_03024_),
    .A1(net6174),
    .A2(net4459));
 sg13g2_a21oi_1 _17681_ (.A1(_02771_),
    .A2(net4459),
    .Y(_00372_),
    .B1(_03024_));
 sg13g2_o21ai_1 _17682_ (.B1(net5604),
    .Y(_03025_),
    .A1(net4022),
    .A2(_02996_));
 sg13g2_a21oi_1 _17683_ (.A1(_02775_),
    .A2(net4460),
    .Y(_00373_),
    .B1(_03025_));
 sg13g2_o21ai_1 _17684_ (.B1(net5604),
    .Y(_03026_),
    .A1(net4043),
    .A2(_02996_));
 sg13g2_a21oi_1 _17685_ (.A1(_02778_),
    .A2(net4459),
    .Y(_00374_),
    .B1(_03026_));
 sg13g2_o21ai_1 _17686_ (.B1(net5604),
    .Y(_03027_),
    .A1(net6111),
    .A2(net4459));
 sg13g2_a21oi_1 _17687_ (.A1(_02781_),
    .A2(net4459),
    .Y(_00375_),
    .B1(_03027_));
 sg13g2_o21ai_1 _17688_ (.B1(net5603),
    .Y(_03028_),
    .A1(net6147),
    .A2(net4459));
 sg13g2_a21oi_1 _17689_ (.A1(_02784_),
    .A2(net4459),
    .Y(_00376_),
    .B1(_03028_));
 sg13g2_and2_1 _17690_ (.A(net3560),
    .B(_10556_),
    .X(_03029_));
 sg13g2_xor2_1 _17691_ (.B(_10557_),
    .A(net3560),
    .X(_00377_));
 sg13g2_nor3_2 _17692_ (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[1] ),
    .B(_08989_),
    .C(_10555_),
    .Y(_03030_));
 sg13g2_xor2_1 _17693_ (.B(_03029_),
    .A(net2062),
    .X(_00378_));
 sg13g2_nand2_1 _17694_ (.Y(_03031_),
    .A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[1] ),
    .B(_10557_));
 sg13g2_nand2_1 _17695_ (.Y(_03032_),
    .A(net2062),
    .B(_03029_));
 sg13g2_nand3_1 _17696_ (.B(_06928_),
    .C(_03029_),
    .A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[1] ),
    .Y(_03033_));
 sg13g2_xnor2_1 _17697_ (.Y(_00379_),
    .A(net3691),
    .B(_03032_));
 sg13g2_nor2_1 _17698_ (.A(_08911_),
    .B(_09617_),
    .Y(_03034_));
 sg13g2_nor2_1 _17699_ (.A(net3627),
    .B(_03034_),
    .Y(_03035_));
 sg13g2_a21oi_1 _17700_ (.A1(net4920),
    .A2(_03034_),
    .Y(_00380_),
    .B1(_03035_));
 sg13g2_a21oi_1 _17701_ (.A1(\fpga_top.io_uart_out.rx_first_read ),
    .A2(_02738_),
    .Y(_03036_),
    .B1(net1405));
 sg13g2_nor2_1 _17702_ (.A(net1387),
    .B(net1406),
    .Y(_00381_));
 sg13g2_a21oi_1 _17703_ (.A1(_06678_),
    .A2(net5328),
    .Y(_00382_),
    .B1(net1387));
 sg13g2_nor2_1 _17704_ (.A(\fpga_top.io_uart_out.rout[0] ),
    .B(net5327),
    .Y(_03037_));
 sg13g2_a21oi_1 _17705_ (.A1(_06866_),
    .A2(net5327),
    .Y(_00383_),
    .B1(_03037_));
 sg13g2_mux2_1 _17706_ (.A0(\fpga_top.io_uart_out.rout[1] ),
    .A1(net3883),
    .S(net5327),
    .X(_00384_));
 sg13g2_mux2_1 _17707_ (.A0(net2852),
    .A1(net3809),
    .S(net5327),
    .X(_00385_));
 sg13g2_mux2_1 _17708_ (.A0(\fpga_top.io_uart_out.rout[3] ),
    .A1(net3815),
    .S(net5327),
    .X(_00386_));
 sg13g2_mux2_1 _17709_ (.A0(net3623),
    .A1(net3925),
    .S(net5328),
    .X(_00387_));
 sg13g2_mux2_1 _17710_ (.A0(\fpga_top.io_uart_out.rout[5] ),
    .A1(net3735),
    .S(net5327),
    .X(_00388_));
 sg13g2_mux2_1 _17711_ (.A0(\fpga_top.io_uart_out.rout[6] ),
    .A1(net3595),
    .S(net5327),
    .X(_00389_));
 sg13g2_nor2_1 _17712_ (.A(\fpga_top.io_uart_out.rout[7] ),
    .B(net5328),
    .Y(_03038_));
 sg13g2_a21oi_1 _17713_ (.A1(_06895_),
    .A2(net5328),
    .Y(_00390_),
    .B1(_03038_));
 sg13g2_or2_1 _17714_ (.X(_03039_),
    .B(_08616_),
    .A(_06769_));
 sg13g2_a221oi_1 _17715_ (.B2(net3681),
    .C1(net4012),
    .B1(_08681_),
    .A1(net3807),
    .Y(_03040_),
    .A2(_08618_));
 sg13g2_a21oi_1 _17716_ (.A1(_03039_),
    .A2(_03040_),
    .Y(_00391_),
    .B1(\fpga_top.cpu_start ));
 sg13g2_nor3_2 _17717_ (.A(_08902_),
    .B(_09617_),
    .C(_10518_),
    .Y(_03041_));
 sg13g2_nor2_1 _17718_ (.A(net6305),
    .B(_03041_),
    .Y(_03042_));
 sg13g2_a21oi_1 _17719_ (.A1(net4921),
    .A2(_03041_),
    .Y(_00392_),
    .B1(_03042_));
 sg13g2_nor2_1 _17720_ (.A(net6302),
    .B(_03041_),
    .Y(_03043_));
 sg13g2_a21oi_1 _17721_ (.A1(net4918),
    .A2(_03041_),
    .Y(_00393_),
    .B1(_03043_));
 sg13g2_nor2_1 _17722_ (.A(net6325),
    .B(_03041_),
    .Y(_03044_));
 sg13g2_a21oi_1 _17723_ (.A1(net4851),
    .A2(_03041_),
    .Y(_00394_),
    .B1(_03044_));
 sg13g2_mux2_1 _17724_ (.A0(net6411),
    .A1(net4842),
    .S(_03041_),
    .X(_00395_));
 sg13g2_nand2_2 _17725_ (.Y(_03045_),
    .A(_08909_),
    .B(_02734_));
 sg13g2_nor2_1 _17726_ (.A(net4560),
    .B(_03045_),
    .Y(_03046_));
 sg13g2_o21ai_1 _17727_ (.B1(\fpga_top.io_frc.frc_cntrl_val ),
    .Y(_03047_),
    .A1(net4560),
    .A2(_03045_));
 sg13g2_nor2_1 _17728_ (.A(net4560),
    .B(_09615_),
    .Y(_03048_));
 sg13g2_inv_1 _17729_ (.Y(_03049_),
    .A(net4503));
 sg13g2_a21oi_2 _17730_ (.B1(net4503),
    .Y(_03050_),
    .A2(net4845),
    .A1(_08912_));
 sg13g2_and2_1 _17731_ (.A(_03047_),
    .B(_03050_),
    .X(_03051_));
 sg13g2_nand2_1 _17732_ (.Y(_03052_),
    .A(_03047_),
    .B(_03050_));
 sg13g2_nor2b_1 _17733_ (.A(net4512),
    .B_N(_03050_),
    .Y(_03053_));
 sg13g2_nand2b_1 _17734_ (.Y(_03054_),
    .B(_03050_),
    .A_N(net4512));
 sg13g2_a221oi_1 _17735_ (.B2(_06685_),
    .C1(net4449),
    .B1(net4442),
    .A1(_10526_),
    .Y(_03055_),
    .A2(net4501));
 sg13g2_a21oi_1 _17736_ (.A1(_06685_),
    .A2(net4449),
    .Y(_00396_),
    .B1(_03055_));
 sg13g2_xor2_1 _17737_ (.B(net6335),
    .A(net6143),
    .X(_03056_));
 sg13g2_a221oi_1 _17738_ (.B2(_03056_),
    .C1(net4449),
    .B1(net4442),
    .A1(net4846),
    .Y(_03057_),
    .A2(net4501));
 sg13g2_a21oi_1 _17739_ (.A1(_06686_),
    .A2(net4449),
    .Y(_00397_),
    .B1(_03057_));
 sg13g2_nand3_1 _17740_ (.B(net6612),
    .C(net3930),
    .A(net6143),
    .Y(_03058_));
 sg13g2_o21ai_1 _17741_ (.B1(_06689_),
    .Y(_03059_),
    .A1(_06685_),
    .A2(_06686_));
 sg13g2_and2_1 _17742_ (.A(_03058_),
    .B(_03059_),
    .X(_03060_));
 sg13g2_a221oi_1 _17743_ (.B2(_03060_),
    .C1(net4451),
    .B1(net4442),
    .A1(_08915_),
    .Y(_03061_),
    .A2(net4501));
 sg13g2_a21oi_1 _17744_ (.A1(_06689_),
    .A2(net4449),
    .Y(_00398_),
    .B1(_03061_));
 sg13g2_nand4_1 _17745_ (.B(\fpga_top.io_frc.frc_cntr_val[1] ),
    .C(\fpga_top.io_frc.frc_cntr_val[3] ),
    .A(net6143),
    .Y(_03062_),
    .D(net3930));
 sg13g2_xnor2_1 _17746_ (.Y(_03063_),
    .A(net6179),
    .B(_03058_));
 sg13g2_a221oi_1 _17747_ (.B2(_03063_),
    .C1(net4449),
    .B1(net4442),
    .A1(net4843),
    .Y(_03064_),
    .A2(net4501));
 sg13g2_a21oi_1 _17748_ (.A1(_06687_),
    .A2(net4449),
    .Y(_00399_),
    .B1(_03064_));
 sg13g2_nor2_2 _17749_ (.A(_06695_),
    .B(_03062_),
    .Y(_03065_));
 sg13g2_xnor2_1 _17750_ (.Y(_03066_),
    .A(net6321),
    .B(_03062_));
 sg13g2_a221oi_1 _17751_ (.B2(_03066_),
    .C1(net4449),
    .B1(net4442),
    .A1(net4839),
    .Y(_03067_),
    .A2(net4501));
 sg13g2_a21oi_1 _17752_ (.A1(_06695_),
    .A2(net4450),
    .Y(_00400_),
    .B1(_03067_));
 sg13g2_xnor2_1 _17753_ (.Y(_03068_),
    .A(_06693_),
    .B(_03065_));
 sg13g2_a221oi_1 _17754_ (.B2(_03068_),
    .C1(net4450),
    .B1(net4442),
    .A1(net4834),
    .Y(_03069_),
    .A2(net4501));
 sg13g2_a21oi_1 _17755_ (.A1(_06693_),
    .A2(net4450),
    .Y(_00401_),
    .B1(_03069_));
 sg13g2_nand3_1 _17756_ (.B(\fpga_top.io_frc.frc_cntr_val[5] ),
    .C(_03065_),
    .A(net4061),
    .Y(_03070_));
 sg13g2_a21o_1 _17757_ (.A2(_03065_),
    .A1(\fpga_top.io_frc.frc_cntr_val[5] ),
    .B1(net4061),
    .X(_03071_));
 sg13g2_and2_1 _17758_ (.A(_03070_),
    .B(_03071_),
    .X(_03072_));
 sg13g2_a22oi_1 _17759_ (.Y(_03073_),
    .B1(net4442),
    .B2(_03072_),
    .A2(net4501),
    .A1(_02756_));
 sg13g2_nor2_1 _17760_ (.A(net4061),
    .B(net4447),
    .Y(_03074_));
 sg13g2_a21oi_1 _17761_ (.A1(net4447),
    .A2(_03073_),
    .Y(_00402_),
    .B1(_03074_));
 sg13g2_and4_1 _17762_ (.A(\fpga_top.io_frc.frc_cntr_val[7] ),
    .B(\fpga_top.io_frc.frc_cntr_val[6] ),
    .C(\fpga_top.io_frc.frc_cntr_val[5] ),
    .D(_03065_),
    .X(_03075_));
 sg13g2_xnor2_1 _17763_ (.Y(_03076_),
    .A(net6197),
    .B(_03070_));
 sg13g2_a221oi_1 _17764_ (.B2(_03076_),
    .C1(net4451),
    .B1(net4442),
    .A1(_02760_),
    .Y(_03077_),
    .A2(net4501));
 sg13g2_a21oi_1 _17765_ (.A1(_06690_),
    .A2(net4451),
    .Y(_00403_),
    .B1(_03077_));
 sg13g2_xnor2_1 _17766_ (.Y(_03078_),
    .A(_06710_),
    .B(_03075_));
 sg13g2_a221oi_1 _17767_ (.B2(_03078_),
    .C1(net4453),
    .B1(net4443),
    .A1(_02764_),
    .Y(_03079_),
    .A2(net4502));
 sg13g2_a21oi_1 _17768_ (.A1(_06710_),
    .A2(net4453),
    .Y(_00404_),
    .B1(_03079_));
 sg13g2_nand3_1 _17769_ (.B(\fpga_top.io_frc.frc_cntr_val[8] ),
    .C(_03075_),
    .A(net4028),
    .Y(_03080_));
 sg13g2_a21o_1 _17770_ (.A2(_03075_),
    .A1(\fpga_top.io_frc.frc_cntr_val[8] ),
    .B1(net4028),
    .X(_03081_));
 sg13g2_and2_1 _17771_ (.A(_03080_),
    .B(_03081_),
    .X(_03082_));
 sg13g2_a221oi_1 _17772_ (.B2(_03082_),
    .C1(net4453),
    .B1(net4443),
    .A1(_02768_),
    .Y(_03083_),
    .A2(net4502));
 sg13g2_a21oi_1 _17773_ (.A1(_06708_),
    .A2(net4453),
    .Y(_00405_),
    .B1(_03083_));
 sg13g2_and4_1 _17774_ (.A(\fpga_top.io_frc.frc_cntr_val[10] ),
    .B(\fpga_top.io_frc.frc_cntr_val[9] ),
    .C(\fpga_top.io_frc.frc_cntr_val[8] ),
    .D(_03075_),
    .X(_03084_));
 sg13g2_xnor2_1 _17775_ (.Y(_03085_),
    .A(net4016),
    .B(_03080_));
 sg13g2_a221oi_1 _17776_ (.B2(_03085_),
    .C1(net4453),
    .B1(net4443),
    .A1(_08981_),
    .Y(_03086_),
    .A2(net4502));
 sg13g2_a21oi_1 _17777_ (.A1(_06706_),
    .A2(net4453),
    .Y(_00406_),
    .B1(_03086_));
 sg13g2_xor2_1 _17778_ (.B(_03084_),
    .A(net4052),
    .X(_03087_));
 sg13g2_nor2_1 _17779_ (.A(_02771_),
    .B(net4467),
    .Y(_03088_));
 sg13g2_a21oi_1 _17780_ (.A1(net4443),
    .A2(_03087_),
    .Y(_03089_),
    .B1(_03088_));
 sg13g2_nor2_1 _17781_ (.A(net4052),
    .B(net4448),
    .Y(_03090_));
 sg13g2_a21oi_1 _17782_ (.A1(net4448),
    .A2(_03089_),
    .Y(_00407_),
    .B1(_03090_));
 sg13g2_nand3_1 _17783_ (.B(\fpga_top.io_frc.frc_cntr_val[11] ),
    .C(_03084_),
    .A(\fpga_top.io_frc.frc_cntr_val[12] ),
    .Y(_03091_));
 sg13g2_a21o_1 _17784_ (.A2(_03084_),
    .A1(\fpga_top.io_frc.frc_cntr_val[11] ),
    .B1(net6250),
    .X(_03092_));
 sg13g2_and2_1 _17785_ (.A(_03091_),
    .B(_03092_),
    .X(_03093_));
 sg13g2_a221oi_1 _17786_ (.B2(_03093_),
    .C1(net4456),
    .B1(net4444),
    .A1(_02774_),
    .Y(_03094_),
    .A2(net4503));
 sg13g2_a21oi_1 _17787_ (.A1(_06703_),
    .A2(net4456),
    .Y(_00408_),
    .B1(_03094_));
 sg13g2_nor2_1 _17788_ (.A(_06701_),
    .B(_03091_),
    .Y(_03095_));
 sg13g2_xnor2_1 _17789_ (.Y(_03096_),
    .A(net3745),
    .B(_03091_));
 sg13g2_o21ai_1 _17790_ (.B1(net4448),
    .Y(_03097_),
    .A1(_02778_),
    .A2(net4467));
 sg13g2_a21oi_1 _17791_ (.A1(net4445),
    .A2(_03096_),
    .Y(_03098_),
    .B1(_03097_));
 sg13g2_a21oi_1 _17792_ (.A1(_06701_),
    .A2(net4457),
    .Y(_00409_),
    .B1(_03098_));
 sg13g2_xnor2_1 _17793_ (.Y(_03099_),
    .A(_06699_),
    .B(_03095_));
 sg13g2_a221oi_1 _17794_ (.B2(_03099_),
    .C1(net4456),
    .B1(net4445),
    .A1(_02782_),
    .Y(_03100_),
    .A2(net4503));
 sg13g2_a21oi_1 _17795_ (.A1(_06699_),
    .A2(net4457),
    .Y(_00410_),
    .B1(_03100_));
 sg13g2_nor4_2 _17796_ (.A(_06697_),
    .B(_06699_),
    .C(_06701_),
    .Y(_03101_),
    .D(_03091_));
 sg13g2_a21oi_1 _17797_ (.A1(\fpga_top.io_frc.frc_cntr_val[14] ),
    .A2(_03095_),
    .Y(_03102_),
    .B1(net3902));
 sg13g2_nor3_1 _17798_ (.A(_03054_),
    .B(_03101_),
    .C(_03102_),
    .Y(_03103_));
 sg13g2_nor2_1 _17799_ (.A(_02784_),
    .B(net4467),
    .Y(_03104_));
 sg13g2_nor3_1 _17800_ (.A(net4456),
    .B(_03103_),
    .C(_03104_),
    .Y(_03105_));
 sg13g2_a21oi_1 _17801_ (.A1(_06697_),
    .A2(net4456),
    .Y(_00411_),
    .B1(_03105_));
 sg13g2_and2_1 _17802_ (.A(net4039),
    .B(_03101_),
    .X(_03106_));
 sg13g2_xnor2_1 _17803_ (.Y(_03107_),
    .A(_06730_),
    .B(_03101_));
 sg13g2_a221oi_1 _17804_ (.B2(_03107_),
    .C1(net4454),
    .B1(net4443),
    .A1(_10594_),
    .Y(_03108_),
    .A2(net4502));
 sg13g2_a21oi_1 _17805_ (.A1(_06730_),
    .A2(net4457),
    .Y(_00412_),
    .B1(_03108_));
 sg13g2_xnor2_1 _17806_ (.Y(_03109_),
    .A(_06729_),
    .B(_03106_));
 sg13g2_a221oi_1 _17807_ (.B2(_03109_),
    .C1(net4454),
    .B1(net4443),
    .A1(_10599_),
    .Y(_03110_),
    .A2(net4502));
 sg13g2_a21oi_1 _17808_ (.A1(_06729_),
    .A2(net4454),
    .Y(_00413_),
    .B1(_03110_));
 sg13g2_nand4_1 _17809_ (.B(\fpga_top.io_frc.frc_cntr_val[16] ),
    .C(\fpga_top.io_frc.frc_cntr_val[18] ),
    .A(\fpga_top.io_frc.frc_cntr_val[17] ),
    .Y(_03111_),
    .D(_03101_));
 sg13g2_a21o_1 _17810_ (.A2(_03106_),
    .A1(\fpga_top.io_frc.frc_cntr_val[17] ),
    .B1(net3949),
    .X(_03112_));
 sg13g2_and2_1 _17811_ (.A(_03111_),
    .B(_03112_),
    .X(_03113_));
 sg13g2_nor2_1 _17812_ (.A(_10603_),
    .B(net4467),
    .Y(_03114_));
 sg13g2_a21oi_1 _17813_ (.A1(net4445),
    .A2(_03113_),
    .Y(_03115_),
    .B1(_03114_));
 sg13g2_nor2_1 _17814_ (.A(net3949),
    .B(net4447),
    .Y(_03116_));
 sg13g2_a21oi_1 _17815_ (.A1(net4448),
    .A2(_03115_),
    .Y(_00414_),
    .B1(_03116_));
 sg13g2_nor2_1 _17816_ (.A(_06731_),
    .B(_03111_),
    .Y(_03117_));
 sg13g2_xnor2_1 _17817_ (.Y(_03118_),
    .A(net3803),
    .B(_03111_));
 sg13g2_o21ai_1 _17818_ (.B1(net4448),
    .Y(_03119_),
    .A1(_02789_),
    .A2(net4467));
 sg13g2_a21oi_1 _17819_ (.A1(net4443),
    .A2(_03118_),
    .Y(_03120_),
    .B1(_03119_));
 sg13g2_a21oi_1 _17820_ (.A1(_06731_),
    .A2(net4453),
    .Y(_00415_),
    .B1(_03120_));
 sg13g2_xnor2_1 _17821_ (.Y(_03121_),
    .A(_06728_),
    .B(_03117_));
 sg13g2_a221oi_1 _17822_ (.B2(_03121_),
    .C1(net4454),
    .B1(net4445),
    .A1(_10606_),
    .Y(_03122_),
    .A2(net4502));
 sg13g2_a21oi_1 _17823_ (.A1(_06728_),
    .A2(net4454),
    .Y(_00416_),
    .B1(_03122_));
 sg13g2_nor4_2 _17824_ (.A(_06726_),
    .B(_06728_),
    .C(_06731_),
    .Y(_03123_),
    .D(_03111_));
 sg13g2_a21oi_1 _17825_ (.A1(net3756),
    .A2(_03117_),
    .Y(_03124_),
    .B1(net3824));
 sg13g2_nor2_1 _17826_ (.A(_03123_),
    .B(_03124_),
    .Y(_03125_));
 sg13g2_o21ai_1 _17827_ (.B1(net4448),
    .Y(_03126_),
    .A1(_10609_),
    .A2(net4467));
 sg13g2_a21oi_1 _17828_ (.A1(net4445),
    .A2(_03125_),
    .Y(_03127_),
    .B1(_03126_));
 sg13g2_a21oi_1 _17829_ (.A1(_06726_),
    .A2(net4454),
    .Y(_00417_),
    .B1(_03127_));
 sg13g2_and2_1 _17830_ (.A(net4072),
    .B(_03123_),
    .X(_03128_));
 sg13g2_xnor2_1 _17831_ (.Y(_03129_),
    .A(_06724_),
    .B(_03123_));
 sg13g2_a221oi_1 _17832_ (.B2(_03129_),
    .C1(net4453),
    .B1(net4443),
    .A1(_10612_),
    .Y(_03130_),
    .A2(net4502));
 sg13g2_a21oi_1 _17833_ (.A1(_06724_),
    .A2(net4454),
    .Y(_00418_),
    .B1(_03130_));
 sg13g2_xnor2_1 _17834_ (.Y(_03131_),
    .A(_06723_),
    .B(_03128_));
 sg13g2_o21ai_1 _17835_ (.B1(net4447),
    .Y(_03132_),
    .A1(_02795_),
    .A2(net4468));
 sg13g2_a21oi_1 _17836_ (.A1(net4444),
    .A2(_03131_),
    .Y(_03133_),
    .B1(_03132_));
 sg13g2_a21oi_1 _17837_ (.A1(_06723_),
    .A2(net4456),
    .Y(_00419_),
    .B1(_03133_));
 sg13g2_nand4_1 _17838_ (.B(\fpga_top.io_frc.frc_cntr_val[23] ),
    .C(\fpga_top.io_frc.frc_cntr_val[22] ),
    .A(\fpga_top.io_frc.frc_cntr_val[24] ),
    .Y(_03134_),
    .D(_03123_));
 sg13g2_a21o_1 _17839_ (.A2(_03128_),
    .A1(\fpga_top.io_frc.frc_cntr_val[23] ),
    .B1(net4005),
    .X(_03135_));
 sg13g2_and2_1 _17840_ (.A(_03134_),
    .B(_03135_),
    .X(_03136_));
 sg13g2_o21ai_1 _17841_ (.B1(net4447),
    .Y(_03137_),
    .A1(_10615_),
    .A2(net4468));
 sg13g2_a21oi_1 _17842_ (.A1(net4444),
    .A2(_03136_),
    .Y(_03138_),
    .B1(_03137_));
 sg13g2_a21oi_1 _17843_ (.A1(_06721_),
    .A2(net4455),
    .Y(_00420_),
    .B1(_03138_));
 sg13g2_nor2_2 _17844_ (.A(_06719_),
    .B(_03134_),
    .Y(_03139_));
 sg13g2_xnor2_1 _17845_ (.Y(_03140_),
    .A(net6181),
    .B(_03134_));
 sg13g2_a221oi_1 _17846_ (.B2(_03140_),
    .C1(net4455),
    .B1(net4444),
    .A1(_10619_),
    .Y(_03141_),
    .A2(net4502));
 sg13g2_a21oi_1 _17847_ (.A1(_06719_),
    .A2(net4455),
    .Y(_00421_),
    .B1(_03141_));
 sg13g2_xnor2_1 _17848_ (.Y(_03142_),
    .A(_06718_),
    .B(_03139_));
 sg13g2_o21ai_1 _17849_ (.B1(net4447),
    .Y(_03143_),
    .A1(_10622_),
    .A2(net4467));
 sg13g2_a21oi_1 _17850_ (.A1(net4444),
    .A2(_03142_),
    .Y(_03144_),
    .B1(_03143_));
 sg13g2_a21oi_1 _17851_ (.A1(_06718_),
    .A2(net4455),
    .Y(_00422_),
    .B1(_03144_));
 sg13g2_nand3_1 _17852_ (.B(net4040),
    .C(_03139_),
    .A(net3862),
    .Y(_03145_));
 sg13g2_a21o_1 _17853_ (.A2(_03139_),
    .A1(\fpga_top.io_frc.frc_cntr_val[26] ),
    .B1(net3862),
    .X(_03146_));
 sg13g2_and2_1 _17854_ (.A(_03145_),
    .B(_03146_),
    .X(_03147_));
 sg13g2_a221oi_1 _17855_ (.B2(_03147_),
    .C1(net4455),
    .B1(net4444),
    .A1(_02802_),
    .Y(_03148_),
    .A2(net4503));
 sg13g2_a21oi_1 _17856_ (.A1(_06717_),
    .A2(net4456),
    .Y(_00423_),
    .B1(_03148_));
 sg13g2_and4_1 _17857_ (.A(\fpga_top.io_frc.frc_cntr_val[28] ),
    .B(\fpga_top.io_frc.frc_cntr_val[27] ),
    .C(\fpga_top.io_frc.frc_cntr_val[26] ),
    .D(_03139_),
    .X(_03149_));
 sg13g2_xnor2_1 _17858_ (.Y(_03150_),
    .A(net6347),
    .B(_03145_));
 sg13g2_o21ai_1 _17859_ (.B1(net4447),
    .Y(_03151_),
    .A1(_02805_),
    .A2(net4467));
 sg13g2_a21oi_1 _17860_ (.A1(net4444),
    .A2(_03150_),
    .Y(_03152_),
    .B1(_03151_));
 sg13g2_a21oi_1 _17861_ (.A1(_06715_),
    .A2(net4455),
    .Y(_00424_),
    .B1(_03152_));
 sg13g2_xnor2_1 _17862_ (.Y(_03153_),
    .A(_06714_),
    .B(_03149_));
 sg13g2_a221oi_1 _17863_ (.B2(_03153_),
    .C1(net4455),
    .B1(net4444),
    .A1(_02808_),
    .Y(_03154_),
    .A2(net4503));
 sg13g2_a21oi_1 _17864_ (.A1(_06714_),
    .A2(net4455),
    .Y(_00425_),
    .B1(_03154_));
 sg13g2_nand3_1 _17865_ (.B(\fpga_top.io_frc.frc_cntr_val[29] ),
    .C(_03149_),
    .A(net4055),
    .Y(_03155_));
 sg13g2_a21o_1 _17866_ (.A2(_03149_),
    .A1(net6610),
    .B1(net4055),
    .X(_03156_));
 sg13g2_and2_1 _17867_ (.A(_03155_),
    .B(_03156_),
    .X(_03157_));
 sg13g2_a221oi_1 _17868_ (.B2(_03157_),
    .C1(net4452),
    .B1(net4446),
    .A1(_02813_),
    .Y(_03158_),
    .A2(net4504));
 sg13g2_a21oi_1 _17869_ (.A1(_06713_),
    .A2(net4452),
    .Y(_00426_),
    .B1(_03158_));
 sg13g2_nor2_1 _17870_ (.A(_06712_),
    .B(_03155_),
    .Y(_03159_));
 sg13g2_xnor2_1 _17871_ (.Y(_03160_),
    .A(net6086),
    .B(_03155_));
 sg13g2_o21ai_1 _17872_ (.B1(net4447),
    .Y(_03161_),
    .A1(_02817_),
    .A2(net4468));
 sg13g2_a21oi_1 _17873_ (.A1(net4446),
    .A2(_03160_),
    .Y(_03162_),
    .B1(_03161_));
 sg13g2_a21oi_1 _17874_ (.A1(_06712_),
    .A2(net4452),
    .Y(_00427_),
    .B1(_03162_));
 sg13g2_nand2_1 _17875_ (.Y(_03163_),
    .A(_08978_),
    .B(_10552_));
 sg13g2_nor3_2 _17876_ (.A(_08902_),
    .B(_10522_),
    .C(_03163_),
    .Y(_03164_));
 sg13g2_nor2_1 _17877_ (.A(net6373),
    .B(_03164_),
    .Y(_03165_));
 sg13g2_a21oi_1 _17878_ (.A1(net4921),
    .A2(_03164_),
    .Y(_00428_),
    .B1(_03165_));
 sg13g2_nor2_1 _17879_ (.A(net6313),
    .B(_03164_),
    .Y(_03166_));
 sg13g2_a21oi_1 _17880_ (.A1(net4918),
    .A2(_03164_),
    .Y(_00429_),
    .B1(_03166_));
 sg13g2_nor2_1 _17881_ (.A(net6360),
    .B(_03164_),
    .Y(_03167_));
 sg13g2_a21oi_1 _17882_ (.A1(net4851),
    .A2(_03164_),
    .Y(_00430_),
    .B1(_03167_));
 sg13g2_mux2_1 _17883_ (.A0(net6418),
    .A1(net4842),
    .S(_03164_),
    .X(_00431_));
 sg13g2_nand3_1 _17884_ (.B(_09664_),
    .C(_09667_),
    .A(_09661_),
    .Y(_03168_));
 sg13g2_nand2_2 _17885_ (.Y(_03169_),
    .A(_09655_),
    .B(_09657_));
 sg13g2_or2_1 _17886_ (.X(_03170_),
    .B(_03169_),
    .A(_03168_));
 sg13g2_mux2_1 _17887_ (.A0(net4361),
    .A1(net2421),
    .S(net4170),
    .X(_00432_));
 sg13g2_mux2_1 _17888_ (.A0(net4357),
    .A1(net2880),
    .S(net4172),
    .X(_00433_));
 sg13g2_mux2_1 _17889_ (.A0(net4350),
    .A1(net2826),
    .S(net4171),
    .X(_00434_));
 sg13g2_mux2_1 _17890_ (.A0(net4346),
    .A1(net3145),
    .S(net4170),
    .X(_00435_));
 sg13g2_mux2_1 _17891_ (.A0(net4340),
    .A1(net3516),
    .S(net4172),
    .X(_00436_));
 sg13g2_mux2_1 _17892_ (.A0(net4196),
    .A1(net2496),
    .S(net4172),
    .X(_00437_));
 sg13g2_mux2_1 _17893_ (.A0(net4334),
    .A1(net3553),
    .S(net4171),
    .X(_00438_));
 sg13g2_mux2_1 _17894_ (.A0(net4330),
    .A1(net3183),
    .S(net4174),
    .X(_00439_));
 sg13g2_mux2_1 _17895_ (.A0(net4325),
    .A1(net2654),
    .S(net4172),
    .X(_00440_));
 sg13g2_mux2_1 _17896_ (.A0(net4320),
    .A1(net2912),
    .S(net4171),
    .X(_00441_));
 sg13g2_mux2_1 _17897_ (.A0(net4191),
    .A1(net3076),
    .S(net4173),
    .X(_00442_));
 sg13g2_mux2_1 _17898_ (.A0(net4185),
    .A1(net2528),
    .S(net4170),
    .X(_00443_));
 sg13g2_mux2_1 _17899_ (.A0(net4313),
    .A1(net3013),
    .S(net4173),
    .X(_00444_));
 sg13g2_mux2_1 _17900_ (.A0(net4307),
    .A1(net3460),
    .S(net4170),
    .X(_00445_));
 sg13g2_mux2_1 _17901_ (.A0(net4302),
    .A1(net3650),
    .S(net4170),
    .X(_00446_));
 sg13g2_mux2_1 _17902_ (.A0(net4297),
    .A1(net3371),
    .S(net4174),
    .X(_00447_));
 sg13g2_mux2_1 _17903_ (.A0(net4291),
    .A1(net3532),
    .S(net4173),
    .X(_00448_));
 sg13g2_mux2_1 _17904_ (.A0(net4286),
    .A1(net2424),
    .S(net4170),
    .X(_00449_));
 sg13g2_mux2_1 _17905_ (.A0(net4280),
    .A1(net3127),
    .S(net4173),
    .X(_00450_));
 sg13g2_mux2_1 _17906_ (.A0(net4276),
    .A1(net2773),
    .S(net4172),
    .X(_00451_));
 sg13g2_mux2_1 _17907_ (.A0(net4269),
    .A1(net3164),
    .S(net4172),
    .X(_00452_));
 sg13g2_mux2_1 _17908_ (.A0(net4264),
    .A1(net2717),
    .S(net4170),
    .X(_00453_));
 sg13g2_mux2_1 _17909_ (.A0(net4261),
    .A1(net3057),
    .S(net4174),
    .X(_00454_));
 sg13g2_mux2_1 _17910_ (.A0(net4254),
    .A1(net3150),
    .S(net4173),
    .X(_00455_));
 sg13g2_mux2_1 _17911_ (.A0(net4404),
    .A1(net3068),
    .S(net4173),
    .X(_00456_));
 sg13g2_mux2_1 _17912_ (.A0(net4399),
    .A1(net3409),
    .S(net4172),
    .X(_00457_));
 sg13g2_mux2_1 _17913_ (.A0(net4393),
    .A1(net3366),
    .S(net4171),
    .X(_00458_));
 sg13g2_mux2_1 _17914_ (.A0(net4392),
    .A1(net2402),
    .S(net4170),
    .X(_00459_));
 sg13g2_mux2_1 _17915_ (.A0(net4385),
    .A1(net3365),
    .S(net4171),
    .X(_00460_));
 sg13g2_mux2_1 _17916_ (.A0(net4378),
    .A1(net2879),
    .S(net4173),
    .X(_00461_));
 sg13g2_mux2_1 _17917_ (.A0(net4376),
    .A1(net2309),
    .S(net4172),
    .X(_00462_));
 sg13g2_mux2_1 _17918_ (.A0(net4367),
    .A1(net3231),
    .S(net4173),
    .X(_00463_));
 sg13g2_or2_1 _17919_ (.X(_03171_),
    .B(_03168_),
    .A(_09805_));
 sg13g2_mux2_1 _17920_ (.A0(net4361),
    .A1(net2845),
    .S(net4165),
    .X(_00464_));
 sg13g2_mux2_1 _17921_ (.A0(net4357),
    .A1(net3578),
    .S(net4167),
    .X(_00465_));
 sg13g2_mux2_1 _17922_ (.A0(net4350),
    .A1(net2914),
    .S(net4166),
    .X(_00466_));
 sg13g2_mux2_1 _17923_ (.A0(net4346),
    .A1(net2771),
    .S(net4165),
    .X(_00467_));
 sg13g2_mux2_1 _17924_ (.A0(net4340),
    .A1(net3462),
    .S(net4167),
    .X(_00468_));
 sg13g2_mux2_1 _17925_ (.A0(net4196),
    .A1(net2334),
    .S(net4167),
    .X(_00469_));
 sg13g2_mux2_1 _17926_ (.A0(net4334),
    .A1(net2519),
    .S(net4166),
    .X(_00470_));
 sg13g2_mux2_1 _17927_ (.A0(net4329),
    .A1(net2788),
    .S(net4169),
    .X(_00471_));
 sg13g2_mux2_1 _17928_ (.A0(net4325),
    .A1(net2557),
    .S(net4167),
    .X(_00472_));
 sg13g2_mux2_1 _17929_ (.A0(net4320),
    .A1(net2518),
    .S(net4166),
    .X(_00473_));
 sg13g2_mux2_1 _17930_ (.A0(net4191),
    .A1(net2677),
    .S(net4168),
    .X(_00474_));
 sg13g2_mux2_1 _17931_ (.A0(net4185),
    .A1(net3086),
    .S(net4165),
    .X(_00475_));
 sg13g2_mux2_1 _17932_ (.A0(net4312),
    .A1(net3049),
    .S(net4168),
    .X(_00476_));
 sg13g2_mux2_1 _17933_ (.A0(net4307),
    .A1(net3456),
    .S(net4165),
    .X(_00477_));
 sg13g2_mux2_1 _17934_ (.A0(net4302),
    .A1(net2672),
    .S(net4165),
    .X(_00478_));
 sg13g2_mux2_1 _17935_ (.A0(net4297),
    .A1(net3066),
    .S(net4169),
    .X(_00479_));
 sg13g2_mux2_1 _17936_ (.A0(net4291),
    .A1(net3588),
    .S(net4168),
    .X(_00480_));
 sg13g2_mux2_1 _17937_ (.A0(net4286),
    .A1(net2743),
    .S(net4165),
    .X(_00481_));
 sg13g2_mux2_1 _17938_ (.A0(net4280),
    .A1(net3535),
    .S(net4168),
    .X(_00482_));
 sg13g2_mux2_1 _17939_ (.A0(net4276),
    .A1(net3159),
    .S(net4167),
    .X(_00483_));
 sg13g2_mux2_1 _17940_ (.A0(net4269),
    .A1(net2240),
    .S(net4167),
    .X(_00484_));
 sg13g2_mux2_1 _17941_ (.A0(net4264),
    .A1(net2593),
    .S(net4165),
    .X(_00485_));
 sg13g2_mux2_1 _17942_ (.A0(net4261),
    .A1(net3376),
    .S(net4169),
    .X(_00486_));
 sg13g2_mux2_1 _17943_ (.A0(net4254),
    .A1(net2341),
    .S(net4168),
    .X(_00487_));
 sg13g2_mux2_1 _17944_ (.A0(net4404),
    .A1(net3103),
    .S(net4168),
    .X(_00488_));
 sg13g2_mux2_1 _17945_ (.A0(net4399),
    .A1(net2897),
    .S(net4167),
    .X(_00489_));
 sg13g2_mux2_1 _17946_ (.A0(net4393),
    .A1(net2745),
    .S(net4166),
    .X(_00490_));
 sg13g2_mux2_1 _17947_ (.A0(net4389),
    .A1(net3069),
    .S(net4165),
    .X(_00491_));
 sg13g2_mux2_1 _17948_ (.A0(net4384),
    .A1(net2355),
    .S(net4166),
    .X(_00492_));
 sg13g2_mux2_1 _17949_ (.A0(net4381),
    .A1(net3457),
    .S(net4168),
    .X(_00493_));
 sg13g2_mux2_1 _17950_ (.A0(net4373),
    .A1(net2868),
    .S(net4167),
    .X(_00494_));
 sg13g2_mux2_1 _17951_ (.A0(net4367),
    .A1(net3078),
    .S(net4168),
    .X(_00495_));
 sg13g2_or2_1 _17952_ (.X(_03172_),
    .B(_03168_),
    .A(_09659_));
 sg13g2_mux2_1 _17953_ (.A0(net4361),
    .A1(net2523),
    .S(net4160),
    .X(_00496_));
 sg13g2_mux2_1 _17954_ (.A0(net4357),
    .A1(net3223),
    .S(net4162),
    .X(_00497_));
 sg13g2_mux2_1 _17955_ (.A0(net4350),
    .A1(net2491),
    .S(net4161),
    .X(_00498_));
 sg13g2_mux2_1 _17956_ (.A0(net4346),
    .A1(net2922),
    .S(net4160),
    .X(_00499_));
 sg13g2_mux2_1 _17957_ (.A0(net4340),
    .A1(net2839),
    .S(net4162),
    .X(_00500_));
 sg13g2_mux2_1 _17958_ (.A0(net4196),
    .A1(net2465),
    .S(net4162),
    .X(_00501_));
 sg13g2_mux2_1 _17959_ (.A0(net4334),
    .A1(net2787),
    .S(net4161),
    .X(_00502_));
 sg13g2_mux2_1 _17960_ (.A0(net4329),
    .A1(net2608),
    .S(net4164),
    .X(_00503_));
 sg13g2_mux2_1 _17961_ (.A0(net4325),
    .A1(net2874),
    .S(net4162),
    .X(_00504_));
 sg13g2_mux2_1 _17962_ (.A0(net4320),
    .A1(net3568),
    .S(net4161),
    .X(_00505_));
 sg13g2_mux2_1 _17963_ (.A0(net4191),
    .A1(net2621),
    .S(net4163),
    .X(_00506_));
 sg13g2_mux2_1 _17964_ (.A0(net4185),
    .A1(net2565),
    .S(net4160),
    .X(_00507_));
 sg13g2_mux2_1 _17965_ (.A0(net4312),
    .A1(net2643),
    .S(net4163),
    .X(_00508_));
 sg13g2_mux2_1 _17966_ (.A0(net4307),
    .A1(net2544),
    .S(net4160),
    .X(_00509_));
 sg13g2_mux2_1 _17967_ (.A0(net4302),
    .A1(net2461),
    .S(net4160),
    .X(_00510_));
 sg13g2_mux2_1 _17968_ (.A0(net4297),
    .A1(net3214),
    .S(net4164),
    .X(_00511_));
 sg13g2_mux2_1 _17969_ (.A0(net4291),
    .A1(net2571),
    .S(net4163),
    .X(_00512_));
 sg13g2_mux2_1 _17970_ (.A0(net4286),
    .A1(net3569),
    .S(net4160),
    .X(_00513_));
 sg13g2_mux2_1 _17971_ (.A0(net4280),
    .A1(net3035),
    .S(net4163),
    .X(_00514_));
 sg13g2_mux2_1 _17972_ (.A0(net4276),
    .A1(net2690),
    .S(net4162),
    .X(_00515_));
 sg13g2_mux2_1 _17973_ (.A0(net4269),
    .A1(net3377),
    .S(net4162),
    .X(_00516_));
 sg13g2_mux2_1 _17974_ (.A0(net4264),
    .A1(net2598),
    .S(net4160),
    .X(_00517_));
 sg13g2_mux2_1 _17975_ (.A0(net4261),
    .A1(net2701),
    .S(net4164),
    .X(_00518_));
 sg13g2_mux2_1 _17976_ (.A0(net4254),
    .A1(net2738),
    .S(net4163),
    .X(_00519_));
 sg13g2_mux2_1 _17977_ (.A0(net4404),
    .A1(net2383),
    .S(net4163),
    .X(_00520_));
 sg13g2_mux2_1 _17978_ (.A0(net4399),
    .A1(net2382),
    .S(net4162),
    .X(_00521_));
 sg13g2_mux2_1 _17979_ (.A0(net4393),
    .A1(net2540),
    .S(net4161),
    .X(_00522_));
 sg13g2_mux2_1 _17980_ (.A0(net4389),
    .A1(net3058),
    .S(net4160),
    .X(_00523_));
 sg13g2_mux2_1 _17981_ (.A0(net4385),
    .A1(net2816),
    .S(net4161),
    .X(_00524_));
 sg13g2_mux2_1 _17982_ (.A0(net4378),
    .A1(net2907),
    .S(net4163),
    .X(_00525_));
 sg13g2_mux2_1 _17983_ (.A0(net4373),
    .A1(net2258),
    .S(net4162),
    .X(_00526_));
 sg13g2_mux2_1 _17984_ (.A0(net4367),
    .A1(net2555),
    .S(net4163),
    .X(_00527_));
 sg13g2_or3_1 _17985_ (.A(net3898),
    .B(net5351),
    .C(_09101_),
    .X(_03173_));
 sg13g2_nand2_1 _17986_ (.Y(_03174_),
    .A(net3898),
    .B(net5353));
 sg13g2_xnor2_1 _17987_ (.Y(_03175_),
    .A(_06675_),
    .B(_03174_));
 sg13g2_nand2_1 _17988_ (.Y(_00528_),
    .A(_03173_),
    .B(_03175_));
 sg13g2_nand3_1 _17989_ (.B(net5353),
    .C(_08918_),
    .A(net3898),
    .Y(_03176_));
 sg13g2_o21ai_1 _17990_ (.B1(net6420),
    .Y(_03177_),
    .A1(\fpga_top.qspi_if.cmd_ofs[0] ),
    .A2(_03174_));
 sg13g2_nand3_1 _17991_ (.B(_03176_),
    .C(net6421),
    .A(_03173_),
    .Y(_00529_));
 sg13g2_xor2_1 _17992_ (.B(_03176_),
    .A(net6503),
    .X(_03178_));
 sg13g2_nand2_1 _17993_ (.Y(_00530_),
    .A(_03173_),
    .B(_03178_));
 sg13g2_and3_2 _17994_ (.X(_03179_),
    .A(_09661_),
    .B(_09664_),
    .C(_09666_));
 sg13g2_nand3_1 _17995_ (.B(_09657_),
    .C(_03179_),
    .A(_09655_),
    .Y(_03180_));
 sg13g2_mux2_1 _17996_ (.A0(net4362),
    .A1(net3210),
    .S(net4249),
    .X(_00531_));
 sg13g2_mux2_1 _17997_ (.A0(net4356),
    .A1(net2577),
    .S(net4251),
    .X(_00532_));
 sg13g2_mux2_1 _17998_ (.A0(net4349),
    .A1(net2895),
    .S(net4250),
    .X(_00533_));
 sg13g2_mux2_1 _17999_ (.A0(net4344),
    .A1(net2475),
    .S(net4249),
    .X(_00534_));
 sg13g2_mux2_1 _18000_ (.A0(net4339),
    .A1(net2262),
    .S(net4251),
    .X(_00535_));
 sg13g2_mux2_1 _18001_ (.A0(net4196),
    .A1(net3551),
    .S(net4251),
    .X(_00536_));
 sg13g2_mux2_1 _18002_ (.A0(net4335),
    .A1(net2568),
    .S(net4250),
    .X(_00537_));
 sg13g2_mux2_1 _18003_ (.A0(net4329),
    .A1(net3372),
    .S(net4252),
    .X(_00538_));
 sg13g2_mux2_1 _18004_ (.A0(net4324),
    .A1(net2827),
    .S(net4251),
    .X(_00539_));
 sg13g2_mux2_1 _18005_ (.A0(net4322),
    .A1(net2888),
    .S(net4250),
    .X(_00540_));
 sg13g2_mux2_1 _18006_ (.A0(net4190),
    .A1(net2674),
    .S(net4252),
    .X(_00541_));
 sg13g2_mux2_1 _18007_ (.A0(net4186),
    .A1(net3561),
    .S(net4249),
    .X(_00542_));
 sg13g2_mux2_1 _18008_ (.A0(net4312),
    .A1(net2522),
    .S(net4252),
    .X(_00543_));
 sg13g2_mux2_1 _18009_ (.A0(net4307),
    .A1(net2324),
    .S(net4249),
    .X(_00544_));
 sg13g2_mux2_1 _18010_ (.A0(net4301),
    .A1(net2861),
    .S(net4249),
    .X(_00545_));
 sg13g2_mux2_1 _18011_ (.A0(net4296),
    .A1(net2376),
    .S(net4252),
    .X(_00546_));
 sg13g2_mux2_1 _18012_ (.A0(net4290),
    .A1(net2661),
    .S(net4252),
    .X(_00547_));
 sg13g2_mux2_1 _18013_ (.A0(net4284),
    .A1(net2885),
    .S(net4249),
    .X(_00548_));
 sg13g2_mux2_1 _18014_ (.A0(net4279),
    .A1(net3656),
    .S(net4253),
    .X(_00549_));
 sg13g2_mux2_1 _18015_ (.A0(net4275),
    .A1(net3186),
    .S(net4251),
    .X(_00550_));
 sg13g2_mux2_1 _18016_ (.A0(net4273),
    .A1(net2488),
    .S(net4251),
    .X(_00551_));
 sg13g2_mux2_1 _18017_ (.A0(net4265),
    .A1(net2663),
    .S(net4249),
    .X(_00552_));
 sg13g2_mux2_1 _18018_ (.A0(net4260),
    .A1(net3527),
    .S(net4253),
    .X(_00553_));
 sg13g2_mux2_1 _18019_ (.A0(net4254),
    .A1(net3117),
    .S(net4252),
    .X(_00554_));
 sg13g2_mux2_1 _18020_ (.A0(net4404),
    .A1(net3427),
    .S(net4252),
    .X(_00555_));
 sg13g2_mux2_1 _18021_ (.A0(net4398),
    .A1(net2502),
    .S(net4251),
    .X(_00556_));
 sg13g2_mux2_1 _18022_ (.A0(net4393),
    .A1(net2812),
    .S(net4250),
    .X(_00557_));
 sg13g2_mux2_1 _18023_ (.A0(net4392),
    .A1(net2368),
    .S(net4249),
    .X(_00558_));
 sg13g2_mux2_1 _18024_ (.A0(net4387),
    .A1(net3663),
    .S(net4250),
    .X(_00559_));
 sg13g2_mux2_1 _18025_ (.A0(net4377),
    .A1(net2264),
    .S(net4252),
    .X(_00560_));
 sg13g2_mux2_1 _18026_ (.A0(net4373),
    .A1(net3360),
    .S(net4251),
    .X(_00561_));
 sg13g2_mux2_1 _18027_ (.A0(net4368),
    .A1(net3655),
    .S(net4253),
    .X(_00562_));
 sg13g2_or2_1 _18028_ (.X(_03181_),
    .B(_03168_),
    .A(_02993_));
 sg13g2_mux2_1 _18029_ (.A0(net4361),
    .A1(net2612),
    .S(net4155),
    .X(_00563_));
 sg13g2_mux2_1 _18030_ (.A0(net4357),
    .A1(net2410),
    .S(net4157),
    .X(_00564_));
 sg13g2_mux2_1 _18031_ (.A0(net4349),
    .A1(net2228),
    .S(net4156),
    .X(_00565_));
 sg13g2_mux2_1 _18032_ (.A0(net4344),
    .A1(net3052),
    .S(net4155),
    .X(_00566_));
 sg13g2_mux2_1 _18033_ (.A0(net4340),
    .A1(net3273),
    .S(net4157),
    .X(_00567_));
 sg13g2_mux2_1 _18034_ (.A0(net4196),
    .A1(net2689),
    .S(net4157),
    .X(_00568_));
 sg13g2_mux2_1 _18035_ (.A0(net4334),
    .A1(net3458),
    .S(net4156),
    .X(_00569_));
 sg13g2_mux2_1 _18036_ (.A0(net4329),
    .A1(net2824),
    .S(net4159),
    .X(_00570_));
 sg13g2_mux2_1 _18037_ (.A0(net4325),
    .A1(net2999),
    .S(net4157),
    .X(_00571_));
 sg13g2_mux2_1 _18038_ (.A0(net4320),
    .A1(net2215),
    .S(net4156),
    .X(_00572_));
 sg13g2_mux2_1 _18039_ (.A0(net4191),
    .A1(net2391),
    .S(net4158),
    .X(_00573_));
 sg13g2_mux2_1 _18040_ (.A0(net4185),
    .A1(net3239),
    .S(net4155),
    .X(_00574_));
 sg13g2_mux2_1 _18041_ (.A0(net4313),
    .A1(net2396),
    .S(net4158),
    .X(_00575_));
 sg13g2_mux2_1 _18042_ (.A0(net4307),
    .A1(net2497),
    .S(net4155),
    .X(_00576_));
 sg13g2_mux2_1 _18043_ (.A0(net4302),
    .A1(net3246),
    .S(net4155),
    .X(_00577_));
 sg13g2_mux2_1 _18044_ (.A0(net4297),
    .A1(net2238),
    .S(net4159),
    .X(_00578_));
 sg13g2_mux2_1 _18045_ (.A0(net4291),
    .A1(net2206),
    .S(net4158),
    .X(_00579_));
 sg13g2_mux2_1 _18046_ (.A0(net4286),
    .A1(net2492),
    .S(net4155),
    .X(_00580_));
 sg13g2_mux2_1 _18047_ (.A0(net4280),
    .A1(net2863),
    .S(net4158),
    .X(_00581_));
 sg13g2_mux2_1 _18048_ (.A0(net4276),
    .A1(net2425),
    .S(net4157),
    .X(_00582_));
 sg13g2_mux2_1 _18049_ (.A0(net4270),
    .A1(net2576),
    .S(net4157),
    .X(_00583_));
 sg13g2_mux2_1 _18050_ (.A0(net4264),
    .A1(net3255),
    .S(net4155),
    .X(_00584_));
 sg13g2_mux2_1 _18051_ (.A0(net4261),
    .A1(net2293),
    .S(net4159),
    .X(_00585_));
 sg13g2_mux2_1 _18052_ (.A0(net4254),
    .A1(net2318),
    .S(net4158),
    .X(_00586_));
 sg13g2_mux2_1 _18053_ (.A0(net4403),
    .A1(net2973),
    .S(net4158),
    .X(_00587_));
 sg13g2_mux2_1 _18054_ (.A0(net4399),
    .A1(net2369),
    .S(net4157),
    .X(_00588_));
 sg13g2_mux2_1 _18055_ (.A0(net4393),
    .A1(net2750),
    .S(net4156),
    .X(_00589_));
 sg13g2_mux2_1 _18056_ (.A0(net4389),
    .A1(net2611),
    .S(net4155),
    .X(_00590_));
 sg13g2_mux2_1 _18057_ (.A0(net4384),
    .A1(net2242),
    .S(net4156),
    .X(_00591_));
 sg13g2_mux2_1 _18058_ (.A0(net4377),
    .A1(net2485),
    .S(net4158),
    .X(_00592_));
 sg13g2_mux2_1 _18059_ (.A0(net4373),
    .A1(net2171),
    .S(net4157),
    .X(_00593_));
 sg13g2_mux2_1 _18060_ (.A0(net4367),
    .A1(net2728),
    .S(net4158),
    .X(_00594_));
 sg13g2_nand3_1 _18061_ (.B(_09804_),
    .C(_03179_),
    .A(_09657_),
    .Y(_03182_));
 sg13g2_mux2_1 _18062_ (.A0(net4362),
    .A1(net2243),
    .S(net4244),
    .X(_00595_));
 sg13g2_mux2_1 _18063_ (.A0(net4356),
    .A1(net2676),
    .S(net4246),
    .X(_00596_));
 sg13g2_mux2_1 _18064_ (.A0(net4349),
    .A1(net3406),
    .S(net4245),
    .X(_00597_));
 sg13g2_mux2_1 _18065_ (.A0(net4344),
    .A1(net2493),
    .S(net4244),
    .X(_00598_));
 sg13g2_mux2_1 _18066_ (.A0(net4339),
    .A1(net2629),
    .S(net4246),
    .X(_00599_));
 sg13g2_mux2_1 _18067_ (.A0(net4196),
    .A1(net2231),
    .S(net4246),
    .X(_00600_));
 sg13g2_mux2_1 _18068_ (.A0(net4334),
    .A1(net3187),
    .S(net4245),
    .X(_00601_));
 sg13g2_mux2_1 _18069_ (.A0(net4329),
    .A1(net3378),
    .S(net4247),
    .X(_00602_));
 sg13g2_mux2_1 _18070_ (.A0(net4324),
    .A1(net3597),
    .S(net4246),
    .X(_00603_));
 sg13g2_mux2_1 _18071_ (.A0(net4322),
    .A1(net2337),
    .S(net4245),
    .X(_00604_));
 sg13g2_mux2_1 _18072_ (.A0(net4190),
    .A1(net3048),
    .S(net4247),
    .X(_00605_));
 sg13g2_mux2_1 _18073_ (.A0(net4185),
    .A1(net3610),
    .S(net4244),
    .X(_00606_));
 sg13g2_mux2_1 _18074_ (.A0(net4312),
    .A1(net2968),
    .S(net4247),
    .X(_00607_));
 sg13g2_mux2_1 _18075_ (.A0(net4307),
    .A1(net3009),
    .S(net4244),
    .X(_00608_));
 sg13g2_mux2_1 _18076_ (.A0(net4301),
    .A1(net3446),
    .S(net4244),
    .X(_00609_));
 sg13g2_mux2_1 _18077_ (.A0(net4296),
    .A1(net2515),
    .S(net4247),
    .X(_00610_));
 sg13g2_mux2_1 _18078_ (.A0(net4290),
    .A1(net3628),
    .S(net4248),
    .X(_00611_));
 sg13g2_mux2_1 _18079_ (.A0(net4284),
    .A1(net3029),
    .S(net4244),
    .X(_00612_));
 sg13g2_mux2_1 _18080_ (.A0(net4279),
    .A1(net3232),
    .S(net4248),
    .X(_00613_));
 sg13g2_mux2_1 _18081_ (.A0(net4275),
    .A1(net3278),
    .S(net4246),
    .X(_00614_));
 sg13g2_mux2_1 _18082_ (.A0(net4269),
    .A1(net3491),
    .S(net4246),
    .X(_00615_));
 sg13g2_mux2_1 _18083_ (.A0(net4265),
    .A1(net3004),
    .S(net4244),
    .X(_00616_));
 sg13g2_mux2_1 _18084_ (.A0(net4260),
    .A1(net3081),
    .S(net4248),
    .X(_00617_));
 sg13g2_mux2_1 _18085_ (.A0(net4254),
    .A1(net3063),
    .S(net4247),
    .X(_00618_));
 sg13g2_mux2_1 _18086_ (.A0(net4404),
    .A1(net3039),
    .S(net4247),
    .X(_00619_));
 sg13g2_mux2_1 _18087_ (.A0(net4398),
    .A1(net3286),
    .S(net4246),
    .X(_00620_));
 sg13g2_mux2_1 _18088_ (.A0(net4393),
    .A1(net2556),
    .S(net4245),
    .X(_00621_));
 sg13g2_mux2_1 _18089_ (.A0(net4389),
    .A1(net3105),
    .S(net4244),
    .X(_00622_));
 sg13g2_mux2_1 _18090_ (.A0(net4386),
    .A1(net3469),
    .S(net4245),
    .X(_00623_));
 sg13g2_mux2_1 _18091_ (.A0(net4378),
    .A1(net3383),
    .S(net4247),
    .X(_00624_));
 sg13g2_mux2_1 _18092_ (.A0(net4372),
    .A1(net2758),
    .S(net4246),
    .X(_00625_));
 sg13g2_mux2_1 _18093_ (.A0(net4367),
    .A1(net3242),
    .S(net4247),
    .X(_00626_));
 sg13g2_or2_1 _18094_ (.X(_03183_),
    .B(_02993_),
    .A(_09668_));
 sg13g2_mux2_1 _18095_ (.A0(net4362),
    .A1(net3112),
    .S(net4150),
    .X(_00627_));
 sg13g2_mux2_1 _18096_ (.A0(net4355),
    .A1(net2656),
    .S(net4152),
    .X(_00628_));
 sg13g2_mux2_1 _18097_ (.A0(net4351),
    .A1(net3119),
    .S(net4151),
    .X(_00629_));
 sg13g2_mux2_1 _18098_ (.A0(net4344),
    .A1(net2742),
    .S(net4150),
    .X(_00630_));
 sg13g2_mux2_1 _18099_ (.A0(net4339),
    .A1(net3328),
    .S(net4152),
    .X(_00631_));
 sg13g2_mux2_1 _18100_ (.A0(net4195),
    .A1(net2248),
    .S(net4152),
    .X(_00632_));
 sg13g2_mux2_1 _18101_ (.A0(net4335),
    .A1(net2818),
    .S(net4151),
    .X(_00633_));
 sg13g2_mux2_1 _18102_ (.A0(net4329),
    .A1(net2817),
    .S(net4154),
    .X(_00634_));
 sg13g2_mux2_1 _18103_ (.A0(net4325),
    .A1(net2808),
    .S(net4152),
    .X(_00635_));
 sg13g2_mux2_1 _18104_ (.A0(net4320),
    .A1(net2599),
    .S(net4151),
    .X(_00636_));
 sg13g2_mux2_1 _18105_ (.A0(net4191),
    .A1(net2162),
    .S(net4153),
    .X(_00637_));
 sg13g2_mux2_1 _18106_ (.A0(net4186),
    .A1(net3521),
    .S(net4150),
    .X(_00638_));
 sg13g2_mux2_1 _18107_ (.A0(net4313),
    .A1(net2872),
    .S(net4153),
    .X(_00639_));
 sg13g2_mux2_1 _18108_ (.A0(net4309),
    .A1(net2838),
    .S(net4150),
    .X(_00640_));
 sg13g2_mux2_1 _18109_ (.A0(net4303),
    .A1(net2564),
    .S(net4150),
    .X(_00641_));
 sg13g2_mux2_1 _18110_ (.A0(net4297),
    .A1(net2900),
    .S(net4153),
    .X(_00642_));
 sg13g2_mux2_1 _18111_ (.A0(net4292),
    .A1(net2859),
    .S(net4153),
    .X(_00643_));
 sg13g2_mux2_1 _18112_ (.A0(net4285),
    .A1(net3031),
    .S(net4150),
    .X(_00644_));
 sg13g2_mux2_1 _18113_ (.A0(net4279),
    .A1(net2413),
    .S(net4153),
    .X(_00645_));
 sg13g2_mux2_1 _18114_ (.A0(net4274),
    .A1(net2514),
    .S(net4152),
    .X(_00646_));
 sg13g2_mux2_1 _18115_ (.A0(net4270),
    .A1(net2446),
    .S(net4152),
    .X(_00647_));
 sg13g2_mux2_1 _18116_ (.A0(net4266),
    .A1(net3190),
    .S(net4150),
    .X(_00648_));
 sg13g2_mux2_1 _18117_ (.A0(net4259),
    .A1(net2998),
    .S(net4154),
    .X(_00649_));
 sg13g2_mux2_1 _18118_ (.A0(net4255),
    .A1(net3482),
    .S(net4153),
    .X(_00650_));
 sg13g2_mux2_1 _18119_ (.A0(net4403),
    .A1(net2744),
    .S(net4153),
    .X(_00651_));
 sg13g2_mux2_1 _18120_ (.A0(net4400),
    .A1(net3096),
    .S(net4152),
    .X(_00652_));
 sg13g2_mux2_1 _18121_ (.A0(net4397),
    .A1(net2219),
    .S(net4151),
    .X(_00653_));
 sg13g2_mux2_1 _18122_ (.A0(net4388),
    .A1(net2623),
    .S(net4150),
    .X(_00654_));
 sg13g2_mux2_1 _18123_ (.A0(net4384),
    .A1(net3222),
    .S(net4151),
    .X(_00655_));
 sg13g2_mux2_1 _18124_ (.A0(net4377),
    .A1(net2209),
    .S(net4154),
    .X(_00656_));
 sg13g2_mux2_1 _18125_ (.A0(net4372),
    .A1(net2441),
    .S(net4152),
    .X(_00657_));
 sg13g2_mux2_1 _18126_ (.A0(net4367),
    .A1(net2429),
    .S(net4153),
    .X(_00658_));
 sg13g2_nand3_1 _18127_ (.B(_09804_),
    .C(_03179_),
    .A(_09658_),
    .Y(_03184_));
 sg13g2_mux2_1 _18128_ (.A0(net4362),
    .A1(net3370),
    .S(net4239),
    .X(_00659_));
 sg13g2_mux2_1 _18129_ (.A0(net4356),
    .A1(net2474),
    .S(net4241),
    .X(_00660_));
 sg13g2_mux2_1 _18130_ (.A0(net4349),
    .A1(net3212),
    .S(net4240),
    .X(_00661_));
 sg13g2_mux2_1 _18131_ (.A0(net4344),
    .A1(net2718),
    .S(net4239),
    .X(_00662_));
 sg13g2_mux2_1 _18132_ (.A0(net4339),
    .A1(net3061),
    .S(net4241),
    .X(_00663_));
 sg13g2_mux2_1 _18133_ (.A0(net4199),
    .A1(net2965),
    .S(net4241),
    .X(_00664_));
 sg13g2_mux2_1 _18134_ (.A0(net4334),
    .A1(net3402),
    .S(net4240),
    .X(_00665_));
 sg13g2_mux2_1 _18135_ (.A0(net4329),
    .A1(net2851),
    .S(net4242),
    .X(_00666_));
 sg13g2_mux2_1 _18136_ (.A0(net4324),
    .A1(net2417),
    .S(net4241),
    .X(_00667_));
 sg13g2_mux2_1 _18137_ (.A0(net4322),
    .A1(net2222),
    .S(net4240),
    .X(_00668_));
 sg13g2_mux2_1 _18138_ (.A0(net4190),
    .A1(net3102),
    .S(net4242),
    .X(_00669_));
 sg13g2_mux2_1 _18139_ (.A0(net4185),
    .A1(net3266),
    .S(net4239),
    .X(_00670_));
 sg13g2_mux2_1 _18140_ (.A0(net4312),
    .A1(net2292),
    .S(net4242),
    .X(_00671_));
 sg13g2_mux2_1 _18141_ (.A0(net4307),
    .A1(net2473),
    .S(net4239),
    .X(_00672_));
 sg13g2_mux2_1 _18142_ (.A0(net4301),
    .A1(net2682),
    .S(net4239),
    .X(_00673_));
 sg13g2_mux2_1 _18143_ (.A0(net4296),
    .A1(net3045),
    .S(net4242),
    .X(_00674_));
 sg13g2_mux2_1 _18144_ (.A0(net4290),
    .A1(net2554),
    .S(net4243),
    .X(_00675_));
 sg13g2_mux2_1 _18145_ (.A0(net4284),
    .A1(net3463),
    .S(net4239),
    .X(_00676_));
 sg13g2_mux2_1 _18146_ (.A0(net4279),
    .A1(net2605),
    .S(net4243),
    .X(_00677_));
 sg13g2_mux2_1 _18147_ (.A0(net4275),
    .A1(net2972),
    .S(net4241),
    .X(_00678_));
 sg13g2_mux2_1 _18148_ (.A0(net4269),
    .A1(net2505),
    .S(net4241),
    .X(_00679_));
 sg13g2_mux2_1 _18149_ (.A0(net4265),
    .A1(net2377),
    .S(net4239),
    .X(_00680_));
 sg13g2_mux2_1 _18150_ (.A0(net4260),
    .A1(net2822),
    .S(net4243),
    .X(_00681_));
 sg13g2_mux2_1 _18151_ (.A0(net4254),
    .A1(net3439),
    .S(net4242),
    .X(_00682_));
 sg13g2_mux2_1 _18152_ (.A0(net4407),
    .A1(net3046),
    .S(net4242),
    .X(_00683_));
 sg13g2_mux2_1 _18153_ (.A0(net4398),
    .A1(net2321),
    .S(net4241),
    .X(_00684_));
 sg13g2_mux2_1 _18154_ (.A0(net4394),
    .A1(net2216),
    .S(net4240),
    .X(_00685_));
 sg13g2_mux2_1 _18155_ (.A0(net4389),
    .A1(net2245),
    .S(net4239),
    .X(_00686_));
 sg13g2_mux2_1 _18156_ (.A0(net4386),
    .A1(net2772),
    .S(net4240),
    .X(_00687_));
 sg13g2_mux2_1 _18157_ (.A0(net4377),
    .A1(net2271),
    .S(net4242),
    .X(_00688_));
 sg13g2_mux2_1 _18158_ (.A0(net4373),
    .A1(net2443),
    .S(net4241),
    .X(_00689_));
 sg13g2_mux2_1 _18159_ (.A0(net4367),
    .A1(net2323),
    .S(net4242),
    .X(_00690_));
 sg13g2_nor3_1 _18160_ (.A(_09661_),
    .B(_09663_),
    .C(_09666_),
    .Y(_03185_));
 sg13g2_nand3_1 _18161_ (.B(_09657_),
    .C(_03185_),
    .A(_09655_),
    .Y(_03186_));
 sg13g2_mux2_1 _18162_ (.A0(net4361),
    .A1(net2727),
    .S(net4234),
    .X(_00691_));
 sg13g2_mux2_1 _18163_ (.A0(net4355),
    .A1(net3467),
    .S(net4236),
    .X(_00692_));
 sg13g2_mux2_1 _18164_ (.A0(net4351),
    .A1(net2471),
    .S(net4234),
    .X(_00693_));
 sg13g2_mux2_1 _18165_ (.A0(net4345),
    .A1(net3602),
    .S(net4236),
    .X(_00694_));
 sg13g2_mux2_1 _18166_ (.A0(net4339),
    .A1(net3325),
    .S(net4236),
    .X(_00695_));
 sg13g2_mux2_1 _18167_ (.A0(net4195),
    .A1(net3090),
    .S(net4236),
    .X(_00696_));
 sg13g2_mux2_1 _18168_ (.A0(_10235_),
    .A1(net2679),
    .S(net4235),
    .X(_00697_));
 sg13g2_mux2_1 _18169_ (.A0(net4331),
    .A1(net2362),
    .S(net4237),
    .X(_00698_));
 sg13g2_mux2_1 _18170_ (.A0(net4324),
    .A1(net2604),
    .S(net4236),
    .X(_00699_));
 sg13g2_mux2_1 _18171_ (.A0(net4321),
    .A1(net2635),
    .S(net4235),
    .X(_00700_));
 sg13g2_mux2_1 _18172_ (.A0(net4190),
    .A1(net3698),
    .S(net4237),
    .X(_00701_));
 sg13g2_mux2_1 _18173_ (.A0(net4186),
    .A1(net3466),
    .S(net4234),
    .X(_00702_));
 sg13g2_mux2_1 _18174_ (.A0(net4314),
    .A1(net3258),
    .S(net4237),
    .X(_00703_));
 sg13g2_mux2_1 _18175_ (.A0(net4308),
    .A1(net3536),
    .S(net4234),
    .X(_00704_));
 sg13g2_mux2_1 _18176_ (.A0(net4304),
    .A1(net2651),
    .S(net4234),
    .X(_00705_));
 sg13g2_mux2_1 _18177_ (.A0(net4296),
    .A1(net2649),
    .S(net4237),
    .X(_00706_));
 sg13g2_mux2_1 _18178_ (.A0(net4290),
    .A1(net3011),
    .S(net4237),
    .X(_00707_));
 sg13g2_mux2_1 _18179_ (.A0(net4284),
    .A1(net3616),
    .S(net4234),
    .X(_00708_));
 sg13g2_mux2_1 _18180_ (.A0(net4279),
    .A1(net3340),
    .S(net4237),
    .X(_00709_));
 sg13g2_mux2_1 _18181_ (.A0(net4274),
    .A1(net3296),
    .S(net4236),
    .X(_00710_));
 sg13g2_mux2_1 _18182_ (.A0(net4270),
    .A1(net3268),
    .S(net4236),
    .X(_00711_));
 sg13g2_mux2_1 _18183_ (.A0(net4268),
    .A1(net3411),
    .S(net4234),
    .X(_00712_));
 sg13g2_mux2_1 _18184_ (.A0(net4259),
    .A1(net2602),
    .S(net4238),
    .X(_00713_));
 sg13g2_mux2_1 _18185_ (.A0(net4256),
    .A1(net3474),
    .S(net4238),
    .X(_00714_));
 sg13g2_mux2_1 _18186_ (.A0(net4403),
    .A1(net3546),
    .S(net4237),
    .X(_00715_));
 sg13g2_mux2_1 _18187_ (.A0(net4398),
    .A1(net3158),
    .S(net4236),
    .X(_00716_));
 sg13g2_mux2_1 _18188_ (.A0(net4394),
    .A1(net3262),
    .S(net4235),
    .X(_00717_));
 sg13g2_mux2_1 _18189_ (.A0(net4388),
    .A1(net3088),
    .S(net4234),
    .X(_00718_));
 sg13g2_mux2_1 _18190_ (.A0(net4384),
    .A1(net2345),
    .S(net4235),
    .X(_00719_));
 sg13g2_mux2_1 _18191_ (.A0(net4377),
    .A1(net3375),
    .S(net4237),
    .X(_00720_));
 sg13g2_mux2_1 _18192_ (.A0(net4372),
    .A1(net2832),
    .S(net4238),
    .X(_00721_));
 sg13g2_mux2_1 _18193_ (.A0(net4368),
    .A1(net2958),
    .S(net4238),
    .X(_00722_));
 sg13g2_nand3_1 _18194_ (.B(_09804_),
    .C(_03185_),
    .A(_09657_),
    .Y(_03187_));
 sg13g2_mux2_1 _18195_ (.A0(net4361),
    .A1(net2606),
    .S(net4229),
    .X(_00723_));
 sg13g2_mux2_1 _18196_ (.A0(net4355),
    .A1(net3254),
    .S(net4231),
    .X(_00724_));
 sg13g2_mux2_1 _18197_ (.A0(net4349),
    .A1(net3188),
    .S(net4229),
    .X(_00725_));
 sg13g2_mux2_1 _18198_ (.A0(net4346),
    .A1(net3001),
    .S(net4231),
    .X(_00726_));
 sg13g2_mux2_1 _18199_ (.A0(net4339),
    .A1(net2619),
    .S(net4231),
    .X(_00727_));
 sg13g2_mux2_1 _18200_ (.A0(net4195),
    .A1(net2464),
    .S(net4231),
    .X(_00728_));
 sg13g2_mux2_1 _18201_ (.A0(net4335),
    .A1(net3016),
    .S(net4230),
    .X(_00729_));
 sg13g2_mux2_1 _18202_ (.A0(net4330),
    .A1(net2911),
    .S(net4232),
    .X(_00730_));
 sg13g2_mux2_1 _18203_ (.A0(net4324),
    .A1(net2173),
    .S(net4231),
    .X(_00731_));
 sg13g2_mux2_1 _18204_ (.A0(net4321),
    .A1(net3319),
    .S(net4230),
    .X(_00732_));
 sg13g2_mux2_1 _18205_ (.A0(net4190),
    .A1(net2904),
    .S(net4232),
    .X(_00733_));
 sg13g2_mux2_1 _18206_ (.A0(net4185),
    .A1(net2706),
    .S(net4229),
    .X(_00734_));
 sg13g2_mux2_1 _18207_ (.A0(net4314),
    .A1(net2609),
    .S(net4232),
    .X(_00735_));
 sg13g2_mux2_1 _18208_ (.A0(net4308),
    .A1(net3471),
    .S(net4229),
    .X(_00736_));
 sg13g2_mux2_1 _18209_ (.A0(net4304),
    .A1(net3177),
    .S(net4229),
    .X(_00737_));
 sg13g2_mux2_1 _18210_ (.A0(net4296),
    .A1(net3272),
    .S(net4232),
    .X(_00738_));
 sg13g2_mux2_1 _18211_ (.A0(net4290),
    .A1(net2908),
    .S(net4232),
    .X(_00739_));
 sg13g2_mux2_1 _18212_ (.A0(net4284),
    .A1(net3549),
    .S(net4229),
    .X(_00740_));
 sg13g2_mux2_1 _18213_ (.A0(net4279),
    .A1(net3279),
    .S(net4232),
    .X(_00741_));
 sg13g2_mux2_1 _18214_ (.A0(net4274),
    .A1(net3136),
    .S(net4231),
    .X(_00742_));
 sg13g2_mux2_1 _18215_ (.A0(net4270),
    .A1(net2754),
    .S(net4231),
    .X(_00743_));
 sg13g2_mux2_1 _18216_ (.A0(net4265),
    .A1(net2939),
    .S(net4229),
    .X(_00744_));
 sg13g2_mux2_1 _18217_ (.A0(net4259),
    .A1(net2332),
    .S(net4233),
    .X(_00745_));
 sg13g2_mux2_1 _18218_ (.A0(net4256),
    .A1(net3065),
    .S(net4233),
    .X(_00746_));
 sg13g2_mux2_1 _18219_ (.A0(net4403),
    .A1(net3217),
    .S(net4232),
    .X(_00747_));
 sg13g2_mux2_1 _18220_ (.A0(net4398),
    .A1(net2354),
    .S(net4231),
    .X(_00748_));
 sg13g2_mux2_1 _18221_ (.A0(net4393),
    .A1(net2960),
    .S(net4230),
    .X(_00749_));
 sg13g2_mux2_1 _18222_ (.A0(net4388),
    .A1(net2597),
    .S(net4229),
    .X(_00750_));
 sg13g2_mux2_1 _18223_ (.A0(net4384),
    .A1(net3226),
    .S(net4230),
    .X(_00751_));
 sg13g2_mux2_1 _18224_ (.A0(net4377),
    .A1(net3342),
    .S(net4232),
    .X(_00752_));
 sg13g2_mux2_1 _18225_ (.A0(net4372),
    .A1(net3563),
    .S(net4233),
    .X(_00753_));
 sg13g2_mux2_1 _18226_ (.A0(net4368),
    .A1(net3299),
    .S(net4233),
    .X(_00754_));
 sg13g2_nand3_1 _18227_ (.B(_09658_),
    .C(_03185_),
    .A(_09655_),
    .Y(_03188_));
 sg13g2_mux2_1 _18228_ (.A0(net4361),
    .A1(net2763),
    .S(net4224),
    .X(_00755_));
 sg13g2_mux2_1 _18229_ (.A0(net4355),
    .A1(net2286),
    .S(net4226),
    .X(_00756_));
 sg13g2_mux2_1 _18230_ (.A0(net4349),
    .A1(net2699),
    .S(net4224),
    .X(_00757_));
 sg13g2_mux2_1 _18231_ (.A0(net4345),
    .A1(net2850),
    .S(net4226),
    .X(_00758_));
 sg13g2_mux2_1 _18232_ (.A0(net4339),
    .A1(net2948),
    .S(net4226),
    .X(_00759_));
 sg13g2_mux2_1 _18233_ (.A0(net4195),
    .A1(net2823),
    .S(net4226),
    .X(_00760_));
 sg13g2_mux2_1 _18234_ (.A0(net4335),
    .A1(net2646),
    .S(net4225),
    .X(_00761_));
 sg13g2_mux2_1 _18235_ (.A0(net4330),
    .A1(net2342),
    .S(net4227),
    .X(_00762_));
 sg13g2_mux2_1 _18236_ (.A0(net4324),
    .A1(net3237),
    .S(net4226),
    .X(_00763_));
 sg13g2_mux2_1 _18237_ (.A0(net4321),
    .A1(net3236),
    .S(net4225),
    .X(_00764_));
 sg13g2_mux2_1 _18238_ (.A0(net4190),
    .A1(net2585),
    .S(net4227),
    .X(_00765_));
 sg13g2_mux2_1 _18239_ (.A0(net4186),
    .A1(net2180),
    .S(net4224),
    .X(_00766_));
 sg13g2_mux2_1 _18240_ (.A0(net4314),
    .A1(net2356),
    .S(net4227),
    .X(_00767_));
 sg13g2_mux2_1 _18241_ (.A0(net4308),
    .A1(net3389),
    .S(net4224),
    .X(_00768_));
 sg13g2_mux2_1 _18242_ (.A0(net4304),
    .A1(net3007),
    .S(net4224),
    .X(_00769_));
 sg13g2_mux2_1 _18243_ (.A0(net4296),
    .A1(net3442),
    .S(net4227),
    .X(_00770_));
 sg13g2_mux2_1 _18244_ (.A0(net4290),
    .A1(net3034),
    .S(net4227),
    .X(_00771_));
 sg13g2_mux2_1 _18245_ (.A0(net4284),
    .A1(net2915),
    .S(net4224),
    .X(_00772_));
 sg13g2_mux2_1 _18246_ (.A0(net4279),
    .A1(net3534),
    .S(net4227),
    .X(_00773_));
 sg13g2_mux2_1 _18247_ (.A0(net4274),
    .A1(net3260),
    .S(net4226),
    .X(_00774_));
 sg13g2_mux2_1 _18248_ (.A0(net4269),
    .A1(net3636),
    .S(net4226),
    .X(_00775_));
 sg13g2_mux2_1 _18249_ (.A0(net4265),
    .A1(net2749),
    .S(net4224),
    .X(_00776_));
 sg13g2_mux2_1 _18250_ (.A0(net4259),
    .A1(net3175),
    .S(net4228),
    .X(_00777_));
 sg13g2_mux2_1 _18251_ (.A0(net4256),
    .A1(net2251),
    .S(net4228),
    .X(_00778_));
 sg13g2_mux2_1 _18252_ (.A0(net4403),
    .A1(net3180),
    .S(net4227),
    .X(_00779_));
 sg13g2_mux2_1 _18253_ (.A0(net4398),
    .A1(net3036),
    .S(net4226),
    .X(_00780_));
 sg13g2_mux2_1 _18254_ (.A0(net4393),
    .A1(net2448),
    .S(net4225),
    .X(_00781_));
 sg13g2_mux2_1 _18255_ (.A0(net4388),
    .A1(net2317),
    .S(net4224),
    .X(_00782_));
 sg13g2_mux2_1 _18256_ (.A0(net4384),
    .A1(net3055),
    .S(net4225),
    .X(_00783_));
 sg13g2_mux2_1 _18257_ (.A0(net4377),
    .A1(net2436),
    .S(net4227),
    .X(_00784_));
 sg13g2_mux2_1 _18258_ (.A0(net4372),
    .A1(net2548),
    .S(net4228),
    .X(_00785_));
 sg13g2_mux2_1 _18259_ (.A0(net4368),
    .A1(net2454),
    .S(net4228),
    .X(_00786_));
 sg13g2_nand3_1 _18260_ (.B(_09804_),
    .C(_03185_),
    .A(_09658_),
    .Y(_03189_));
 sg13g2_mux2_1 _18261_ (.A0(net4361),
    .A1(net3432),
    .S(net4219),
    .X(_00787_));
 sg13g2_mux2_1 _18262_ (.A0(net4355),
    .A1(net2340),
    .S(net4221),
    .X(_00788_));
 sg13g2_mux2_1 _18263_ (.A0(net4349),
    .A1(net2253),
    .S(net4219),
    .X(_00789_));
 sg13g2_mux2_1 _18264_ (.A0(net4345),
    .A1(net3333),
    .S(net4221),
    .X(_00790_));
 sg13g2_mux2_1 _18265_ (.A0(net4339),
    .A1(net2632),
    .S(net4221),
    .X(_00791_));
 sg13g2_mux2_1 _18266_ (.A0(net4195),
    .A1(net3292),
    .S(net4221),
    .X(_00792_));
 sg13g2_mux2_1 _18267_ (.A0(net4334),
    .A1(net3358),
    .S(net4220),
    .X(_00793_));
 sg13g2_mux2_1 _18268_ (.A0(net4330),
    .A1(net2930),
    .S(net4222),
    .X(_00794_));
 sg13g2_mux2_1 _18269_ (.A0(net4324),
    .A1(net2926),
    .S(net4221),
    .X(_00795_));
 sg13g2_mux2_1 _18270_ (.A0(net4321),
    .A1(net2587),
    .S(net4220),
    .X(_00796_));
 sg13g2_mux2_1 _18271_ (.A0(net4190),
    .A1(net2669),
    .S(net4222),
    .X(_00797_));
 sg13g2_mux2_1 _18272_ (.A0(net4186),
    .A1(net2378),
    .S(net4219),
    .X(_00798_));
 sg13g2_mux2_1 _18273_ (.A0(net4314),
    .A1(net2862),
    .S(net4222),
    .X(_00799_));
 sg13g2_mux2_1 _18274_ (.A0(net4308),
    .A1(net2833),
    .S(net4219),
    .X(_00800_));
 sg13g2_mux2_1 _18275_ (.A0(net4304),
    .A1(net2702),
    .S(net4219),
    .X(_00801_));
 sg13g2_mux2_1 _18276_ (.A0(net4296),
    .A1(net2358),
    .S(net4222),
    .X(_00802_));
 sg13g2_mux2_1 _18277_ (.A0(net4290),
    .A1(net2394),
    .S(net4222),
    .X(_00803_));
 sg13g2_mux2_1 _18278_ (.A0(net4284),
    .A1(net2588),
    .S(net4219),
    .X(_00804_));
 sg13g2_mux2_1 _18279_ (.A0(net4280),
    .A1(net3459),
    .S(net4222),
    .X(_00805_));
 sg13g2_mux2_1 _18280_ (.A0(net4276),
    .A1(net2444),
    .S(net4221),
    .X(_00806_));
 sg13g2_mux2_1 _18281_ (.A0(net4269),
    .A1(net3199),
    .S(net4221),
    .X(_00807_));
 sg13g2_mux2_1 _18282_ (.A0(_10490_),
    .A1(net2236),
    .S(net4219),
    .X(_00808_));
 sg13g2_mux2_1 _18283_ (.A0(net4259),
    .A1(net3479),
    .S(net4223),
    .X(_00809_));
 sg13g2_mux2_1 _18284_ (.A0(net4256),
    .A1(net2828),
    .S(net4223),
    .X(_00810_));
 sg13g2_mux2_1 _18285_ (.A0(net4404),
    .A1(net3355),
    .S(net4222),
    .X(_00811_));
 sg13g2_mux2_1 _18286_ (.A0(net4398),
    .A1(net2495),
    .S(net4221),
    .X(_00812_));
 sg13g2_mux2_1 _18287_ (.A0(net4394),
    .A1(net2199),
    .S(net4220),
    .X(_00813_));
 sg13g2_mux2_1 _18288_ (.A0(net4388),
    .A1(net3295),
    .S(net4219),
    .X(_00814_));
 sg13g2_mux2_1 _18289_ (.A0(net4384),
    .A1(net2275),
    .S(net4220),
    .X(_00815_));
 sg13g2_mux2_1 _18290_ (.A0(net4377),
    .A1(net2266),
    .S(net4222),
    .X(_00816_));
 sg13g2_mux2_1 _18291_ (.A0(net4372),
    .A1(net2405),
    .S(net4223),
    .X(_00817_));
 sg13g2_mux2_1 _18292_ (.A0(net4368),
    .A1(net3335),
    .S(net4223),
    .X(_00818_));
 sg13g2_or2_1 _18293_ (.X(_03190_),
    .B(_03169_),
    .A(_09668_));
 sg13g2_mux2_1 _18294_ (.A0(net4363),
    .A1(net2730),
    .S(net4145),
    .X(_00819_));
 sg13g2_mux2_1 _18295_ (.A0(net4355),
    .A1(net2534),
    .S(net4147),
    .X(_00820_));
 sg13g2_mux2_1 _18296_ (.A0(net4351),
    .A1(net2986),
    .S(net4146),
    .X(_00821_));
 sg13g2_mux2_1 _18297_ (.A0(net4345),
    .A1(net3307),
    .S(net4145),
    .X(_00822_));
 sg13g2_mux2_1 _18298_ (.A0(net4343),
    .A1(net2847),
    .S(net4147),
    .X(_00823_));
 sg13g2_mux2_1 _18299_ (.A0(net4195),
    .A1(net3520),
    .S(net4147),
    .X(_00824_));
 sg13g2_mux2_1 _18300_ (.A0(net4335),
    .A1(net3194),
    .S(net4146),
    .X(_00825_));
 sg13g2_mux2_1 _18301_ (.A0(net4331),
    .A1(net3373),
    .S(net4149),
    .X(_00826_));
 sg13g2_mux2_1 _18302_ (.A0(net4325),
    .A1(net2974),
    .S(net4147),
    .X(_00827_));
 sg13g2_mux2_1 _18303_ (.A0(net4320),
    .A1(net3073),
    .S(net4146),
    .X(_00828_));
 sg13g2_mux2_1 _18304_ (.A0(net4191),
    .A1(net2889),
    .S(net4148),
    .X(_00829_));
 sg13g2_mux2_1 _18305_ (.A0(net4187),
    .A1(net2642),
    .S(net4145),
    .X(_00830_));
 sg13g2_mux2_1 _18306_ (.A0(net4313),
    .A1(net3570),
    .S(net4148),
    .X(_00831_));
 sg13g2_mux2_1 _18307_ (.A0(net4309),
    .A1(net3477),
    .S(net4145),
    .X(_00832_));
 sg13g2_mux2_1 _18308_ (.A0(net4303),
    .A1(net3129),
    .S(net4145),
    .X(_00833_));
 sg13g2_mux2_1 _18309_ (.A0(net4297),
    .A1(net3582),
    .S(net4148),
    .X(_00834_));
 sg13g2_mux2_1 _18310_ (.A0(net4292),
    .A1(net2336),
    .S(net4148),
    .X(_00835_));
 sg13g2_mux2_1 _18311_ (.A0(net4285),
    .A1(net3677),
    .S(net4145),
    .X(_00836_));
 sg13g2_mux2_1 _18312_ (.A0(net4283),
    .A1(net2821),
    .S(net4148),
    .X(_00837_));
 sg13g2_mux2_1 _18313_ (.A0(net4274),
    .A1(net2731),
    .S(net4147),
    .X(_00838_));
 sg13g2_mux2_1 _18314_ (.A0(net4270),
    .A1(net3475),
    .S(net4147),
    .X(_00839_));
 sg13g2_mux2_1 _18315_ (.A0(net4266),
    .A1(net3483),
    .S(net4145),
    .X(_00840_));
 sg13g2_mux2_1 _18316_ (.A0(net4259),
    .A1(net3531),
    .S(net4149),
    .X(_00841_));
 sg13g2_mux2_1 _18317_ (.A0(net4255),
    .A1(net3092),
    .S(net4148),
    .X(_00842_));
 sg13g2_mux2_1 _18318_ (.A0(net4403),
    .A1(net2811),
    .S(net4148),
    .X(_00843_));
 sg13g2_mux2_1 _18319_ (.A0(net4400),
    .A1(net2359),
    .S(net4147),
    .X(_00844_));
 sg13g2_mux2_1 _18320_ (.A0(net4397),
    .A1(net2607),
    .S(net4146),
    .X(_00845_));
 sg13g2_mux2_1 _18321_ (.A0(net4388),
    .A1(net3008),
    .S(net4145),
    .X(_00846_));
 sg13g2_mux2_1 _18322_ (.A0(net4385),
    .A1(net3132),
    .S(net4146),
    .X(_00847_));
 sg13g2_mux2_1 _18323_ (.A0(net4378),
    .A1(net3470),
    .S(net4149),
    .X(_00848_));
 sg13g2_mux2_1 _18324_ (.A0(net4373),
    .A1(net2570),
    .S(net4147),
    .X(_00849_));
 sg13g2_mux2_1 _18325_ (.A0(net4368),
    .A1(net3334),
    .S(net4148),
    .X(_00850_));
 sg13g2_nand3_1 _18326_ (.B(_09663_),
    .C(_09667_),
    .A(_09661_),
    .Y(_03191_));
 sg13g2_or2_1 _18327_ (.X(_03192_),
    .B(_03191_),
    .A(_03169_));
 sg13g2_mux2_1 _18328_ (.A0(net4365),
    .A1(net3329),
    .S(net4140),
    .X(_00851_));
 sg13g2_mux2_1 _18329_ (.A0(net4358),
    .A1(net2989),
    .S(net4142),
    .X(_00852_));
 sg13g2_mux2_1 _18330_ (.A0(net4352),
    .A1(net3601),
    .S(net4141),
    .X(_00853_));
 sg13g2_mux2_1 _18331_ (.A0(net4347),
    .A1(net2966),
    .S(net4141),
    .X(_00854_));
 sg13g2_mux2_1 _18332_ (.A0(net4342),
    .A1(net3541),
    .S(net4142),
    .X(_00855_));
 sg13g2_mux2_1 _18333_ (.A0(net4198),
    .A1(net2675),
    .S(net4144),
    .X(_00856_));
 sg13g2_mux2_1 _18334_ (.A0(net4337),
    .A1(net3399),
    .S(net4141),
    .X(_00857_));
 sg13g2_mux2_1 _18335_ (.A0(net4332),
    .A1(net2916),
    .S(net4143),
    .X(_00858_));
 sg13g2_mux2_1 _18336_ (.A0(net4326),
    .A1(net3116),
    .S(net4142),
    .X(_00859_));
 sg13g2_mux2_1 _18337_ (.A0(net4318),
    .A1(net2633),
    .S(net4140),
    .X(_00860_));
 sg13g2_mux2_1 _18338_ (.A0(net4193),
    .A1(net3461),
    .S(net4143),
    .X(_00861_));
 sg13g2_mux2_1 _18339_ (.A0(net4188),
    .A1(net3301),
    .S(net4140),
    .X(_00862_));
 sg13g2_mux2_1 _18340_ (.A0(net4315),
    .A1(net2813),
    .S(net4143),
    .X(_00863_));
 sg13g2_mux2_1 _18341_ (.A0(net4310),
    .A1(net2600),
    .S(net4140),
    .X(_00864_));
 sg13g2_mux2_1 _18342_ (.A0(net4305),
    .A1(net2765),
    .S(net4140),
    .X(_00865_));
 sg13g2_mux2_1 _18343_ (.A0(net4298),
    .A1(net3284),
    .S(net4142),
    .X(_00866_));
 sg13g2_mux2_1 _18344_ (.A0(net4293),
    .A1(net2622),
    .S(net4143),
    .X(_00867_));
 sg13g2_mux2_1 _18345_ (.A0(net4287),
    .A1(net2734),
    .S(net4140),
    .X(_00868_));
 sg13g2_mux2_1 _18346_ (.A0(net4281),
    .A1(net3620),
    .S(net4143),
    .X(_00869_));
 sg13g2_mux2_1 _18347_ (.A0(net4277),
    .A1(net2647),
    .S(net4141),
    .X(_00870_));
 sg13g2_mux2_1 _18348_ (.A0(net4272),
    .A1(net2586),
    .S(net4142),
    .X(_00871_));
 sg13g2_mux2_1 _18349_ (.A0(net4266),
    .A1(net2653),
    .S(net4140),
    .X(_00872_));
 sg13g2_mux2_1 _18350_ (.A0(net4263),
    .A1(net3361),
    .S(net4142),
    .X(_00873_));
 sg13g2_mux2_1 _18351_ (.A0(net4257),
    .A1(net3243),
    .S(net4144),
    .X(_00874_));
 sg13g2_mux2_1 _18352_ (.A0(net4405),
    .A1(net3353),
    .S(net4143),
    .X(_00875_));
 sg13g2_mux2_1 _18353_ (.A0(net4402),
    .A1(net3093),
    .S(net4142),
    .X(_00876_));
 sg13g2_mux2_1 _18354_ (.A0(net4395),
    .A1(net2639),
    .S(net4141),
    .X(_00877_));
 sg13g2_mux2_1 _18355_ (.A0(net4391),
    .A1(net3431),
    .S(net4141),
    .X(_00878_));
 sg13g2_mux2_1 _18356_ (.A0(net4386),
    .A1(net3104),
    .S(net4140),
    .X(_00879_));
 sg13g2_mux2_1 _18357_ (.A0(net4379),
    .A1(net3426),
    .S(net4143),
    .X(_00880_));
 sg13g2_mux2_1 _18358_ (.A0(net4374),
    .A1(net2239),
    .S(net4142),
    .X(_00881_));
 sg13g2_mux2_1 _18359_ (.A0(net4370),
    .A1(net2815),
    .S(net4143),
    .X(_00882_));
 sg13g2_or2_1 _18360_ (.X(_03193_),
    .B(_03191_),
    .A(_09659_));
 sg13g2_mux2_1 _18361_ (.A0(net4365),
    .A1(net3010),
    .S(net4135),
    .X(_00883_));
 sg13g2_mux2_1 _18362_ (.A0(net4358),
    .A1(net3006),
    .S(net4137),
    .X(_00884_));
 sg13g2_mux2_1 _18363_ (.A0(net4352),
    .A1(net3302),
    .S(net4136),
    .X(_00885_));
 sg13g2_mux2_1 _18364_ (.A0(net4347),
    .A1(net2601),
    .S(net4136),
    .X(_00886_));
 sg13g2_mux2_1 _18365_ (.A0(net4342),
    .A1(net3577),
    .S(net4137),
    .X(_00887_));
 sg13g2_mux2_1 _18366_ (.A0(net4197),
    .A1(net2415),
    .S(net4139),
    .X(_00888_));
 sg13g2_mux2_1 _18367_ (.A0(net4337),
    .A1(net2678),
    .S(net4136),
    .X(_00889_));
 sg13g2_mux2_1 _18368_ (.A0(net4332),
    .A1(net3267),
    .S(net4138),
    .X(_00890_));
 sg13g2_mux2_1 _18369_ (.A0(net4326),
    .A1(net2618),
    .S(net4137),
    .X(_00891_));
 sg13g2_mux2_1 _18370_ (.A0(net4318),
    .A1(net2395),
    .S(net4135),
    .X(_00892_));
 sg13g2_mux2_1 _18371_ (.A0(net4193),
    .A1(net3379),
    .S(net4138),
    .X(_00893_));
 sg13g2_mux2_1 _18372_ (.A0(net4188),
    .A1(net2709),
    .S(net4135),
    .X(_00894_));
 sg13g2_mux2_1 _18373_ (.A0(net4315),
    .A1(net3413),
    .S(net4138),
    .X(_00895_));
 sg13g2_mux2_1 _18374_ (.A0(net4310),
    .A1(net2178),
    .S(net4135),
    .X(_00896_));
 sg13g2_mux2_1 _18375_ (.A0(net4305),
    .A1(net3097),
    .S(net4135),
    .X(_00897_));
 sg13g2_mux2_1 _18376_ (.A0(net4299),
    .A1(net2698),
    .S(net4137),
    .X(_00898_));
 sg13g2_mux2_1 _18377_ (.A0(net4293),
    .A1(net2963),
    .S(net4138),
    .X(_00899_));
 sg13g2_mux2_1 _18378_ (.A0(net4287),
    .A1(net3331),
    .S(net4135),
    .X(_00900_));
 sg13g2_mux2_1 _18379_ (.A0(net4281),
    .A1(net2829),
    .S(net4138),
    .X(_00901_));
 sg13g2_mux2_1 _18380_ (.A0(net4277),
    .A1(net2146),
    .S(net4136),
    .X(_00902_));
 sg13g2_mux2_1 _18381_ (.A0(net4272),
    .A1(net3091),
    .S(net4137),
    .X(_00903_));
 sg13g2_mux2_1 _18382_ (.A0(net4267),
    .A1(net2710),
    .S(net4135),
    .X(_00904_));
 sg13g2_mux2_1 _18383_ (.A0(net4263),
    .A1(net2404),
    .S(net4137),
    .X(_00905_));
 sg13g2_mux2_1 _18384_ (.A0(net4257),
    .A1(net2416),
    .S(net4139),
    .X(_00906_));
 sg13g2_mux2_1 _18385_ (.A0(net4405),
    .A1(net3005),
    .S(net4138),
    .X(_00907_));
 sg13g2_mux2_1 _18386_ (.A0(net4402),
    .A1(net2761),
    .S(net4137),
    .X(_00908_));
 sg13g2_mux2_1 _18387_ (.A0(net4395),
    .A1(net2792),
    .S(net4136),
    .X(_00909_));
 sg13g2_mux2_1 _18388_ (.A0(net4391),
    .A1(net2780),
    .S(net4136),
    .X(_00910_));
 sg13g2_mux2_1 _18389_ (.A0(net4386),
    .A1(net2614),
    .S(net4135),
    .X(_00911_));
 sg13g2_mux2_1 _18390_ (.A0(net4379),
    .A1(net2645),
    .S(net4138),
    .X(_00912_));
 sg13g2_mux2_1 _18391_ (.A0(net4374),
    .A1(net2257),
    .S(net4137),
    .X(_00913_));
 sg13g2_mux2_1 _18392_ (.A0(net4369),
    .A1(net3015),
    .S(net4138),
    .X(_00914_));
 sg13g2_nor2_1 _18393_ (.A(net3203),
    .B(net4462),
    .Y(_03194_));
 sg13g2_a21oi_1 _18394_ (.A1(net4461),
    .A2(net4920),
    .Y(_00915_),
    .B1(_03194_));
 sg13g2_nor2_1 _18395_ (.A(net3805),
    .B(net4462),
    .Y(_03195_));
 sg13g2_a21oi_1 _18396_ (.A1(net4462),
    .A2(net4918),
    .Y(_00916_),
    .B1(_03195_));
 sg13g2_nor2_1 _18397_ (.A(net3144),
    .B(net4462),
    .Y(_03196_));
 sg13g2_a21oi_1 _18398_ (.A1(net4852),
    .A2(net4462),
    .Y(_00917_),
    .B1(_03196_));
 sg13g2_mux2_1 _18399_ (.A0(net3854),
    .A1(net4844),
    .S(net4462),
    .X(_00918_));
 sg13g2_mux2_1 _18400_ (.A0(net3881),
    .A1(net4839),
    .S(net4461),
    .X(_00919_));
 sg13g2_nor2_1 _18401_ (.A(net3171),
    .B(net4461),
    .Y(_03197_));
 sg13g2_a21oi_1 _18402_ (.A1(net4461),
    .A2(net4836),
    .Y(_00920_),
    .B1(_03197_));
 sg13g2_nor2_1 _18403_ (.A(net3120),
    .B(net4461),
    .Y(_03198_));
 sg13g2_a21oi_1 _18404_ (.A1(net4461),
    .A2(net4833),
    .Y(_00921_),
    .B1(_03198_));
 sg13g2_nor2_1 _18405_ (.A(net3382),
    .B(net4461),
    .Y(_03199_));
 sg13g2_a21oi_1 _18406_ (.A1(net4461),
    .A2(net4831),
    .Y(_00922_),
    .B1(_03199_));
 sg13g2_nor2_2 _18407_ (.A(_08845_),
    .B(net4941),
    .Y(_03200_));
 sg13g2_nand2b_2 _18408_ (.Y(_03201_),
    .B(_09559_),
    .A_N(_08845_));
 sg13g2_nor2_1 _18409_ (.A(net5624),
    .B(_09559_),
    .Y(_03202_));
 sg13g2_a22oi_1 _18410_ (.Y(_03203_),
    .B1(net4911),
    .B2(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .A2(net4555),
    .A1(net6227));
 sg13g2_o21ai_1 _18411_ (.B1(net6228),
    .Y(_00923_),
    .A1(_06562_),
    .A2(net4541));
 sg13g2_a22oi_1 _18412_ (.Y(_03204_),
    .B1(net4913),
    .B2(\fpga_top.cpu_top.csr_wdata_mon[1] ),
    .A2(net4555),
    .A1(net6134));
 sg13g2_o21ai_1 _18413_ (.B1(net6135),
    .Y(_00924_),
    .A1(_06561_),
    .A2(net4541));
 sg13g2_nand2_1 _18414_ (.Y(_03205_),
    .A(net2796),
    .B(net4550));
 sg13g2_a22oi_1 _18415_ (.Y(_03206_),
    .B1(net4911),
    .B2(net5664),
    .A2(net4549),
    .A1(\fpga_top.bus_gather.d_write_data[2] ));
 sg13g2_nand2_1 _18416_ (.Y(_00925_),
    .A(_03205_),
    .B(_03206_));
 sg13g2_a22oi_1 _18417_ (.Y(_03207_),
    .B1(net4912),
    .B2(net5662),
    .A2(net4556),
    .A1(net6160));
 sg13g2_o21ai_1 _18418_ (.B1(net6161),
    .Y(_00926_),
    .A1(_06570_),
    .A2(net4542));
 sg13g2_a22oi_1 _18419_ (.Y(_03208_),
    .B1(net4913),
    .B2(net5660),
    .A2(net4556),
    .A1(net4053));
 sg13g2_o21ai_1 _18420_ (.B1(net4054),
    .Y(_00927_),
    .A1(_06577_),
    .A2(net4542));
 sg13g2_a22oi_1 _18421_ (.Y(_03209_),
    .B1(net4911),
    .B2(net5658),
    .A2(net4550),
    .A1(net6230));
 sg13g2_o21ai_1 _18422_ (.B1(_03209_),
    .Y(_00928_),
    .A1(_06586_),
    .A2(net4541));
 sg13g2_nand2_1 _18423_ (.Y(_03210_),
    .A(net1782),
    .B(net4550));
 sg13g2_a22oi_1 _18424_ (.Y(_03211_),
    .B1(net4913),
    .B2(\fpga_top.cpu_start_adr[6] ),
    .A2(net4549),
    .A1(\fpga_top.bus_gather.d_write_data[6] ));
 sg13g2_nand2_1 _18425_ (.Y(_00929_),
    .A(_03210_),
    .B(_03211_));
 sg13g2_nand2_1 _18426_ (.Y(_03212_),
    .A(net1904),
    .B(net4550));
 sg13g2_a22oi_1 _18427_ (.Y(_03213_),
    .B1(net4913),
    .B2(net5656),
    .A2(net4549),
    .A1(\fpga_top.bus_gather.d_write_data[7] ));
 sg13g2_nand2_1 _18428_ (.Y(_00930_),
    .A(_03212_),
    .B(_03213_));
 sg13g2_nand2_1 _18429_ (.Y(_03214_),
    .A(net1838),
    .B(net4550));
 sg13g2_a22oi_1 _18430_ (.Y(_03215_),
    .B1(net4911),
    .B2(net5654),
    .A2(net4549),
    .A1(\fpga_top.bus_gather.d_write_data[8] ));
 sg13g2_nand2_1 _18431_ (.Y(_00931_),
    .A(_03214_),
    .B(_03215_));
 sg13g2_nand2_1 _18432_ (.Y(_03216_),
    .A(net1667),
    .B(net4550));
 sg13g2_a22oi_1 _18433_ (.Y(_03217_),
    .B1(net4911),
    .B2(net5653),
    .A2(net4549),
    .A1(\fpga_top.bus_gather.d_write_data[9] ));
 sg13g2_nand2_1 _18434_ (.Y(_00932_),
    .A(_03216_),
    .B(_03217_));
 sg13g2_a22oi_1 _18435_ (.Y(_03218_),
    .B1(net4912),
    .B2(net5652),
    .A2(net4556),
    .A1(net6191));
 sg13g2_o21ai_1 _18436_ (.B1(_03218_),
    .Y(_00933_),
    .A1(_06593_),
    .A2(net4542));
 sg13g2_nand2_1 _18437_ (.Y(_03219_),
    .A(net2115),
    .B(net4556));
 sg13g2_a22oi_1 _18438_ (.Y(_03220_),
    .B1(net4914),
    .B2(net5651),
    .A2(net4549),
    .A1(\fpga_top.bus_gather.d_write_data[11] ));
 sg13g2_nand2_1 _18439_ (.Y(_00934_),
    .A(_03219_),
    .B(_03220_));
 sg13g2_a22oi_1 _18440_ (.Y(_03221_),
    .B1(net4912),
    .B2(\fpga_top.cpu_start_adr[12] ),
    .A2(net4556),
    .A1(net6243));
 sg13g2_o21ai_1 _18441_ (.B1(net6244),
    .Y(_00935_),
    .A1(_06598_),
    .A2(net4542));
 sg13g2_a22oi_1 _18442_ (.Y(_03222_),
    .B1(net4913),
    .B2(\fpga_top.cpu_start_adr[13] ),
    .A2(net4556),
    .A1(net6235));
 sg13g2_o21ai_1 _18443_ (.B1(net6236),
    .Y(_00936_),
    .A1(_06600_),
    .A2(net4541));
 sg13g2_a22oi_1 _18444_ (.Y(_03223_),
    .B1(net4914),
    .B2(net5650),
    .A2(net4557),
    .A1(net6183));
 sg13g2_o21ai_1 _18445_ (.B1(net6184),
    .Y(_00937_),
    .A1(_06602_),
    .A2(net4544));
 sg13g2_a22oi_1 _18446_ (.Y(_03224_),
    .B1(net4914),
    .B2(\fpga_top.cpu_start_adr[15] ),
    .A2(net4557),
    .A1(net6138));
 sg13g2_o21ai_1 _18447_ (.B1(net6139),
    .Y(_00938_),
    .A1(_06604_),
    .A2(net4544));
 sg13g2_a22oi_1 _18448_ (.Y(_03225_),
    .B1(net4911),
    .B2(net5649),
    .A2(net4559),
    .A1(net6251));
 sg13g2_o21ai_1 _18449_ (.B1(net6252),
    .Y(_00939_),
    .A1(_06606_),
    .A2(net4541));
 sg13g2_a22oi_1 _18450_ (.Y(_03226_),
    .B1(net4911),
    .B2(net5648),
    .A2(net4555),
    .A1(net6222));
 sg13g2_o21ai_1 _18451_ (.B1(_03226_),
    .Y(_00940_),
    .A1(_06610_),
    .A2(net4543));
 sg13g2_a22oi_1 _18452_ (.Y(_03227_),
    .B1(net4914),
    .B2(net5647),
    .A2(net4557),
    .A1(net6126));
 sg13g2_o21ai_1 _18453_ (.B1(net6127),
    .Y(_00941_),
    .A1(_06612_),
    .A2(net4544));
 sg13g2_a22oi_1 _18454_ (.Y(_03228_),
    .B1(net4914),
    .B2(\fpga_top.cpu_start_adr[19] ),
    .A2(net4557),
    .A1(net4030));
 sg13g2_o21ai_1 _18455_ (.B1(net4031),
    .Y(_00942_),
    .A1(_06616_),
    .A2(net4544));
 sg13g2_a22oi_1 _18456_ (.Y(_03229_),
    .B1(net4912),
    .B2(net5646),
    .A2(net4555),
    .A1(net6187));
 sg13g2_o21ai_1 _18457_ (.B1(_03229_),
    .Y(_00943_),
    .A1(_06619_),
    .A2(net4543));
 sg13g2_a22oi_1 _18458_ (.Y(_03230_),
    .B1(net4912),
    .B2(net5644),
    .A2(net4555),
    .A1(net3962));
 sg13g2_o21ai_1 _18459_ (.B1(_03230_),
    .Y(_00944_),
    .A1(_06622_),
    .A2(net4542));
 sg13g2_a22oi_1 _18460_ (.Y(_03231_),
    .B1(net4915),
    .B2(net5643),
    .A2(net4558),
    .A1(net3990));
 sg13g2_o21ai_1 _18461_ (.B1(net3991),
    .Y(_00945_),
    .A1(_06624_),
    .A2(net4545));
 sg13g2_a22oi_1 _18462_ (.Y(_03232_),
    .B1(net4914),
    .B2(net5642),
    .A2(net4557),
    .A1(net4058));
 sg13g2_o21ai_1 _18463_ (.B1(net4059),
    .Y(_00946_),
    .A1(_06625_),
    .A2(net4545));
 sg13g2_a22oi_1 _18464_ (.Y(_03233_),
    .B1(net4915),
    .B2(\fpga_top.cpu_start_adr[24] ),
    .A2(net4557),
    .A1(net6103));
 sg13g2_o21ai_1 _18465_ (.B1(net6104),
    .Y(_00947_),
    .A1(_06628_),
    .A2(net4544));
 sg13g2_a22oi_1 _18466_ (.Y(_03234_),
    .B1(net4915),
    .B2(\fpga_top.cpu_start_adr[25] ),
    .A2(net4558),
    .A1(net6144));
 sg13g2_o21ai_1 _18467_ (.B1(net6145),
    .Y(_00948_),
    .A1(_06630_),
    .A2(net4544));
 sg13g2_a22oi_1 _18468_ (.Y(_03235_),
    .B1(net4914),
    .B2(\fpga_top.cpu_start_adr[26] ),
    .A2(net4556),
    .A1(net4062));
 sg13g2_o21ai_1 _18469_ (.B1(net4063),
    .Y(_00949_),
    .A1(_06633_),
    .A2(net4544));
 sg13g2_a22oi_1 _18470_ (.Y(_03236_),
    .B1(net4911),
    .B2(net5640),
    .A2(net4550),
    .A1(net3983));
 sg13g2_o21ai_1 _18471_ (.B1(_03236_),
    .Y(_00950_),
    .A1(_06635_),
    .A2(net4541));
 sg13g2_a22oi_1 _18472_ (.Y(_03237_),
    .B1(net4912),
    .B2(net5638),
    .A2(net4555),
    .A1(net4070));
 sg13g2_o21ai_1 _18473_ (.B1(_03237_),
    .Y(_00951_),
    .A1(_06639_),
    .A2(net4542));
 sg13g2_a22oi_1 _18474_ (.Y(_03238_),
    .B1(net4912),
    .B2(net5637),
    .A2(net4555),
    .A1(net6177));
 sg13g2_o21ai_1 _18475_ (.B1(_03238_),
    .Y(_00952_),
    .A1(_06640_),
    .A2(net4541));
 sg13g2_a22oi_1 _18476_ (.Y(_03239_),
    .B1(net4912),
    .B2(net5635),
    .A2(net4555),
    .A1(net6113));
 sg13g2_o21ai_1 _18477_ (.B1(_03239_),
    .Y(_00953_),
    .A1(_06642_),
    .A2(net4541));
 sg13g2_a22oi_1 _18478_ (.Y(_03240_),
    .B1(net4914),
    .B2(net2221),
    .A2(net4557),
    .A1(net3876));
 sg13g2_o21ai_1 _18479_ (.B1(_03240_),
    .Y(_00954_),
    .A1(_06645_),
    .A2(net4544));
 sg13g2_nor2b_2 _18480_ (.A(net4535),
    .B_N(net4558),
    .Y(_03241_));
 sg13g2_inv_1 _18481_ (.Y(_03242_),
    .A(_03241_));
 sg13g2_a21oi_2 _18482_ (.B1(_09551_),
    .Y(_03243_),
    .A2(net4941),
    .A1(net4570));
 sg13g2_a21oi_1 _18483_ (.A1(_08845_),
    .A2(net4570),
    .Y(_03244_),
    .B1(_07606_));
 sg13g2_a22oi_1 _18484_ (.Y(_00955_),
    .B1(_03243_),
    .B2(_03244_),
    .A2(_03241_),
    .A1(_06815_));
 sg13g2_a21oi_1 _18485_ (.A1(_08845_),
    .A2(net4570),
    .Y(_03245_),
    .B1(net5343));
 sg13g2_o21ai_1 _18486_ (.B1(_03243_),
    .Y(_03246_),
    .A1(net6327),
    .A2(_03242_));
 sg13g2_nor2_1 _18487_ (.A(_03245_),
    .B(_03246_),
    .Y(_00956_));
 sg13g2_nand2b_1 _18488_ (.Y(_03247_),
    .B(_09099_),
    .A_N(_09096_));
 sg13g2_nor2b_1 _18489_ (.A(\fpga_top.qspi_if.qspi_state[11] ),
    .B_N(_09088_),
    .Y(_03248_));
 sg13g2_nand2b_1 _18490_ (.Y(_03249_),
    .B(_03248_),
    .A_N(_03247_));
 sg13g2_inv_1 _18491_ (.Y(_03250_),
    .A(net4755));
 sg13g2_nand2_1 _18492_ (.Y(_03251_),
    .A(_08870_),
    .B(net4755));
 sg13g2_nand2_1 _18493_ (.Y(_03252_),
    .A(\fpga_top.qspi_if.rdedge[2] ),
    .B(_00089_));
 sg13g2_o21ai_1 _18494_ (.B1(_00090_),
    .Y(_03253_),
    .A1(_00095_),
    .A2(_03252_));
 sg13g2_and3_1 _18495_ (.X(_03254_),
    .A(_00123_),
    .B(_06676_),
    .C(net4948));
 sg13g2_nor2b_1 _18496_ (.A(_00115_),
    .B_N(_00107_),
    .Y(_03255_));
 sg13g2_and2_1 _18497_ (.A(\fpga_top.qspi_if.rdedge[2] ),
    .B(_00087_),
    .X(_03256_));
 sg13g2_a22oi_1 _18498_ (.Y(_03257_),
    .B1(_03256_),
    .B2(_06930_),
    .A2(_03255_),
    .A1(_06676_));
 sg13g2_a21oi_1 _18499_ (.A1(_06500_),
    .A2(_03257_),
    .Y(_03258_),
    .B1(\fpga_top.qspi_if.rdedge[0] ));
 sg13g2_o21ai_1 _18500_ (.B1(_03258_),
    .Y(_03259_),
    .A1(_03253_),
    .A2(_03254_));
 sg13g2_nor2b_1 _18501_ (.A(_00107_),
    .B_N(_00095_),
    .Y(_03260_));
 sg13g2_nor2_1 _18502_ (.A(_00123_),
    .B(_06500_),
    .Y(_03261_));
 sg13g2_a221oi_1 _18503_ (.B2(_00115_),
    .C1(\fpga_top.qspi_if.rdedge[2] ),
    .B1(_03261_),
    .A1(_06500_),
    .Y(_03262_),
    .A2(_03260_));
 sg13g2_nand2_1 _18504_ (.Y(_03263_),
    .A(_06500_),
    .B(_00086_));
 sg13g2_nor3_1 _18505_ (.A(_06500_),
    .B(_06930_),
    .C(_00089_),
    .Y(_03264_));
 sg13g2_o21ai_1 _18506_ (.B1(\fpga_top.qspi_if.rdedge[2] ),
    .Y(_03265_),
    .A1(_00087_),
    .A2(_03263_));
 sg13g2_o21ai_1 _18507_ (.B1(\fpga_top.qspi_if.rdedge[0] ),
    .Y(_03266_),
    .A1(_03264_),
    .A2(_03265_));
 sg13g2_o21ai_1 _18508_ (.B1(_03259_),
    .Y(_03267_),
    .A1(_03262_),
    .A2(_03266_));
 sg13g2_nand2_2 _18509_ (.Y(_03268_),
    .A(_03251_),
    .B(_03267_));
 sg13g2_mux2_1 _18510_ (.A0(net3737),
    .A1(\fpga_top.qspi_if.word_data[0] ),
    .S(net4710),
    .X(_00957_));
 sg13g2_mux2_1 _18511_ (.A0(net3765),
    .A1(\fpga_top.qspi_if.word_data[1] ),
    .S(net4710),
    .X(_00958_));
 sg13g2_mux2_1 _18512_ (.A0(net1629),
    .A1(\fpga_top.qspi_if.word_data[2] ),
    .S(net4710),
    .X(_00959_));
 sg13g2_mux2_1 _18513_ (.A0(net3743),
    .A1(\fpga_top.qspi_if.word_data[3] ),
    .S(net4710),
    .X(_00960_));
 sg13g2_nand2_1 _18514_ (.Y(_03269_),
    .A(\fpga_top.qspi_if.word_data[0] ),
    .B(net4750));
 sg13g2_nand2_1 _18515_ (.Y(_03270_),
    .A(net3288),
    .B(net4702));
 sg13g2_o21ai_1 _18516_ (.B1(_03270_),
    .Y(_00961_),
    .A1(net4702),
    .A2(_03269_));
 sg13g2_nand2_1 _18517_ (.Y(_03271_),
    .A(\fpga_top.qspi_if.word_data[1] ),
    .B(net4752));
 sg13g2_nand2_1 _18518_ (.Y(_03272_),
    .A(net2095),
    .B(net4705));
 sg13g2_o21ai_1 _18519_ (.B1(_03272_),
    .Y(_00962_),
    .A1(net4705),
    .A2(_03271_));
 sg13g2_nand2_1 _18520_ (.Y(_03273_),
    .A(\fpga_top.qspi_if.word_data[2] ),
    .B(net4753));
 sg13g2_nand2_1 _18521_ (.Y(_03274_),
    .A(net3879),
    .B(net4706));
 sg13g2_o21ai_1 _18522_ (.B1(_03274_),
    .Y(_00963_),
    .A1(net4705),
    .A2(_03273_));
 sg13g2_nand2_1 _18523_ (.Y(_03275_),
    .A(\fpga_top.qspi_if.word_data[3] ),
    .B(net4750));
 sg13g2_nand2_1 _18524_ (.Y(_03276_),
    .A(net3790),
    .B(net4703));
 sg13g2_o21ai_1 _18525_ (.B1(_03276_),
    .Y(_00964_),
    .A1(net4702),
    .A2(_03275_));
 sg13g2_nand2_1 _18526_ (.Y(_03277_),
    .A(net3288),
    .B(net4751));
 sg13g2_nand2_1 _18527_ (.Y(_03278_),
    .A(net3837),
    .B(net4701));
 sg13g2_o21ai_1 _18528_ (.B1(_03278_),
    .Y(_00965_),
    .A1(net4701),
    .A2(_03277_));
 sg13g2_nand2_1 _18529_ (.Y(_03279_),
    .A(net2095),
    .B(net4753));
 sg13g2_nand2_1 _18530_ (.Y(_03280_),
    .A(net2241),
    .B(net4705));
 sg13g2_o21ai_1 _18531_ (.B1(_03280_),
    .Y(_00966_),
    .A1(net4705),
    .A2(_03279_));
 sg13g2_nand2_1 _18532_ (.Y(_03281_),
    .A(\fpga_top.qspi_if.word_data[6] ),
    .B(net4752));
 sg13g2_nand2_1 _18533_ (.Y(_03282_),
    .A(net1863),
    .B(net4706));
 sg13g2_o21ai_1 _18534_ (.B1(_03282_),
    .Y(_00967_),
    .A1(net4705),
    .A2(_03281_));
 sg13g2_nand2_1 _18535_ (.Y(_03283_),
    .A(\fpga_top.qspi_if.word_data[7] ),
    .B(net4750));
 sg13g2_nand2_1 _18536_ (.Y(_03284_),
    .A(net1999),
    .B(net4702));
 sg13g2_o21ai_1 _18537_ (.B1(_03284_),
    .Y(_00968_),
    .A1(net4702),
    .A2(_03283_));
 sg13g2_nand2_1 _18538_ (.Y(_03285_),
    .A(\fpga_top.qspi_if.word_data[8] ),
    .B(net4750));
 sg13g2_nand2_1 _18539_ (.Y(_03286_),
    .A(net3728),
    .B(net4700));
 sg13g2_o21ai_1 _18540_ (.B1(_03286_),
    .Y(_00969_),
    .A1(net4700),
    .A2(_03285_));
 sg13g2_nand2_1 _18541_ (.Y(_03287_),
    .A(\fpga_top.qspi_if.word_data[9] ),
    .B(net4753));
 sg13g2_nand2_1 _18542_ (.Y(_03288_),
    .A(net1718),
    .B(net4705));
 sg13g2_o21ai_1 _18543_ (.B1(_03288_),
    .Y(_00970_),
    .A1(net4705),
    .A2(_03287_));
 sg13g2_nand2_1 _18544_ (.Y(_03289_),
    .A(net1863),
    .B(net4753));
 sg13g2_nand2_1 _18545_ (.Y(_03290_),
    .A(net3207),
    .B(net4704));
 sg13g2_o21ai_1 _18546_ (.B1(_03290_),
    .Y(_00971_),
    .A1(net4704),
    .A2(_03289_));
 sg13g2_nand2_1 _18547_ (.Y(_03291_),
    .A(\fpga_top.qspi_if.word_data[11] ),
    .B(net4750));
 sg13g2_nand2_1 _18548_ (.Y(_03292_),
    .A(net1910),
    .B(net4701));
 sg13g2_o21ai_1 _18549_ (.B1(_03292_),
    .Y(_00972_),
    .A1(net4700),
    .A2(_03291_));
 sg13g2_nand2_1 _18550_ (.Y(_03293_),
    .A(\fpga_top.qspi_if.word_data[12] ),
    .B(net4750));
 sg13g2_nand2_1 _18551_ (.Y(_03294_),
    .A(net2006),
    .B(net4702));
 sg13g2_o21ai_1 _18552_ (.B1(_03294_),
    .Y(_00973_),
    .A1(net4700),
    .A2(_03293_));
 sg13g2_nand2_1 _18553_ (.Y(_03295_),
    .A(\fpga_top.qspi_if.word_data[13] ),
    .B(net4752));
 sg13g2_nand2_1 _18554_ (.Y(_03296_),
    .A(net1610),
    .B(net4707));
 sg13g2_o21ai_1 _18555_ (.B1(_03296_),
    .Y(_00974_),
    .A1(net4708),
    .A2(_03295_));
 sg13g2_nand2_1 _18556_ (.Y(_03297_),
    .A(\fpga_top.qspi_if.word_data[14] ),
    .B(net4753));
 sg13g2_nand2_1 _18557_ (.Y(_03298_),
    .A(net1784),
    .B(net4706));
 sg13g2_o21ai_1 _18558_ (.B1(_03298_),
    .Y(_00975_),
    .A1(net4706),
    .A2(_03297_));
 sg13g2_nand2_1 _18559_ (.Y(_03299_),
    .A(\fpga_top.qspi_if.word_data[15] ),
    .B(net4751));
 sg13g2_nand2_1 _18560_ (.Y(_03300_),
    .A(net1846),
    .B(net4704));
 sg13g2_o21ai_1 _18561_ (.B1(_03300_),
    .Y(_00976_),
    .A1(net4703),
    .A2(_03299_));
 sg13g2_nand2_1 _18562_ (.Y(_03301_),
    .A(\fpga_top.qspi_if.word_data[16] ),
    .B(net4751));
 sg13g2_nand2_1 _18563_ (.Y(_03302_),
    .A(net1657),
    .B(net4703));
 sg13g2_o21ai_1 _18564_ (.B1(_03302_),
    .Y(_00977_),
    .A1(net4703),
    .A2(_03301_));
 sg13g2_nand2_1 _18565_ (.Y(_03303_),
    .A(net1610),
    .B(net4753));
 sg13g2_nand2_1 _18566_ (.Y(_03304_),
    .A(net1660),
    .B(net4707));
 sg13g2_o21ai_1 _18567_ (.B1(_03304_),
    .Y(_00978_),
    .A1(net4707),
    .A2(_03303_));
 sg13g2_nand2_1 _18568_ (.Y(_03305_),
    .A(\fpga_top.qspi_if.word_data[18] ),
    .B(net4752));
 sg13g2_nand2_1 _18569_ (.Y(_03306_),
    .A(net1669),
    .B(net4708));
 sg13g2_o21ai_1 _18570_ (.B1(_03306_),
    .Y(_00979_),
    .A1(net4708),
    .A2(_03305_));
 sg13g2_nand2_1 _18571_ (.Y(_03307_),
    .A(net1846),
    .B(net4753));
 sg13g2_nand2_1 _18572_ (.Y(_03308_),
    .A(net2042),
    .B(net4704));
 sg13g2_o21ai_1 _18573_ (.B1(_03308_),
    .Y(_00980_),
    .A1(net4704),
    .A2(_03307_));
 sg13g2_nand2_1 _18574_ (.Y(_03309_),
    .A(net1657),
    .B(net4751));
 sg13g2_nand2_1 _18575_ (.Y(_03310_),
    .A(net1927),
    .B(net4700));
 sg13g2_o21ai_1 _18576_ (.B1(_03310_),
    .Y(_00981_),
    .A1(net4700),
    .A2(_03309_));
 sg13g2_nand2_1 _18577_ (.Y(_03311_),
    .A(net1660),
    .B(net4752));
 sg13g2_nand2_1 _18578_ (.Y(_03312_),
    .A(net1858),
    .B(net4707));
 sg13g2_o21ai_1 _18579_ (.B1(_03312_),
    .Y(_00982_),
    .A1(net4708),
    .A2(_03311_));
 sg13g2_nand2_1 _18580_ (.Y(_03313_),
    .A(net1669),
    .B(net4752));
 sg13g2_nand2_1 _18581_ (.Y(_03314_),
    .A(net1715),
    .B(net4707));
 sg13g2_o21ai_1 _18582_ (.B1(_03314_),
    .Y(_00983_),
    .A1(net4707),
    .A2(_03313_));
 sg13g2_nand2_1 _18583_ (.Y(_03315_),
    .A(\fpga_top.qspi_if.word_data[23] ),
    .B(net4753));
 sg13g2_nand2_1 _18584_ (.Y(_03316_),
    .A(net1683),
    .B(net4704));
 sg13g2_o21ai_1 _18585_ (.B1(_03316_),
    .Y(_00984_),
    .A1(net4709),
    .A2(_03315_));
 sg13g2_nand2_1 _18586_ (.Y(_03317_),
    .A(\fpga_top.qspi_if.word_data[24] ),
    .B(net4750));
 sg13g2_nand2_1 _18587_ (.Y(_03318_),
    .A(net1497),
    .B(net4700));
 sg13g2_o21ai_1 _18588_ (.B1(_03318_),
    .Y(_00985_),
    .A1(net4700),
    .A2(_03317_));
 sg13g2_nand2_1 _18589_ (.Y(_03319_),
    .A(\fpga_top.qspi_if.word_data[25] ),
    .B(net4752));
 sg13g2_nand2_1 _18590_ (.Y(_03320_),
    .A(net1615),
    .B(net4707));
 sg13g2_o21ai_1 _18591_ (.B1(_03320_),
    .Y(_00986_),
    .A1(net4707),
    .A2(_03319_));
 sg13g2_nand2_1 _18592_ (.Y(_03321_),
    .A(\fpga_top.qspi_if.word_data[26] ),
    .B(net4752));
 sg13g2_nand2_1 _18593_ (.Y(_03322_),
    .A(net1442),
    .B(net4708));
 sg13g2_o21ai_1 _18594_ (.B1(_03322_),
    .Y(_00987_),
    .A1(net4708),
    .A2(_03321_));
 sg13g2_nand2_1 _18595_ (.Y(_03323_),
    .A(\fpga_top.qspi_if.word_data[27] ),
    .B(net4750));
 sg13g2_nand2_1 _18596_ (.Y(_03324_),
    .A(net1402),
    .B(net4702));
 sg13g2_o21ai_1 _18597_ (.B1(_03324_),
    .Y(_00988_),
    .A1(net4702),
    .A2(_03323_));
 sg13g2_nand2_1 _18598_ (.Y(_03325_),
    .A(net1597),
    .B(_03241_));
 sg13g2_nand2b_1 _18599_ (.Y(_03326_),
    .B(_03243_),
    .A_N(_09902_));
 sg13g2_o21ai_1 _18600_ (.B1(_03325_),
    .Y(_00989_),
    .A1(_03241_),
    .A2(_03326_));
 sg13g2_nand2_1 _18601_ (.Y(_03327_),
    .A(net1633),
    .B(_03241_));
 sg13g2_nand2b_1 _18602_ (.Y(_03328_),
    .B(_03243_),
    .A_N(_09978_));
 sg13g2_o21ai_1 _18603_ (.B1(_03327_),
    .Y(_00990_),
    .A1(_03241_),
    .A2(_03328_));
 sg13g2_nand2_1 _18604_ (.Y(_03329_),
    .A(net5616),
    .B(net5622));
 sg13g2_o21ai_1 _18605_ (.B1(_03329_),
    .Y(_03330_),
    .A1(net5622),
    .A2(_06665_));
 sg13g2_a21oi_1 _18606_ (.A1(net4941),
    .A2(_03330_),
    .Y(_03331_),
    .B1(net4535));
 sg13g2_a22oi_1 _18607_ (.Y(_03332_),
    .B1(_03200_),
    .B2(_08159_),
    .A2(net4557),
    .A1(net6295));
 sg13g2_a21oi_1 _18608_ (.A1(\fpga_top.bus_gather.i_read_adr[2] ),
    .A2(net5167),
    .Y(_03333_),
    .B1(net4568));
 sg13g2_o21ai_1 _18609_ (.B1(_03333_),
    .Y(_03334_),
    .A1(_08158_),
    .A2(net5168));
 sg13g2_o21ai_1 _18610_ (.B1(_03334_),
    .Y(_03335_),
    .A1(net5616),
    .A2(_09548_));
 sg13g2_a22oi_1 _18611_ (.Y(_00991_),
    .B1(_03335_),
    .B2(net4535),
    .A2(_03332_),
    .A1(_03331_));
 sg13g2_nand2_1 _18612_ (.Y(_03336_),
    .A(net5615),
    .B(net5624));
 sg13g2_o21ai_1 _18613_ (.B1(_03336_),
    .Y(_03337_),
    .A1(net5622),
    .A2(_06666_));
 sg13g2_a21oi_1 _18614_ (.A1(net4941),
    .A2(_03337_),
    .Y(_03338_),
    .B1(net4535));
 sg13g2_a22oi_1 _18615_ (.Y(_03339_),
    .B1(_03200_),
    .B2(_08192_),
    .A2(net4553),
    .A1(net6248));
 sg13g2_nor2_1 _18616_ (.A(_08191_),
    .B(net5168),
    .Y(_03340_));
 sg13g2_a21oi_1 _18617_ (.A1(\fpga_top.bus_gather.i_read_adr[3] ),
    .A2(net5167),
    .Y(_03341_),
    .B1(_03340_));
 sg13g2_nor2_1 _18618_ (.A(net4569),
    .B(_03341_),
    .Y(_03342_));
 sg13g2_a21oi_1 _18619_ (.A1(net5615),
    .A2(net4569),
    .Y(_03343_),
    .B1(_03342_));
 sg13g2_a22oi_1 _18620_ (.Y(_00992_),
    .B1(_03343_),
    .B2(net4535),
    .A2(_03339_),
    .A1(_03338_));
 sg13g2_mux2_1 _18621_ (.A0(\fpga_top.cpu_top.csr_wadr_mon[2] ),
    .A1(\fpga_top.bus_gather.u_read_adr[4] ),
    .S(net5623),
    .X(_03344_));
 sg13g2_a22oi_1 _18622_ (.Y(_03345_),
    .B1(_03344_),
    .B2(net4941),
    .A2(net4553),
    .A1(net6277));
 sg13g2_a21oi_1 _18623_ (.A1(_08222_),
    .A2(net4547),
    .Y(_03346_),
    .B1(net4533));
 sg13g2_nand2_1 _18624_ (.Y(_03347_),
    .A(_08222_),
    .B(net5163));
 sg13g2_nand2_1 _18625_ (.Y(_03348_),
    .A(net5597),
    .B(net5168));
 sg13g2_a21oi_1 _18626_ (.A1(_03347_),
    .A2(_03348_),
    .Y(_03349_),
    .B1(net4569));
 sg13g2_a21oi_1 _18627_ (.A1(\fpga_top.bus_gather.u_read_adr[4] ),
    .A2(net4569),
    .Y(_03350_),
    .B1(_03349_));
 sg13g2_a22oi_1 _18628_ (.Y(_00993_),
    .B1(_03350_),
    .B2(net4535),
    .A2(_03346_),
    .A1(_03345_));
 sg13g2_nand2b_1 _18629_ (.Y(_03351_),
    .B(net4549),
    .A_N(_08101_));
 sg13g2_mux2_1 _18630_ (.A0(\fpga_top.cpu_top.csr_wadr_mon[3] ),
    .A1(\fpga_top.bus_gather.u_read_adr[5] ),
    .S(net5622),
    .X(_03352_));
 sg13g2_a221oi_1 _18631_ (.B2(net4939),
    .C1(net4529),
    .B1(_03352_),
    .A1(net6453),
    .Y(_03353_),
    .A2(net4554));
 sg13g2_nor2_1 _18632_ (.A(_08101_),
    .B(net5168),
    .Y(_03354_));
 sg13g2_a21oi_1 _18633_ (.A1(\fpga_top.bus_gather.i_read_adr[5] ),
    .A2(net5165),
    .Y(_03355_),
    .B1(_03354_));
 sg13g2_nor2_1 _18634_ (.A(net4564),
    .B(_03355_),
    .Y(_03356_));
 sg13g2_a21oi_1 _18635_ (.A1(net6303),
    .A2(net4569),
    .Y(_03357_),
    .B1(_03356_));
 sg13g2_a22oi_1 _18636_ (.Y(_00994_),
    .B1(_03357_),
    .B2(net4529),
    .A2(_03353_),
    .A1(_03351_));
 sg13g2_nand2b_1 _18637_ (.Y(_03358_),
    .B(net4547),
    .A_N(_08247_));
 sg13g2_nand2_1 _18638_ (.Y(_03359_),
    .A(net6315),
    .B(net5623));
 sg13g2_o21ai_1 _18639_ (.B1(_03359_),
    .Y(_03360_),
    .A1(net5622),
    .A2(_06667_));
 sg13g2_a221oi_1 _18640_ (.B2(net4939),
    .C1(net4533),
    .B1(_03360_),
    .A1(net6443),
    .Y(_03361_),
    .A2(net4553));
 sg13g2_nor2_1 _18641_ (.A(_08247_),
    .B(net5165),
    .Y(_03362_));
 sg13g2_a21oi_1 _18642_ (.A1(net5596),
    .A2(net5167),
    .Y(_03363_),
    .B1(_03362_));
 sg13g2_nor2_1 _18643_ (.A(net4564),
    .B(_03363_),
    .Y(_03364_));
 sg13g2_a21oi_1 _18644_ (.A1(net6315),
    .A2(net4564),
    .Y(_03365_),
    .B1(_03364_));
 sg13g2_a22oi_1 _18645_ (.Y(_00995_),
    .B1(_03365_),
    .B2(net4533),
    .A2(_03361_),
    .A1(_03358_));
 sg13g2_nand2b_1 _18646_ (.Y(_03366_),
    .B(net4547),
    .A_N(_08073_));
 sg13g2_nand2_1 _18647_ (.Y(_03367_),
    .A(net6149),
    .B(net5622));
 sg13g2_o21ai_1 _18648_ (.B1(_03367_),
    .Y(_03368_),
    .A1(net5622),
    .A2(_06668_));
 sg13g2_a221oi_1 _18649_ (.B2(net4940),
    .C1(net4529),
    .B1(_03368_),
    .A1(net6267),
    .Y(_03369_),
    .A2(net4554));
 sg13g2_nor2_1 _18650_ (.A(_08073_),
    .B(net5165),
    .Y(_03370_));
 sg13g2_a21oi_1 _18651_ (.A1(\fpga_top.bus_gather.i_read_adr[7] ),
    .A2(net5165),
    .Y(_03371_),
    .B1(_03370_));
 sg13g2_nor2_1 _18652_ (.A(net4564),
    .B(_03371_),
    .Y(_03372_));
 sg13g2_a21oi_1 _18653_ (.A1(net6149),
    .A2(net4564),
    .Y(_03373_),
    .B1(_03372_));
 sg13g2_a22oi_1 _18654_ (.Y(_00996_),
    .B1(_03373_),
    .B2(net4533),
    .A2(_03369_),
    .A1(_03366_));
 sg13g2_mux2_1 _18655_ (.A0(\fpga_top.cpu_top.csr_wadr_mon[6] ),
    .A1(net6364),
    .S(net5623),
    .X(_03374_));
 sg13g2_a22oi_1 _18656_ (.Y(_03375_),
    .B1(_03374_),
    .B2(net4940),
    .A2(net4553),
    .A1(net6412));
 sg13g2_a21oi_1 _18657_ (.A1(_08129_),
    .A2(net4547),
    .Y(_03376_),
    .B1(net4533));
 sg13g2_nor2_1 _18658_ (.A(_08128_),
    .B(net5167),
    .Y(_03377_));
 sg13g2_a21oi_1 _18659_ (.A1(net5595),
    .A2(net5167),
    .Y(_03378_),
    .B1(_03377_));
 sg13g2_nor2_1 _18660_ (.A(net4564),
    .B(_03378_),
    .Y(_03379_));
 sg13g2_a21oi_1 _18661_ (.A1(net6364),
    .A2(net4564),
    .Y(_03380_),
    .B1(_03379_));
 sg13g2_a22oi_1 _18662_ (.Y(_00997_),
    .B1(_03380_),
    .B2(net4534),
    .A2(_03376_),
    .A1(_03375_));
 sg13g2_nor2_1 _18663_ (.A(_08313_),
    .B(net4543),
    .Y(_03381_));
 sg13g2_mux2_1 _18664_ (.A0(\fpga_top.cpu_top.csr_wadr_mon[7] ),
    .A1(net6119),
    .S(net5622),
    .X(_03382_));
 sg13g2_a21oi_1 _18665_ (.A1(net4940),
    .A2(_03382_),
    .Y(_03383_),
    .B1(net4529));
 sg13g2_a21oi_1 _18666_ (.A1(net6253),
    .A2(net4554),
    .Y(_03384_),
    .B1(_03381_));
 sg13g2_a21oi_1 _18667_ (.A1(\fpga_top.bus_gather.i_read_adr[9] ),
    .A2(net5165),
    .Y(_03385_),
    .B1(net4564));
 sg13g2_o21ai_1 _18668_ (.B1(_03385_),
    .Y(_03386_),
    .A1(_08313_),
    .A2(net5165));
 sg13g2_o21ai_1 _18669_ (.B1(_03386_),
    .Y(_03387_),
    .A1(net6119),
    .A2(_09548_));
 sg13g2_a22oi_1 _18670_ (.Y(_00998_),
    .B1(_03387_),
    .B2(net4529),
    .A2(_03384_),
    .A1(_03383_));
 sg13g2_nand2b_1 _18671_ (.Y(_03388_),
    .B(net4549),
    .A_N(_08012_));
 sg13g2_mux2_1 _18672_ (.A0(net6433),
    .A1(net6341),
    .S(net5617),
    .X(_03389_));
 sg13g2_a221oi_1 _18673_ (.B2(net4940),
    .C1(net4528),
    .B1(_03389_),
    .A1(net6461),
    .Y(_03390_),
    .A2(net4554));
 sg13g2_a21oi_1 _18674_ (.A1(\fpga_top.bus_gather.i_read_adr[10] ),
    .A2(net5164),
    .Y(_03391_),
    .B1(net4563));
 sg13g2_o21ai_1 _18675_ (.B1(_03391_),
    .Y(_03392_),
    .A1(_08012_),
    .A2(net5164));
 sg13g2_o21ai_1 _18676_ (.B1(_03392_),
    .Y(_03393_),
    .A1(net6341),
    .A2(_09548_));
 sg13g2_a22oi_1 _18677_ (.Y(_00999_),
    .B1(_03393_),
    .B2(net4528),
    .A2(_03390_),
    .A1(_03388_));
 sg13g2_nand2_1 _18678_ (.Y(_03394_),
    .A(_08278_),
    .B(net4548));
 sg13g2_nand2_1 _18679_ (.Y(_03395_),
    .A(net6214),
    .B(net5617));
 sg13g2_o21ai_1 _18680_ (.B1(_03395_),
    .Y(_03396_),
    .A1(net5621),
    .A2(_06669_));
 sg13g2_a221oi_1 _18681_ (.B2(net4939),
    .C1(net4528),
    .B1(_03396_),
    .A1(net6451),
    .Y(_03397_),
    .A2(net4554));
 sg13g2_a21oi_1 _18682_ (.A1(\fpga_top.bus_gather.i_read_adr[11] ),
    .A2(net5164),
    .Y(_03398_),
    .B1(net4565));
 sg13g2_o21ai_1 _18683_ (.B1(_03398_),
    .Y(_03399_),
    .A1(_08279_),
    .A2(net5164));
 sg13g2_o21ai_1 _18684_ (.B1(_03399_),
    .Y(_03400_),
    .A1(net6214),
    .A2(_09548_));
 sg13g2_a22oi_1 _18685_ (.Y(_01000_),
    .B1(_03400_),
    .B2(net4528),
    .A2(_03397_),
    .A1(_03394_));
 sg13g2_nand2_1 _18686_ (.Y(_03401_),
    .A(net3173),
    .B(net4551));
 sg13g2_nand2_1 _18687_ (.Y(_03402_),
    .A(\fpga_top.bus_gather.u_read_adr[12] ),
    .B(net5617));
 sg13g2_o21ai_1 _18688_ (.B1(_03402_),
    .Y(_03403_),
    .A1(net5617),
    .A2(_06670_));
 sg13g2_a221oi_1 _18689_ (.B2(net4939),
    .C1(net4528),
    .B1(_03403_),
    .A1(_08345_),
    .Y(_03404_),
    .A2(net4548));
 sg13g2_nand2b_1 _18690_ (.Y(_03405_),
    .B(net5161),
    .A_N(_08345_));
 sg13g2_a21oi_1 _18691_ (.A1(_06599_),
    .A2(net5164),
    .Y(_03406_),
    .B1(net4563));
 sg13g2_a22oi_1 _18692_ (.Y(_03407_),
    .B1(_03405_),
    .B2(_03406_),
    .A2(net4563),
    .A1(\fpga_top.bus_gather.u_read_adr[12] ));
 sg13g2_a22oi_1 _18693_ (.Y(_01001_),
    .B1(_03407_),
    .B2(net4530),
    .A2(_03404_),
    .A1(_03401_));
 sg13g2_mux2_1 _18694_ (.A0(\fpga_top.cpu_top.csr_wadr_mon[11] ),
    .A1(\fpga_top.bus_gather.u_read_adr[13] ),
    .S(net5621),
    .X(_03408_));
 sg13g2_a22oi_1 _18695_ (.Y(_03409_),
    .B1(net4548),
    .B2(_07970_),
    .A2(net4551),
    .A1(net6130));
 sg13g2_o21ai_1 _18696_ (.B1(_09548_),
    .Y(_03410_),
    .A1(_07970_),
    .A2(net5164));
 sg13g2_a21oi_1 _18697_ (.A1(_06601_),
    .A2(net5164),
    .Y(_03411_),
    .B1(_03410_));
 sg13g2_a21oi_1 _18698_ (.A1(\fpga_top.bus_gather.u_read_adr[13] ),
    .A2(net4563),
    .Y(_03412_),
    .B1(_03411_));
 sg13g2_a21oi_1 _18699_ (.A1(net4939),
    .A2(_03408_),
    .Y(_03413_),
    .B1(net4528));
 sg13g2_a22oi_1 _18700_ (.Y(_01002_),
    .B1(_03413_),
    .B2(_03409_),
    .A2(_03412_),
    .A1(net4528));
 sg13g2_mux2_1 _18701_ (.A0(\fpga_top.dma_io_wadr_u[14] ),
    .A1(net6257),
    .S(net5617),
    .X(_03414_));
 sg13g2_a22oi_1 _18702_ (.Y(_03415_),
    .B1(net4548),
    .B2(_07944_),
    .A2(net4551),
    .A1(net6271));
 sg13g2_nand2b_1 _18703_ (.Y(_03416_),
    .B(net5161),
    .A_N(_07944_));
 sg13g2_a21oi_1 _18704_ (.A1(_06603_),
    .A2(net5164),
    .Y(_03417_),
    .B1(net4567));
 sg13g2_a22oi_1 _18705_ (.Y(_03418_),
    .B1(_03416_),
    .B2(_03417_),
    .A2(net4563),
    .A1(net6257));
 sg13g2_a21oi_1 _18706_ (.A1(net4939),
    .A2(_03414_),
    .Y(_03419_),
    .B1(net4533));
 sg13g2_a22oi_1 _18707_ (.Y(_01003_),
    .B1(_03419_),
    .B2(_03415_),
    .A2(_03418_),
    .A1(net4530));
 sg13g2_nand2b_1 _18708_ (.Y(_03420_),
    .B(net5161),
    .A_N(_08548_));
 sg13g2_a21oi_1 _18709_ (.A1(_06605_),
    .A2(net5166),
    .Y(_03421_),
    .B1(net4567));
 sg13g2_a22oi_1 _18710_ (.Y(_03422_),
    .B1(_03420_),
    .B2(_03421_),
    .A2(net4563),
    .A1(net6224));
 sg13g2_nand2b_1 _18711_ (.Y(_03423_),
    .B(net4546),
    .A_N(_08548_));
 sg13g2_nor2b_1 _18712_ (.A(net5617),
    .B_N(net6365),
    .Y(_03424_));
 sg13g2_a21oi_1 _18713_ (.A1(net6224),
    .A2(net5620),
    .Y(_03425_),
    .B1(_03424_));
 sg13g2_a22oi_1 _18714_ (.Y(_03426_),
    .B1(_03425_),
    .B2(net4940),
    .A2(net4551),
    .A1(_06827_));
 sg13g2_a21oi_1 _18715_ (.A1(_03423_),
    .A2(_03426_),
    .Y(_03427_),
    .B1(net4530));
 sg13g2_a21oi_1 _18716_ (.A1(net4530),
    .A2(_03422_),
    .Y(_01004_),
    .B1(_03427_));
 sg13g2_nand2_1 _18717_ (.Y(_03428_),
    .A(net6231),
    .B(net5620));
 sg13g2_o21ai_1 _18718_ (.B1(_03428_),
    .Y(_03429_),
    .A1(net5620),
    .A2(_06829_));
 sg13g2_a22oi_1 _18719_ (.Y(_03430_),
    .B1(net4547),
    .B2(_08038_),
    .A2(net4552),
    .A1(net6261));
 sg13g2_nand2_1 _18720_ (.Y(_03431_),
    .A(_08038_),
    .B(net5162));
 sg13g2_nand2_1 _18721_ (.Y(_03432_),
    .A(net5593),
    .B(net5167));
 sg13g2_a21oi_1 _18722_ (.A1(_03431_),
    .A2(_03432_),
    .Y(_03433_),
    .B1(net4567));
 sg13g2_a21oi_1 _18723_ (.A1(net6231),
    .A2(net4567),
    .Y(_03434_),
    .B1(_03433_));
 sg13g2_a21oi_1 _18724_ (.A1(net4940),
    .A2(_03429_),
    .Y(_03435_),
    .B1(net4532));
 sg13g2_a22oi_1 _18725_ (.Y(_01005_),
    .B1(_03435_),
    .B2(_03430_),
    .A2(_03434_),
    .A1(net4532));
 sg13g2_nor2b_1 _18726_ (.A(net5618),
    .B_N(net6169),
    .Y(_03436_));
 sg13g2_a21oi_1 _18727_ (.A1(net6255),
    .A2(net5618),
    .Y(_03437_),
    .B1(_03436_));
 sg13g2_a22oi_1 _18728_ (.Y(_03438_),
    .B1(net4546),
    .B2(_08377_),
    .A2(net4551),
    .A1(net6566));
 sg13g2_o21ai_1 _18729_ (.B1(_03438_),
    .Y(_03439_),
    .A1(_09559_),
    .A2(_03437_));
 sg13g2_nand2_1 _18730_ (.Y(_03440_),
    .A(_08377_),
    .B(net5161));
 sg13g2_a21oi_1 _18731_ (.A1(\fpga_top.bus_gather.i_read_adr[17] ),
    .A2(net5166),
    .Y(_03441_),
    .B1(net4566));
 sg13g2_a22oi_1 _18732_ (.Y(_03442_),
    .B1(_03440_),
    .B2(_03441_),
    .A2(net4565),
    .A1(_06515_));
 sg13g2_mux2_1 _18733_ (.A0(_03439_),
    .A1(_03442_),
    .S(net4531),
    .X(_01006_));
 sg13g2_mux2_1 _18734_ (.A0(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[18] ),
    .A1(\fpga_top.bus_gather.u_read_adr[18] ),
    .S(net5618),
    .X(_03443_));
 sg13g2_nor2_1 _18735_ (.A(_08526_),
    .B(net4545),
    .Y(_03444_));
 sg13g2_a221oi_1 _18736_ (.B2(net4941),
    .C1(_03444_),
    .B1(_03443_),
    .A1(net6436),
    .Y(_03445_),
    .A2(net4553));
 sg13g2_nand2_1 _18737_ (.Y(_03446_),
    .A(_06529_),
    .B(net4565));
 sg13g2_a21oi_1 _18738_ (.A1(\fpga_top.bus_gather.i_read_adr[18] ),
    .A2(net5166),
    .Y(_03447_),
    .B1(net4566));
 sg13g2_o21ai_1 _18739_ (.B1(_03447_),
    .Y(_03448_),
    .A1(_08526_),
    .A2(net5166));
 sg13g2_nand3_1 _18740_ (.B(_03446_),
    .C(_03448_),
    .A(net4531),
    .Y(_03449_));
 sg13g2_o21ai_1 _18741_ (.B1(_03449_),
    .Y(_01007_),
    .A1(net4534),
    .A2(net6437));
 sg13g2_nor2b_1 _18742_ (.A(net5618),
    .B_N(net6140),
    .Y(_03450_));
 sg13g2_a21oi_1 _18743_ (.A1(net6264),
    .A2(net5618),
    .Y(_03451_),
    .B1(_03450_));
 sg13g2_nor2_1 _18744_ (.A(_09559_),
    .B(_03451_),
    .Y(_03452_));
 sg13g2_a221oi_1 _18745_ (.B2(_08405_),
    .C1(_03452_),
    .B1(net4546),
    .A1(net6448),
    .Y(_03453_),
    .A2(net4552));
 sg13g2_nand2_1 _18746_ (.Y(_03454_),
    .A(_08405_),
    .B(net5162));
 sg13g2_a21oi_1 _18747_ (.A1(\fpga_top.bus_gather.i_read_adr[19] ),
    .A2(net5166),
    .Y(_03455_),
    .B1(net4566));
 sg13g2_a22oi_1 _18748_ (.Y(_03456_),
    .B1(_03454_),
    .B2(_03455_),
    .A2(net4565),
    .A1(_06527_));
 sg13g2_nand2_1 _18749_ (.Y(_03457_),
    .A(net4531),
    .B(_03456_));
 sg13g2_o21ai_1 _18750_ (.B1(_03457_),
    .Y(_01008_),
    .A1(net4532),
    .A2(_03453_));
 sg13g2_mux2_1 _18751_ (.A0(net6186),
    .A1(\fpga_top.bus_gather.u_read_adr[20] ),
    .S(net5619),
    .X(_03458_));
 sg13g2_a21oi_1 _18752_ (.A1(net4941),
    .A2(_03458_),
    .Y(_03459_),
    .B1(net4531));
 sg13g2_a22oi_1 _18753_ (.Y(_03460_),
    .B1(net4546),
    .B2(_08428_),
    .A2(net4552),
    .A1(net6397));
 sg13g2_nand2_1 _18754_ (.Y(_03461_),
    .A(_08427_),
    .B(net5162));
 sg13g2_a21oi_1 _18755_ (.A1(_06620_),
    .A2(net5167),
    .Y(_03462_),
    .B1(net4566));
 sg13g2_a22oi_1 _18756_ (.Y(_03463_),
    .B1(_03461_),
    .B2(_03462_),
    .A2(net4566),
    .A1(net6291));
 sg13g2_a22oi_1 _18757_ (.Y(_01009_),
    .B1(_03463_),
    .B2(net4532),
    .A2(_03460_),
    .A1(_03459_));
 sg13g2_nor2b_1 _18758_ (.A(net5618),
    .B_N(net6115),
    .Y(_03464_));
 sg13g2_a21oi_1 _18759_ (.A1(\fpga_top.bus_gather.u_read_adr[21] ),
    .A2(net5618),
    .Y(_03465_),
    .B1(_03464_));
 sg13g2_nor2_1 _18760_ (.A(_09559_),
    .B(_03465_),
    .Y(_03466_));
 sg13g2_a221oi_1 _18761_ (.B2(_07867_),
    .C1(_03466_),
    .B1(net4546),
    .A1(net6500),
    .Y(_03467_),
    .A2(net4552));
 sg13g2_nand2_1 _18762_ (.Y(_03468_),
    .A(_07867_),
    .B(net5161));
 sg13g2_a21oi_1 _18763_ (.A1(\fpga_top.bus_gather.i_read_adr[21] ),
    .A2(net5166),
    .Y(_03469_),
    .B1(net4566));
 sg13g2_a22oi_1 _18764_ (.Y(_03470_),
    .B1(_03468_),
    .B2(_03469_),
    .A2(net4566),
    .A1(_06525_));
 sg13g2_nand2_1 _18765_ (.Y(_03471_),
    .A(net4531),
    .B(_03470_));
 sg13g2_o21ai_1 _18766_ (.B1(_03471_),
    .Y(_01010_),
    .A1(net4531),
    .A2(net6501));
 sg13g2_nand2b_1 _18767_ (.Y(_03472_),
    .B(net4546),
    .A_N(_07837_));
 sg13g2_mux2_1 _18768_ (.A0(net6108),
    .A1(net6494),
    .S(net5618),
    .X(_03473_));
 sg13g2_a221oi_1 _18769_ (.B2(net4940),
    .C1(net4531),
    .B1(_03473_),
    .A1(net6485),
    .Y(_03474_),
    .A2(net4552));
 sg13g2_nand2b_1 _18770_ (.Y(_03475_),
    .B(net5166),
    .A_N(net5591));
 sg13g2_a21oi_1 _18771_ (.A1(_07837_),
    .A2(net5161),
    .Y(_03476_),
    .B1(net4565));
 sg13g2_a22oi_1 _18772_ (.Y(_03477_),
    .B1(_03475_),
    .B2(_03476_),
    .A2(net4565),
    .A1(net6233));
 sg13g2_a22oi_1 _18773_ (.Y(_01011_),
    .B1(_03477_),
    .B2(net4531),
    .A2(_03474_),
    .A1(_03472_));
 sg13g2_nor2b_1 _18774_ (.A(net5619),
    .B_N(net6082),
    .Y(_03478_));
 sg13g2_a21oi_1 _18775_ (.A1(net3901),
    .A2(net5619),
    .Y(_03479_),
    .B1(_03478_));
 sg13g2_a22oi_1 _18776_ (.Y(_03480_),
    .B1(net4546),
    .B2(_08475_),
    .A2(net4551),
    .A1(net6513));
 sg13g2_o21ai_1 _18777_ (.B1(_03480_),
    .Y(_03481_),
    .A1(_09559_),
    .A2(_03479_));
 sg13g2_nand2_1 _18778_ (.Y(_03482_),
    .A(_08475_),
    .B(net5161));
 sg13g2_a21oi_1 _18779_ (.A1(\fpga_top.bus_gather.i_read_adr[23] ),
    .A2(net5166),
    .Y(_03483_),
    .B1(net4566));
 sg13g2_a22oi_1 _18780_ (.Y(_03484_),
    .B1(_03482_),
    .B2(_03483_),
    .A2(net4563),
    .A1(_06532_));
 sg13g2_mux2_1 _18781_ (.A0(_03481_),
    .A1(_03484_),
    .S(net4530),
    .X(_01012_));
 sg13g2_a21oi_1 _18782_ (.A1(_07907_),
    .A2(net5162),
    .Y(_03485_),
    .B1(net4565));
 sg13g2_o21ai_1 _18783_ (.B1(_03485_),
    .Y(_03486_),
    .A1(_06629_),
    .A2(net5162));
 sg13g2_o21ai_1 _18784_ (.B1(_03486_),
    .Y(_03487_),
    .A1(net6319),
    .A2(_09548_));
 sg13g2_nand2_1 _18785_ (.Y(_03488_),
    .A(_07907_),
    .B(net4546));
 sg13g2_mux2_1 _18786_ (.A0(net6162),
    .A1(net6319),
    .S(net5617),
    .X(_03489_));
 sg13g2_a221oi_1 _18787_ (.B2(net4939),
    .C1(net4528),
    .B1(_03489_),
    .A1(net6529),
    .Y(_03490_),
    .A2(net4551));
 sg13g2_a22oi_1 _18788_ (.Y(_01013_),
    .B1(_03488_),
    .B2(_03490_),
    .A2(_03487_),
    .A1(net4530));
 sg13g2_mux2_1 _18789_ (.A0(net6213),
    .A1(net6239),
    .S(net5617),
    .X(_03491_));
 sg13g2_a21oi_1 _18790_ (.A1(net4939),
    .A2(_03491_),
    .Y(_03492_),
    .B1(net4530));
 sg13g2_a22oi_1 _18791_ (.Y(_03493_),
    .B1(net4548),
    .B2(_08500_),
    .A2(net4551),
    .A1(net6262));
 sg13g2_nand2b_1 _18792_ (.Y(_03494_),
    .B(net5161),
    .A_N(_08500_));
 sg13g2_a21oi_1 _18793_ (.A1(_06631_),
    .A2(net5165),
    .Y(_03495_),
    .B1(net4565));
 sg13g2_a22oi_1 _18794_ (.Y(_03496_),
    .B1(_03494_),
    .B2(_03495_),
    .A2(net4563),
    .A1(net6239));
 sg13g2_a22oi_1 _18795_ (.Y(_01014_),
    .B1(_03496_),
    .B2(net4530),
    .A2(_03493_),
    .A1(_03492_));
 sg13g2_nor2_1 _18796_ (.A(net3944),
    .B(_08726_),
    .Y(_03497_));
 sg13g2_a21oi_1 _18797_ (.A1(_03267_),
    .A2(_03497_),
    .Y(_03498_),
    .B1(_03250_));
 sg13g2_o21ai_1 _18798_ (.B1(_03498_),
    .Y(_01015_),
    .A1(_06545_),
    .A2(_03267_));
 sg13g2_xnor2_1 _18799_ (.Y(_03499_),
    .A(\fpga_top.qspi_if.read_cntr[0] ),
    .B(net3911));
 sg13g2_nand4_1 _18800_ (.B(net4755),
    .C(_03267_),
    .A(_08727_),
    .Y(_03500_),
    .D(_03499_));
 sg13g2_nor2_1 _18801_ (.A(_03250_),
    .B(_03267_),
    .Y(_03501_));
 sg13g2_o21ai_1 _18802_ (.B1(_03500_),
    .Y(_03502_),
    .A1(net5331),
    .A2(net4755));
 sg13g2_a21o_1 _18803_ (.A2(_03501_),
    .A1(net3911),
    .B1(_03502_),
    .X(_01016_));
 sg13g2_o21ai_1 _18804_ (.B1(net4067),
    .Y(_03503_),
    .A1(net3944),
    .A2(net3911));
 sg13g2_nand2_1 _18805_ (.Y(_03504_),
    .A(net1489),
    .B(net4755));
 sg13g2_nand2_1 _18806_ (.Y(_03505_),
    .A(net1489),
    .B(_08725_));
 sg13g2_nand2_1 _18807_ (.Y(_03506_),
    .A(_03503_),
    .B(_03505_));
 sg13g2_nand3_1 _18808_ (.B(_03267_),
    .C(_03506_),
    .A(net4755),
    .Y(_03507_));
 sg13g2_a22oi_1 _18809_ (.Y(_03508_),
    .B1(_03501_),
    .B2(net4067),
    .A2(_03250_),
    .A1(net5709));
 sg13g2_nand2_1 _18810_ (.Y(_01017_),
    .A(_03507_),
    .B(net4068));
 sg13g2_a21oi_1 _18811_ (.A1(_08725_),
    .A2(_03267_),
    .Y(_01018_),
    .B1(_03504_));
 sg13g2_nor3_1 _18812_ (.A(net6247),
    .B(net5352),
    .C(_08862_),
    .Y(_03509_));
 sg13g2_a21oi_1 _18813_ (.A1(net6247),
    .A2(net5352),
    .Y(_03510_),
    .B1(_03509_));
 sg13g2_nor3_2 _18814_ (.A(net3762),
    .B(_09094_),
    .C(_03247_),
    .Y(_03511_));
 sg13g2_nor2_2 _18815_ (.A(_06947_),
    .B(_06949_),
    .Y(_03512_));
 sg13g2_nand2_1 _18816_ (.Y(_03513_),
    .A(net3913),
    .B(_03512_));
 sg13g2_a22oi_1 _18817_ (.Y(_03514_),
    .B1(_06949_),
    .B2(net3832),
    .A2(_06947_),
    .A1(net3888));
 sg13g2_nand2_1 _18818_ (.Y(_03515_),
    .A(_03513_),
    .B(_03514_));
 sg13g2_nand2_1 _18819_ (.Y(_03516_),
    .A(_03511_),
    .B(_03515_));
 sg13g2_o21ai_1 _18820_ (.B1(_03516_),
    .Y(_01019_),
    .A1(_03510_),
    .A2(_03511_));
 sg13g2_nor2_1 _18821_ (.A(net5355),
    .B(_03511_),
    .Y(_03517_));
 sg13g2_xor2_1 _18822_ (.B(net6351),
    .A(net6247),
    .X(_03518_));
 sg13g2_nor4_1 _18823_ (.A(net5352),
    .B(_08862_),
    .C(_03511_),
    .D(_03518_),
    .Y(_03519_));
 sg13g2_nand2_1 _18824_ (.Y(_03520_),
    .A(net3750),
    .B(_03512_));
 sg13g2_a22oi_1 _18825_ (.Y(_03521_),
    .B1(_06949_),
    .B2(net3818),
    .A2(_06947_),
    .A1(net3961));
 sg13g2_nand2_1 _18826_ (.Y(_03522_),
    .A(_03520_),
    .B(_03521_));
 sg13g2_a221oi_1 _18827_ (.B2(_03511_),
    .C1(_03519_),
    .B1(_03522_),
    .A1(net6351),
    .Y(_03523_),
    .A2(_03517_));
 sg13g2_inv_1 _18828_ (.Y(_01020_),
    .A(_03523_));
 sg13g2_o21ai_1 _18829_ (.B1(net6473),
    .Y(_03524_),
    .A1(net5352),
    .A2(_08860_));
 sg13g2_nand2_1 _18830_ (.Y(_03525_),
    .A(net2398),
    .B(net5355));
 sg13g2_o21ai_1 _18831_ (.B1(net6474),
    .Y(_03526_),
    .A1(_08861_),
    .A2(_03525_));
 sg13g2_nand2_1 _18832_ (.Y(_03527_),
    .A(net3742),
    .B(_03512_));
 sg13g2_a22oi_1 _18833_ (.Y(_03528_),
    .B1(_06949_),
    .B2(net3819),
    .A2(_06947_),
    .A1(net3947));
 sg13g2_nand2_1 _18834_ (.Y(_03529_),
    .A(_03527_),
    .B(_03528_));
 sg13g2_mux2_1 _18835_ (.A0(_03526_),
    .A1(_03529_),
    .S(_03511_),
    .X(_01021_));
 sg13g2_nand2_1 _18836_ (.Y(_03530_),
    .A(net2398),
    .B(_03517_));
 sg13g2_nand2b_1 _18837_ (.Y(_03531_),
    .B(_08861_),
    .A_N(_03525_));
 sg13g2_nand2_1 _18838_ (.Y(_03532_),
    .A(\fpga_top.qspi_if.read_latency_0[3] ),
    .B(_03512_));
 sg13g2_a22oi_1 _18839_ (.Y(_03533_),
    .B1(_06949_),
    .B2(\fpga_top.qspi_if.read_latency_1[3] ),
    .A2(_06947_),
    .A1(\fpga_top.qspi_if.read_latency_2[3] ));
 sg13g2_and3_1 _18840_ (.X(_03534_),
    .A(_03511_),
    .B(_03532_),
    .C(_03533_));
 sg13g2_nor2b_1 _18841_ (.A(_03511_),
    .B_N(_03531_),
    .Y(_03535_));
 sg13g2_o21ai_1 _18842_ (.B1(_03530_),
    .Y(_01022_),
    .A1(_03534_),
    .A2(_03535_));
 sg13g2_nand3b_1 _18843_ (.B(_08909_),
    .C(_08900_),
    .Y(_03536_),
    .A_N(_08901_));
 sg13g2_nand2_2 _18844_ (.Y(_03537_),
    .A(_08891_),
    .B(_09616_));
 sg13g2_nand2_2 _18845_ (.Y(_03538_),
    .A(_08891_),
    .B(_10521_));
 sg13g2_nor3_2 _18846_ (.A(_02733_),
    .B(_03536_),
    .C(_03538_),
    .Y(_03539_));
 sg13g2_nor2_1 _18847_ (.A(net3600),
    .B(_03539_),
    .Y(_03540_));
 sg13g2_a21oi_1 _18848_ (.A1(net4919),
    .A2(_03539_),
    .Y(_01023_),
    .B1(_03540_));
 sg13g2_nor2_1 _18849_ (.A(net3500),
    .B(net4441),
    .Y(_03541_));
 sg13g2_a21oi_1 _18850_ (.A1(net4845),
    .A2(net4441),
    .Y(_01024_),
    .B1(_03541_));
 sg13g2_nor2_1 _18851_ (.A(net6099),
    .B(net4441),
    .Y(_03542_));
 sg13g2_a21oi_1 _18852_ (.A1(net4850),
    .A2(_03539_),
    .Y(_01025_),
    .B1(_03542_));
 sg13g2_mux2_1 _18853_ (.A0(net6323),
    .A1(net4838),
    .S(net4441),
    .X(_01026_));
 sg13g2_nor2_1 _18854_ (.A(net3849),
    .B(net4441),
    .Y(_03543_));
 sg13g2_a21oi_1 _18855_ (.A1(net4834),
    .A2(net4441),
    .Y(_01027_),
    .B1(_03543_));
 sg13g2_nor2_1 _18856_ (.A(net3347),
    .B(net4441),
    .Y(_03544_));
 sg13g2_a21oi_1 _18857_ (.A1(net4833),
    .A2(net4441),
    .Y(_01028_),
    .B1(_03544_));
 sg13g2_or3_1 _18858_ (.A(_08898_),
    .B(_03536_),
    .C(net4466),
    .X(_03545_));
 sg13g2_and2_1 _18859_ (.A(net5599),
    .B(_03545_),
    .X(_03546_));
 sg13g2_nand2b_1 _18860_ (.Y(_03547_),
    .B(net3),
    .A_N(net5600));
 sg13g2_o21ai_1 _18861_ (.B1(_03547_),
    .Y(_03548_),
    .A1(_02999_),
    .A2(_03545_));
 sg13g2_a21o_1 _18862_ (.A2(_03546_),
    .A1(net3772),
    .B1(_03548_),
    .X(_01029_));
 sg13g2_o21ai_1 _18863_ (.B1(_03547_),
    .Y(_03549_),
    .A1(_03002_),
    .A2(_03545_));
 sg13g2_a21o_1 _18864_ (.A2(_03546_),
    .A1(net3813),
    .B1(_03549_),
    .X(_01030_));
 sg13g2_nand2_1 _18865_ (.Y(_03550_),
    .A(net3661),
    .B(_03546_));
 sg13g2_nand2_1 _18866_ (.Y(_03551_),
    .A(net5599),
    .B(_08915_));
 sg13g2_o21ai_1 _18867_ (.B1(_03550_),
    .Y(_01031_),
    .A1(_03545_),
    .A2(_03551_));
 sg13g2_nand2_1 _18868_ (.Y(_03552_),
    .A(net3708),
    .B(_03546_));
 sg13g2_o21ai_1 _18869_ (.B1(_03552_),
    .Y(_01032_),
    .A1(_03008_),
    .A2(_03545_));
 sg13g2_nand2_1 _18870_ (.Y(_03553_),
    .A(net5688),
    .B(_03546_));
 sg13g2_o21ai_1 _18871_ (.B1(_03553_),
    .Y(_01033_),
    .A1(_03012_),
    .A2(_03545_));
 sg13g2_nand2_1 _18872_ (.Y(_03554_),
    .A(net2357),
    .B(_03546_));
 sg13g2_o21ai_1 _18873_ (.B1(_03554_),
    .Y(_01034_),
    .A1(_03015_),
    .A2(_03545_));
 sg13g2_nor2_1 _18874_ (.A(_08910_),
    .B(net4466),
    .Y(_03555_));
 sg13g2_nor3_2 _18875_ (.A(_08910_),
    .B(_08983_),
    .C(net4466),
    .Y(_03556_));
 sg13g2_nor2_1 _18876_ (.A(net3933),
    .B(net4440),
    .Y(_03557_));
 sg13g2_a21oi_1 _18877_ (.A1(net4919),
    .A2(net4440),
    .Y(_01035_),
    .B1(_03557_));
 sg13g2_nor2_1 _18878_ (.A(net3751),
    .B(net4439),
    .Y(_03558_));
 sg13g2_a21oi_1 _18879_ (.A1(net4917),
    .A2(net4439),
    .Y(_01036_),
    .B1(_03558_));
 sg13g2_nor2_1 _18880_ (.A(net3701),
    .B(net4440),
    .Y(_03559_));
 sg13g2_a21oi_1 _18881_ (.A1(net4849),
    .A2(net4440),
    .Y(_01037_),
    .B1(_03559_));
 sg13g2_nor2_1 _18882_ (.A(net3678),
    .B(net4440),
    .Y(_03560_));
 sg13g2_a21oi_1 _18883_ (.A1(net4843),
    .A2(net4440),
    .Y(_01038_),
    .B1(_03560_));
 sg13g2_nor2_1 _18884_ (.A(net3715),
    .B(net4439),
    .Y(_03561_));
 sg13g2_a21oi_1 _18885_ (.A1(net4838),
    .A2(net4439),
    .Y(_01039_),
    .B1(_03561_));
 sg13g2_nor2_1 _18886_ (.A(net3683),
    .B(net4440),
    .Y(_03562_));
 sg13g2_a21oi_1 _18887_ (.A1(net4834),
    .A2(net4440),
    .Y(_01040_),
    .B1(_03562_));
 sg13g2_nor2_1 _18888_ (.A(net3795),
    .B(net4439),
    .Y(_03563_));
 sg13g2_a21oi_1 _18889_ (.A1(net4833),
    .A2(net4439),
    .Y(_01041_),
    .B1(_03563_));
 sg13g2_nor2_1 _18890_ (.A(net3492),
    .B(net4439),
    .Y(_03564_));
 sg13g2_a21oi_1 _18891_ (.A1(net4831),
    .A2(net4439),
    .Y(_01042_),
    .B1(_03564_));
 sg13g2_nor2_1 _18892_ (.A(_06661_),
    .B(net5354),
    .Y(_03565_));
 sg13g2_nand2_1 _18893_ (.Y(_03566_),
    .A(net5683),
    .B(_08854_));
 sg13g2_o21ai_1 _18894_ (.B1(_03566_),
    .Y(_01043_),
    .A1(net5683),
    .A2(_03565_));
 sg13g2_nand3b_1 _18895_ (.B(_09106_),
    .C(net5629),
    .Y(_03567_),
    .A_N(_08851_));
 sg13g2_o21ai_1 _18896_ (.B1(_08854_),
    .Y(_03568_),
    .A1(net5629),
    .A2(net5331));
 sg13g2_a22oi_1 _18897_ (.Y(_03569_),
    .B1(_03567_),
    .B2(_03568_),
    .A2(_03565_),
    .A1(net6195));
 sg13g2_inv_1 _18898_ (.Y(_01044_),
    .A(net6196));
 sg13g2_a21oi_1 _18899_ (.A1(net5354),
    .A2(_08851_),
    .Y(_03570_),
    .B1(_06661_));
 sg13g2_a22oi_1 _18900_ (.Y(_03571_),
    .B1(_03570_),
    .B2(net5682),
    .A2(net5699),
    .A1(_06661_));
 sg13g2_nand2_1 _18901_ (.Y(_01045_),
    .A(_08856_),
    .B(net6546));
 sg13g2_and2_1 _18902_ (.A(_10552_),
    .B(_03555_),
    .X(_03572_));
 sg13g2_nor2_1 _18903_ (.A(net3703),
    .B(net4420),
    .Y(_03573_));
 sg13g2_a21oi_1 _18904_ (.A1(net4919),
    .A2(net4419),
    .Y(_01046_),
    .B1(_03573_));
 sg13g2_nor2_1 _18905_ (.A(net3724),
    .B(net4419),
    .Y(_03574_));
 sg13g2_a21oi_1 _18906_ (.A1(net4917),
    .A2(net4420),
    .Y(_01047_),
    .B1(_03574_));
 sg13g2_nor2_1 _18907_ (.A(net3796),
    .B(net4420),
    .Y(_03575_));
 sg13g2_a21oi_1 _18908_ (.A1(net4849),
    .A2(net4420),
    .Y(_01048_),
    .B1(_03575_));
 sg13g2_nor2_1 _18909_ (.A(net3830),
    .B(net4420),
    .Y(_03576_));
 sg13g2_a21oi_1 _18910_ (.A1(net4843),
    .A2(net4420),
    .Y(_01049_),
    .B1(_03576_));
 sg13g2_nor2_1 _18911_ (.A(net3486),
    .B(net4419),
    .Y(_03577_));
 sg13g2_a21oi_1 _18912_ (.A1(net4838),
    .A2(net4419),
    .Y(_01050_),
    .B1(_03577_));
 sg13g2_nor2_1 _18913_ (.A(net3012),
    .B(_03572_),
    .Y(_03578_));
 sg13g2_a21oi_1 _18914_ (.A1(_02752_),
    .A2(net4420),
    .Y(_01051_),
    .B1(_03578_));
 sg13g2_nor2_1 _18915_ (.A(net3764),
    .B(net4419),
    .Y(_03579_));
 sg13g2_a21oi_1 _18916_ (.A1(net4833),
    .A2(net4419),
    .Y(_01052_),
    .B1(_03579_));
 sg13g2_nor2_1 _18917_ (.A(net3712),
    .B(net4419),
    .Y(_03580_));
 sg13g2_a21oi_1 _18918_ (.A1(net4831),
    .A2(net4419),
    .Y(_01053_),
    .B1(_03580_));
 sg13g2_nor3_1 _18919_ (.A(_08910_),
    .B(_02733_),
    .C(net4466),
    .Y(_03581_));
 sg13g2_nor2_1 _18920_ (.A(net3644),
    .B(net4438),
    .Y(_03582_));
 sg13g2_a21oi_1 _18921_ (.A1(_10526_),
    .A2(net4437),
    .Y(_01054_),
    .B1(_03582_));
 sg13g2_nor2_1 _18922_ (.A(net3801),
    .B(net4436),
    .Y(_03583_));
 sg13g2_a21oi_1 _18923_ (.A1(net4845),
    .A2(net4437),
    .Y(_01055_),
    .B1(_03583_));
 sg13g2_nor2_1 _18924_ (.A(net1733),
    .B(net4436),
    .Y(_03584_));
 sg13g2_a21oi_1 _18925_ (.A1(net4850),
    .A2(net4436),
    .Y(_01056_),
    .B1(_03584_));
 sg13g2_nor2_1 _18926_ (.A(net3021),
    .B(net4438),
    .Y(_03585_));
 sg13g2_a21oi_1 _18927_ (.A1(net4843),
    .A2(net4438),
    .Y(_01057_),
    .B1(_03585_));
 sg13g2_mux2_1 _18928_ (.A0(net3891),
    .A1(net4838),
    .S(net4436),
    .X(_01058_));
 sg13g2_nor2_1 _18929_ (.A(net3643),
    .B(net4436),
    .Y(_03586_));
 sg13g2_a21oi_1 _18930_ (.A1(_02752_),
    .A2(net4436),
    .Y(_01059_),
    .B1(_03586_));
 sg13g2_nor2_1 _18931_ (.A(net3825),
    .B(net4437),
    .Y(_03587_));
 sg13g2_a21oi_1 _18932_ (.A1(_02756_),
    .A2(net4437),
    .Y(_01060_),
    .B1(_03587_));
 sg13g2_nor2_1 _18933_ (.A(net3785),
    .B(net4436),
    .Y(_03588_));
 sg13g2_a21oi_1 _18934_ (.A1(net4831),
    .A2(net4436),
    .Y(_01061_),
    .B1(_03588_));
 sg13g2_nor2_1 _18935_ (.A(_08911_),
    .B(net4466),
    .Y(_03589_));
 sg13g2_nor2_1 _18936_ (.A(net3653),
    .B(net4435),
    .Y(_03590_));
 sg13g2_a21oi_1 _18937_ (.A1(_10526_),
    .A2(net4435),
    .Y(_01062_),
    .B1(_03590_));
 sg13g2_nor2_1 _18938_ (.A(net3517),
    .B(net4435),
    .Y(_03591_));
 sg13g2_a21oi_1 _18939_ (.A1(net4845),
    .A2(net4435),
    .Y(_01063_),
    .B1(_03591_));
 sg13g2_nor2_1 _18940_ (.A(net3840),
    .B(net4434),
    .Y(_03592_));
 sg13g2_a21oi_1 _18941_ (.A1(net4850),
    .A2(net4434),
    .Y(_01064_),
    .B1(_03592_));
 sg13g2_nor2_1 _18942_ (.A(net3802),
    .B(net4435),
    .Y(_03593_));
 sg13g2_a21oi_1 _18943_ (.A1(net4843),
    .A2(net4435),
    .Y(_01065_),
    .B1(_03593_));
 sg13g2_mux2_1 _18944_ (.A0(net3910),
    .A1(net4838),
    .S(net4435),
    .X(_01066_));
 sg13g2_nor2_1 _18945_ (.A(net3204),
    .B(net4434),
    .Y(_03594_));
 sg13g2_a21oi_1 _18946_ (.A1(net4834),
    .A2(net4434),
    .Y(_01067_),
    .B1(_03594_));
 sg13g2_nor2_1 _18947_ (.A(net3936),
    .B(net4434),
    .Y(_03595_));
 sg13g2_a21oi_1 _18948_ (.A1(_02756_),
    .A2(net4434),
    .Y(_01068_),
    .B1(_03595_));
 sg13g2_nor2_1 _18949_ (.A(net3905),
    .B(net4434),
    .Y(_03596_));
 sg13g2_a21oi_1 _18950_ (.A1(_02760_),
    .A2(net4434),
    .Y(_01069_),
    .B1(_03596_));
 sg13g2_nor2_1 _18951_ (.A(_02740_),
    .B(net4466),
    .Y(_03597_));
 sg13g2_nor2_1 _18952_ (.A(net3326),
    .B(net4432),
    .Y(_03598_));
 sg13g2_a21oi_1 _18953_ (.A1(_10595_),
    .A2(net4432),
    .Y(_01070_),
    .B1(_03598_));
 sg13g2_nor2_1 _18954_ (.A(net6194),
    .B(net4430),
    .Y(_03599_));
 sg13g2_a21oi_1 _18955_ (.A1(_10600_),
    .A2(net4430),
    .Y(_01071_),
    .B1(_03599_));
 sg13g2_nor2_1 _18956_ (.A(net3773),
    .B(net4430),
    .Y(_03600_));
 sg13g2_a21oi_1 _18957_ (.A1(_10603_),
    .A2(net4431),
    .Y(_01072_),
    .B1(_03600_));
 sg13g2_nor2_1 _18958_ (.A(net3690),
    .B(net4430),
    .Y(_03601_));
 sg13g2_a21oi_1 _18959_ (.A1(_02789_),
    .A2(net4430),
    .Y(_01073_),
    .B1(_03601_));
 sg13g2_nor2_1 _18960_ (.A(net6210),
    .B(net4432),
    .Y(_03602_));
 sg13g2_a21oi_1 _18961_ (.A1(_10605_),
    .A2(net4432),
    .Y(_01074_),
    .B1(_03602_));
 sg13g2_nor2_1 _18962_ (.A(net3681),
    .B(net4430),
    .Y(_03603_));
 sg13g2_a21oi_1 _18963_ (.A1(_10609_),
    .A2(net4430),
    .Y(_01075_),
    .B1(_03603_));
 sg13g2_nor2_1 _18964_ (.A(net3839),
    .B(net4430),
    .Y(_03604_));
 sg13g2_a21oi_1 _18965_ (.A1(_10611_),
    .A2(net4431),
    .Y(_01076_),
    .B1(_03604_));
 sg13g2_nor2_1 _18966_ (.A(net3807),
    .B(net4431),
    .Y(_03605_));
 sg13g2_a21oi_1 _18967_ (.A1(_02795_),
    .A2(net4431),
    .Y(_01077_),
    .B1(_03605_));
 sg13g2_nor2_1 _18968_ (.A(net3697),
    .B(net4427),
    .Y(_03606_));
 sg13g2_a21oi_1 _18969_ (.A1(_10526_),
    .A2(net4428),
    .Y(_01078_),
    .B1(_03606_));
 sg13g2_nor2_1 _18970_ (.A(net3666),
    .B(net4428),
    .Y(_03607_));
 sg13g2_a21oi_1 _18971_ (.A1(net4916),
    .A2(net4428),
    .Y(_01079_),
    .B1(_03607_));
 sg13g2_nor2_1 _18972_ (.A(net3147),
    .B(net4429),
    .Y(_03608_));
 sg13g2_a21oi_1 _18973_ (.A1(net4850),
    .A2(net4429),
    .Y(_01080_),
    .B1(_03608_));
 sg13g2_nand2_1 _18974_ (.Y(_03609_),
    .A(net4842),
    .B(net4428));
 sg13g2_o21ai_1 _18975_ (.B1(_03609_),
    .Y(_01081_),
    .A1(_06653_),
    .A2(net4428));
 sg13g2_mux2_1 _18976_ (.A0(net3906),
    .A1(net4840),
    .S(net4427),
    .X(_01082_));
 sg13g2_nor2_1 _18977_ (.A(net2126),
    .B(net4427),
    .Y(_03610_));
 sg13g2_a21oi_1 _18978_ (.A1(net4835),
    .A2(net4427),
    .Y(_01083_),
    .B1(_03610_));
 sg13g2_nor2_1 _18979_ (.A(net3614),
    .B(net4427),
    .Y(_03611_));
 sg13g2_a21oi_1 _18980_ (.A1(net4832),
    .A2(net4427),
    .Y(_01084_),
    .B1(_03611_));
 sg13g2_nor2_1 _18981_ (.A(net3429),
    .B(net4427),
    .Y(_03612_));
 sg13g2_a21oi_1 _18982_ (.A1(net4830),
    .A2(net4427),
    .Y(_01085_),
    .B1(_03612_));
 sg13g2_nor2_1 _18983_ (.A(net3853),
    .B(net4433),
    .Y(_03613_));
 sg13g2_a21oi_1 _18984_ (.A1(_02763_),
    .A2(net4433),
    .Y(_01086_),
    .B1(_03613_));
 sg13g2_nor2_1 _18985_ (.A(net4056),
    .B(net4433),
    .Y(_03614_));
 sg13g2_a21oi_1 _18986_ (.A1(_02767_),
    .A2(net4433),
    .Y(_01087_),
    .B1(_03614_));
 sg13g2_o21ai_1 _18987_ (.B1(net5603),
    .Y(_03615_),
    .A1(_02995_),
    .A2(net4466));
 sg13g2_o21ai_1 _18988_ (.B1(_02999_),
    .Y(_03616_),
    .A1(net4),
    .A2(net5600));
 sg13g2_nand2_1 _18989_ (.Y(_03617_),
    .A(_03615_),
    .B(_03616_));
 sg13g2_o21ai_1 _18990_ (.B1(_03617_),
    .Y(_01088_),
    .A1(_06830_),
    .A2(_03615_));
 sg13g2_xnor2_1 _18991_ (.Y(_03618_),
    .A(net5),
    .B(net4));
 sg13g2_nor2_1 _18992_ (.A(net5600),
    .B(_03618_),
    .Y(_03619_));
 sg13g2_a21oi_1 _18993_ (.A1(net5599),
    .A2(net4916),
    .Y(_03620_),
    .B1(_03619_));
 sg13g2_mux2_1 _18994_ (.A0(net3961),
    .A1(_03620_),
    .S(_03615_),
    .X(_01089_));
 sg13g2_a21oi_1 _18995_ (.A1(net5599),
    .A2(net4850),
    .Y(_03621_),
    .B1(_03619_));
 sg13g2_mux2_1 _18996_ (.A0(net3947),
    .A1(_03621_),
    .S(_03615_),
    .X(_01090_));
 sg13g2_o21ai_1 _18997_ (.B1(_03008_),
    .Y(_03622_),
    .A1(net5599),
    .A2(_03618_));
 sg13g2_mux2_1 _18998_ (.A0(net3917),
    .A1(_03622_),
    .S(_03615_),
    .X(_01091_));
 sg13g2_o21ai_1 _18999_ (.B1(net5603),
    .Y(_03623_),
    .A1(_03045_),
    .A2(net4466));
 sg13g2_mux2_1 _19000_ (.A0(net3832),
    .A1(_03616_),
    .S(_03623_),
    .X(_01092_));
 sg13g2_mux2_1 _19001_ (.A0(net3818),
    .A1(_03620_),
    .S(_03623_),
    .X(_01093_));
 sg13g2_mux2_1 _19002_ (.A0(net3819),
    .A1(_03621_),
    .S(_03623_),
    .X(_01094_));
 sg13g2_mux2_1 _19003_ (.A0(net3793),
    .A1(_03622_),
    .S(_03623_),
    .X(_01095_));
 sg13g2_o21ai_1 _19004_ (.B1(net5604),
    .Y(_03624_),
    .A1(_09615_),
    .A2(_03537_));
 sg13g2_mux2_1 _19005_ (.A0(net3913),
    .A1(_03616_),
    .S(_03624_),
    .X(_01096_));
 sg13g2_mux2_1 _19006_ (.A0(net3750),
    .A1(_03620_),
    .S(_03624_),
    .X(_01097_));
 sg13g2_mux2_1 _19007_ (.A0(net3742),
    .A1(_03621_),
    .S(_03624_),
    .X(_01098_));
 sg13g2_mux2_1 _19008_ (.A0(net3700),
    .A1(_03622_),
    .S(_03624_),
    .X(_01099_));
 sg13g2_a21oi_1 _19009_ (.A1(net5681),
    .A2(net5351),
    .Y(_03625_),
    .B1(net5378));
 sg13g2_o21ai_1 _19010_ (.B1(_03625_),
    .Y(_01100_),
    .A1(net5681),
    .A2(net5352));
 sg13g2_nand2_1 _19011_ (.Y(_03626_),
    .A(net5354),
    .B(_08865_));
 sg13g2_o21ai_1 _19012_ (.B1(net6157),
    .Y(_03627_),
    .A1(net5681),
    .A2(net5352));
 sg13g2_a21oi_1 _19013_ (.A1(_03626_),
    .A2(net6158),
    .Y(_01101_),
    .B1(net5377));
 sg13g2_a21oi_1 _19014_ (.A1(net5680),
    .A2(_03626_),
    .Y(_03628_),
    .B1(net5377));
 sg13g2_o21ai_1 _19015_ (.B1(_03628_),
    .Y(_01102_),
    .A1(net5680),
    .A2(_03626_));
 sg13g2_nand2_1 _19016_ (.Y(_03629_),
    .A(_09093_),
    .B(_09096_));
 sg13g2_nor4_2 _19017_ (.A(net1400),
    .B(_08930_),
    .C(_09099_),
    .Y(_03630_),
    .D(_03629_));
 sg13g2_nor4_1 _19018_ (.A(net3870),
    .B(net3524),
    .C(net3589),
    .D(net3788),
    .Y(_03631_));
 sg13g2_xnor2_1 _19019_ (.Y(_03632_),
    .A(net3870),
    .B(net5355));
 sg13g2_nor3_1 _19020_ (.A(_03630_),
    .B(_03631_),
    .C(_03632_),
    .Y(_01103_));
 sg13g2_nand2_1 _19021_ (.Y(_03633_),
    .A(net3524),
    .B(_06942_));
 sg13g2_or2_1 _19022_ (.X(_03634_),
    .B(_03631_),
    .A(_06944_));
 sg13g2_a21oi_1 _19023_ (.A1(net3525),
    .A2(_03634_),
    .Y(_01104_),
    .B1(_03630_));
 sg13g2_nand2_1 _19024_ (.Y(_03635_),
    .A(net3788),
    .B(_06944_));
 sg13g2_nor2_1 _19025_ (.A(net3788),
    .B(_06944_),
    .Y(_03636_));
 sg13g2_nand2_1 _19026_ (.Y(_03637_),
    .A(net3589),
    .B(_03636_));
 sg13g2_a21oi_1 _19027_ (.A1(_03635_),
    .A2(_03637_),
    .Y(_01105_),
    .B1(_03630_));
 sg13g2_o21ai_1 _19028_ (.B1(net3589),
    .Y(_03638_),
    .A1(\fpga_top.qspi_if.rst_cntr[2] ),
    .A2(_06944_));
 sg13g2_nand2b_1 _19029_ (.Y(_01106_),
    .B(net3590),
    .A_N(_03630_));
 sg13g2_nand4_1 _19030_ (.B(_09287_),
    .C(_09290_),
    .A(_09277_),
    .Y(_03639_),
    .D(_09291_));
 sg13g2_nor2_2 _19031_ (.A(_09541_),
    .B(net6600),
    .Y(_03640_));
 sg13g2_xor2_1 _19032_ (.B(_03640_),
    .A(net1519),
    .X(_01107_));
 sg13g2_and2_1 _19033_ (.A(net1519),
    .B(_03640_),
    .X(_03641_));
 sg13g2_nand2_1 _19034_ (.Y(_03642_),
    .A(net1909),
    .B(_03641_));
 sg13g2_xor2_1 _19035_ (.B(_03641_),
    .A(net1909),
    .X(_01108_));
 sg13g2_nor2_2 _19036_ (.A(net5668),
    .B(_03642_),
    .Y(_03643_));
 sg13g2_xnor2_1 _19037_ (.Y(_01109_),
    .A(net5668),
    .B(_03642_));
 sg13g2_nand2_1 _19038_ (.Y(_03644_),
    .A(net1370),
    .B(\fpga_top.uart_top.rx_fifo_dvalid ));
 sg13g2_xnor2_1 _19039_ (.Y(_01110_),
    .A(net1370),
    .B(net5338));
 sg13g2_nand3_1 _19040_ (.B(net1367),
    .C(\fpga_top.uart_top.rx_fifo_dvalid ),
    .A(net1370),
    .Y(_03645_));
 sg13g2_xnor2_1 _19041_ (.Y(_01111_),
    .A(net1367),
    .B(_03644_));
 sg13g2_xnor2_1 _19042_ (.Y(_01112_),
    .A(net1364),
    .B(_03645_));
 sg13g2_xnor2_1 _19043_ (.Y(_03646_),
    .A(\fpga_top.uart_top.rx_fifo_dvalid ),
    .B(_03640_));
 sg13g2_xnor2_1 _19044_ (.Y(_01113_),
    .A(net1614),
    .B(_03646_));
 sg13g2_or3_1 _19045_ (.A(net1390),
    .B(net1614),
    .C(_03640_),
    .X(_03647_));
 sg13g2_o21ai_1 _19046_ (.B1(net1390),
    .Y(_03648_),
    .A1(net1614),
    .A2(_03640_));
 sg13g2_o21ai_1 _19047_ (.B1(_03648_),
    .Y(_01114_),
    .A1(_08872_),
    .A2(_03647_));
 sg13g2_and2_1 _19048_ (.A(net2176),
    .B(_03647_),
    .X(_03649_));
 sg13g2_nor2_1 _19049_ (.A(net2176),
    .B(_03647_),
    .Y(_03650_));
 sg13g2_a21o_1 _19050_ (.A2(_03650_),
    .A1(net1897),
    .B1(_03649_),
    .X(_01115_));
 sg13g2_nor2b_1 _19051_ (.A(_03650_),
    .B_N(net1897),
    .Y(_01116_));
 sg13g2_nand2_1 _19052_ (.Y(_03651_),
    .A(net5666),
    .B(_09905_));
 sg13g2_nor2_1 _19053_ (.A(\fpga_top.uart_top.uart_send_char.send_cntr[4] ),
    .B(net5712),
    .Y(_03652_));
 sg13g2_a21oi_2 _19054_ (.B1(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[3] ),
    .Y(_03653_),
    .A2(_03652_),
    .A1(_03651_));
 sg13g2_inv_1 _19055_ (.Y(_03654_),
    .A(_03653_));
 sg13g2_nand2_2 _19056_ (.Y(_03655_),
    .A(net3032),
    .B(net5146));
 sg13g2_xor2_1 _19057_ (.B(net6118),
    .A(net3032),
    .X(_01117_));
 sg13g2_nand3_1 _19058_ (.B(net3889),
    .C(_03653_),
    .A(net3032),
    .Y(_03656_));
 sg13g2_xnor2_1 _19059_ (.Y(_01118_),
    .A(net3889),
    .B(_03655_));
 sg13g2_nor2_1 _19060_ (.A(net6592),
    .B(_03656_),
    .Y(_03657_));
 sg13g2_xnor2_1 _19061_ (.Y(_01119_),
    .A(net3356),
    .B(_03656_));
 sg13g2_xor2_1 _19062_ (.B(net1393),
    .A(net1368),
    .X(_01120_));
 sg13g2_a21oi_1 _19063_ (.A1(net1368),
    .A2(net1393),
    .Y(_03658_),
    .B1(net1365));
 sg13g2_nand3_1 _19064_ (.B(net1365),
    .C(net1393),
    .A(net1368),
    .Y(_03659_));
 sg13g2_nor2b_1 _19065_ (.A(_03658_),
    .B_N(_03659_),
    .Y(_01121_));
 sg13g2_xnor2_1 _19066_ (.Y(_01122_),
    .A(net1362),
    .B(_03659_));
 sg13g2_xnor2_1 _19067_ (.Y(_03660_),
    .A(_09519_),
    .B(net5146));
 sg13g2_xnor2_1 _19068_ (.Y(_01123_),
    .A(net1536),
    .B(_03660_));
 sg13g2_xnor2_1 _19069_ (.Y(_03661_),
    .A(net3855),
    .B(net5146));
 sg13g2_nand2_1 _19070_ (.Y(_03662_),
    .A(net1536),
    .B(_03661_));
 sg13g2_or2_1 _19071_ (.X(_03663_),
    .B(_03661_),
    .A(net1536));
 sg13g2_a21oi_1 _19072_ (.A1(_03662_),
    .A2(_03663_),
    .Y(_03664_),
    .B1(_03660_));
 sg13g2_a21oi_1 _19073_ (.A1(_06502_),
    .A2(_03660_),
    .Y(_01124_),
    .B1(_03664_));
 sg13g2_xnor2_1 _19074_ (.Y(_03665_),
    .A(net3386),
    .B(net5146));
 sg13g2_o21ai_1 _19075_ (.B1(_03662_),
    .Y(_03666_),
    .A1(_06502_),
    .A2(net5146));
 sg13g2_a21oi_1 _19076_ (.A1(_03665_),
    .A2(_03666_),
    .Y(_03667_),
    .B1(_03660_));
 sg13g2_o21ai_1 _19077_ (.B1(_03667_),
    .Y(_03668_),
    .A1(_03665_),
    .A2(_03666_));
 sg13g2_nand2_1 _19078_ (.Y(_03669_),
    .A(net3386),
    .B(_03660_));
 sg13g2_nand2_1 _19079_ (.Y(_01125_),
    .A(_03668_),
    .B(_03669_));
 sg13g2_a21oi_1 _19080_ (.A1(_09520_),
    .A2(net5146),
    .Y(_03670_),
    .B1(net6117));
 sg13g2_o21ai_1 _19081_ (.B1(_03667_),
    .Y(_03671_),
    .A1(_06503_),
    .A2(net5146));
 sg13g2_xor2_1 _19082_ (.B(_03671_),
    .A(_03670_),
    .X(_01126_));
 sg13g2_and2_1 _19083_ (.A(_06674_),
    .B(_09346_),
    .X(_03672_));
 sg13g2_nor2_1 _19084_ (.A(_06674_),
    .B(_09345_),
    .Y(_03673_));
 sg13g2_nor3_1 _19085_ (.A(_09335_),
    .B(_03672_),
    .C(net6284),
    .Y(_01127_));
 sg13g2_nor2_1 _19086_ (.A(\fpga_top.uart_top.uart_if.tx_out_cntr[1] ),
    .B(_09518_),
    .Y(_03674_));
 sg13g2_inv_1 _19087_ (.Y(_03675_),
    .A(_03674_));
 sg13g2_xnor2_1 _19088_ (.Y(_03676_),
    .A(net6348),
    .B(_09517_));
 sg13g2_o21ai_1 _19089_ (.B1(net5284),
    .Y(_01128_),
    .A1(net1393),
    .A2(net6349));
 sg13g2_nand2_1 _19090_ (.Y(_03677_),
    .A(net3443),
    .B(_03675_));
 sg13g2_nand3b_1 _19091_ (.B(_03674_),
    .C(net1392),
    .Y(_03678_),
    .A_N(net3443));
 sg13g2_a21oi_1 _19092_ (.A1(_03677_),
    .A2(_03678_),
    .Y(_01129_),
    .B1(net3731));
 sg13g2_o21ai_1 _19093_ (.B1(net1392),
    .Y(_03679_),
    .A1(net3443),
    .A2(_03675_));
 sg13g2_nand2_1 _19094_ (.Y(_01130_),
    .A(net5284),
    .B(net3444));
 sg13g2_a21oi_1 _19095_ (.A1(_00121_),
    .A2(_09346_),
    .Y(_03680_),
    .B1(_09335_));
 sg13g2_o21ai_1 _19096_ (.B1(_03680_),
    .Y(_01131_),
    .A1(net1385),
    .A2(_09346_));
 sg13g2_mux4_1 _19097_ (.S0(net5413),
    .A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][0] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][0] ),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][0] ),
    .A3(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][0] ),
    .S1(net5410),
    .X(_03681_));
 sg13g2_mux2_1 _19098_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][0] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][0] ),
    .S(net5413),
    .X(_03682_));
 sg13g2_nor2b_1 _19099_ (.A(net1431),
    .B_N(net5413),
    .Y(_03683_));
 sg13g2_o21ai_1 _19100_ (.B1(net5410),
    .Y(_03684_),
    .A1(net5413),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][0] ));
 sg13g2_o21ai_1 _19101_ (.B1(net5407),
    .Y(_03685_),
    .A1(_03683_),
    .A2(_03684_));
 sg13g2_a21oi_1 _19102_ (.A1(_06848_),
    .A2(_03682_),
    .Y(_03686_),
    .B1(_03685_));
 sg13g2_nor2_1 _19103_ (.A(net5284),
    .B(_03686_),
    .Y(_03687_));
 sg13g2_o21ai_1 _19104_ (.B1(_03687_),
    .Y(_03688_),
    .A1(net5407),
    .A2(_03681_));
 sg13g2_o21ai_1 _19105_ (.B1(net5282),
    .Y(_03689_),
    .A1(net1631),
    .A2(_09346_));
 sg13g2_a22oi_1 _19106_ (.Y(_01132_),
    .B1(_03688_),
    .B2(_03689_),
    .A2(net4945),
    .A1(_06847_));
 sg13g2_nor2b_1 _19107_ (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][1] ),
    .B_N(net5418),
    .Y(_03690_));
 sg13g2_nor2_1 _19108_ (.A(net5420),
    .B(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][1] ),
    .Y(_03691_));
 sg13g2_nor3_1 _19109_ (.A(net5409),
    .B(_03690_),
    .C(_03691_),
    .Y(_03692_));
 sg13g2_nor2b_1 _19110_ (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][1] ),
    .B_N(net5419),
    .Y(_03693_));
 sg13g2_o21ai_1 _19111_ (.B1(net5412),
    .Y(_03694_),
    .A1(net5419),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][1] ));
 sg13g2_o21ai_1 _19112_ (.B1(net5406),
    .Y(_03695_),
    .A1(_03693_),
    .A2(_03694_));
 sg13g2_a21oi_1 _19113_ (.A1(net5415),
    .A2(_06850_),
    .Y(_03696_),
    .B1(net5411));
 sg13g2_o21ai_1 _19114_ (.B1(_03696_),
    .Y(_03697_),
    .A1(net5415),
    .A2(net1693));
 sg13g2_o21ai_1 _19115_ (.B1(net5410),
    .Y(_03698_),
    .A1(net5413),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][1] ));
 sg13g2_a21oi_1 _19116_ (.A1(net5413),
    .A2(_06851_),
    .Y(_03699_),
    .B1(_03698_));
 sg13g2_nor2_1 _19117_ (.A(net5407),
    .B(_03699_),
    .Y(_03700_));
 sg13g2_a21oi_1 _19118_ (.A1(net1694),
    .A2(_03700_),
    .Y(_03701_),
    .B1(net5284));
 sg13g2_o21ai_1 _19119_ (.B1(_03701_),
    .Y(_03702_),
    .A1(_03692_),
    .A2(_03695_));
 sg13g2_o21ai_1 _19120_ (.B1(net5283),
    .Y(_03703_),
    .A1(net1491),
    .A2(_09346_));
 sg13g2_a22oi_1 _19121_ (.Y(_01133_),
    .B1(net1695),
    .B2(_03703_),
    .A2(net4946),
    .A1(_06849_));
 sg13g2_nor2b_1 _19122_ (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][2] ),
    .B_N(net5419),
    .Y(_03704_));
 sg13g2_nor2_1 _19123_ (.A(net5420),
    .B(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][2] ),
    .Y(_03705_));
 sg13g2_nor3_1 _19124_ (.A(net5412),
    .B(_03704_),
    .C(_03705_),
    .Y(_03706_));
 sg13g2_nor2b_1 _19125_ (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][2] ),
    .B_N(net5419),
    .Y(_03707_));
 sg13g2_o21ai_1 _19126_ (.B1(net5412),
    .Y(_03708_),
    .A1(net5419),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][2] ));
 sg13g2_o21ai_1 _19127_ (.B1(_00013_),
    .Y(_03709_),
    .A1(_03707_),
    .A2(_03708_));
 sg13g2_or2_1 _19128_ (.X(_03710_),
    .B(_03709_),
    .A(_03706_));
 sg13g2_a21oi_1 _19129_ (.A1(net5415),
    .A2(_06852_),
    .Y(_03711_),
    .B1(net5411));
 sg13g2_o21ai_1 _19130_ (.B1(_03711_),
    .Y(_03712_),
    .A1(net5419),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][2] ));
 sg13g2_o21ai_1 _19131_ (.B1(net5412),
    .Y(_03713_),
    .A1(net5415),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][2] ));
 sg13g2_a21oi_1 _19132_ (.A1(net5419),
    .A2(_06853_),
    .Y(_03714_),
    .B1(_03713_));
 sg13g2_nor2_1 _19133_ (.A(net5407),
    .B(_03714_),
    .Y(_03715_));
 sg13g2_a21oi_1 _19134_ (.A1(_03712_),
    .A2(_03715_),
    .Y(_03716_),
    .B1(net5283));
 sg13g2_a22oi_1 _19135_ (.Y(_03717_),
    .B1(_03710_),
    .B2(_03716_),
    .A2(net5283),
    .A1(\fpga_top.uart_top.uart_if.tx_out_data[4] ));
 sg13g2_nand2_1 _19136_ (.Y(_03718_),
    .A(net1491),
    .B(net4946));
 sg13g2_o21ai_1 _19137_ (.B1(_03718_),
    .Y(_01134_),
    .A1(net4945),
    .A2(_03717_));
 sg13g2_a21oi_1 _19138_ (.A1(net5418),
    .A2(_06855_),
    .Y(_03719_),
    .B1(net5408));
 sg13g2_o21ai_1 _19139_ (.B1(_03719_),
    .Y(_03720_),
    .A1(net5418),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][3] ));
 sg13g2_o21ai_1 _19140_ (.B1(net5408),
    .Y(_03721_),
    .A1(net5418),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][3] ));
 sg13g2_a21oi_1 _19141_ (.A1(net5418),
    .A2(_06856_),
    .Y(_03722_),
    .B1(_03721_));
 sg13g2_nor2_1 _19142_ (.A(net5406),
    .B(_03722_),
    .Y(_03723_));
 sg13g2_nor2b_1 _19143_ (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][3] ),
    .B_N(net5417),
    .Y(_03724_));
 sg13g2_nor2_1 _19144_ (.A(net5417),
    .B(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][3] ),
    .Y(_03725_));
 sg13g2_nor3_1 _19145_ (.A(net5408),
    .B(_03724_),
    .C(_03725_),
    .Y(_03726_));
 sg13g2_nor2b_1 _19146_ (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][3] ),
    .B_N(net5417),
    .Y(_03727_));
 sg13g2_o21ai_1 _19147_ (.B1(net5409),
    .Y(_03728_),
    .A1(net5418),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][3] ));
 sg13g2_o21ai_1 _19148_ (.B1(net5406),
    .Y(_03729_),
    .A1(_03727_),
    .A2(_03728_));
 sg13g2_a21oi_1 _19149_ (.A1(_03720_),
    .A2(_03723_),
    .Y(_03730_),
    .B1(net5282));
 sg13g2_o21ai_1 _19150_ (.B1(_03730_),
    .Y(_03731_),
    .A1(_03726_),
    .A2(_03729_));
 sg13g2_o21ai_1 _19151_ (.B1(net5283),
    .Y(_03732_),
    .A1(net1514),
    .A2(_09346_));
 sg13g2_a22oi_1 _19152_ (.Y(_01135_),
    .B1(_03731_),
    .B2(_03732_),
    .A2(net4945),
    .A1(_06854_));
 sg13g2_nand2b_1 _19153_ (.Y(_03733_),
    .B(net5415),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][4] ));
 sg13g2_o21ai_1 _19154_ (.B1(_03733_),
    .Y(_03734_),
    .A1(net5415),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][4] ));
 sg13g2_mux2_1 _19155_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][4] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][4] ),
    .S(net5414),
    .X(_03735_));
 sg13g2_o21ai_1 _19156_ (.B1(net5407),
    .Y(_03736_),
    .A1(net5411),
    .A2(_03734_));
 sg13g2_a21oi_1 _19157_ (.A1(net5411),
    .A2(_03735_),
    .Y(_03737_),
    .B1(_03736_));
 sg13g2_nand2b_1 _19158_ (.Y(_03738_),
    .B(net5414),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][4] ));
 sg13g2_o21ai_1 _19159_ (.B1(_03738_),
    .Y(_03739_),
    .A1(net5415),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][4] ));
 sg13g2_mux2_1 _19160_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][4] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][4] ),
    .S(net5419),
    .X(_03740_));
 sg13g2_a21oi_1 _19161_ (.A1(net5412),
    .A2(_03740_),
    .Y(_03741_),
    .B1(net5406));
 sg13g2_o21ai_1 _19162_ (.B1(_03741_),
    .Y(_03742_),
    .A1(net5412),
    .A2(_03739_));
 sg13g2_nor2_1 _19163_ (.A(net5284),
    .B(_03737_),
    .Y(_03743_));
 sg13g2_a22oi_1 _19164_ (.Y(_03744_),
    .B1(_03742_),
    .B2(_03743_),
    .A2(net5283),
    .A1(\fpga_top.uart_top.uart_if.tx_out_data[6] ));
 sg13g2_nand2_1 _19165_ (.Y(_03745_),
    .A(net1514),
    .B(net4946));
 sg13g2_o21ai_1 _19166_ (.B1(_03745_),
    .Y(_01136_),
    .A1(net4946),
    .A2(_03744_));
 sg13g2_nand2b_1 _19167_ (.Y(_03746_),
    .B(net5413),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][5] ));
 sg13g2_o21ai_1 _19168_ (.B1(_03746_),
    .Y(_03747_),
    .A1(net5413),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][5] ));
 sg13g2_mux2_1 _19169_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][5] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][5] ),
    .S(net5416),
    .X(_03748_));
 sg13g2_o21ai_1 _19170_ (.B1(net5406),
    .Y(_03749_),
    .A1(net5410),
    .A2(_03747_));
 sg13g2_a21oi_1 _19171_ (.A1(net5408),
    .A2(_03748_),
    .Y(_03750_),
    .B1(_03749_));
 sg13g2_nand2b_1 _19172_ (.Y(_03751_),
    .B(net5420),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][5] ));
 sg13g2_o21ai_1 _19173_ (.B1(_03751_),
    .Y(_03752_),
    .A1(net5420),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][5] ));
 sg13g2_mux2_1 _19174_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][5] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][5] ),
    .S(net5418),
    .X(_03753_));
 sg13g2_a21oi_1 _19175_ (.A1(net5409),
    .A2(_03753_),
    .Y(_03754_),
    .B1(net5406));
 sg13g2_o21ai_1 _19176_ (.B1(_03754_),
    .Y(_03755_),
    .A1(net5409),
    .A2(_03752_));
 sg13g2_nor2_1 _19177_ (.A(net5282),
    .B(_03750_),
    .Y(_03756_));
 sg13g2_a22oi_1 _19178_ (.Y(_03757_),
    .B1(_03755_),
    .B2(_03756_),
    .A2(net5282),
    .A1(net1411));
 sg13g2_nand2_1 _19179_ (.Y(_03758_),
    .A(net1576),
    .B(net4946));
 sg13g2_o21ai_1 _19180_ (.B1(_03758_),
    .Y(_01137_),
    .A1(net4946),
    .A2(_03757_));
 sg13g2_nand2b_1 _19181_ (.Y(_03759_),
    .B(net5414),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][6] ));
 sg13g2_o21ai_1 _19182_ (.B1(_03759_),
    .Y(_03760_),
    .A1(net5414),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][6] ));
 sg13g2_mux2_1 _19183_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][6] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][6] ),
    .S(net5414),
    .X(_03761_));
 sg13g2_o21ai_1 _19184_ (.B1(net5407),
    .Y(_03762_),
    .A1(net5411),
    .A2(_03760_));
 sg13g2_a21oi_1 _19185_ (.A1(net5411),
    .A2(_03761_),
    .Y(_03763_),
    .B1(_03762_));
 sg13g2_nand2b_1 _19186_ (.Y(_03764_),
    .B(net5414),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][6] ));
 sg13g2_o21ai_1 _19187_ (.B1(_03764_),
    .Y(_03765_),
    .A1(net5414),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][6] ));
 sg13g2_mux2_1 _19188_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][6] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][6] ),
    .S(net5414),
    .X(_03766_));
 sg13g2_a21oi_1 _19189_ (.A1(net5411),
    .A2(_03766_),
    .Y(_03767_),
    .B1(net5407));
 sg13g2_o21ai_1 _19190_ (.B1(_03767_),
    .Y(_03768_),
    .A1(net5411),
    .A2(_03765_));
 sg13g2_nor2_1 _19191_ (.A(net5284),
    .B(_03763_),
    .Y(_03769_));
 sg13g2_a22oi_1 _19192_ (.Y(_03770_),
    .B1(_03768_),
    .B2(_03769_),
    .A2(net5284),
    .A1(\fpga_top.uart_top.uart_if.tx_out_data[8] ));
 sg13g2_nand2_1 _19193_ (.Y(_03771_),
    .A(net1411),
    .B(net4945));
 sg13g2_o21ai_1 _19194_ (.B1(_03771_),
    .Y(_01138_),
    .A1(net4945),
    .A2(_03770_));
 sg13g2_nand2b_1 _19195_ (.Y(_03772_),
    .B(net5417),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][7] ));
 sg13g2_o21ai_1 _19196_ (.B1(_03772_),
    .Y(_03773_),
    .A1(net5417),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][7] ));
 sg13g2_mux2_1 _19197_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][7] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][7] ),
    .S(net5417),
    .X(_03774_));
 sg13g2_o21ai_1 _19198_ (.B1(net5406),
    .Y(_03775_),
    .A1(net5408),
    .A2(_03773_));
 sg13g2_a21oi_1 _19199_ (.A1(net5408),
    .A2(_03774_),
    .Y(_03776_),
    .B1(_03775_));
 sg13g2_nand2b_1 _19200_ (.Y(_03777_),
    .B(net5421),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][7] ));
 sg13g2_o21ai_1 _19201_ (.B1(_03777_),
    .Y(_03778_),
    .A1(net5417),
    .A2(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][7] ));
 sg13g2_mux2_1 _19202_ (.A0(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][7] ),
    .A1(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][7] ),
    .S(net5417),
    .X(_03779_));
 sg13g2_a21oi_1 _19203_ (.A1(net5408),
    .A2(_03779_),
    .Y(_03780_),
    .B1(net5406));
 sg13g2_o21ai_1 _19204_ (.B1(_03780_),
    .Y(_03781_),
    .A1(net5408),
    .A2(_03778_));
 sg13g2_nor2_1 _19205_ (.A(net5282),
    .B(_03776_),
    .Y(_03782_));
 sg13g2_a22oi_1 _19206_ (.Y(_03783_),
    .B1(_03781_),
    .B2(_03782_),
    .A2(net5282),
    .A1(net1596));
 sg13g2_nand2_1 _19207_ (.Y(_03784_),
    .A(net1604),
    .B(net4945));
 sg13g2_o21ai_1 _19208_ (.B1(_03784_),
    .Y(_01139_),
    .A1(net4945),
    .A2(_03783_));
 sg13g2_nand2b_1 _19209_ (.Y(_01140_),
    .B(net4945),
    .A_N(net1596));
 sg13g2_xor2_1 _19210_ (.B(net4948),
    .A(net2105),
    .X(_01141_));
 sg13g2_nor2_1 _19211_ (.A(\fpga_top.bus_gather.u_read_adr[30] ),
    .B(_09563_),
    .Y(_03785_));
 sg13g2_or2_1 _19212_ (.X(_03786_),
    .B(_09563_),
    .A(\fpga_top.bus_gather.u_read_adr[30] ));
 sg13g2_nand2_1 _19213_ (.Y(_03787_),
    .A(\fpga_top.bus_gather.u_read_adr[5] ),
    .B(net5065));
 sg13g2_and2_1 _19214_ (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[31] ),
    .B(_09651_),
    .X(_03788_));
 sg13g2_nand2_2 _19215_ (.Y(_03789_),
    .A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[31] ),
    .B(_09651_));
 sg13g2_nor2_1 _19216_ (.A(\fpga_top.cpu_top.csr_wadr_mon[3] ),
    .B(_03789_),
    .Y(_03790_));
 sg13g2_o21ai_1 _19217_ (.B1(_03786_),
    .Y(_03791_),
    .A1(\fpga_top.cpu_top.alui_shamt[3] ),
    .A2(net4908));
 sg13g2_o21ai_1 _19218_ (.B1(_03787_),
    .Y(_03792_),
    .A1(_03790_),
    .A2(_03791_));
 sg13g2_nand2_1 _19219_ (.Y(_03793_),
    .A(\fpga_top.bus_gather.u_read_adr[4] ),
    .B(net5065));
 sg13g2_nor2_1 _19220_ (.A(\fpga_top.cpu_top.csr_wadr_mon[2] ),
    .B(_03789_),
    .Y(_03794_));
 sg13g2_o21ai_1 _19221_ (.B1(_03786_),
    .Y(_03795_),
    .A1(\fpga_top.cpu_top.alui_shamt[2] ),
    .A2(net4908));
 sg13g2_o21ai_1 _19222_ (.B1(_03793_),
    .Y(_03796_),
    .A1(_03794_),
    .A2(_03795_));
 sg13g2_nor2_2 _19223_ (.A(_03792_),
    .B(_03796_),
    .Y(_03797_));
 sg13g2_o21ai_1 _19224_ (.B1(_03786_),
    .Y(_03798_),
    .A1(net5573),
    .A2(net4908));
 sg13g2_a21oi_1 _19225_ (.A1(_06665_),
    .A2(net4908),
    .Y(_03799_),
    .B1(_03798_));
 sg13g2_a21oi_2 _19226_ (.B1(_03799_),
    .Y(_03800_),
    .A2(net5065),
    .A1(net5616));
 sg13g2_inv_1 _19227_ (.Y(_03801_),
    .A(_03800_));
 sg13g2_nand2_1 _19228_ (.Y(_03802_),
    .A(\fpga_top.cpu_top.alui_shamt[1] ),
    .B(_03789_));
 sg13g2_a21oi_1 _19229_ (.A1(\fpga_top.cpu_top.csr_wadr_mon[1] ),
    .A2(_03788_),
    .Y(_03803_),
    .B1(net5066));
 sg13g2_a22oi_1 _19230_ (.Y(_03804_),
    .B1(_03802_),
    .B2(_03803_),
    .A2(net5066),
    .A1(_06505_));
 sg13g2_nor2_2 _19231_ (.A(_03801_),
    .B(_03804_),
    .Y(_03805_));
 sg13g2_nand2_2 _19232_ (.Y(_03806_),
    .A(_03797_),
    .B(_03805_));
 sg13g2_nand2_1 _19233_ (.Y(_03807_),
    .A(_06509_),
    .B(_06513_));
 sg13g2_nor4_2 _19234_ (.A(\fpga_top.bus_gather.u_read_adr[13] ),
    .B(\fpga_top.bus_gather.u_read_adr[12] ),
    .C(_06523_),
    .Y(_03808_),
    .D(_03807_));
 sg13g2_nand2b_1 _19235_ (.Y(_03809_),
    .B(\fpga_top.cpu_top.csr_wadr_mon[8] ),
    .A_N(\fpga_top.cpu_top.csr_wadr_mon[11] ));
 sg13g2_nor4_2 _19236_ (.A(\fpga_top.cpu_top.csr_wadr_mon[5] ),
    .B(\fpga_top.cpu_top.csr_wadr_mon[7] ),
    .C(\fpga_top.cpu_top.csr_wadr_mon[10] ),
    .Y(_03810_),
    .D(_03809_));
 sg13g2_nand2_1 _19237_ (.Y(_03811_),
    .A(net4908),
    .B(_03810_));
 sg13g2_nor2b_1 _19238_ (.A(\fpga_top.cpu_top.br_ofs[10] ),
    .B_N(\fpga_top.cpu_top.br_ofs[8] ),
    .Y(_03812_));
 sg13g2_nand4_1 _19239_ (.B(_07288_),
    .C(_03789_),
    .A(_06558_),
    .Y(_03813_),
    .D(_03812_));
 sg13g2_nand3_1 _19240_ (.B(_03811_),
    .C(_03813_),
    .A(_03786_),
    .Y(_03814_));
 sg13g2_o21ai_1 _19241_ (.B1(_03814_),
    .Y(_03815_),
    .A1(_03786_),
    .A2(_03808_));
 sg13g2_nand2_1 _19242_ (.Y(_03816_),
    .A(_06669_),
    .B(net4908));
 sg13g2_a21oi_1 _19243_ (.A1(_06556_),
    .A2(_03789_),
    .Y(_03817_),
    .B1(net5065));
 sg13g2_a22oi_1 _19244_ (.Y(_03818_),
    .B1(_03816_),
    .B2(_03817_),
    .A2(net5065),
    .A1(\fpga_top.bus_gather.u_read_adr[11] ));
 sg13g2_inv_4 _19245_ (.A(_03818_),
    .Y(_03819_));
 sg13g2_nand2_1 _19246_ (.Y(_03820_),
    .A(net5571),
    .B(_03789_));
 sg13g2_a21oi_1 _19247_ (.A1(\fpga_top.cpu_top.csr_wadr_mon[6] ),
    .A2(net4908),
    .Y(_03821_),
    .B1(net5065));
 sg13g2_a22oi_1 _19248_ (.Y(_03822_),
    .B1(_03820_),
    .B2(_03821_),
    .A2(net5065),
    .A1(_06511_));
 sg13g2_inv_1 _19249_ (.Y(_03823_),
    .A(_03822_));
 sg13g2_or4_1 _19250_ (.A(_03806_),
    .B(_03815_),
    .C(_03818_),
    .D(_03822_),
    .X(_03824_));
 sg13g2_nand2_1 _19251_ (.Y(_03825_),
    .A(\fpga_top.bus_gather.u_read_adr[6] ),
    .B(net5065));
 sg13g2_nor2_1 _19252_ (.A(\fpga_top.cpu_top.csr_wadr_mon[4] ),
    .B(_03789_),
    .Y(_03826_));
 sg13g2_o21ai_1 _19253_ (.B1(_03786_),
    .Y(_03827_),
    .A1(\fpga_top.cpu_top.alui_shamt[4] ),
    .A2(net4908));
 sg13g2_o21ai_1 _19254_ (.B1(_03825_),
    .Y(_03828_),
    .A1(_03826_),
    .A2(_03827_));
 sg13g2_nor2b_2 _19255_ (.A(_03824_),
    .B_N(_03828_),
    .Y(_03829_));
 sg13g2_nor2_2 _19256_ (.A(net5193),
    .B(_09459_),
    .Y(_03830_));
 sg13g2_nand3_1 _19257_ (.B(net5293),
    .C(_09445_),
    .A(net6533),
    .Y(_03831_));
 sg13g2_nor2_2 _19258_ (.A(_03788_),
    .B(net5050),
    .Y(_03832_));
 sg13g2_nand2_1 _19259_ (.Y(_03833_),
    .A(_03789_),
    .B(net5136));
 sg13g2_and2_1 _19260_ (.A(net4629),
    .B(net4829),
    .X(_03834_));
 sg13g2_nand2_2 _19261_ (.Y(_03835_),
    .A(net4628),
    .B(net4828));
 sg13g2_and2_1 _19262_ (.A(net4631),
    .B(net5059),
    .X(_03836_));
 sg13g2_nand2_2 _19263_ (.Y(_03837_),
    .A(net4629),
    .B(net5048));
 sg13g2_nor2_2 _19264_ (.A(net5343),
    .B(_07606_),
    .Y(_03838_));
 sg13g2_or2_1 _19265_ (.X(_03839_),
    .B(_07606_),
    .A(net5343));
 sg13g2_mux2_1 _19266_ (.A0(net5825),
    .A1(\fpga_top.cpu_top.csr_uimm[0] ),
    .S(net5576),
    .X(_03840_));
 sg13g2_nor2_1 _19267_ (.A(net5385),
    .B(_03840_),
    .Y(_03841_));
 sg13g2_nor3_1 _19268_ (.A(_03815_),
    .B(_03823_),
    .C(_03828_),
    .Y(_03842_));
 sg13g2_and2_1 _19269_ (.A(_03819_),
    .B(_03842_),
    .X(_03843_));
 sg13g2_nand3_1 _19270_ (.B(_03804_),
    .C(_03843_),
    .A(_03797_),
    .Y(_03844_));
 sg13g2_nor2_2 _19271_ (.A(_03800_),
    .B(_03844_),
    .Y(_03845_));
 sg13g2_nor2_2 _19272_ (.A(_03801_),
    .B(_03844_),
    .Y(_03846_));
 sg13g2_inv_4 _19273_ (.A(net4670),
    .Y(_03847_));
 sg13g2_a22oi_1 _19274_ (.Y(_03848_),
    .B1(net4670),
    .B2(net3493),
    .A2(net4673),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[0] ));
 sg13g2_nand3_1 _19275_ (.B(_03805_),
    .C(_03842_),
    .A(_03797_),
    .Y(_03849_));
 sg13g2_nor2_2 _19276_ (.A(_03819_),
    .B(_03849_),
    .Y(_03850_));
 sg13g2_a22oi_1 _19277_ (.Y(_03851_),
    .B1(net4666),
    .B2(net2147),
    .A2(net4629),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[0] ));
 sg13g2_nor2_2 _19278_ (.A(_03818_),
    .B(_03849_),
    .Y(_03852_));
 sg13g2_or4_1 _19279_ (.A(_03815_),
    .B(_03818_),
    .C(_03822_),
    .D(_03828_),
    .X(_03853_));
 sg13g2_nor2_2 _19280_ (.A(_03800_),
    .B(_03804_),
    .Y(_03854_));
 sg13g2_or2_1 _19281_ (.X(_03855_),
    .B(_03804_),
    .A(_03800_));
 sg13g2_nand2b_2 _19282_ (.Y(_03856_),
    .B(_03796_),
    .A_N(_03792_));
 sg13g2_inv_1 _19283_ (.Y(_03857_),
    .A(_03856_));
 sg13g2_nor3_2 _19284_ (.A(_03853_),
    .B(_03855_),
    .C(_03856_),
    .Y(_03858_));
 sg13g2_nand3b_1 _19285_ (.B(_03854_),
    .C(_03857_),
    .Y(_03859_),
    .A_N(_03853_));
 sg13g2_a22oi_1 _19286_ (.Y(_03860_),
    .B1(net4699),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[0] ),
    .A2(net4664),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[0] ));
 sg13g2_nand3_1 _19287_ (.B(_03851_),
    .C(_03860_),
    .A(_03848_),
    .Y(_03861_));
 sg13g2_nor2_2 _19288_ (.A(_03853_),
    .B(_03856_),
    .Y(_03862_));
 sg13g2_nor3_2 _19289_ (.A(_03853_),
    .B(_03855_),
    .C(_03856_),
    .Y(_03863_));
 sg13g2_nand2_2 _19290_ (.Y(_03864_),
    .A(_03854_),
    .B(_03862_));
 sg13g2_nor2b_1 _19291_ (.A(_03806_),
    .B_N(_03843_),
    .Y(_03865_));
 sg13g2_a22oi_1 _19292_ (.Y(_03866_),
    .B1(_03841_),
    .B2(_03861_),
    .A2(_03840_),
    .A1(net5129));
 sg13g2_nor2_2 _19293_ (.A(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .B(net5048),
    .Y(_03867_));
 sg13g2_a21oi_1 _19294_ (.A1(_03836_),
    .A2(_03866_),
    .Y(_03868_),
    .B1(_03867_));
 sg13g2_mux2_1 _19295_ (.A0(net3298),
    .A1(_03868_),
    .S(net4587),
    .X(_01142_));
 sg13g2_nor2_1 _19296_ (.A(net5576),
    .B(net5824),
    .Y(_03869_));
 sg13g2_a21oi_2 _19297_ (.B1(_03869_),
    .Y(_03870_),
    .A2(_06608_),
    .A1(net5576));
 sg13g2_nor2_1 _19298_ (.A(net5381),
    .B(_03870_),
    .Y(_03871_));
 sg13g2_nor2_2 _19299_ (.A(_03806_),
    .B(_03853_),
    .Y(_03872_));
 sg13g2_or2_1 _19300_ (.X(_03873_),
    .B(_03828_),
    .A(_03824_));
 sg13g2_a22oi_1 _19301_ (.Y(_03874_),
    .B1(net4660),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[1] ),
    .A2(net4665),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[1] ));
 sg13g2_nand2_1 _19302_ (.Y(_03875_),
    .A(_03824_),
    .B(_03874_));
 sg13g2_o21ai_1 _19303_ (.B1(_03875_),
    .Y(_03876_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[1] ),
    .A2(_03824_));
 sg13g2_a21o_1 _19304_ (.A2(net4671),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[1] ),
    .B1(net4658),
    .X(_03877_));
 sg13g2_a221oi_1 _19305_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[1] ),
    .C1(_03877_),
    .B1(net4692),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mcause[1] ),
    .Y(_03878_),
    .A2(net4670));
 sg13g2_a22oi_1 _19306_ (.Y(_03879_),
    .B1(_03876_),
    .B2(_03878_),
    .A2(net4658),
    .A1(_06878_));
 sg13g2_a22oi_1 _19307_ (.Y(_03880_),
    .B1(_03871_),
    .B2(_03879_),
    .A2(_03870_),
    .A1(net5129));
 sg13g2_nand2_1 _19308_ (.Y(_03881_),
    .A(net5047),
    .B(_03880_));
 sg13g2_o21ai_1 _19309_ (.B1(_03881_),
    .Y(_03882_),
    .A1(\fpga_top.cpu_top.csr_wdata_mon[1] ),
    .A2(net5047));
 sg13g2_nand2_1 _19310_ (.Y(_03883_),
    .A(net1451),
    .B(net4581));
 sg13g2_o21ai_1 _19311_ (.B1(_03883_),
    .Y(_01143_),
    .A1(net4581),
    .A2(_03882_));
 sg13g2_nor2_1 _19312_ (.A(net1951),
    .B(net4587),
    .Y(_03884_));
 sg13g2_mux2_1 _19313_ (.A0(net5821),
    .A1(\fpga_top.cpu_top.csr_uimm[2] ),
    .S(net5576),
    .X(_03885_));
 sg13g2_nand2_1 _19314_ (.Y(_03886_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[2] ),
    .B(net4664));
 sg13g2_a22oi_1 _19315_ (.Y(_03887_),
    .B1(net4666),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[2] ),
    .A2(net4629),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[2] ));
 sg13g2_a21oi_1 _19316_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[2] ),
    .A2(net4673),
    .Y(_03888_),
    .B1(_03846_));
 sg13g2_nand3_1 _19317_ (.B(_03887_),
    .C(_03888_),
    .A(_03886_),
    .Y(_03889_));
 sg13g2_o21ai_1 _19318_ (.B1(_03889_),
    .Y(_03890_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mcause[2] ),
    .A2(_03847_));
 sg13g2_and2_1 _19319_ (.A(_03797_),
    .B(_03854_),
    .X(_03891_));
 sg13g2_and2_1 _19320_ (.A(_03843_),
    .B(_03891_),
    .X(_03892_));
 sg13g2_a21oi_1 _19321_ (.A1(\fpga_top.cpu_top.csr_mepc_ex[2] ),
    .A2(net4686),
    .Y(_03893_),
    .B1(net4699));
 sg13g2_and3_2 _19322_ (.X(_03894_),
    .A(_03819_),
    .B(_03842_),
    .C(_03891_));
 sg13g2_a22oi_1 _19323_ (.Y(_03895_),
    .B1(_03890_),
    .B2(_03893_),
    .A2(net4693),
    .A1(_06882_));
 sg13g2_nor2_1 _19324_ (.A(net5381),
    .B(_03885_),
    .Y(_03896_));
 sg13g2_a22oi_1 _19325_ (.Y(_03897_),
    .B1(_03895_),
    .B2(_03896_),
    .A2(_03885_),
    .A1(net5129));
 sg13g2_nand2_1 _19326_ (.Y(_03898_),
    .A(net5048),
    .B(_03897_));
 sg13g2_o21ai_1 _19327_ (.B1(_03898_),
    .Y(_03899_),
    .A1(net5664),
    .A2(net5048));
 sg13g2_a21oi_1 _19328_ (.A1(_03834_),
    .A2(_03899_),
    .Y(_01144_),
    .B1(_03884_));
 sg13g2_nand2_1 _19329_ (.Y(_03900_),
    .A(net1511),
    .B(net4581));
 sg13g2_mux2_1 _19330_ (.A0(net5818),
    .A1(\fpga_top.cpu_top.csr_uimm[3] ),
    .S(net5577),
    .X(_03901_));
 sg13g2_nand2_1 _19331_ (.Y(_03902_),
    .A(_03805_),
    .B(_03857_));
 sg13g2_nand3_1 _19332_ (.B(_03843_),
    .C(_03857_),
    .A(_03805_),
    .Y(_03903_));
 sg13g2_inv_1 _19333_ (.Y(_03904_),
    .A(_03903_));
 sg13g2_nor2b_2 _19334_ (.A(_07039_),
    .B_N(_07297_),
    .Y(_03905_));
 sg13g2_nor3_1 _19335_ (.A(net5308),
    .B(_07289_),
    .C(_03905_),
    .Y(_03906_));
 sg13g2_nor2_1 _19336_ (.A(net5571),
    .B(net5570),
    .Y(_03907_));
 sg13g2_and4_1 _19337_ (.A(\fpga_top.cpu_top.br_ofs[5] ),
    .B(_07288_),
    .C(_03812_),
    .D(_03907_),
    .X(_03908_));
 sg13g2_a221oi_1 _19338_ (.B2(_03908_),
    .C1(net5293),
    .B1(_07575_),
    .A1(_07293_),
    .Y(_03909_),
    .A2(_07296_));
 sg13g2_nor2_1 _19339_ (.A(\fpga_top.cpu_top.br_ofs[2] ),
    .B(\fpga_top.cpu_top.br_ofs[1] ),
    .Y(_03910_));
 sg13g2_nor3_1 _19340_ (.A(\fpga_top.cpu_top.br_ofs[11] ),
    .B(\fpga_top.cpu_top.br_ofs[3] ),
    .C(\fpga_top.cpu_top.br_ofs[4] ),
    .Y(_03911_));
 sg13g2_nand3_1 _19341_ (.B(_03910_),
    .C(_03911_),
    .A(_07037_),
    .Y(_03912_));
 sg13g2_nor4_2 _19342_ (.A(_07295_),
    .B(_07576_),
    .C(_10624_),
    .Y(_03913_),
    .D(_03912_));
 sg13g2_nor2_1 _19343_ (.A(\fpga_top.cpu_top.alui_shamt[2] ),
    .B(\fpga_top.cpu_top.alui_shamt[3] ),
    .Y(_03914_));
 sg13g2_nand3_1 _19344_ (.B(_06575_),
    .C(_03914_),
    .A(_06559_),
    .Y(_03915_));
 sg13g2_nor4_1 _19345_ (.A(\fpga_top.cpu_top.alui_shamt[2] ),
    .B(\fpga_top.cpu_top.alui_shamt[1] ),
    .C(net5572),
    .D(\fpga_top.cpu_top.alui_shamt[3] ),
    .Y(_03916_));
 sg13g2_nor2_2 _19346_ (.A(net5572),
    .B(_03915_),
    .Y(_03917_));
 sg13g2_nor4_1 _19347_ (.A(\fpga_top.cpu_top.br_ofs[8] ),
    .B(\fpga_top.cpu_top.br_ofs[9] ),
    .C(\fpga_top.cpu_top.br_ofs[10] ),
    .D(net5569),
    .Y(_03918_));
 sg13g2_nand2b_1 _19348_ (.Y(_03919_),
    .B(_03918_),
    .A_N(_07078_));
 sg13g2_nor4_1 _19349_ (.A(_07031_),
    .B(_10624_),
    .C(_03912_),
    .D(_03919_),
    .Y(_03920_));
 sg13g2_nor3_1 _19350_ (.A(_07295_),
    .B(_10624_),
    .C(_03912_),
    .Y(_03921_));
 sg13g2_nor3_1 _19351_ (.A(\fpga_top.cpu_top.br_ofs[3] ),
    .B(\fpga_top.cpu_top.alui_shamt[4] ),
    .C(\fpga_top.cpu_top.br_ofs[4] ),
    .Y(_03922_));
 sg13g2_nor3_1 _19352_ (.A(net5571),
    .B(\fpga_top.cpu_top.br_ofs[5] ),
    .C(\fpga_top.cpu_top.br_ofs[11] ),
    .Y(_03923_));
 sg13g2_nand3_1 _19353_ (.B(_03910_),
    .C(_03923_),
    .A(_06554_),
    .Y(_03924_));
 sg13g2_nand4_1 _19354_ (.B(_03916_),
    .C(_03918_),
    .A(_07037_),
    .Y(_03925_),
    .D(_03922_));
 sg13g2_nor4_1 _19355_ (.A(_07301_),
    .B(_10624_),
    .C(_03924_),
    .D(_03925_),
    .Y(_03926_));
 sg13g2_nor4_2 _19356_ (.A(_08276_),
    .B(_03913_),
    .C(_03920_),
    .Y(_03927_),
    .D(_03926_));
 sg13g2_and4_1 _19357_ (.A(net5207),
    .B(net5205),
    .C(_03906_),
    .D(_03909_),
    .X(_03928_));
 sg13g2_nand2_2 _19358_ (.Y(_03929_),
    .A(_03927_),
    .B(_03928_));
 sg13g2_nor2_1 _19359_ (.A(_03903_),
    .B(_03929_),
    .Y(_03930_));
 sg13g2_a21oi_1 _19360_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[3] ),
    .A2(net4628),
    .Y(_03931_),
    .B1(_03930_));
 sg13g2_nor2_1 _19361_ (.A(_03853_),
    .B(_03902_),
    .Y(_03932_));
 sg13g2_nor2b_2 _19362_ (.A(_03853_),
    .B_N(_03891_),
    .Y(_03933_));
 sg13g2_or2_1 _19363_ (.X(_03934_),
    .B(_03933_),
    .A(net4659));
 sg13g2_a22oi_1 _19364_ (.Y(_03935_),
    .B1(net4660),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[3] ),
    .A2(net4665),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[3] ));
 sg13g2_and2_1 _19365_ (.A(_03805_),
    .B(_03862_),
    .X(_03936_));
 sg13g2_nand2_1 _19366_ (.Y(_03937_),
    .A(\fpga_top.cpu_top.csr_msie ),
    .B(_03936_));
 sg13g2_a21oi_1 _19367_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[3] ),
    .A2(net4671),
    .Y(_03938_),
    .B1(net4670));
 sg13g2_nand4_1 _19368_ (.B(_03935_),
    .C(_03937_),
    .A(_03931_),
    .Y(_03939_),
    .D(_03938_));
 sg13g2_o21ai_1 _19369_ (.B1(_03939_),
    .Y(_03940_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mcause[3] ),
    .A2(_03847_));
 sg13g2_a21oi_1 _19370_ (.A1(\fpga_top.cpu_top.csr_mepc_ex[3] ),
    .A2(_03894_),
    .Y(_03941_),
    .B1(net4692));
 sg13g2_a221oi_1 _19371_ (.B2(_03941_),
    .C1(_03934_),
    .B1(_03940_),
    .A1(_06884_),
    .Y(_03942_),
    .A2(net4692));
 sg13g2_a21oi_2 _19372_ (.B1(_03942_),
    .Y(_03943_),
    .A2(net4659),
    .A1(\fpga_top.cpu_top.csr_rmie ));
 sg13g2_nor3_1 _19373_ (.A(net5381),
    .B(_03901_),
    .C(_03943_),
    .Y(_03944_));
 sg13g2_a21o_2 _19374_ (.A2(_03901_),
    .A1(net5129),
    .B1(_03944_),
    .X(_03945_));
 sg13g2_inv_1 _19375_ (.Y(_03946_),
    .A(_03945_));
 sg13g2_nand2_2 _19376_ (.Y(_03947_),
    .A(_06789_),
    .B(net5134));
 sg13g2_o21ai_1 _19377_ (.B1(_03947_),
    .Y(_03948_),
    .A1(_03837_),
    .A2(_03945_));
 sg13g2_o21ai_1 _19378_ (.B1(_03900_),
    .Y(_01145_),
    .A1(net4581),
    .A2(_03948_));
 sg13g2_nand2_1 _19379_ (.Y(_03949_),
    .A(net1571),
    .B(net4581));
 sg13g2_nand3_1 _19380_ (.B(net5809),
    .C(net5129),
    .A(net5379),
    .Y(_03950_));
 sg13g2_a21o_1 _19381_ (.A2(net5809),
    .A1(net5379),
    .B1(net5381),
    .X(_03951_));
 sg13g2_nand2_1 _19382_ (.Y(_03952_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[6] ),
    .B(net4665));
 sg13g2_a22oi_1 _19383_ (.Y(_03953_),
    .B1(net4686),
    .B2(\fpga_top.cpu_top.csr_mepc_ex[6] ),
    .A2(net4664),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[6] ));
 sg13g2_a221oi_1 _19384_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_mtval[6] ),
    .C1(net4699),
    .B1(net4671),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[6] ),
    .Y(_03954_),
    .A2(net4628));
 sg13g2_nand3_1 _19385_ (.B(_03953_),
    .C(_03954_),
    .A(_03952_),
    .Y(_03955_));
 sg13g2_o21ai_1 _19386_ (.B1(_03955_),
    .Y(_03956_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[6] ),
    .A2(net4695));
 sg13g2_o21ai_1 _19387_ (.B1(_03950_),
    .Y(_03957_),
    .A1(_03951_),
    .A2(_03956_));
 sg13g2_inv_1 _19388_ (.Y(_03958_),
    .A(_03957_));
 sg13g2_nand2_2 _19389_ (.Y(_03959_),
    .A(_06790_),
    .B(net5134));
 sg13g2_o21ai_1 _19390_ (.B1(_03959_),
    .Y(_03960_),
    .A1(_03837_),
    .A2(_03957_));
 sg13g2_o21ai_1 _19391_ (.B1(_03949_),
    .Y(_01146_),
    .A1(net4581),
    .A2(_03960_));
 sg13g2_nand2_1 _19392_ (.Y(_03961_),
    .A(net5379),
    .B(net5805));
 sg13g2_a22oi_1 _19393_ (.Y(_03962_),
    .B1(net4660),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[7] ),
    .A2(net4665),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[7] ));
 sg13g2_a221oi_1 _19394_ (.B2(\fpga_top.cpu_top.csr_mtie ),
    .C1(net4628),
    .B1(_03932_),
    .A1(\fpga_top.cpu_top.execution.csr_array.frc_cntr_val_leq ),
    .Y(_03963_),
    .A2(_03904_));
 sg13g2_a22oi_1 _19395_ (.Y(_03964_),
    .B1(_03962_),
    .B2(_03963_),
    .A2(net4628),
    .A1(_06893_));
 sg13g2_nand2b_1 _19396_ (.Y(_03965_),
    .B(net4671),
    .A_N(\fpga_top.cpu_top.execution.csr_array.csr_mtval[7] ));
 sg13g2_o21ai_1 _19397_ (.B1(_03965_),
    .Y(_03966_),
    .A1(net4671),
    .A2(_03964_));
 sg13g2_a21oi_1 _19398_ (.A1(\fpga_top.cpu_top.csr_mepc_ex[7] ),
    .A2(net4686),
    .Y(_03967_),
    .B1(net4692));
 sg13g2_a22oi_1 _19399_ (.Y(_03968_),
    .B1(_03966_),
    .B2(_03967_),
    .A2(net4692),
    .A1(_06894_));
 sg13g2_a21o_2 _19400_ (.A2(net4658),
    .A1(net2066),
    .B1(_03968_),
    .X(_03969_));
 sg13g2_nand3_1 _19401_ (.B(_03961_),
    .C(_03969_),
    .A(net5581),
    .Y(_03970_));
 sg13g2_o21ai_1 _19402_ (.B1(_03970_),
    .Y(_03971_),
    .A1(_03838_),
    .A2(_03961_));
 sg13g2_inv_1 _19403_ (.Y(_03972_),
    .A(_03971_));
 sg13g2_a221oi_1 _19404_ (.B2(_03971_),
    .C1(net4581),
    .B1(_03836_),
    .A1(net5657),
    .Y(_03973_),
    .A2(net5134));
 sg13g2_a21oi_1 _19405_ (.A1(_06893_),
    .A2(net4582),
    .Y(_01147_),
    .B1(_03973_));
 sg13g2_nor2_2 _19406_ (.A(net5577),
    .B(_06566_),
    .Y(_03974_));
 sg13g2_nor2_1 _19407_ (.A(net5381),
    .B(_03974_),
    .Y(_03975_));
 sg13g2_a21oi_1 _19408_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[8] ),
    .A2(net4628),
    .Y(_03976_),
    .B1(net4672));
 sg13g2_a22oi_1 _19409_ (.Y(_03977_),
    .B1(net4660),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[8] ),
    .A2(net4666),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[8] ));
 sg13g2_a22oi_1 _19410_ (.Y(_03978_),
    .B1(_03976_),
    .B2(_03977_),
    .A2(net4672),
    .A1(_06899_));
 sg13g2_a21oi_1 _19411_ (.A1(\fpga_top.cpu_top.csr_mepc_ex[8] ),
    .A2(_03894_),
    .Y(_03979_),
    .B1(_03978_));
 sg13g2_a21oi_1 _19412_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[8] ),
    .A2(net4692),
    .Y(_03980_),
    .B1(_03934_));
 sg13g2_a22oi_1 _19413_ (.Y(_03981_),
    .B1(_03979_),
    .B2(_03980_),
    .A2(net4659),
    .A1(_06901_));
 sg13g2_a22oi_1 _19414_ (.Y(_03982_),
    .B1(_03975_),
    .B2(_03981_),
    .A2(_03974_),
    .A1(net5129));
 sg13g2_nand2_2 _19415_ (.Y(_03983_),
    .A(net5047),
    .B(_03982_));
 sg13g2_nand2b_2 _19416_ (.Y(_03984_),
    .B(net5136),
    .A_N(net5655));
 sg13g2_nand3_1 _19417_ (.B(_03983_),
    .C(_03984_),
    .A(net4587),
    .Y(_03985_));
 sg13g2_o21ai_1 _19418_ (.B1(_03985_),
    .Y(_01148_),
    .A1(_06898_),
    .A2(net4587));
 sg13g2_nand2_1 _19419_ (.Y(_03986_),
    .A(net1450),
    .B(net4582));
 sg13g2_o21ai_1 _19420_ (.B1(net4587),
    .Y(_03987_),
    .A1(net5653),
    .A2(net5049));
 sg13g2_nand2_2 _19421_ (.Y(_03988_),
    .A(net5380),
    .B(net5801));
 sg13g2_nor2_1 _19422_ (.A(_03838_),
    .B(_03988_),
    .Y(_03989_));
 sg13g2_nand2_1 _19423_ (.Y(_03990_),
    .A(net5582),
    .B(_03988_));
 sg13g2_nand2_1 _19424_ (.Y(_03991_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[9] ),
    .B(net4669));
 sg13g2_a22oi_1 _19425_ (.Y(_03992_),
    .B1(_03892_),
    .B2(\fpga_top.cpu_top.csr_mepc_ex[9] ),
    .A2(net4664),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[9] ));
 sg13g2_a221oi_1 _19426_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_mtval[9] ),
    .C1(net4699),
    .B1(net4673),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[9] ),
    .Y(_03993_),
    .A2(net4629));
 sg13g2_nand3_1 _19427_ (.B(_03992_),
    .C(_03993_),
    .A(_03991_),
    .Y(_03994_));
 sg13g2_o21ai_1 _19428_ (.B1(_03994_),
    .Y(_03995_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[9] ),
    .A2(net4695));
 sg13g2_nor2_1 _19429_ (.A(_03990_),
    .B(_03995_),
    .Y(_03996_));
 sg13g2_nor2_1 _19430_ (.A(_03989_),
    .B(_03996_),
    .Y(_03997_));
 sg13g2_or2_1 _19431_ (.X(_03998_),
    .B(_03996_),
    .A(_03989_));
 sg13g2_nor2_1 _19432_ (.A(net5139),
    .B(_03998_),
    .Y(_03999_));
 sg13g2_o21ai_1 _19433_ (.B1(_03986_),
    .Y(_01149_),
    .A1(_03987_),
    .A2(_03999_));
 sg13g2_nor2_2 _19434_ (.A(net5575),
    .B(_06571_),
    .Y(_04000_));
 sg13g2_nand2_1 _19435_ (.Y(_04001_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[10] ),
    .B(net4630));
 sg13g2_a22oi_1 _19436_ (.Y(_04002_),
    .B1(net4662),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[10] ),
    .A2(net4667),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[10] ));
 sg13g2_a221oi_1 _19437_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[10] ),
    .C1(net4696),
    .B1(net4687),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[10] ),
    .Y(_04003_),
    .A2(net4674));
 sg13g2_nand3_1 _19438_ (.B(_04002_),
    .C(_04003_),
    .A(_04001_),
    .Y(_04004_));
 sg13g2_o21ai_1 _19439_ (.B1(_04004_),
    .Y(_04005_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[10] ),
    .A2(net4695));
 sg13g2_nor3_1 _19440_ (.A(net5382),
    .B(_04000_),
    .C(_04005_),
    .Y(_04006_));
 sg13g2_a21oi_2 _19441_ (.B1(_04006_),
    .Y(_04007_),
    .A2(_04000_),
    .A1(net5130));
 sg13g2_and2_1 _19442_ (.A(net5059),
    .B(_04007_),
    .X(_04008_));
 sg13g2_nor2_2 _19443_ (.A(\fpga_top.cpu_start_adr[10] ),
    .B(net5059),
    .Y(_04009_));
 sg13g2_nor3_1 _19444_ (.A(net4585),
    .B(_04008_),
    .C(_04009_),
    .Y(_04010_));
 sg13g2_a21o_1 _19445_ (.A2(net4583),
    .A1(net2343),
    .B1(_04010_),
    .X(_01150_));
 sg13g2_nand2_1 _19446_ (.Y(_04011_),
    .A(net5379),
    .B(net5797));
 sg13g2_a22oi_1 _19447_ (.Y(_04012_),
    .B1(net4660),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[11] ),
    .A2(net4665),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[11] ));
 sg13g2_a221oi_1 _19448_ (.B2(\fpga_top.cpu_top.csr_meie ),
    .C1(net4628),
    .B1(_03932_),
    .A1(\fpga_top.cpu_top.execution.csr_array.g_interrupt ),
    .Y(_04013_),
    .A2(_03904_));
 sg13g2_a22oi_1 _19449_ (.Y(_04014_),
    .B1(_04012_),
    .B2(_04013_),
    .A2(net4628),
    .A1(_06904_));
 sg13g2_nand2b_1 _19450_ (.Y(_04015_),
    .B(net4671),
    .A_N(\fpga_top.cpu_top.execution.csr_array.csr_mtval[11] ));
 sg13g2_o21ai_1 _19451_ (.B1(_04015_),
    .Y(_04016_),
    .A1(net4671),
    .A2(_04014_));
 sg13g2_a21oi_1 _19452_ (.A1(\fpga_top.cpu_top.csr_mepc_ex[11] ),
    .A2(net4686),
    .Y(_04017_),
    .B1(net4693));
 sg13g2_a22oi_1 _19453_ (.Y(_04018_),
    .B1(_04016_),
    .B2(_04017_),
    .A2(net4693),
    .A1(_06905_));
 sg13g2_a21oi_2 _19454_ (.B1(_04018_),
    .Y(_04019_),
    .A2(net4658),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mpp[0] ));
 sg13g2_nand3b_1 _19455_ (.B(net5581),
    .C(_04011_),
    .Y(_04020_),
    .A_N(_04019_));
 sg13g2_o21ai_1 _19456_ (.B1(_04020_),
    .Y(_04021_),
    .A1(_03838_),
    .A2(_04011_));
 sg13g2_inv_1 _19457_ (.Y(_04022_),
    .A(_04021_));
 sg13g2_a221oi_1 _19458_ (.B2(_04021_),
    .C1(net4581),
    .B1(_03836_),
    .A1(\fpga_top.cpu_start_adr[11] ),
    .Y(_04023_),
    .A2(net5134));
 sg13g2_a21oi_1 _19459_ (.A1(_06904_),
    .A2(net4582),
    .Y(_01151_),
    .B1(_04023_));
 sg13g2_nor2_1 _19460_ (.A(net1796),
    .B(net4587),
    .Y(_04024_));
 sg13g2_nor2b_1 _19461_ (.A(net5576),
    .B_N(net5795),
    .Y(_04025_));
 sg13g2_or2_1 _19462_ (.X(_04026_),
    .B(_03824_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[12] ));
 sg13g2_nand2_1 _19463_ (.Y(_04027_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[12] ),
    .B(net4664));
 sg13g2_nand2_1 _19464_ (.Y(_04028_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[12] ),
    .B(net4665));
 sg13g2_nand3_1 _19465_ (.B(_04027_),
    .C(_04028_),
    .A(_03824_),
    .Y(_04029_));
 sg13g2_a22oi_1 _19466_ (.Y(_04030_),
    .B1(_04026_),
    .B2(_04029_),
    .A2(net4672),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[12] ));
 sg13g2_a21oi_1 _19467_ (.A1(\fpga_top.cpu_top.csr_mepc_ex[12] ),
    .A2(net4686),
    .Y(_04031_),
    .B1(net4699));
 sg13g2_a221oi_1 _19468_ (.B2(_04031_),
    .C1(net4659),
    .B1(_04030_),
    .A1(_06906_),
    .Y(_04032_),
    .A2(net4699));
 sg13g2_a21oi_2 _19469_ (.B1(_04032_),
    .Y(_04033_),
    .A2(net4658),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mpp[1] ));
 sg13g2_nor3_1 _19470_ (.A(net5382),
    .B(_04025_),
    .C(_04033_),
    .Y(_04034_));
 sg13g2_a21oi_2 _19471_ (.B1(_04034_),
    .Y(_04035_),
    .A2(_04025_),
    .A1(net5130));
 sg13g2_nor2_1 _19472_ (.A(_03837_),
    .B(_04035_),
    .Y(_04036_));
 sg13g2_a21oi_1 _19473_ (.A1(\fpga_top.cpu_start_adr[12] ),
    .A2(net5135),
    .Y(_04037_),
    .B1(_04036_));
 sg13g2_a21oi_1 _19474_ (.A1(net4587),
    .A2(_04037_),
    .Y(_01152_),
    .B1(_04024_));
 sg13g2_a21oi_1 _19475_ (.A1(\fpga_top.cpu_start_adr[13] ),
    .A2(net5140),
    .Y(_04038_),
    .B1(net4586));
 sg13g2_nor2b_1 _19476_ (.A(net5580),
    .B_N(net5792),
    .Y(_04039_));
 sg13g2_nand2_1 _19477_ (.Y(_04040_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[13] ),
    .B(net4664));
 sg13g2_a22oi_1 _19478_ (.Y(_04041_),
    .B1(net4669),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[13] ),
    .A2(net4632),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[13] ));
 sg13g2_a221oi_1 _19479_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[13] ),
    .C1(net4699),
    .B1(net4686),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[13] ),
    .Y(_04042_),
    .A2(net4676));
 sg13g2_nand3_1 _19480_ (.B(_04041_),
    .C(_04042_),
    .A(_04040_),
    .Y(_04043_));
 sg13g2_o21ai_1 _19481_ (.B1(_04043_),
    .Y(_04044_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[13] ),
    .A2(_03864_));
 sg13g2_nor3_1 _19482_ (.A(net5382),
    .B(_04039_),
    .C(_04044_),
    .Y(_04045_));
 sg13g2_a21oi_2 _19483_ (.B1(_04045_),
    .Y(_04046_),
    .A2(_04039_),
    .A1(net5130));
 sg13g2_o21ai_1 _19484_ (.B1(_04038_),
    .Y(_04047_),
    .A1(net5140),
    .A2(_04046_));
 sg13g2_o21ai_1 _19485_ (.B1(_04047_),
    .Y(_04048_),
    .A1(net3820),
    .A2(net4589));
 sg13g2_inv_1 _19486_ (.Y(_01153_),
    .A(_04048_));
 sg13g2_nand2_1 _19487_ (.Y(_04049_),
    .A(net1479),
    .B(net4582));
 sg13g2_o21ai_1 _19488_ (.B1(net4587),
    .Y(_04050_),
    .A1(net5650),
    .A2(net5049));
 sg13g2_nand2_2 _19489_ (.Y(_04051_),
    .A(net5380),
    .B(net5790));
 sg13g2_nor2_1 _19490_ (.A(_03838_),
    .B(_04051_),
    .Y(_04052_));
 sg13g2_nand2_1 _19491_ (.Y(_04053_),
    .A(net5582),
    .B(_04051_));
 sg13g2_nand2_1 _19492_ (.Y(_04054_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[14] ),
    .B(net4664));
 sg13g2_a22oi_1 _19493_ (.Y(_04055_),
    .B1(net4686),
    .B2(\fpga_top.cpu_top.csr_mepc_ex[14] ),
    .A2(net4666),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[14] ));
 sg13g2_a221oi_1 _19494_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_mtval[14] ),
    .C1(net4699),
    .B1(net4673),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[14] ),
    .Y(_04056_),
    .A2(net4629));
 sg13g2_nand3_1 _19495_ (.B(_04055_),
    .C(_04056_),
    .A(_04054_),
    .Y(_04057_));
 sg13g2_o21ai_1 _19496_ (.B1(_04057_),
    .Y(_04058_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[14] ),
    .A2(net4695));
 sg13g2_nor2_1 _19497_ (.A(_04053_),
    .B(_04058_),
    .Y(_04059_));
 sg13g2_nor2_2 _19498_ (.A(_04052_),
    .B(_04059_),
    .Y(_04060_));
 sg13g2_nor3_1 _19499_ (.A(net5139),
    .B(_04052_),
    .C(_04059_),
    .Y(_04061_));
 sg13g2_o21ai_1 _19500_ (.B1(_04049_),
    .Y(_01154_),
    .A1(_04050_),
    .A2(_04061_));
 sg13g2_nor2b_1 _19501_ (.A(net5580),
    .B_N(net5789),
    .Y(_04062_));
 sg13g2_nand2_1 _19502_ (.Y(_04063_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[15] ),
    .B(net4632));
 sg13g2_a22oi_1 _19503_ (.Y(_04064_),
    .B1(net4663),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[15] ),
    .A2(net4669),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[15] ));
 sg13g2_a221oi_1 _19504_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[15] ),
    .C1(net4698),
    .B1(net4689),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[15] ),
    .Y(_04065_),
    .A2(net4676));
 sg13g2_nand3_1 _19505_ (.B(_04064_),
    .C(_04065_),
    .A(_04063_),
    .Y(_04066_));
 sg13g2_o21ai_1 _19506_ (.B1(_04066_),
    .Y(_04067_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[15] ),
    .A2(_03859_));
 sg13g2_nor3_1 _19507_ (.A(net5381),
    .B(_04062_),
    .C(_04067_),
    .Y(_04068_));
 sg13g2_a21oi_2 _19508_ (.B1(_04068_),
    .Y(_04069_),
    .A2(_04062_),
    .A1(net5130));
 sg13g2_o21ai_1 _19509_ (.B1(net4589),
    .Y(_04070_),
    .A1(\fpga_top.cpu_start_adr[15] ),
    .A2(net5055));
 sg13g2_a21oi_1 _19510_ (.A1(net5055),
    .A2(_04069_),
    .Y(_04071_),
    .B1(_04070_));
 sg13g2_a21o_1 _19511_ (.A2(net4586),
    .A1(net1950),
    .B1(_04071_),
    .X(_01155_));
 sg13g2_nand2_1 _19512_ (.Y(_04072_),
    .A(net1437),
    .B(net4586));
 sg13g2_o21ai_1 _19513_ (.B1(net4589),
    .Y(_04073_),
    .A1(net5649),
    .A2(net5055));
 sg13g2_nand2_1 _19514_ (.Y(_04074_),
    .A(net5380),
    .B(net5786));
 sg13g2_nor2_1 _19515_ (.A(_03838_),
    .B(_04074_),
    .Y(_04075_));
 sg13g2_and2_1 _19516_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[16] ),
    .B(net4663),
    .X(_04076_));
 sg13g2_a221oi_1 _19517_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[16] ),
    .C1(_04076_),
    .B1(net4689),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[16] ),
    .Y(_04077_),
    .A2(net4632));
 sg13g2_a221oi_1 _19518_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[16] ),
    .C1(net4698),
    .B1(net4669),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[16] ),
    .Y(_04078_),
    .A2(net4676));
 sg13g2_a22oi_1 _19519_ (.Y(_04079_),
    .B1(_04077_),
    .B2(_04078_),
    .A2(net4694),
    .A1(_06909_));
 sg13g2_and3_1 _19520_ (.X(_04080_),
    .A(net5582),
    .B(_04074_),
    .C(_04079_));
 sg13g2_or2_1 _19521_ (.X(_04081_),
    .B(_04080_),
    .A(_04075_));
 sg13g2_nor2_1 _19522_ (.A(net5141),
    .B(_04081_),
    .Y(_04082_));
 sg13g2_o21ai_1 _19523_ (.B1(_04072_),
    .Y(_01156_),
    .A1(_04073_),
    .A2(_04082_));
 sg13g2_nand2_1 _19524_ (.Y(_04083_),
    .A(net1436),
    .B(net4585));
 sg13g2_o21ai_1 _19525_ (.B1(net4588),
    .Y(_04084_),
    .A1(net5648),
    .A2(net5058));
 sg13g2_nor2b_1 _19526_ (.A(net5578),
    .B_N(net5785),
    .Y(_04085_));
 sg13g2_and2_1 _19527_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[17] ),
    .B(net4667),
    .X(_04086_));
 sg13g2_a221oi_1 _19528_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[17] ),
    .C1(_04086_),
    .B1(net4662),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[17] ),
    .Y(_04087_),
    .A2(net4630));
 sg13g2_a221oi_1 _19529_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[17] ),
    .C1(net4696),
    .B1(net4689),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[17] ),
    .Y(_04088_),
    .A2(net4674));
 sg13g2_a22oi_1 _19530_ (.Y(_04089_),
    .B1(_04087_),
    .B2(_04088_),
    .A2(net4694),
    .A1(_06911_));
 sg13g2_nor2_1 _19531_ (.A(net5383),
    .B(_04085_),
    .Y(_04090_));
 sg13g2_a22oi_1 _19532_ (.Y(_04091_),
    .B1(_04089_),
    .B2(_04090_),
    .A2(_04085_),
    .A1(net5131));
 sg13g2_and2_1 _19533_ (.A(net5060),
    .B(_04091_),
    .X(_04092_));
 sg13g2_o21ai_1 _19534_ (.B1(_04083_),
    .Y(_01157_),
    .A1(_04084_),
    .A2(_04092_));
 sg13g2_nor2b_1 _19535_ (.A(net5578),
    .B_N(\fpga_top.cpu_top.execution.csr_array.rs1_sel[18] ),
    .Y(_04093_));
 sg13g2_and2_1 _19536_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[18] ),
    .B(net4669),
    .X(_04094_));
 sg13g2_a221oi_1 _19537_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[18] ),
    .C1(_04094_),
    .B1(net4689),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[18] ),
    .Y(_04095_),
    .A2(net4632));
 sg13g2_a221oi_1 _19538_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[18] ),
    .C1(net4698),
    .B1(net4663),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[18] ),
    .Y(_04096_),
    .A2(net4676));
 sg13g2_a22oi_1 _19539_ (.Y(_04097_),
    .B1(_04095_),
    .B2(_04096_),
    .A2(net4694),
    .A1(_06912_));
 sg13g2_nor2_1 _19540_ (.A(net5383),
    .B(_04093_),
    .Y(_04098_));
 sg13g2_a22oi_1 _19541_ (.Y(_04099_),
    .B1(_04097_),
    .B2(_04098_),
    .A2(_04093_),
    .A1(net5133));
 sg13g2_o21ai_1 _19542_ (.B1(net4588),
    .Y(_04100_),
    .A1(net5647),
    .A2(net5055));
 sg13g2_a21oi_1 _19543_ (.A1(net5055),
    .A2(_04099_),
    .Y(_04101_),
    .B1(_04100_));
 sg13g2_a21o_1 _19544_ (.A2(net4586),
    .A1(net1985),
    .B1(_04101_),
    .X(_01158_));
 sg13g2_nor2b_1 _19545_ (.A(net5579),
    .B_N(net5780),
    .Y(_04102_));
 sg13g2_nand2_1 _19546_ (.Y(_04103_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[19] ),
    .B(net4630));
 sg13g2_a22oi_1 _19547_ (.Y(_04104_),
    .B1(net4662),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[19] ),
    .A2(net4667),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[19] ));
 sg13g2_a221oi_1 _19548_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[19] ),
    .C1(net4697),
    .B1(net4688),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[19] ),
    .Y(_04105_),
    .A2(net4674));
 sg13g2_nand3_1 _19549_ (.B(_04104_),
    .C(_04105_),
    .A(_04103_),
    .Y(_04106_));
 sg13g2_o21ai_1 _19550_ (.B1(_04106_),
    .Y(_04107_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[19] ),
    .A2(net4695));
 sg13g2_nor3_1 _19551_ (.A(net5384),
    .B(_04102_),
    .C(_04107_),
    .Y(_04108_));
 sg13g2_a21oi_2 _19552_ (.B1(_04108_),
    .Y(_04109_),
    .A2(_04102_),
    .A1(net5131));
 sg13g2_nand2_2 _19553_ (.Y(_04110_),
    .A(net5056),
    .B(_04109_));
 sg13g2_nor2_2 _19554_ (.A(\fpga_top.cpu_start_adr[19] ),
    .B(net5058),
    .Y(_04111_));
 sg13g2_nor2_1 _19555_ (.A(net4583),
    .B(_04111_),
    .Y(_04112_));
 sg13g2_a22oi_1 _19556_ (.Y(_04113_),
    .B1(_04110_),
    .B2(_04112_),
    .A2(net4583),
    .A1(net3098));
 sg13g2_inv_1 _19557_ (.Y(_01159_),
    .A(_04113_));
 sg13g2_a21oi_1 _19558_ (.A1(net5646),
    .A2(net5142),
    .Y(_04114_),
    .B1(net4585));
 sg13g2_nor2_1 _19559_ (.A(net5579),
    .B(_06578_),
    .Y(_04115_));
 sg13g2_nand2_1 _19560_ (.Y(_04116_),
    .A(\fpga_top.cpu_top.csr_mepc_ex[20] ),
    .B(net4687));
 sg13g2_a22oi_1 _19561_ (.Y(_04117_),
    .B1(net4662),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[20] ),
    .A2(net4631),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[20] ));
 sg13g2_a221oi_1 _19562_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[20] ),
    .C1(net4696),
    .B1(net4668),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[20] ),
    .Y(_04118_),
    .A2(net4674));
 sg13g2_nand3_1 _19563_ (.B(_04117_),
    .C(_04118_),
    .A(_04116_),
    .Y(_04119_));
 sg13g2_o21ai_1 _19564_ (.B1(_04119_),
    .Y(_04120_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[20] ),
    .A2(net4695));
 sg13g2_nor3_1 _19565_ (.A(net5383),
    .B(_04115_),
    .C(_04120_),
    .Y(_04121_));
 sg13g2_a21oi_2 _19566_ (.B1(_04121_),
    .Y(_04122_),
    .A2(_04115_),
    .A1(net5131));
 sg13g2_o21ai_1 _19567_ (.B1(_04114_),
    .Y(_04123_),
    .A1(net5142),
    .A2(_04122_));
 sg13g2_o21ai_1 _19568_ (.B1(_04123_),
    .Y(_04124_),
    .A1(net3810),
    .A2(net4589));
 sg13g2_inv_1 _19569_ (.Y(_01160_),
    .A(_04124_));
 sg13g2_nor2b_1 _19570_ (.A(net5578),
    .B_N(net5776),
    .Y(_04125_));
 sg13g2_nand2_1 _19571_ (.Y(_04126_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[21] ),
    .B(net4662));
 sg13g2_a22oi_1 _19572_ (.Y(_04127_),
    .B1(net4688),
    .B2(\fpga_top.cpu_top.csr_mepc_ex[21] ),
    .A2(net4630),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[21] ));
 sg13g2_a221oi_1 _19573_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[21] ),
    .C1(net4697),
    .B1(net4667),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[21] ),
    .Y(_04128_),
    .A2(net4675));
 sg13g2_nand3_1 _19574_ (.B(_04127_),
    .C(_04128_),
    .A(_04126_),
    .Y(_04129_));
 sg13g2_o21ai_1 _19575_ (.B1(_04129_),
    .Y(_04130_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ),
    .A2(_03859_));
 sg13g2_nor3_1 _19576_ (.A(net5384),
    .B(_04125_),
    .C(_04130_),
    .Y(_04131_));
 sg13g2_a21oi_2 _19577_ (.B1(_04131_),
    .Y(_04132_),
    .A2(_04125_),
    .A1(net5132));
 sg13g2_and2_1 _19578_ (.A(net5060),
    .B(_04132_),
    .X(_04133_));
 sg13g2_nor2_2 _19579_ (.A(net5645),
    .B(net5060),
    .Y(_04134_));
 sg13g2_nor3_1 _19580_ (.A(net4583),
    .B(_04133_),
    .C(_04134_),
    .Y(_04135_));
 sg13g2_a21o_1 _19581_ (.A2(net4583),
    .A1(net2214),
    .B1(_04135_),
    .X(_01161_));
 sg13g2_a21oi_1 _19582_ (.A1(net5643),
    .A2(net5142),
    .Y(_04136_),
    .B1(net4585));
 sg13g2_nor2_1 _19583_ (.A(net5578),
    .B(_06579_),
    .Y(_04137_));
 sg13g2_nand2_1 _19584_ (.Y(_04138_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[22] ),
    .B(net4631));
 sg13g2_a22oi_1 _19585_ (.Y(_04139_),
    .B1(net4661),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[22] ),
    .A2(net4668),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[22] ));
 sg13g2_a221oi_1 _19586_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[22] ),
    .C1(net4696),
    .B1(net4687),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[22] ),
    .Y(_04140_),
    .A2(net4675));
 sg13g2_nand3_1 _19587_ (.B(_04139_),
    .C(_04140_),
    .A(_04138_),
    .Y(_04141_));
 sg13g2_o21ai_1 _19588_ (.B1(_04141_),
    .Y(_04142_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[22] ),
    .A2(_03864_));
 sg13g2_nor3_1 _19589_ (.A(net5383),
    .B(_04137_),
    .C(_04142_),
    .Y(_04143_));
 sg13g2_a21oi_2 _19590_ (.B1(_04143_),
    .Y(_04144_),
    .A2(_04137_),
    .A1(net5131));
 sg13g2_o21ai_1 _19591_ (.B1(_04136_),
    .Y(_04145_),
    .A1(_03837_),
    .A2(_04144_));
 sg13g2_o21ai_1 _19592_ (.B1(_04145_),
    .Y(_04146_),
    .A1(net3767),
    .A2(net4588));
 sg13g2_inv_1 _19593_ (.Y(_01162_),
    .A(_04146_));
 sg13g2_nor2b_1 _19594_ (.A(net5578),
    .B_N(net5773),
    .Y(_04147_));
 sg13g2_nand2_1 _19595_ (.Y(_04148_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[23] ),
    .B(net4631));
 sg13g2_a22oi_1 _19596_ (.Y(_04149_),
    .B1(net4661),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[23] ),
    .A2(net4667),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[23] ));
 sg13g2_a221oi_1 _19597_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[23] ),
    .C1(net4696),
    .B1(net4687),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[23] ),
    .Y(_04150_),
    .A2(net4675));
 sg13g2_nand3_1 _19598_ (.B(_04149_),
    .C(_04150_),
    .A(_04148_),
    .Y(_04151_));
 sg13g2_o21ai_1 _19599_ (.B1(_04151_),
    .Y(_04152_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[23] ),
    .A2(_03864_));
 sg13g2_nor3_1 _19600_ (.A(net5383),
    .B(_04147_),
    .C(_04152_),
    .Y(_04153_));
 sg13g2_a21oi_2 _19601_ (.B1(_04153_),
    .Y(_04154_),
    .A2(_04147_),
    .A1(net5132));
 sg13g2_and2_1 _19602_ (.A(net5056),
    .B(_04154_),
    .X(_04155_));
 sg13g2_nor2_2 _19603_ (.A(\fpga_top.cpu_start_adr[23] ),
    .B(net5056),
    .Y(_04156_));
 sg13g2_nor3_1 _19604_ (.A(net4584),
    .B(_04155_),
    .C(_04156_),
    .Y(_04157_));
 sg13g2_a21o_1 _19605_ (.A2(net4584),
    .A1(net1983),
    .B1(_04157_),
    .X(_01163_));
 sg13g2_a21oi_1 _19606_ (.A1(\fpga_top.cpu_start_adr[24] ),
    .A2(net5141),
    .Y(_04158_),
    .B1(net4586));
 sg13g2_nor2b_1 _19607_ (.A(net5578),
    .B_N(\fpga_top.cpu_top.execution.csr_array.rs1_sel[24] ),
    .Y(_04159_));
 sg13g2_nand2_1 _19608_ (.Y(_04160_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[24] ),
    .B(net4632));
 sg13g2_a22oi_1 _19609_ (.Y(_04161_),
    .B1(net4661),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[24] ),
    .A2(net4669),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[24] ));
 sg13g2_a221oi_1 _19610_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[24] ),
    .C1(net4698),
    .B1(net4689),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[24] ),
    .Y(_04162_),
    .A2(net4676));
 sg13g2_nand3_1 _19611_ (.B(_04161_),
    .C(_04162_),
    .A(_04160_),
    .Y(_04163_));
 sg13g2_o21ai_1 _19612_ (.B1(_04163_),
    .Y(_04164_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[24] ),
    .A2(_03864_));
 sg13g2_nor3_1 _19613_ (.A(net5385),
    .B(_04159_),
    .C(_04164_),
    .Y(_04165_));
 sg13g2_a21oi_2 _19614_ (.B1(_04165_),
    .Y(_04166_),
    .A2(_04159_),
    .A1(net5133));
 sg13g2_o21ai_1 _19615_ (.B1(_04158_),
    .Y(_04167_),
    .A1(_03837_),
    .A2(_04166_));
 sg13g2_o21ai_1 _19616_ (.B1(_04167_),
    .Y(_04168_),
    .A1(net3812),
    .A2(net4589));
 sg13g2_inv_1 _19617_ (.Y(_01164_),
    .A(_04168_));
 sg13g2_a21oi_1 _19618_ (.A1(net6618),
    .A2(net5143),
    .Y(_04169_),
    .B1(net4586));
 sg13g2_nor2b_1 _19619_ (.A(net5578),
    .B_N(net5768),
    .Y(_04170_));
 sg13g2_and2_1 _19620_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[25] ),
    .B(net4663),
    .X(_04171_));
 sg13g2_a221oi_1 _19621_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[25] ),
    .C1(_04171_),
    .B1(net4689),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[25] ),
    .Y(_04172_),
    .A2(net4632));
 sg13g2_a221oi_1 _19622_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[25] ),
    .C1(net4698),
    .B1(net4669),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[25] ),
    .Y(_04173_),
    .A2(net4676));
 sg13g2_a22oi_1 _19623_ (.Y(_04174_),
    .B1(_04172_),
    .B2(_04173_),
    .A2(net4694),
    .A1(_06918_));
 sg13g2_nor2_1 _19624_ (.A(net5383),
    .B(_04170_),
    .Y(_04175_));
 sg13g2_a22oi_1 _19625_ (.Y(_04176_),
    .B1(_04174_),
    .B2(_04175_),
    .A2(_04170_),
    .A1(net5131));
 sg13g2_o21ai_1 _19626_ (.B1(_04169_),
    .Y(_04177_),
    .A1(net5141),
    .A2(_04176_));
 sg13g2_o21ai_1 _19627_ (.B1(_04177_),
    .Y(_04178_),
    .A1(net3845),
    .A2(net4588));
 sg13g2_inv_1 _19628_ (.Y(_01165_),
    .A(_04178_));
 sg13g2_nor2b_1 _19629_ (.A(net5579),
    .B_N(\fpga_top.cpu_top.execution.csr_array.rs1_sel[26] ),
    .Y(_04179_));
 sg13g2_nand2_1 _19630_ (.Y(_04180_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[26] ),
    .B(net4630));
 sg13g2_a22oi_1 _19631_ (.Y(_04181_),
    .B1(net4661),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[26] ),
    .A2(net4667),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[26] ));
 sg13g2_a221oi_1 _19632_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[26] ),
    .C1(net4697),
    .B1(net4688),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[26] ),
    .Y(_04182_),
    .A2(net4674));
 sg13g2_nand3_1 _19633_ (.B(_04181_),
    .C(_04182_),
    .A(_04180_),
    .Y(_04183_));
 sg13g2_o21ai_1 _19634_ (.B1(_04183_),
    .Y(_04184_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[26] ),
    .A2(_03864_));
 sg13g2_nor3_1 _19635_ (.A(net5384),
    .B(_04179_),
    .C(_04184_),
    .Y(_04185_));
 sg13g2_a21oi_2 _19636_ (.B1(_04185_),
    .Y(_04186_),
    .A2(_04179_),
    .A1(net5132));
 sg13g2_and2_1 _19637_ (.A(net5056),
    .B(_04186_),
    .X(_04187_));
 sg13g2_nor2_2 _19638_ (.A(\fpga_top.cpu_start_adr[26] ),
    .B(net5056),
    .Y(_04188_));
 sg13g2_nor3_1 _19639_ (.A(net4584),
    .B(_04187_),
    .C(_04188_),
    .Y(_04189_));
 sg13g2_a21o_1 _19640_ (.A2(net4583),
    .A1(net2102),
    .B1(_04189_),
    .X(_01166_));
 sg13g2_nand2_1 _19641_ (.Y(_04190_),
    .A(net5380),
    .B(net5763));
 sg13g2_inv_1 _19642_ (.Y(_04191_),
    .A(_04190_));
 sg13g2_and2_1 _19643_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[27] ),
    .B(net4667),
    .X(_04192_));
 sg13g2_a221oi_1 _19644_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[27] ),
    .C1(_04192_),
    .B1(net4687),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[27] ),
    .Y(_04193_),
    .A2(net4630));
 sg13g2_a221oi_1 _19645_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[27] ),
    .C1(net4696),
    .B1(net4662),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[27] ),
    .Y(_04194_),
    .A2(net4674));
 sg13g2_a22oi_1 _19646_ (.Y(_04195_),
    .B1(_04193_),
    .B2(_04194_),
    .A2(net4694),
    .A1(_06919_));
 sg13g2_nor2_1 _19647_ (.A(net5384),
    .B(_04191_),
    .Y(_04196_));
 sg13g2_a22oi_1 _19648_ (.Y(_04197_),
    .B1(_04195_),
    .B2(_04196_),
    .A2(_04191_),
    .A1(net5131));
 sg13g2_and2_1 _19649_ (.A(net5057),
    .B(_04197_),
    .X(_04198_));
 sg13g2_o21ai_1 _19650_ (.B1(net4588),
    .Y(_04199_),
    .A1(net5641),
    .A2(net5057));
 sg13g2_nand2_1 _19651_ (.Y(_04200_),
    .A(net1560),
    .B(net4583));
 sg13g2_o21ai_1 _19652_ (.B1(_04200_),
    .Y(_01167_),
    .A1(_04198_),
    .A2(_04199_));
 sg13g2_nand2_1 _19653_ (.Y(_04201_),
    .A(net1457),
    .B(net4585));
 sg13g2_o21ai_1 _19654_ (.B1(net4588),
    .Y(_04202_),
    .A1(net5638),
    .A2(net5058));
 sg13g2_nor2_1 _19655_ (.A(net5579),
    .B(_06580_),
    .Y(_04203_));
 sg13g2_nand2_1 _19656_ (.Y(_04204_),
    .A(\fpga_top.cpu_top.csr_mepc_ex[28] ),
    .B(net4687));
 sg13g2_a22oi_1 _19657_ (.Y(_04205_),
    .B1(net4667),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[28] ),
    .A2(net4630),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[28] ));
 sg13g2_a221oi_1 _19658_ (.B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[28] ),
    .C1(net4697),
    .B1(net4662),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[28] ),
    .Y(_04206_),
    .A2(net4675));
 sg13g2_nand3_1 _19659_ (.B(_04205_),
    .C(_04206_),
    .A(_04204_),
    .Y(_04207_));
 sg13g2_o21ai_1 _19660_ (.B1(_04207_),
    .Y(_04208_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[28] ),
    .A2(net4695));
 sg13g2_nor3_1 _19661_ (.A(net5384),
    .B(_04203_),
    .C(_04208_),
    .Y(_04209_));
 sg13g2_a21oi_2 _19662_ (.B1(_04209_),
    .Y(_04210_),
    .A2(_04203_),
    .A1(net5131));
 sg13g2_and2_1 _19663_ (.A(net5057),
    .B(_04210_),
    .X(_04211_));
 sg13g2_o21ai_1 _19664_ (.B1(_04201_),
    .Y(_01168_),
    .A1(_04202_),
    .A2(_04211_));
 sg13g2_nor2b_1 _19665_ (.A(net5578),
    .B_N(net5759),
    .Y(_04212_));
 sg13g2_nand2_1 _19666_ (.Y(_04213_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[29] ),
    .B(net4663));
 sg13g2_a22oi_1 _19667_ (.Y(_04214_),
    .B1(net4668),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[29] ),
    .A2(net4630),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[29] ));
 sg13g2_a221oi_1 _19668_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[29] ),
    .C1(net4696),
    .B1(net4688),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[29] ),
    .Y(_04215_),
    .A2(net4674));
 sg13g2_nand3_1 _19669_ (.B(_04214_),
    .C(_04215_),
    .A(_04213_),
    .Y(_04216_));
 sg13g2_o21ai_1 _19670_ (.B1(_04216_),
    .Y(_04217_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[29] ),
    .A2(_03864_));
 sg13g2_nor3_1 _19671_ (.A(net5383),
    .B(_04212_),
    .C(_04217_),
    .Y(_04218_));
 sg13g2_a21oi_2 _19672_ (.B1(_04218_),
    .Y(_04219_),
    .A2(_04212_),
    .A1(net5132));
 sg13g2_and2_1 _19673_ (.A(net5056),
    .B(_04219_),
    .X(_04220_));
 sg13g2_nor2_2 _19674_ (.A(net5637),
    .B(net5056),
    .Y(_04221_));
 sg13g2_nor3_1 _19675_ (.A(net4584),
    .B(_04220_),
    .C(_04221_),
    .Y(_04222_));
 sg13g2_a21o_1 _19676_ (.A2(net4583),
    .A1(net1933),
    .B1(_04222_),
    .X(_01169_));
 sg13g2_nor2_1 _19677_ (.A(net5579),
    .B(_06581_),
    .Y(_04223_));
 sg13g2_nand2_1 _19678_ (.Y(_04224_),
    .A(net5131),
    .B(_04223_));
 sg13g2_nand2_1 _19679_ (.Y(_04225_),
    .A(net1482),
    .B(net4668));
 sg13g2_a22oi_1 _19680_ (.Y(_04226_),
    .B1(net4662),
    .B2(net1595),
    .A2(net4631),
    .A1(net1826));
 sg13g2_a21o_1 _19681_ (.A2(net4696),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[30] ),
    .B1(_03933_),
    .X(_04227_));
 sg13g2_a221oi_1 _19682_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[30] ),
    .C1(_04227_),
    .B1(net4687),
    .A1(net1410),
    .Y(_04228_),
    .A2(net4674));
 sg13g2_and3_2 _19683_ (.X(_04229_),
    .A(_04225_),
    .B(_04226_),
    .C(_04228_));
 sg13g2_or3_1 _19684_ (.A(net5383),
    .B(_04223_),
    .C(_04229_),
    .X(_04230_));
 sg13g2_and2_1 _19685_ (.A(_04224_),
    .B(_04230_),
    .X(_04231_));
 sg13g2_nand2_2 _19686_ (.Y(_04232_),
    .A(_04224_),
    .B(_04230_));
 sg13g2_nor2_1 _19687_ (.A(net1826),
    .B(net4588),
    .Y(_04233_));
 sg13g2_a22oi_1 _19688_ (.Y(_04234_),
    .B1(_03836_),
    .B2(_04232_),
    .A2(net5142),
    .A1(net5635));
 sg13g2_a21oi_1 _19689_ (.A1(net4588),
    .A2(_04234_),
    .Y(_01170_),
    .B1(_04233_));
 sg13g2_nor2_1 _19690_ (.A(net5580),
    .B(_06582_),
    .Y(_04235_));
 sg13g2_nor2_1 _19691_ (.A(net5385),
    .B(_04235_),
    .Y(_04236_));
 sg13g2_nand2_1 _19692_ (.Y(_04237_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[31] ),
    .B(net4666));
 sg13g2_a22oi_1 _19693_ (.Y(_04238_),
    .B1(net4661),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[31] ),
    .A2(net4629),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[31] ));
 sg13g2_a21oi_1 _19694_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[31] ),
    .A2(net4673),
    .Y(_04239_),
    .B1(_03846_));
 sg13g2_nand3_1 _19695_ (.B(_04238_),
    .C(_04239_),
    .A(_04237_),
    .Y(_04240_));
 sg13g2_o21ai_1 _19696_ (.B1(_04240_),
    .Y(_04241_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mcause[6] ),
    .A2(_03847_));
 sg13g2_a21oi_1 _19697_ (.A1(\fpga_top.cpu_top.csr_mepc_ex[31] ),
    .A2(_03894_),
    .Y(_04242_),
    .B1(net4694));
 sg13g2_a22oi_1 _19698_ (.Y(_04243_),
    .B1(_04241_),
    .B2(_04242_),
    .A2(_03863_),
    .A1(_06923_));
 sg13g2_a22oi_1 _19699_ (.Y(_04244_),
    .B1(_04236_),
    .B2(_04243_),
    .A2(_04235_),
    .A1(net5129));
 sg13g2_nand2_2 _19700_ (.Y(_04245_),
    .A(net5049),
    .B(_04244_));
 sg13g2_nor2_1 _19701_ (.A(net6588),
    .B(net5049),
    .Y(_04246_));
 sg13g2_nor2_1 _19702_ (.A(net4582),
    .B(_04246_),
    .Y(_04247_));
 sg13g2_a22oi_1 _19703_ (.Y(_04248_),
    .B1(_04245_),
    .B2(_04247_),
    .A2(net4582),
    .A1(net3109));
 sg13g2_inv_1 _19704_ (.Y(_01171_),
    .A(_04248_));
 sg13g2_or2_1 _19705_ (.X(_04249_),
    .B(_03169_),
    .A(_09803_));
 sg13g2_mux2_1 _19706_ (.A0(net4364),
    .A1(net3705),
    .S(net4130),
    .X(_01172_));
 sg13g2_mux2_1 _19707_ (.A0(net4358),
    .A1(net3455),
    .S(net4132),
    .X(_01173_));
 sg13g2_mux2_1 _19708_ (.A0(net4354),
    .A1(net3552),
    .S(net4131),
    .X(_01174_));
 sg13g2_mux2_1 _19709_ (.A0(net4347),
    .A1(net3193),
    .S(net4130),
    .X(_01175_));
 sg13g2_mux2_1 _19710_ (.A0(net4341),
    .A1(net3075),
    .S(net4132),
    .X(_01176_));
 sg13g2_mux2_1 _19711_ (.A0(net4197),
    .A1(net2379),
    .S(net4132),
    .X(_01177_));
 sg13g2_mux2_1 _19712_ (.A0(net4336),
    .A1(net2858),
    .S(net4130),
    .X(_01178_));
 sg13g2_mux2_1 _19713_ (.A0(net4332),
    .A1(net2363),
    .S(net4133),
    .X(_01179_));
 sg13g2_mux2_1 _19714_ (.A0(net4328),
    .A1(net3123),
    .S(net4132),
    .X(_01180_));
 sg13g2_mux2_1 _19715_ (.A0(net4318),
    .A1(net2388),
    .S(net4131),
    .X(_01181_));
 sg13g2_mux2_1 _19716_ (.A0(net4193),
    .A1(net2442),
    .S(net4133),
    .X(_01182_));
 sg13g2_mux2_1 _19717_ (.A0(net4189),
    .A1(net3702),
    .S(net4131),
    .X(_01183_));
 sg13g2_mux2_1 _19718_ (.A0(net4315),
    .A1(net2300),
    .S(net4133),
    .X(_01184_));
 sg13g2_mux2_1 _19719_ (.A0(net4311),
    .A1(net3192),
    .S(net4131),
    .X(_01185_));
 sg13g2_mux2_1 _19720_ (.A0(net4303),
    .A1(net3554),
    .S(net4130),
    .X(_01186_));
 sg13g2_mux2_1 _19721_ (.A0(net4299),
    .A1(net3605),
    .S(net4133),
    .X(_01187_));
 sg13g2_mux2_1 _19722_ (.A0(net4293),
    .A1(net2834),
    .S(net4133),
    .X(_01188_));
 sg13g2_mux2_1 _19723_ (.A0(net4288),
    .A1(net2494),
    .S(net4130),
    .X(_01189_));
 sg13g2_mux2_1 _19724_ (.A0(net4282),
    .A1(net2901),
    .S(net4133),
    .X(_01190_));
 sg13g2_mux2_1 _19725_ (.A0(net4277),
    .A1(net3530),
    .S(net4130),
    .X(_01191_));
 sg13g2_mux2_1 _19726_ (.A0(net4271),
    .A1(net2776),
    .S(net4132),
    .X(_01192_));
 sg13g2_mux2_1 _19727_ (.A0(net4264),
    .A1(net2894),
    .S(net4130),
    .X(_01193_));
 sg13g2_mux2_1 _19728_ (.A0(net4262),
    .A1(net3160),
    .S(net4134),
    .X(_01194_));
 sg13g2_mux2_1 _19729_ (.A0(net4258),
    .A1(net3437),
    .S(net4133),
    .X(_01195_));
 sg13g2_mux2_1 _19730_ (.A0(net4406),
    .A1(net2463),
    .S(net4134),
    .X(_01196_));
 sg13g2_mux2_1 _19731_ (.A0(net4401),
    .A1(net2810),
    .S(net4132),
    .X(_01197_));
 sg13g2_mux2_1 _19732_ (.A0(net4396),
    .A1(net2959),
    .S(net4131),
    .X(_01198_));
 sg13g2_mux2_1 _19733_ (.A0(net4390),
    .A1(net3684),
    .S(net4131),
    .X(_01199_));
 sg13g2_mux2_1 _19734_ (.A0(net4382),
    .A1(net2695),
    .S(net4130),
    .X(_01200_));
 sg13g2_mux2_1 _19735_ (.A0(net4380),
    .A1(net3354),
    .S(net4133),
    .X(_01201_));
 sg13g2_mux2_1 _19736_ (.A0(net4374),
    .A1(net3401),
    .S(net4132),
    .X(_01202_));
 sg13g2_mux2_1 _19737_ (.A0(net4371),
    .A1(net3253),
    .S(net4132),
    .X(_01203_));
 sg13g2_a21oi_2 _19738_ (.B1(_06546_),
    .Y(_04250_),
    .A2(_07015_),
    .A1(_07002_));
 sg13g2_nor2_2 _19739_ (.A(_08874_),
    .B(_09555_),
    .Y(_04251_));
 sg13g2_or2_1 _19740_ (.X(_04252_),
    .B(_09555_),
    .A(_08874_));
 sg13g2_nor2_2 _19741_ (.A(net5126),
    .B(net5044),
    .Y(_04253_));
 sg13g2_a21oi_1 _19742_ (.A1(net5665),
    .A2(net5046),
    .Y(_04254_),
    .B1(net5127));
 sg13g2_a21oi_1 _19743_ (.A1(net5664),
    .A2(net5127),
    .Y(_04255_),
    .B1(_04254_));
 sg13g2_nor3_1 _19744_ (.A(net5665),
    .B(net5127),
    .C(net5046),
    .Y(_04256_));
 sg13g2_nor2_1 _19745_ (.A(_04255_),
    .B(_04256_),
    .Y(_01204_));
 sg13g2_nand2_1 _19746_ (.Y(_04257_),
    .A(net5662),
    .B(net5127));
 sg13g2_a21oi_1 _19747_ (.A1(net5665),
    .A2(net6402),
    .Y(_04258_),
    .B1(net5128));
 sg13g2_nor2_1 _19748_ (.A(_04253_),
    .B(_04258_),
    .Y(_04259_));
 sg13g2_a22oi_1 _19749_ (.Y(_01205_),
    .B1(_04257_),
    .B2(_04259_),
    .A2(_04254_),
    .A1(_06666_));
 sg13g2_nand2_1 _19750_ (.Y(_04260_),
    .A(net5660),
    .B(net5127));
 sg13g2_nand4_1 _19751_ (.B(net6402),
    .C(net6434),
    .A(net5665),
    .Y(_04261_),
    .D(net5046));
 sg13g2_nand2b_1 _19752_ (.Y(_04262_),
    .B(_04261_),
    .A_N(net5127));
 sg13g2_nor2_1 _19753_ (.A(net6434),
    .B(_04259_),
    .Y(_04263_));
 sg13g2_a21oi_1 _19754_ (.A1(_04260_),
    .A2(_04262_),
    .Y(_01206_),
    .B1(_04263_));
 sg13g2_and4_1 _19755_ (.A(net5665),
    .B(\fpga_top.cpu_top.csr_wadr_mon[1] ),
    .C(\fpga_top.cpu_top.csr_wadr_mon[2] ),
    .D(\fpga_top.cpu_top.csr_wadr_mon[3] ),
    .X(_04264_));
 sg13g2_a21oi_1 _19756_ (.A1(net5046),
    .A2(_04264_),
    .Y(_04265_),
    .B1(net5127));
 sg13g2_a21oi_1 _19757_ (.A1(net5658),
    .A2(net5127),
    .Y(_04266_),
    .B1(_04265_));
 sg13g2_nor2_1 _19758_ (.A(net6386),
    .B(_04262_),
    .Y(_04267_));
 sg13g2_nor2_1 _19759_ (.A(_04266_),
    .B(net6387),
    .Y(_01207_));
 sg13g2_and2_1 _19760_ (.A(\fpga_top.cpu_top.csr_wadr_mon[4] ),
    .B(_04264_),
    .X(_04268_));
 sg13g2_a21oi_1 _19761_ (.A1(_04252_),
    .A2(_04268_),
    .Y(_04269_),
    .B1(net5128));
 sg13g2_a21oi_1 _19762_ (.A1(\fpga_top.cpu_start_adr[6] ),
    .A2(net5128),
    .Y(_04270_),
    .B1(_04269_));
 sg13g2_a21oi_1 _19763_ (.A1(_06667_),
    .A2(_04265_),
    .Y(_01208_),
    .B1(_04270_));
 sg13g2_and2_1 _19764_ (.A(\fpga_top.cpu_top.csr_wadr_mon[5] ),
    .B(_04268_),
    .X(_04271_));
 sg13g2_nand2_1 _19765_ (.Y(_04272_),
    .A(net3937),
    .B(_04268_));
 sg13g2_nor2_1 _19766_ (.A(_04251_),
    .B(_04272_),
    .Y(_04273_));
 sg13g2_nor2_1 _19767_ (.A(net5123),
    .B(_04273_),
    .Y(_04274_));
 sg13g2_a21oi_1 _19768_ (.A1(net5656),
    .A2(net5128),
    .Y(_04275_),
    .B1(_04274_));
 sg13g2_a21oi_1 _19769_ (.A1(_06668_),
    .A2(_04269_),
    .Y(_01209_),
    .B1(_04275_));
 sg13g2_nand2_1 _19770_ (.Y(_04276_),
    .A(net5654),
    .B(net5123));
 sg13g2_and3_1 _19771_ (.X(_04277_),
    .A(\fpga_top.cpu_top.csr_wadr_mon[6] ),
    .B(net5045),
    .C(_04271_));
 sg13g2_or2_1 _19772_ (.X(_04278_),
    .B(_04277_),
    .A(net5123));
 sg13g2_nor2_1 _19773_ (.A(net6440),
    .B(_04273_),
    .Y(_04279_));
 sg13g2_o21ai_1 _19774_ (.B1(_04276_),
    .Y(_01210_),
    .A1(_04278_),
    .A2(_04279_));
 sg13g2_nand2_1 _19775_ (.Y(_04280_),
    .A(net6374),
    .B(_04277_));
 sg13g2_o21ai_1 _19776_ (.B1(_04280_),
    .Y(_04281_),
    .A1(net6374),
    .A2(_04278_));
 sg13g2_a21oi_1 _19777_ (.A1(_06792_),
    .A2(net5123),
    .Y(_01211_),
    .B1(_04281_));
 sg13g2_and2_1 _19778_ (.A(\fpga_top.cpu_top.csr_wadr_mon[7] ),
    .B(net6480),
    .X(_04282_));
 sg13g2_nand4_1 _19779_ (.B(\fpga_top.cpu_top.csr_wadr_mon[7] ),
    .C(net6480),
    .A(\fpga_top.cpu_top.csr_wadr_mon[6] ),
    .Y(_04283_),
    .D(_04271_));
 sg13g2_a21oi_1 _19780_ (.A1(_04277_),
    .A2(_04282_),
    .Y(_04284_),
    .B1(net5123));
 sg13g2_nor2_1 _19781_ (.A(net6433),
    .B(_04280_),
    .Y(_04285_));
 sg13g2_a221oi_1 _19782_ (.B2(net6433),
    .C1(_04285_),
    .B1(_04284_),
    .A1(net5652),
    .Y(_04286_),
    .A2(net5123));
 sg13g2_inv_1 _19783_ (.Y(_01212_),
    .A(_04286_));
 sg13g2_nand2_1 _19784_ (.Y(_04287_),
    .A(net5651),
    .B(net5124));
 sg13g2_nand2_1 _19785_ (.Y(_04288_),
    .A(\fpga_top.cpu_top.csr_wadr_mon[9] ),
    .B(_04282_));
 sg13g2_nor2_1 _19786_ (.A(net6238),
    .B(net5123),
    .Y(_04289_));
 sg13g2_nor2_1 _19787_ (.A(_04284_),
    .B(_04289_),
    .Y(_04290_));
 sg13g2_a22oi_1 _19788_ (.Y(_01213_),
    .B1(_04287_),
    .B2(_04290_),
    .A2(_04284_),
    .A1(_06669_));
 sg13g2_nor2_1 _19789_ (.A(net4035),
    .B(_04290_),
    .Y(_04291_));
 sg13g2_nor3_2 _19790_ (.A(_06669_),
    .B(_06670_),
    .C(_04283_),
    .Y(_04292_));
 sg13g2_and2_1 _19791_ (.A(net5045),
    .B(_04292_),
    .X(_04293_));
 sg13g2_a221oi_1 _19792_ (.B2(_04292_),
    .C1(net4036),
    .B1(net5045),
    .A1(net5375),
    .Y(_01214_),
    .A2(net5123));
 sg13g2_nor2_1 _19793_ (.A(net6274),
    .B(net5122),
    .Y(_04294_));
 sg13g2_a21oi_1 _19794_ (.A1(net5374),
    .A2(net5122),
    .Y(_04295_),
    .B1(_04294_));
 sg13g2_nor2_1 _19795_ (.A(_04293_),
    .B(_04295_),
    .Y(_04296_));
 sg13g2_nand2_1 _19796_ (.Y(_04297_),
    .A(net6274),
    .B(_04293_));
 sg13g2_nor2b_1 _19797_ (.A(_04296_),
    .B_N(_04297_),
    .Y(_01215_));
 sg13g2_nor2_1 _19798_ (.A(\fpga_top.dma_io_wadr_u[14] ),
    .B(net5122),
    .Y(_04298_));
 sg13g2_and4_1 _19799_ (.A(net6274),
    .B(\fpga_top.dma_io_wadr_u[14] ),
    .C(net5045),
    .D(_04292_),
    .X(_04299_));
 sg13g2_a221oi_1 _19800_ (.B2(_04298_),
    .C1(_04299_),
    .B1(_04297_),
    .A1(_06796_),
    .Y(_01216_),
    .A2(net5122));
 sg13g2_nand3_1 _19801_ (.B(\fpga_top.dma_io_wadr_u[14] ),
    .C(\fpga_top.dma_io_wadr_u[15] ),
    .A(\fpga_top.cpu_top.csr_wadr_mon[6] ),
    .Y(_04300_));
 sg13g2_xnor2_1 _19802_ (.Y(_04301_),
    .A(net6365),
    .B(_04299_));
 sg13g2_nand2_1 _19803_ (.Y(_04302_),
    .A(\fpga_top.cpu_start_adr[15] ),
    .B(net5125));
 sg13g2_o21ai_1 _19804_ (.B1(_04302_),
    .Y(_01217_),
    .A1(net5122),
    .A2(net6366));
 sg13g2_nor4_1 _19805_ (.A(_08881_),
    .B(_04272_),
    .C(_04288_),
    .D(_04300_),
    .Y(_04303_));
 sg13g2_nand4_1 _19806_ (.B(\fpga_top.dma_io_wadr_u[14] ),
    .C(\fpga_top.dma_io_wadr_u[15] ),
    .A(\fpga_top.cpu_top.csr_wadr_mon[11] ),
    .Y(_04304_),
    .D(_04292_));
 sg13g2_o21ai_1 _19807_ (.B1(net5044),
    .Y(_04305_),
    .A1(net6151),
    .A2(_04303_));
 sg13g2_nor2_1 _19808_ (.A(_06829_),
    .B(_04304_),
    .Y(_04306_));
 sg13g2_a22oi_1 _19809_ (.Y(_04307_),
    .B1(net4906),
    .B2(net6151),
    .A2(net5126),
    .A1(net5649));
 sg13g2_o21ai_1 _19810_ (.B1(_04307_),
    .Y(_01218_),
    .A1(_04305_),
    .A2(_04306_));
 sg13g2_o21ai_1 _19811_ (.B1(net5046),
    .Y(_04308_),
    .A1(net6169),
    .A2(_04306_));
 sg13g2_and2_1 _19812_ (.A(net6169),
    .B(_04306_),
    .X(_04309_));
 sg13g2_a22oi_1 _19813_ (.Y(_04310_),
    .B1(net4906),
    .B2(net6169),
    .A2(net5126),
    .A1(net5648));
 sg13g2_o21ai_1 _19814_ (.B1(_04310_),
    .Y(_01219_),
    .A1(_04308_),
    .A2(_04309_));
 sg13g2_o21ai_1 _19815_ (.B1(net5046),
    .Y(_04311_),
    .A1(net6094),
    .A2(_04309_));
 sg13g2_and4_1 _19816_ (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[16] ),
    .B(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[17] ),
    .C(net6094),
    .D(_04303_),
    .X(_04312_));
 sg13g2_a22oi_1 _19817_ (.Y(_04313_),
    .B1(net4906),
    .B2(net6094),
    .A2(net5126),
    .A1(net5647));
 sg13g2_o21ai_1 _19818_ (.B1(net6095),
    .Y(_01220_),
    .A1(_04311_),
    .A2(_04312_));
 sg13g2_o21ai_1 _19819_ (.B1(net5044),
    .Y(_04314_),
    .A1(net6140),
    .A2(_04312_));
 sg13g2_and3_1 _19820_ (.X(_04315_),
    .A(net6094),
    .B(net6140),
    .C(_04309_));
 sg13g2_a22oi_1 _19821_ (.Y(_04316_),
    .B1(_04253_),
    .B2(net6140),
    .A2(net5125),
    .A1(\fpga_top.cpu_start_adr[19] ));
 sg13g2_o21ai_1 _19822_ (.B1(net6141),
    .Y(_01221_),
    .A1(_04314_),
    .A2(_04315_));
 sg13g2_o21ai_1 _19823_ (.B1(net5044),
    .Y(_04317_),
    .A1(net6186),
    .A2(_04315_));
 sg13g2_and2_1 _19824_ (.A(net6186),
    .B(_04315_),
    .X(_04318_));
 sg13g2_a22oi_1 _19825_ (.Y(_04319_),
    .B1(net4907),
    .B2(net6186),
    .A2(net5125),
    .A1(net5646));
 sg13g2_o21ai_1 _19826_ (.B1(_04319_),
    .Y(_01222_),
    .A1(_04317_),
    .A2(_04318_));
 sg13g2_o21ai_1 _19827_ (.B1(net5044),
    .Y(_04320_),
    .A1(net6115),
    .A2(_04318_));
 sg13g2_and4_1 _19828_ (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[19] ),
    .B(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[20] ),
    .C(net6115),
    .D(_04312_),
    .X(_04321_));
 sg13g2_a22oi_1 _19829_ (.Y(_04322_),
    .B1(net4906),
    .B2(net6115),
    .A2(net5126),
    .A1(net5644));
 sg13g2_o21ai_1 _19830_ (.B1(_04322_),
    .Y(_01223_),
    .A1(_04320_),
    .A2(_04321_));
 sg13g2_o21ai_1 _19831_ (.B1(net5044),
    .Y(_04323_),
    .A1(net6108),
    .A2(_04321_));
 sg13g2_and3_1 _19832_ (.X(_04324_),
    .A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[21] ),
    .B(net6108),
    .C(_04318_));
 sg13g2_a22oi_1 _19833_ (.Y(_04325_),
    .B1(net4906),
    .B2(net6108),
    .A2(net5125),
    .A1(net5643));
 sg13g2_o21ai_1 _19834_ (.B1(net6109),
    .Y(_01224_),
    .A1(_04323_),
    .A2(_04324_));
 sg13g2_o21ai_1 _19835_ (.B1(net5044),
    .Y(_04326_),
    .A1(net6082),
    .A2(_04324_));
 sg13g2_and2_1 _19836_ (.A(net6082),
    .B(_04324_),
    .X(_04327_));
 sg13g2_a22oi_1 _19837_ (.Y(_04328_),
    .B1(net4906),
    .B2(net6082),
    .A2(net5126),
    .A1(net5642));
 sg13g2_o21ai_1 _19838_ (.B1(_04328_),
    .Y(_01225_),
    .A1(_04326_),
    .A2(_04327_));
 sg13g2_nor2_1 _19839_ (.A(net6162),
    .B(_04327_),
    .Y(_04329_));
 sg13g2_and4_1 _19840_ (.A(net6108),
    .B(net6082),
    .C(net6162),
    .D(_04321_),
    .X(_04330_));
 sg13g2_or2_1 _19841_ (.X(_04331_),
    .B(_04330_),
    .A(_04251_));
 sg13g2_a22oi_1 _19842_ (.Y(_04332_),
    .B1(net4907),
    .B2(net6162),
    .A2(net5125),
    .A1(\fpga_top.cpu_start_adr[24] ));
 sg13g2_o21ai_1 _19843_ (.B1(net6163),
    .Y(_01226_),
    .A1(_04329_),
    .A2(_04331_));
 sg13g2_and3_1 _19844_ (.X(_04333_),
    .A(net6162),
    .B(net6213),
    .C(_04327_));
 sg13g2_o21ai_1 _19845_ (.B1(net5044),
    .Y(_04334_),
    .A1(net6213),
    .A2(_04330_));
 sg13g2_a22oi_1 _19846_ (.Y(_04335_),
    .B1(net4906),
    .B2(net6213),
    .A2(net5125),
    .A1(net6587));
 sg13g2_o21ai_1 _19847_ (.B1(_04335_),
    .Y(_01227_),
    .A1(_04333_),
    .A2(_04334_));
 sg13g2_and2_1 _19848_ (.A(net4049),
    .B(_04333_),
    .X(_04336_));
 sg13g2_o21ai_1 _19849_ (.B1(net5045),
    .Y(_04337_),
    .A1(net4049),
    .A2(_04333_));
 sg13g2_a22oi_1 _19850_ (.Y(_04338_),
    .B1(net4907),
    .B2(net4049),
    .A2(net5125),
    .A1(\fpga_top.cpu_start_adr[26] ));
 sg13g2_o21ai_1 _19851_ (.B1(_04338_),
    .Y(_01228_),
    .A1(_04336_),
    .A2(_04337_));
 sg13g2_and4_1 _19852_ (.A(net6213),
    .B(net4049),
    .C(net4007),
    .D(_04330_),
    .X(_04339_));
 sg13g2_and2_1 _19853_ (.A(net4007),
    .B(_04336_),
    .X(_04340_));
 sg13g2_o21ai_1 _19854_ (.B1(net5045),
    .Y(_04341_),
    .A1(net4007),
    .A2(_04336_));
 sg13g2_a22oi_1 _19855_ (.Y(_04342_),
    .B1(net4907),
    .B2(net4007),
    .A2(net5122),
    .A1(net5640));
 sg13g2_o21ai_1 _19856_ (.B1(_04342_),
    .Y(_01229_),
    .A1(_04340_),
    .A2(_04341_));
 sg13g2_a21oi_1 _19857_ (.A1(net6246),
    .A2(_04339_),
    .Y(_04343_),
    .B1(_04251_));
 sg13g2_o21ai_1 _19858_ (.B1(_04343_),
    .Y(_04344_),
    .A1(net6246),
    .A2(_04339_));
 sg13g2_a22oi_1 _19859_ (.Y(_04345_),
    .B1(net4907),
    .B2(net6246),
    .A2(net5122),
    .A1(net5638));
 sg13g2_nand2_1 _19860_ (.Y(_01230_),
    .A(_04344_),
    .B(_04345_));
 sg13g2_a21oi_1 _19861_ (.A1(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[28] ),
    .A2(_04339_),
    .Y(_04346_),
    .B1(net4074));
 sg13g2_nand3_1 _19862_ (.B(net4074),
    .C(_04339_),
    .A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[28] ),
    .Y(_04347_));
 sg13g2_nand2_1 _19863_ (.Y(_04348_),
    .A(net5045),
    .B(_04347_));
 sg13g2_a22oi_1 _19864_ (.Y(_04349_),
    .B1(net4907),
    .B2(net4074),
    .A2(net5124),
    .A1(net5637));
 sg13g2_o21ai_1 _19865_ (.B1(_04349_),
    .Y(_01231_),
    .A1(_04346_),
    .A2(_04348_));
 sg13g2_and2_1 _19866_ (.A(_06664_),
    .B(_04347_),
    .X(_04350_));
 sg13g2_o21ai_1 _19867_ (.B1(net5045),
    .Y(_04351_),
    .A1(_06664_),
    .A2(_04347_));
 sg13g2_nand4_1 _19868_ (.B(net6246),
    .C(net4074),
    .A(net3981),
    .Y(_04352_),
    .D(_04340_));
 sg13g2_a22oi_1 _19869_ (.Y(_04353_),
    .B1(net4907),
    .B2(net3981),
    .A2(net5122),
    .A1(net5635));
 sg13g2_o21ai_1 _19870_ (.B1(_04353_),
    .Y(_01232_),
    .A1(_04350_),
    .A2(_04351_));
 sg13g2_xor2_1 _19871_ (.B(_04352_),
    .A(net6424),
    .X(_04354_));
 sg13g2_a22oi_1 _19872_ (.Y(_04355_),
    .B1(net4906),
    .B2(net6424),
    .A2(net5125),
    .A1(net2221));
 sg13g2_o21ai_1 _19873_ (.B1(_04355_),
    .Y(_01233_),
    .A1(_04251_),
    .A2(_04354_));
 sg13g2_nand2_1 _19874_ (.Y(_04356_),
    .A(_08704_),
    .B(_09627_));
 sg13g2_nand2_2 _19875_ (.Y(_04357_),
    .A(net5633),
    .B(_04356_));
 sg13g2_a22oi_1 _19876_ (.Y(_04358_),
    .B1(_04357_),
    .B2(net6091),
    .A2(_07009_),
    .A1(net5633));
 sg13g2_inv_1 _19877_ (.Y(_01234_),
    .A(net6092));
 sg13g2_o21ai_1 _19878_ (.B1(_06542_),
    .Y(_04359_),
    .A1(net5628),
    .A2(net5627));
 sg13g2_nor3_1 _19879_ (.A(net5626),
    .B(_06957_),
    .C(_04359_),
    .Y(_04360_));
 sg13g2_o21ai_1 _19880_ (.B1(net3885),
    .Y(_04361_),
    .A1(_09630_),
    .A2(_09631_));
 sg13g2_nand2b_2 _19881_ (.Y(_04362_),
    .B(_04361_),
    .A_N(_04360_));
 sg13g2_mux2_1 _19882_ (.A0(net6581),
    .A1(_04362_),
    .S(net4711),
    .X(_01235_));
 sg13g2_a21oi_2 _19883_ (.B1(_09634_),
    .Y(_04363_),
    .A2(_09630_),
    .A1(\fpga_top.uart_top.uart_rec_char.pdata[1] ));
 sg13g2_nor2_1 _19884_ (.A(net6486),
    .B(net4712),
    .Y(_04364_));
 sg13g2_a21oi_1 _19885_ (.A1(net4712),
    .A2(_04363_),
    .Y(_01236_),
    .B1(_04364_));
 sg13g2_o21ai_1 _19886_ (.B1(net2232),
    .Y(_04365_),
    .A1(_09630_),
    .A2(_09634_));
 sg13g2_nor2b_2 _19887_ (.A(_09633_),
    .B_N(_04365_),
    .Y(_04366_));
 sg13g2_nor2_1 _19888_ (.A(net5664),
    .B(net4713),
    .Y(_04367_));
 sg13g2_a21oi_1 _19889_ (.A1(net4712),
    .A2(_04366_),
    .Y(_01237_),
    .B1(_04367_));
 sg13g2_nor2_1 _19890_ (.A(net5662),
    .B(net4712),
    .Y(_04368_));
 sg13g2_a21oi_1 _19891_ (.A1(_09635_),
    .A2(net4712),
    .Y(_01238_),
    .B1(_04368_));
 sg13g2_mux2_1 _19892_ (.A0(net5660),
    .A1(net3798),
    .S(net4711),
    .X(_01239_));
 sg13g2_mux2_1 _19893_ (.A0(net5658),
    .A1(net1865),
    .S(net4711),
    .X(_01240_));
 sg13g2_nand2_1 _19894_ (.Y(_04369_),
    .A(net1855),
    .B(net4715));
 sg13g2_o21ai_1 _19895_ (.B1(_04369_),
    .Y(_01241_),
    .A1(_06790_),
    .A2(net4715));
 sg13g2_nand2_1 _19896_ (.Y(_04370_),
    .A(net2282),
    .B(net4715));
 sg13g2_o21ai_1 _19897_ (.B1(_04370_),
    .Y(_01242_),
    .A1(_06791_),
    .A2(net4715));
 sg13g2_mux2_1 _19898_ (.A0(net5654),
    .A1(net2085),
    .S(net4711),
    .X(_01243_));
 sg13g2_nand2_1 _19899_ (.Y(_04371_),
    .A(net1931),
    .B(net4711));
 sg13g2_o21ai_1 _19900_ (.B1(_04371_),
    .Y(_01244_),
    .A1(_06792_),
    .A2(net4711));
 sg13g2_nand2_1 _19901_ (.Y(_04372_),
    .A(net1736),
    .B(net4713));
 sg13g2_o21ai_1 _19902_ (.B1(_04372_),
    .Y(_01245_),
    .A1(_06679_),
    .A2(net4713));
 sg13g2_nand2_1 _19903_ (.Y(_04373_),
    .A(net2129),
    .B(net4714));
 sg13g2_o21ai_1 _19904_ (.B1(_04373_),
    .Y(_01246_),
    .A1(_06793_),
    .A2(net4714));
 sg13g2_nand2_1 _19905_ (.Y(_04374_),
    .A(net1548),
    .B(net4711));
 sg13g2_o21ai_1 _19906_ (.B1(_04374_),
    .Y(_01247_),
    .A1(net5375),
    .A2(net4711));
 sg13g2_nand2_1 _19907_ (.Y(_04375_),
    .A(net1659),
    .B(net4713));
 sg13g2_o21ai_1 _19908_ (.B1(_04375_),
    .Y(_01248_),
    .A1(net5374),
    .A2(net4718));
 sg13g2_nand2_1 _19909_ (.Y(_04376_),
    .A(net2014),
    .B(net4714));
 sg13g2_o21ai_1 _19910_ (.B1(_04376_),
    .Y(_01249_),
    .A1(_06796_),
    .A2(net4714));
 sg13g2_nand2_1 _19911_ (.Y(_04377_),
    .A(net1724),
    .B(net4715));
 sg13g2_o21ai_1 _19912_ (.B1(_04377_),
    .Y(_01250_),
    .A1(net5373),
    .A2(net4715));
 sg13g2_nand2_1 _19913_ (.Y(_04378_),
    .A(net2071),
    .B(net4712));
 sg13g2_o21ai_1 _19914_ (.B1(_04378_),
    .Y(_01251_),
    .A1(_06798_),
    .A2(net4712));
 sg13g2_nand2_1 _19915_ (.Y(_04379_),
    .A(net1692),
    .B(net4713));
 sg13g2_o21ai_1 _19916_ (.B1(_04379_),
    .Y(_01252_),
    .A1(_06799_),
    .A2(net4713));
 sg13g2_nand2_1 _19917_ (.Y(_04380_),
    .A(net1779),
    .B(net4717));
 sg13g2_o21ai_1 _19918_ (.B1(_04380_),
    .Y(_01253_),
    .A1(_06800_),
    .A2(net4717));
 sg13g2_nand2_1 _19919_ (.Y(_04381_),
    .A(net1647),
    .B(net4714));
 sg13g2_o21ai_1 _19920_ (.B1(_04381_),
    .Y(_01254_),
    .A1(_06801_),
    .A2(net4715));
 sg13g2_nand2_1 _19921_ (.Y(_04382_),
    .A(net1737),
    .B(net4718));
 sg13g2_o21ai_1 _19922_ (.B1(_04382_),
    .Y(_01255_),
    .A1(_06802_),
    .A2(net4713));
 sg13g2_mux2_1 _19923_ (.A0(net5644),
    .A1(net3206),
    .S(net4717),
    .X(_01256_));
 sg13g2_nand2_1 _19924_ (.Y(_04383_),
    .A(net1812),
    .B(net4716));
 sg13g2_o21ai_1 _19925_ (.B1(_04383_),
    .Y(_01257_),
    .A1(_06803_),
    .A2(net4717));
 sg13g2_nand2_1 _19926_ (.Y(_04384_),
    .A(net3629),
    .B(net4717));
 sg13g2_o21ai_1 _19927_ (.B1(_04384_),
    .Y(_01258_),
    .A1(_06804_),
    .A2(net4717));
 sg13g2_nand2_1 _19928_ (.Y(_04385_),
    .A(net1835),
    .B(net4714));
 sg13g2_o21ai_1 _19929_ (.B1(_04385_),
    .Y(_01259_),
    .A1(_06805_),
    .A2(net4714));
 sg13g2_nand2_1 _19930_ (.Y(_04386_),
    .A(net2117),
    .B(net4716));
 sg13g2_o21ai_1 _19931_ (.B1(_04386_),
    .Y(_01260_),
    .A1(_06806_),
    .A2(net4716));
 sg13g2_nand2_1 _19932_ (.Y(_04387_),
    .A(net1578),
    .B(net4716));
 sg13g2_o21ai_1 _19933_ (.B1(_04387_),
    .Y(_01261_),
    .A1(_06807_),
    .A2(net4716));
 sg13g2_mux2_1 _19934_ (.A0(net5640),
    .A1(net3424),
    .S(net4716),
    .X(_01262_));
 sg13g2_mux2_1 _19935_ (.A0(net5638),
    .A1(net1678),
    .S(net4714),
    .X(_01263_));
 sg13g2_mux2_1 _19936_ (.A0(net5637),
    .A1(net1887),
    .S(net4717),
    .X(_01264_));
 sg13g2_mux2_1 _19937_ (.A0(net5635),
    .A1(net1824),
    .S(net4716),
    .X(_01265_));
 sg13g2_mux2_1 _19938_ (.A0(net2221),
    .A1(net1598),
    .S(net4716),
    .X(_01266_));
 sg13g2_nand2_1 _19939_ (.Y(_04388_),
    .A(net2069),
    .B(net4820));
 sg13g2_o21ai_1 _19940_ (.B1(_04388_),
    .Y(_01267_),
    .A1(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .A2(net4821));
 sg13g2_nand2_1 _19941_ (.Y(_04389_),
    .A(net2137),
    .B(net4818));
 sg13g2_o21ai_1 _19942_ (.B1(_04389_),
    .Y(_01268_),
    .A1(_06684_),
    .A2(net4821));
 sg13g2_nand2_1 _19943_ (.Y(_04390_),
    .A(net1959),
    .B(net4820));
 sg13g2_o21ai_1 _19944_ (.B1(_04390_),
    .Y(_01269_),
    .A1(_06789_),
    .A2(net4820));
 sg13g2_mux2_1 _19945_ (.A0(net5660),
    .A1(net3959),
    .S(net4820),
    .X(_01270_));
 sg13g2_mux2_1 _19946_ (.A0(net5659),
    .A1(net4045),
    .S(net4826),
    .X(_01271_));
 sg13g2_nand2_1 _19947_ (.Y(_04391_),
    .A(net2099),
    .B(net4826));
 sg13g2_o21ai_1 _19948_ (.B1(_04391_),
    .Y(_01272_),
    .A1(_06790_),
    .A2(net4826));
 sg13g2_nand2_1 _19949_ (.Y(_04392_),
    .A(net1970),
    .B(net4820));
 sg13g2_o21ai_1 _19950_ (.B1(_04392_),
    .Y(_01273_),
    .A1(_06791_),
    .A2(net4820));
 sg13g2_nor2_1 _19951_ (.A(net5654),
    .B(net4821),
    .Y(_04393_));
 sg13g2_a21oi_1 _19952_ (.A1(_06591_),
    .A2(net4821),
    .Y(_01274_),
    .B1(_04393_));
 sg13g2_nand2_1 _19953_ (.Y(_04394_),
    .A(net2230),
    .B(net4818));
 sg13g2_o21ai_1 _19954_ (.B1(_04394_),
    .Y(_01275_),
    .A1(_06792_),
    .A2(net4819));
 sg13g2_nor2_1 _19955_ (.A(net5652),
    .B(net4825),
    .Y(_04395_));
 sg13g2_a21oi_1 _19956_ (.A1(_06595_),
    .A2(net4825),
    .Y(_01276_),
    .B1(_04395_));
 sg13g2_nand2_1 _19957_ (.Y(_04396_),
    .A(net3198),
    .B(net4822));
 sg13g2_o21ai_1 _19958_ (.B1(_04396_),
    .Y(_01277_),
    .A1(_06793_),
    .A2(net4818));
 sg13g2_nand2_1 _19959_ (.Y(_04397_),
    .A(net3441),
    .B(net4824));
 sg13g2_o21ai_1 _19960_ (.B1(_04397_),
    .Y(_01278_),
    .A1(net5375),
    .A2(net4824));
 sg13g2_nand2_1 _19961_ (.Y(_04398_),
    .A(net2866),
    .B(net4819));
 sg13g2_o21ai_1 _19962_ (.B1(_04398_),
    .Y(_01279_),
    .A1(net5374),
    .A2(net4819));
 sg13g2_nand2_1 _19963_ (.Y(_04399_),
    .A(net2143),
    .B(net4825));
 sg13g2_o21ai_1 _19964_ (.B1(_04399_),
    .Y(_01280_),
    .A1(_06796_),
    .A2(net4827));
 sg13g2_nand2_1 _19965_ (.Y(_04400_),
    .A(net2139),
    .B(net4824));
 sg13g2_o21ai_1 _19966_ (.B1(_04400_),
    .Y(_01281_),
    .A1(net5373),
    .A2(net4822));
 sg13g2_nor2_1 _19967_ (.A(net5649),
    .B(net4822),
    .Y(_04401_));
 sg13g2_a21oi_1 _19968_ (.A1(_06609_),
    .A2(net4822),
    .Y(_01282_),
    .B1(_04401_));
 sg13g2_nand2_1 _19969_ (.Y(_04402_),
    .A(net2109),
    .B(net4818));
 sg13g2_o21ai_1 _19970_ (.B1(_04402_),
    .Y(_01283_),
    .A1(_06799_),
    .A2(net4818));
 sg13g2_nor2_1 _19971_ (.A(net5647),
    .B(net4822),
    .Y(_04403_));
 sg13g2_a21oi_1 _19972_ (.A1(_06615_),
    .A2(net4822),
    .Y(_01284_),
    .B1(_04403_));
 sg13g2_nand2_1 _19973_ (.Y(_04404_),
    .A(net2087),
    .B(net4823));
 sg13g2_o21ai_1 _19974_ (.B1(_04404_),
    .Y(_01285_),
    .A1(_06801_),
    .A2(net4823));
 sg13g2_nor2_1 _19975_ (.A(net5646),
    .B(net4825),
    .Y(_04405_));
 sg13g2_a21oi_1 _19976_ (.A1(_06621_),
    .A2(net4825),
    .Y(_01286_),
    .B1(_04405_));
 sg13g2_mux2_1 _19977_ (.A0(net5644),
    .A1(net4025),
    .S(net4819),
    .X(_01287_));
 sg13g2_nand2_1 _19978_ (.Y(_04406_),
    .A(net2875),
    .B(net4818));
 sg13g2_o21ai_1 _19979_ (.B1(_04406_),
    .Y(_01288_),
    .A1(_06803_),
    .A2(net4818));
 sg13g2_nor2_1 _19980_ (.A(net5642),
    .B(net4823),
    .Y(_04407_));
 sg13g2_a21oi_1 _19981_ (.A1(_06627_),
    .A2(net4823),
    .Y(_01289_),
    .B1(_04407_));
 sg13g2_nand2_1 _19982_ (.Y(_04408_),
    .A(net2008),
    .B(net4825));
 sg13g2_o21ai_1 _19983_ (.B1(_04408_),
    .Y(_01290_),
    .A1(_06805_),
    .A2(net4825));
 sg13g2_nand2_1 _19984_ (.Y(_04409_),
    .A(net2891),
    .B(net4818));
 sg13g2_o21ai_1 _19985_ (.B1(_04409_),
    .Y(_01291_),
    .A1(_06806_),
    .A2(net4819));
 sg13g2_nand2_1 _19986_ (.Y(_04410_),
    .A(net1860),
    .B(net4826));
 sg13g2_o21ai_1 _19987_ (.B1(_04410_),
    .Y(_01292_),
    .A1(_06807_),
    .A2(net4826));
 sg13g2_nor2_1 _19988_ (.A(net5640),
    .B(net4827),
    .Y(_04411_));
 sg13g2_a21oi_1 _19989_ (.A1(_06637_),
    .A2(net4826),
    .Y(_01293_),
    .B1(_04411_));
 sg13g2_nand2_1 _19990_ (.Y(_04412_),
    .A(net2024),
    .B(net4820));
 sg13g2_o21ai_1 _19991_ (.B1(_04412_),
    .Y(_01294_),
    .A1(_06808_),
    .A2(net4820));
 sg13g2_nand2_1 _19992_ (.Y(_04413_),
    .A(net2432),
    .B(net4822));
 sg13g2_o21ai_1 _19993_ (.B1(_04413_),
    .Y(_01295_),
    .A1(_06809_),
    .A2(net4822));
 sg13g2_nor2_1 _19994_ (.A(net5635),
    .B(net4827),
    .Y(_04414_));
 sg13g2_a21oi_1 _19995_ (.A1(_06644_),
    .A2(net4827),
    .Y(_01296_),
    .B1(_04414_));
 sg13g2_nand2_1 _19996_ (.Y(_04415_),
    .A(net1981),
    .B(net4826));
 sg13g2_o21ai_1 _19997_ (.B1(_04415_),
    .Y(_01297_),
    .A1(_06811_),
    .A2(net4826));
 sg13g2_nor2_1 _19998_ (.A(_07027_),
    .B(\fpga_top.uart_top.uart_rec_char.next_cmd_status[1] ),
    .Y(_04416_));
 sg13g2_or2_1 _19999_ (.X(_04417_),
    .B(\fpga_top.uart_top.uart_rec_char.next_cmd_status[3] ),
    .A(\fpga_top.uart_top.uart_rec_char.next_cmd_status[2] ));
 sg13g2_nand2b_1 _20000_ (.Y(_04418_),
    .B(_08751_),
    .A_N(_04417_));
 sg13g2_nand2b_1 _20001_ (.Y(_04419_),
    .B(_04418_),
    .A_N(\fpga_top.uart_top.uart_rec_char.next_cmd_status[2] ));
 sg13g2_a21oi_1 _20002_ (.A1(\fpga_top.uart_top.uart_rec_char.next_cmd_status[3] ),
    .A2(_08836_),
    .Y(_04420_),
    .B1(_04419_));
 sg13g2_a21oi_1 _20003_ (.A1(\fpga_top.uart_top.uart_rec_char.next_cmd_status[4] ),
    .A2(_04417_),
    .Y(_04421_),
    .B1(_06955_));
 sg13g2_o21ai_1 _20004_ (.B1(_04421_),
    .Y(_04422_),
    .A1(_04416_),
    .A2(_04420_));
 sg13g2_nor2_1 _20005_ (.A(net1396),
    .B(net5228),
    .Y(_04423_));
 sg13g2_nor2_2 _20006_ (.A(net5228),
    .B(_09637_),
    .Y(_04424_));
 sg13g2_inv_1 _20007_ (.Y(_04425_),
    .A(_04424_));
 sg13g2_nor2_1 _20008_ (.A(net1396),
    .B(_04425_),
    .Y(_04426_));
 sg13g2_nand3_1 _20009_ (.B(_04422_),
    .C(_04426_),
    .A(net3513),
    .Y(_04427_));
 sg13g2_o21ai_1 _20010_ (.B1(_04422_),
    .Y(_04428_),
    .A1(net1396),
    .A2(_04425_));
 sg13g2_nand2b_1 _20011_ (.Y(_04429_),
    .B(_04423_),
    .A_N(net3513));
 sg13g2_o21ai_1 _20012_ (.B1(_04427_),
    .Y(_01298_),
    .A1(_04428_),
    .A2(_04429_));
 sg13g2_nand3_1 _20013_ (.B(_04422_),
    .C(_04426_),
    .A(net2790),
    .Y(_04430_));
 sg13g2_or2_1 _20014_ (.X(_04431_),
    .B(\fpga_top.uart_top.uart_rec_char.data_cntr[0] ),
    .A(net2790));
 sg13g2_nand3_1 _20015_ (.B(_04423_),
    .C(_04431_),
    .A(_09639_),
    .Y(_04432_));
 sg13g2_o21ai_1 _20016_ (.B1(_04430_),
    .Y(_01299_),
    .A1(_04428_),
    .A2(_04432_));
 sg13g2_nand3_1 _20017_ (.B(_04422_),
    .C(_04426_),
    .A(net2141),
    .Y(_04433_));
 sg13g2_nand2b_1 _20018_ (.Y(_04434_),
    .B(_09639_),
    .A_N(net2141));
 sg13g2_nand3_1 _20019_ (.B(_04423_),
    .C(_04434_),
    .A(_09640_),
    .Y(_04435_));
 sg13g2_o21ai_1 _20020_ (.B1(_04433_),
    .Y(_01300_),
    .A1(_04428_),
    .A2(_04435_));
 sg13g2_mux2_1 _20021_ (.A0(_04362_),
    .A1(net3798),
    .S(net4745),
    .X(_01302_));
 sg13g2_nand2_1 _20022_ (.Y(_04436_),
    .A(net1865),
    .B(net4745));
 sg13g2_o21ai_1 _20023_ (.B1(_04436_),
    .Y(_01303_),
    .A1(_04363_),
    .A2(net4745));
 sg13g2_nand2_1 _20024_ (.Y(_04437_),
    .A(net1855),
    .B(net4747));
 sg13g2_o21ai_1 _20025_ (.B1(_04437_),
    .Y(_01304_),
    .A1(_04366_),
    .A2(net4747));
 sg13g2_nand2_1 _20026_ (.Y(_04438_),
    .A(net2282),
    .B(net4745));
 sg13g2_o21ai_1 _20027_ (.B1(_04438_),
    .Y(_01305_),
    .A1(_09635_),
    .A2(net4745));
 sg13g2_a22oi_1 _20028_ (.Y(_04439_),
    .B1(net4745),
    .B2(net2085),
    .A2(net4780),
    .A1(\fpga_top.uart_top.uart_rec_char.data_word[0] ));
 sg13g2_inv_1 _20029_ (.Y(_01306_),
    .A(net2086));
 sg13g2_a22oi_1 _20030_ (.Y(_04440_),
    .B1(net4746),
    .B2(net1931),
    .A2(net4780),
    .A1(net1865));
 sg13g2_inv_1 _20031_ (.Y(_01307_),
    .A(_04440_));
 sg13g2_a22oi_1 _20032_ (.Y(_04441_),
    .B1(net4747),
    .B2(net1736),
    .A2(net4780),
    .A1(net1855));
 sg13g2_inv_1 _20033_ (.Y(_01308_),
    .A(_04441_));
 sg13g2_a22oi_1 _20034_ (.Y(_04442_),
    .B1(net4749),
    .B2(net2129),
    .A2(net4782),
    .A1(net2282));
 sg13g2_inv_1 _20035_ (.Y(_01309_),
    .A(_04442_));
 sg13g2_a22oi_1 _20036_ (.Y(_04443_),
    .B1(net4745),
    .B2(net1548),
    .A2(net4780),
    .A1(net2085));
 sg13g2_inv_1 _20037_ (.Y(_01310_),
    .A(_04443_));
 sg13g2_a22oi_1 _20038_ (.Y(_04444_),
    .B1(net4746),
    .B2(net1659),
    .A2(net4780),
    .A1(net1931));
 sg13g2_inv_1 _20039_ (.Y(_01311_),
    .A(_04444_));
 sg13g2_a22oi_1 _20040_ (.Y(_04445_),
    .B1(net4749),
    .B2(net2014),
    .A2(net4780),
    .A1(net1736));
 sg13g2_inv_1 _20041_ (.Y(_01312_),
    .A(_04445_));
 sg13g2_a22oi_1 _20042_ (.Y(_04446_),
    .B1(net4749),
    .B2(net1724),
    .A2(net4782),
    .A1(net2129));
 sg13g2_inv_1 _20043_ (.Y(_01313_),
    .A(_04446_));
 sg13g2_a22oi_1 _20044_ (.Y(_04447_),
    .B1(net4745),
    .B2(net2071),
    .A2(net4780),
    .A1(net1548));
 sg13g2_inv_1 _20045_ (.Y(_01314_),
    .A(_04447_));
 sg13g2_a22oi_1 _20046_ (.Y(_04448_),
    .B1(net4747),
    .B2(net1692),
    .A2(net4783),
    .A1(net1659));
 sg13g2_inv_1 _20047_ (.Y(_01315_),
    .A(_04448_));
 sg13g2_a22oi_1 _20048_ (.Y(_04449_),
    .B1(net4748),
    .B2(net1779),
    .A2(net4781),
    .A1(net2014));
 sg13g2_inv_1 _20049_ (.Y(_01316_),
    .A(_04449_));
 sg13g2_a22oi_1 _20050_ (.Y(_04450_),
    .B1(net4749),
    .B2(net1647),
    .A2(net4782),
    .A1(net1724));
 sg13g2_inv_1 _20051_ (.Y(_01317_),
    .A(_04450_));
 sg13g2_a22oi_1 _20052_ (.Y(_04451_),
    .B1(net4746),
    .B2(net1737),
    .A2(net4780),
    .A1(net2071));
 sg13g2_inv_1 _20053_ (.Y(_01318_),
    .A(_04451_));
 sg13g2_a22oi_1 _20054_ (.Y(_04452_),
    .B1(net4749),
    .B2(net3206),
    .A2(net4782),
    .A1(net1692));
 sg13g2_inv_1 _20055_ (.Y(_01319_),
    .A(_04452_));
 sg13g2_a22oi_1 _20056_ (.Y(_04453_),
    .B1(net4748),
    .B2(net1812),
    .A2(net4781),
    .A1(net1779));
 sg13g2_inv_1 _20057_ (.Y(_01320_),
    .A(_04453_));
 sg13g2_a22oi_1 _20058_ (.Y(_04454_),
    .B1(net4748),
    .B2(net3629),
    .A2(net4781),
    .A1(net1647));
 sg13g2_inv_1 _20059_ (.Y(_01321_),
    .A(_04454_));
 sg13g2_a22oi_1 _20060_ (.Y(_04455_),
    .B1(net4747),
    .B2(net1835),
    .A2(net4783),
    .A1(net1737));
 sg13g2_inv_1 _20061_ (.Y(_01322_),
    .A(_04455_));
 sg13g2_a22oi_1 _20062_ (.Y(_04456_),
    .B1(net4748),
    .B2(net2117),
    .A2(net4781),
    .A1(net3206));
 sg13g2_inv_1 _20063_ (.Y(_01323_),
    .A(_04456_));
 sg13g2_a22oi_1 _20064_ (.Y(_04457_),
    .B1(net4748),
    .B2(net1578),
    .A2(net4781),
    .A1(net1812));
 sg13g2_inv_1 _20065_ (.Y(_01324_),
    .A(_04457_));
 sg13g2_a22oi_1 _20066_ (.Y(_04458_),
    .B1(net4748),
    .B2(net3424),
    .A2(net4781),
    .A1(\fpga_top.uart_top.uart_rec_char.data_word[19] ));
 sg13g2_inv_1 _20067_ (.Y(_01325_),
    .A(net3425));
 sg13g2_a22oi_1 _20068_ (.Y(_04459_),
    .B1(net4749),
    .B2(net1678),
    .A2(net4782),
    .A1(\fpga_top.uart_top.uart_rec_char.data_word[20] ));
 sg13g2_inv_1 _20069_ (.Y(_01326_),
    .A(net1679));
 sg13g2_a22oi_1 _20070_ (.Y(_04460_),
    .B1(net4749),
    .B2(net1887),
    .A2(net4782),
    .A1(\fpga_top.uart_top.uart_rec_char.data_word[21] ));
 sg13g2_inv_1 _20071_ (.Y(_01327_),
    .A(net1888));
 sg13g2_a22oi_1 _20072_ (.Y(_04461_),
    .B1(net4748),
    .B2(net1824),
    .A2(net4781),
    .A1(net1578));
 sg13g2_inv_1 _20073_ (.Y(_01328_),
    .A(_04461_));
 sg13g2_a22oi_1 _20074_ (.Y(_04462_),
    .B1(net4748),
    .B2(net1598),
    .A2(net4781),
    .A1(\fpga_top.uart_top.uart_rec_char.data_word[23] ));
 sg13g2_inv_1 _20075_ (.Y(_01329_),
    .A(net1599));
 sg13g2_nand2_1 _20076_ (.Y(_04463_),
    .A(net5667),
    .B(net2724));
 sg13g2_o21ai_1 _20077_ (.B1(net2725),
    .Y(_01330_),
    .A1(_06542_),
    .A2(net5667));
 sg13g2_mux2_1 _20078_ (.A0(net5628),
    .A1(net3914),
    .S(net5666),
    .X(_01331_));
 sg13g2_nand2_1 _20079_ (.Y(_04464_),
    .A(net5666),
    .B(net2852));
 sg13g2_o21ai_1 _20080_ (.B1(net2853),
    .Y(_01332_),
    .A1(_06543_),
    .A2(net5667));
 sg13g2_mux2_1 _20081_ (.A0(net3918),
    .A1(\fpga_top.io_uart_out.rout[3] ),
    .S(net5666),
    .X(_01333_));
 sg13g2_nand2_1 _20082_ (.Y(_04465_),
    .A(net5666),
    .B(net3623));
 sg13g2_o21ai_1 _20083_ (.B1(net3624),
    .Y(_01334_),
    .A1(_06544_),
    .A2(net5667));
 sg13g2_mux2_1 _20084_ (.A0(net3985),
    .A1(\fpga_top.io_uart_out.rout[5] ),
    .S(net5666),
    .X(_01335_));
 sg13g2_mux2_1 _20085_ (.A0(net4020),
    .A1(\fpga_top.io_uart_out.rout[6] ),
    .S(net5667),
    .X(_01336_));
 sg13g2_mux2_1 _20086_ (.A0(net4033),
    .A1(\fpga_top.io_uart_out.rout[7] ),
    .S(net5666),
    .X(_01337_));
 sg13g2_nand2_1 _20087_ (.Y(_04466_),
    .A(_08714_),
    .B(_08750_));
 sg13g2_nor2_1 _20088_ (.A(net2101),
    .B(net4902),
    .Y(_04467_));
 sg13g2_a21oi_1 _20089_ (.A1(_06684_),
    .A2(net4902),
    .Y(_01338_),
    .B1(_04467_));
 sg13g2_nor2_1 _20090_ (.A(net3027),
    .B(net4903),
    .Y(_04468_));
 sg13g2_a21oi_1 _20091_ (.A1(_06789_),
    .A2(net4903),
    .Y(_01339_),
    .B1(_04468_));
 sg13g2_mux2_1 _20092_ (.A0(net3822),
    .A1(net5660),
    .S(net4903),
    .X(_01340_));
 sg13g2_nand2_1 _20093_ (.Y(_04469_),
    .A(net5658),
    .B(net4902));
 sg13g2_o21ai_1 _20094_ (.B1(_04469_),
    .Y(_01341_),
    .A1(_06506_),
    .A2(net4902));
 sg13g2_nor2_1 _20095_ (.A(net2278),
    .B(net4902),
    .Y(_04470_));
 sg13g2_a21oi_1 _20096_ (.A1(_06790_),
    .A2(net4902),
    .Y(_01342_),
    .B1(_04470_));
 sg13g2_nor2_1 _20097_ (.A(net3537),
    .B(net4902),
    .Y(_04471_));
 sg13g2_a21oi_1 _20098_ (.A1(_06791_),
    .A2(net4902),
    .Y(_01343_),
    .B1(_04471_));
 sg13g2_nand2_1 _20099_ (.Y(_04472_),
    .A(net5654),
    .B(net4904));
 sg13g2_o21ai_1 _20100_ (.B1(_04472_),
    .Y(_01344_),
    .A1(_06510_),
    .A2(net4904));
 sg13g2_nor2_1 _20101_ (.A(net2759),
    .B(net4904),
    .Y(_04473_));
 sg13g2_a21oi_1 _20102_ (.A1(_06792_),
    .A2(net4904),
    .Y(_01345_),
    .B1(_04473_));
 sg13g2_nor2_1 _20103_ (.A(net2197),
    .B(net4897),
    .Y(_04474_));
 sg13g2_a21oi_1 _20104_ (.A1(_06679_),
    .A2(net4897),
    .Y(_01346_),
    .B1(_04474_));
 sg13g2_nor2_1 _20105_ (.A(net2414),
    .B(net4897),
    .Y(_04475_));
 sg13g2_a21oi_1 _20106_ (.A1(_06793_),
    .A2(net4897),
    .Y(_01347_),
    .B1(_04475_));
 sg13g2_nor2_1 _20107_ (.A(net3676),
    .B(net4897),
    .Y(_04476_));
 sg13g2_a21oi_1 _20108_ (.A1(net5375),
    .A2(net4897),
    .Y(_01348_),
    .B1(_04476_));
 sg13g2_nor2_1 _20109_ (.A(net3581),
    .B(net4901),
    .Y(_04477_));
 sg13g2_a21oi_1 _20110_ (.A1(net5374),
    .A2(net4897),
    .Y(_01349_),
    .B1(_04477_));
 sg13g2_nor2_1 _20111_ (.A(net2559),
    .B(net4901),
    .Y(_04478_));
 sg13g2_a21oi_1 _20112_ (.A1(_06796_),
    .A2(net4901),
    .Y(_01350_),
    .B1(_04478_));
 sg13g2_nor2_1 _20113_ (.A(net2170),
    .B(net4901),
    .Y(_04479_));
 sg13g2_a21oi_1 _20114_ (.A1(net5373),
    .A2(net4901),
    .Y(_01351_),
    .B1(_04479_));
 sg13g2_nor2_1 _20115_ (.A(net1802),
    .B(net4900),
    .Y(_04480_));
 sg13g2_a21oi_1 _20116_ (.A1(_06798_),
    .A2(net4900),
    .Y(_01352_),
    .B1(_04480_));
 sg13g2_nor2_1 _20117_ (.A(net2896),
    .B(net4900),
    .Y(_04481_));
 sg13g2_a21oi_1 _20118_ (.A1(_06799_),
    .A2(net4900),
    .Y(_01353_),
    .B1(_04481_));
 sg13g2_nor2_1 _20119_ (.A(net2419),
    .B(net4898),
    .Y(_04482_));
 sg13g2_a21oi_1 _20120_ (.A1(_06800_),
    .A2(net4898),
    .Y(_01354_),
    .B1(_04482_));
 sg13g2_nor2_1 _20121_ (.A(net1948),
    .B(net4900),
    .Y(_04483_));
 sg13g2_a21oi_1 _20122_ (.A1(_06801_),
    .A2(net4898),
    .Y(_01355_),
    .B1(_04483_));
 sg13g2_nor2_1 _20123_ (.A(net3197),
    .B(net4898),
    .Y(_04484_));
 sg13g2_a21oi_1 _20124_ (.A1(_06802_),
    .A2(net4899),
    .Y(_01356_),
    .B1(_04484_));
 sg13g2_nand2_1 _20125_ (.Y(_04485_),
    .A(net5644),
    .B(net4898));
 sg13g2_o21ai_1 _20126_ (.B1(_04485_),
    .Y(_01357_),
    .A1(_06524_),
    .A2(net4898));
 sg13g2_nor2_1 _20127_ (.A(net1873),
    .B(net4898),
    .Y(_04486_));
 sg13g2_a21oi_1 _20128_ (.A1(_06803_),
    .A2(net4898),
    .Y(_01358_),
    .B1(_04486_));
 sg13g2_nor2_1 _20129_ (.A(net3548),
    .B(net4899),
    .Y(_04487_));
 sg13g2_a21oi_1 _20130_ (.A1(_06804_),
    .A2(net4899),
    .Y(_01359_),
    .B1(_04487_));
 sg13g2_nor2_1 _20131_ (.A(net3433),
    .B(net4901),
    .Y(_04488_));
 sg13g2_a21oi_1 _20132_ (.A1(_06805_),
    .A2(net4901),
    .Y(_01360_),
    .B1(_04488_));
 sg13g2_nor2_1 _20133_ (.A(net2268),
    .B(net4899),
    .Y(_04489_));
 sg13g2_a21oi_1 _20134_ (.A1(_06806_),
    .A2(net4899),
    .Y(_01361_),
    .B1(_04489_));
 sg13g2_nor2_1 _20135_ (.A(net2327),
    .B(net4896),
    .Y(_04490_));
 sg13g2_a21oi_1 _20136_ (.A1(_06807_),
    .A2(net4896),
    .Y(_01362_),
    .B1(_04490_));
 sg13g2_nand2_1 _20137_ (.Y(_04491_),
    .A(net5640),
    .B(net4896));
 sg13g2_o21ai_1 _20138_ (.B1(_04491_),
    .Y(_01363_),
    .A1(_06537_),
    .A2(net4896));
 sg13g2_nor2_1 _20139_ (.A(net3567),
    .B(net4896),
    .Y(_04492_));
 sg13g2_a21oi_1 _20140_ (.A1(_06808_),
    .A2(net4896),
    .Y(_01364_),
    .B1(_04492_));
 sg13g2_nor2_1 _20141_ (.A(net3748),
    .B(net4896),
    .Y(_04493_));
 sg13g2_a21oi_1 _20142_ (.A1(_06809_),
    .A2(net4896),
    .Y(_01365_),
    .B1(_04493_));
 sg13g2_nor2_1 _20143_ (.A(net1688),
    .B(net4904),
    .Y(_04494_));
 sg13g2_a21oi_1 _20144_ (.A1(_06810_),
    .A2(net4904),
    .Y(_01366_),
    .B1(_04494_));
 sg13g2_nor2_1 _20145_ (.A(net2500),
    .B(net4904),
    .Y(_04495_));
 sg13g2_a21oi_1 _20146_ (.A1(_06811_),
    .A2(net4904),
    .Y(_01367_),
    .B1(_04495_));
 sg13g2_and3_2 _20147_ (.X(_04496_),
    .A(\fpga_top.bus_gather.u_read_adr[31] ),
    .B(net5613),
    .C(\fpga_top.uart_top.uart_logics.dma_io_data_en ));
 sg13g2_nand3_1 _20148_ (.B(net5613),
    .C(\fpga_top.uart_top.uart_logics.dma_io_data_en ),
    .A(\fpga_top.bus_gather.u_read_adr[31] ),
    .Y(_04497_));
 sg13g2_and2_1 _20149_ (.A(\fpga_top.uart_top.uart_logics.dma_io_data_en ),
    .B(_09396_),
    .X(_04498_));
 sg13g2_nand2_2 _20150_ (.Y(_04499_),
    .A(\fpga_top.uart_top.uart_logics.dma_io_data_en ),
    .B(_09396_));
 sg13g2_nand2_2 _20151_ (.Y(_04500_),
    .A(net5317),
    .B(net5257));
 sg13g2_nor2_1 _20152_ (.A(net5066),
    .B(_04500_),
    .Y(_04501_));
 sg13g2_nor2_2 _20153_ (.A(net5092),
    .B(_04501_),
    .Y(_04502_));
 sg13g2_o21ai_1 _20154_ (.B1(net5174),
    .Y(_04503_),
    .A1(net5066),
    .A2(_04500_));
 sg13g2_o21ai_1 _20155_ (.B1(net5318),
    .Y(_04504_),
    .A1(_10642_),
    .A2(_04499_));
 sg13g2_a21o_2 _20156_ (.A2(net5258),
    .A1(_03861_),
    .B1(_04504_),
    .X(_04505_));
 sg13g2_o21ai_1 _20157_ (.B1(_04505_),
    .Y(_04506_),
    .A1(_09959_),
    .A2(net5316));
 sg13g2_nor3_1 _20158_ (.A(net5092),
    .B(net5066),
    .C(_04500_),
    .Y(_04507_));
 sg13g2_nand2_1 _20159_ (.Y(_04508_),
    .A(net5174),
    .B(_04501_));
 sg13g2_a22oi_1 _20160_ (.Y(_04509_),
    .B1(net4890),
    .B2(net4069),
    .A2(_09809_),
    .A1(net5097));
 sg13g2_o21ai_1 _20161_ (.B1(_04509_),
    .Y(_01368_),
    .A1(net4895),
    .A2(_04506_));
 sg13g2_nand2_1 _20162_ (.Y(_04510_),
    .A(_10024_),
    .B(net5319));
 sg13g2_a21oi_1 _20163_ (.A1(_10660_),
    .A2(net5264),
    .Y(_04511_),
    .B1(net5324));
 sg13g2_o21ai_1 _20164_ (.B1(_04511_),
    .Y(_04512_),
    .A1(_03879_),
    .A2(net5263));
 sg13g2_nand3_1 _20165_ (.B(_04510_),
    .C(_04512_),
    .A(net5174),
    .Y(_04513_));
 sg13g2_a21oi_1 _20166_ (.A1(net5098),
    .A2(_09963_),
    .Y(_04514_),
    .B1(net4891));
 sg13g2_a22oi_1 _20167_ (.Y(_04515_),
    .B1(_04513_),
    .B2(_04514_),
    .A2(net4891),
    .A1(net3638));
 sg13g2_inv_1 _20168_ (.Y(_01369_),
    .A(_04515_));
 sg13g2_a21oi_1 _20169_ (.A1(_10678_),
    .A2(net5264),
    .Y(_04516_),
    .B1(net5324));
 sg13g2_o21ai_1 _20170_ (.B1(_04516_),
    .Y(_04517_),
    .A1(_03895_),
    .A2(net5264));
 sg13g2_a21oi_1 _20171_ (.A1(_10078_),
    .A2(net5319),
    .Y(_04518_),
    .B1(net5093));
 sg13g2_a221oi_1 _20172_ (.B2(_04518_),
    .C1(net4890),
    .B1(_04517_),
    .A1(net5098),
    .Y(_04519_),
    .A2(_10028_));
 sg13g2_a21o_1 _20173_ (.A2(net4891),
    .A1(net2179),
    .B1(_04519_),
    .X(_01370_));
 sg13g2_nand2_1 _20174_ (.Y(_04520_),
    .A(_03943_),
    .B(net5257));
 sg13g2_a21oi_1 _20175_ (.A1(_10696_),
    .A2(net5263),
    .Y(_04521_),
    .B1(_04496_));
 sg13g2_a221oi_1 _20176_ (.B2(_04521_),
    .C1(net5095),
    .B1(_04520_),
    .A1(_10121_),
    .Y(_04522_),
    .A2(net5320));
 sg13g2_a21oi_1 _20177_ (.A1(net5096),
    .A2(_10082_),
    .Y(_04523_),
    .B1(_04522_));
 sg13g2_mux2_1 _20178_ (.A0(net3225),
    .A1(_04523_),
    .S(net4816),
    .X(_01371_));
 sg13g2_a22oi_1 _20179_ (.Y(_04524_),
    .B1(net4661),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[4] ),
    .A2(net4666),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[4] ));
 sg13g2_a21oi_1 _20180_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtval[4] ),
    .A2(net4673),
    .Y(_04525_),
    .B1(net4670));
 sg13g2_a22oi_1 _20181_ (.Y(_04526_),
    .B1(_04524_),
    .B2(_04525_),
    .A2(_03846_),
    .A1(_06886_));
 sg13g2_a221oi_1 _20182_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[4] ),
    .C1(_04526_),
    .B1(_03894_),
    .A1(_03854_),
    .Y(_04527_),
    .A2(_03862_));
 sg13g2_a21oi_2 _20183_ (.B1(_04527_),
    .Y(_04528_),
    .A2(net4693),
    .A1(_06887_));
 sg13g2_a21oi_1 _20184_ (.A1(_10714_),
    .A2(net5264),
    .Y(_04529_),
    .B1(net5324));
 sg13g2_o21ai_1 _20185_ (.B1(_04529_),
    .Y(_04530_),
    .A1(net5264),
    .A2(_04528_));
 sg13g2_nor2_1 _20186_ (.A(_10160_),
    .B(net5316),
    .Y(_04531_));
 sg13g2_nor2_1 _20187_ (.A(net5094),
    .B(_04531_),
    .Y(_04532_));
 sg13g2_nand2_1 _20188_ (.Y(_04533_),
    .A(_10126_),
    .B(net4816));
 sg13g2_a22oi_1 _20189_ (.Y(_04534_),
    .B1(_04533_),
    .B2(net4895),
    .A2(_04532_),
    .A1(_04530_));
 sg13g2_a21o_1 _20190_ (.A2(net4891),
    .A1(net1978),
    .B1(_04534_),
    .X(_01372_));
 sg13g2_nand2_1 _20191_ (.Y(_04535_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[5] ),
    .B(net4672));
 sg13g2_a22oi_1 _20192_ (.Y(_04536_),
    .B1(net4660),
    .B2(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[5] ),
    .A2(net4666),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[5] ));
 sg13g2_nand2_1 _20193_ (.Y(_04537_),
    .A(_04535_),
    .B(_04536_));
 sg13g2_a221oi_1 _20194_ (.B2(\fpga_top.cpu_top.csr_mepc_ex[5] ),
    .C1(_04537_),
    .B1(_03894_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mcause[5] ),
    .Y(_04538_),
    .A2(net4670));
 sg13g2_a21oi_1 _20195_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[5] ),
    .A2(net4692),
    .Y(_04539_),
    .B1(net4659));
 sg13g2_a22oi_1 _20196_ (.Y(_04540_),
    .B1(_04538_),
    .B2(_04539_),
    .A2(net4659),
    .A1(_06890_));
 sg13g2_a21oi_1 _20197_ (.A1(_10732_),
    .A2(net5265),
    .Y(_04541_),
    .B1(net5326));
 sg13g2_o21ai_1 _20198_ (.B1(_04541_),
    .Y(_04542_),
    .A1(net5264),
    .A2(_04540_));
 sg13g2_o21ai_1 _20199_ (.B1(_04542_),
    .Y(_04543_),
    .A1(_10197_),
    .A2(net5317));
 sg13g2_nand2_1 _20200_ (.Y(_04544_),
    .A(net6441),
    .B(net4891));
 sg13g2_o21ai_1 _20201_ (.B1(_04544_),
    .Y(_04545_),
    .A1(net5174),
    .A2(_10165_));
 sg13g2_a21o_1 _20202_ (.A2(_04543_),
    .A1(_04502_),
    .B1(_04545_),
    .X(_01373_));
 sg13g2_nand2_1 _20203_ (.Y(_04546_),
    .A(_03956_),
    .B(net5258));
 sg13g2_a21oi_1 _20204_ (.A1(_10750_),
    .A2(net5262),
    .Y(_04547_),
    .B1(net5324));
 sg13g2_a221oi_1 _20205_ (.B2(_04547_),
    .C1(net4894),
    .B1(_04546_),
    .A1(_10233_),
    .Y(_04548_),
    .A2(net5320));
 sg13g2_a221oi_1 _20206_ (.B2(_06860_),
    .C1(_04548_),
    .B1(net4892),
    .A1(net5095),
    .Y(_01374_),
    .A2(_10202_));
 sg13g2_o21ai_1 _20207_ (.B1(net5317),
    .Y(_04549_),
    .A1(_10768_),
    .A2(net5258));
 sg13g2_a21oi_1 _20208_ (.A1(_03969_),
    .A2(net5258),
    .Y(_04550_),
    .B1(_04549_));
 sg13g2_o21ai_1 _20209_ (.B1(_04502_),
    .Y(_04551_),
    .A1(_10267_),
    .A2(net5316));
 sg13g2_a22oi_1 _20210_ (.Y(_04552_),
    .B1(net4890),
    .B2(net3680),
    .A2(_09672_),
    .A1(net5093));
 sg13g2_o21ai_1 _20211_ (.B1(_04552_),
    .Y(_01375_),
    .A1(_04550_),
    .A2(_04551_));
 sg13g2_a21oi_1 _20212_ (.A1(_10784_),
    .A2(net5265),
    .Y(_04553_),
    .B1(net5326));
 sg13g2_o21ai_1 _20213_ (.B1(_04553_),
    .Y(_04554_),
    .A1(_03981_),
    .A2(net5264));
 sg13g2_nor2_1 _20214_ (.A(_10298_),
    .B(net5316),
    .Y(_04555_));
 sg13g2_nor2_1 _20215_ (.A(net5092),
    .B(_04555_),
    .Y(_04556_));
 sg13g2_a221oi_1 _20216_ (.B2(_04556_),
    .C1(net4893),
    .B1(_04554_),
    .A1(net5094),
    .Y(_04557_),
    .A2(_10272_));
 sg13g2_a21o_1 _20217_ (.A2(net4891),
    .A1(net1932),
    .B1(_04557_),
    .X(_01376_));
 sg13g2_nand2_1 _20218_ (.Y(_04558_),
    .A(_03995_),
    .B(net5258));
 sg13g2_a21oi_1 _20219_ (.A1(_10802_),
    .A2(net5263),
    .Y(_04559_),
    .B1(net5322));
 sg13g2_a221oi_1 _20220_ (.B2(_04559_),
    .C1(net4895),
    .B1(_04558_),
    .A1(_10321_),
    .Y(_04560_),
    .A2(net5323));
 sg13g2_a221oi_1 _20221_ (.B2(_06858_),
    .C1(_04560_),
    .B1(net4892),
    .A1(net5098),
    .Y(_01377_),
    .A2(_10301_));
 sg13g2_nand2_1 _20222_ (.Y(_04561_),
    .A(_04005_),
    .B(net5257));
 sg13g2_a21oi_1 _20223_ (.A1(_10820_),
    .A2(net5263),
    .Y(_04562_),
    .B1(net5324));
 sg13g2_a221oi_1 _20224_ (.B2(_04562_),
    .C1(net5095),
    .B1(_04561_),
    .A1(_10336_),
    .Y(_04563_),
    .A2(net5321));
 sg13g2_a21oi_1 _20225_ (.A1(net5096),
    .A2(_10324_),
    .Y(_04564_),
    .B1(_04563_));
 sg13g2_mux2_1 _20226_ (.A0(net2825),
    .A1(_04564_),
    .S(net4816),
    .X(_01378_));
 sg13g2_nand2_1 _20227_ (.Y(_04565_),
    .A(_04019_),
    .B(net5257));
 sg13g2_a21oi_1 _20228_ (.A1(_10838_),
    .A2(net5262),
    .Y(_04566_),
    .B1(net5324));
 sg13g2_a221oi_1 _20229_ (.B2(_04566_),
    .C1(net5096),
    .B1(_04565_),
    .A1(_10350_),
    .Y(_04567_),
    .A2(net5322));
 sg13g2_a21oi_1 _20230_ (.A1(net5096),
    .A2(_10340_),
    .Y(_04568_),
    .B1(_04567_));
 sg13g2_mux2_1 _20231_ (.A0(net3593),
    .A1(_04568_),
    .S(net4816),
    .X(_01379_));
 sg13g2_nand2_1 _20232_ (.Y(_04569_),
    .A(_04033_),
    .B(net5257));
 sg13g2_a21oi_1 _20233_ (.A1(_10856_),
    .A2(net5263),
    .Y(_04570_),
    .B1(net5324));
 sg13g2_a221oi_1 _20234_ (.B2(_04570_),
    .C1(net5095),
    .B1(_04569_),
    .A1(_10364_),
    .Y(_04571_),
    .A2(net5320));
 sg13g2_a21oi_1 _20235_ (.A1(net5097),
    .A2(_10354_),
    .Y(_04572_),
    .B1(_04571_));
 sg13g2_mux2_1 _20236_ (.A0(net3687),
    .A1(_04572_),
    .S(net4816),
    .X(_01380_));
 sg13g2_nand2_1 _20237_ (.Y(_04573_),
    .A(_04044_),
    .B(net5257));
 sg13g2_a21oi_1 _20238_ (.A1(_10874_),
    .A2(net5262),
    .Y(_04574_),
    .B1(net5322));
 sg13g2_a221oi_1 _20239_ (.B2(_04574_),
    .C1(net4894),
    .B1(_04573_),
    .A1(_10377_),
    .Y(_04575_),
    .A2(net5321));
 sg13g2_a221oi_1 _20240_ (.B2(_06859_),
    .C1(_04575_),
    .B1(net4892),
    .A1(net5097),
    .Y(_01381_),
    .A2(_10367_));
 sg13g2_nor2_1 _20241_ (.A(_10892_),
    .B(net5261),
    .Y(_04576_));
 sg13g2_nor2_1 _20242_ (.A(net5325),
    .B(_04576_),
    .Y(_04577_));
 sg13g2_o21ai_1 _20243_ (.B1(_04577_),
    .Y(_04578_),
    .A1(_04058_),
    .A2(net5267));
 sg13g2_a21oi_1 _20244_ (.A1(_10390_),
    .A2(net5321),
    .Y(_04579_),
    .B1(net4894));
 sg13g2_nor2_1 _20245_ (.A(net5174),
    .B(_10381_),
    .Y(_04580_));
 sg13g2_a221oi_1 _20246_ (.B2(_04579_),
    .C1(_04580_),
    .B1(_04578_),
    .A1(net6279),
    .Y(_04581_),
    .A2(net4892));
 sg13g2_inv_1 _20247_ (.Y(_01382_),
    .A(_04581_));
 sg13g2_nand2_1 _20248_ (.Y(_04582_),
    .A(_04067_),
    .B(net5257));
 sg13g2_a21oi_1 _20249_ (.A1(_10910_),
    .A2(net5262),
    .Y(_04583_),
    .B1(net5320));
 sg13g2_a221oi_1 _20250_ (.B2(_04583_),
    .C1(net4894),
    .B1(_04582_),
    .A1(_10402_),
    .Y(_04584_),
    .A2(net5320));
 sg13g2_a221oi_1 _20251_ (.B2(_06857_),
    .C1(_04584_),
    .B1(net4892),
    .A1(net5095),
    .Y(_01383_),
    .A2(_09675_));
 sg13g2_a21oi_1 _20252_ (.A1(_10928_),
    .A2(net5266),
    .Y(_04585_),
    .B1(net5325));
 sg13g2_o21ai_1 _20253_ (.B1(_04585_),
    .Y(_04586_),
    .A1(_04079_),
    .A2(net5267));
 sg13g2_a21oi_1 _20254_ (.A1(_10418_),
    .A2(net5319),
    .Y(_04587_),
    .B1(net4895));
 sg13g2_nor2_1 _20255_ (.A(net1986),
    .B(net4817),
    .Y(_04588_));
 sg13g2_a221oi_1 _20256_ (.B2(_04587_),
    .C1(_04588_),
    .B1(_04586_),
    .A1(net5093),
    .Y(_01384_),
    .A2(_10405_));
 sg13g2_a21oi_1 _20257_ (.A1(_10944_),
    .A2(net5266),
    .Y(_04589_),
    .B1(net5325));
 sg13g2_o21ai_1 _20258_ (.B1(_04589_),
    .Y(_04590_),
    .A1(_04089_),
    .A2(net5266));
 sg13g2_nor2_1 _20259_ (.A(_10432_),
    .B(net5316),
    .Y(_04591_));
 sg13g2_nor2_1 _20260_ (.A(net5093),
    .B(_04591_),
    .Y(_04592_));
 sg13g2_a22oi_1 _20261_ (.Y(_04593_),
    .B1(_04590_),
    .B2(_04592_),
    .A2(_10421_),
    .A1(net5093));
 sg13g2_mux2_1 _20262_ (.A0(net3336),
    .A1(_04593_),
    .S(net4817),
    .X(_01385_));
 sg13g2_o21ai_1 _20263_ (.B1(net5318),
    .Y(_04594_),
    .A1(_10962_),
    .A2(net5261));
 sg13g2_a21oi_2 _20264_ (.B1(_04594_),
    .Y(_04595_),
    .A2(net5261),
    .A1(_04097_));
 sg13g2_o21ai_1 _20265_ (.B1(_04502_),
    .Y(_04596_),
    .A1(_10447_),
    .A2(net5316));
 sg13g2_a22oi_1 _20266_ (.Y(_04597_),
    .B1(net4890),
    .B2(net3707),
    .A2(_10436_),
    .A1(net5092));
 sg13g2_o21ai_1 _20267_ (.B1(_04597_),
    .Y(_01386_),
    .A1(_04595_),
    .A2(_04596_));
 sg13g2_nand2_2 _20268_ (.Y(_04598_),
    .A(_04107_),
    .B(net5259));
 sg13g2_a21oi_2 _20269_ (.B1(net5325),
    .Y(_04599_),
    .A2(net5266),
    .A1(_10980_));
 sg13g2_a221oi_1 _20270_ (.B2(_04599_),
    .C1(net4894),
    .B1(_04598_),
    .A1(_10460_),
    .Y(_04600_),
    .A2(net5320));
 sg13g2_nor2_1 _20271_ (.A(net3856),
    .B(net4816),
    .Y(_04601_));
 sg13g2_nor2_1 _20272_ (.A(net5174),
    .B(_10450_),
    .Y(_04602_));
 sg13g2_nor3_1 _20273_ (.A(_04600_),
    .B(_04601_),
    .C(_04602_),
    .Y(_01387_));
 sg13g2_nand2_1 _20274_ (.Y(_04603_),
    .A(_04120_),
    .B(net5259));
 sg13g2_a21oi_1 _20275_ (.A1(_10998_),
    .A2(net5266),
    .Y(_04604_),
    .B1(net5325));
 sg13g2_o21ai_1 _20276_ (.B1(net5174),
    .Y(_04605_),
    .A1(_10474_),
    .A2(net5316));
 sg13g2_a21oi_2 _20277_ (.B1(_04605_),
    .Y(_04606_),
    .A2(_04604_),
    .A1(_04603_));
 sg13g2_a21oi_1 _20278_ (.A1(net5098),
    .A2(_10463_),
    .Y(_04607_),
    .B1(_04606_));
 sg13g2_mux2_1 _20279_ (.A0(net2562),
    .A1(_04607_),
    .S(net4817),
    .X(_01388_));
 sg13g2_nand2_1 _20280_ (.Y(_04608_),
    .A(_04130_),
    .B(net5260));
 sg13g2_a21oi_1 _20281_ (.A1(_02553_),
    .A2(net5267),
    .Y(_04609_),
    .B1(net5325));
 sg13g2_o21ai_1 _20282_ (.B1(_04502_),
    .Y(_04610_),
    .A1(_10488_),
    .A2(net5316));
 sg13g2_a21oi_2 _20283_ (.B1(_04610_),
    .Y(_04611_),
    .A2(_04609_),
    .A1(_04608_));
 sg13g2_nor2_1 _20284_ (.A(net2507),
    .B(_04508_),
    .Y(_04612_));
 sg13g2_nor2_1 _20285_ (.A(net5175),
    .B(_10477_),
    .Y(_04613_));
 sg13g2_nor3_1 _20286_ (.A(_04611_),
    .B(_04612_),
    .C(_04613_),
    .Y(_01389_));
 sg13g2_nand2_1 _20287_ (.Y(_04614_),
    .A(_04142_),
    .B(net5259));
 sg13g2_a21oi_1 _20288_ (.A1(_02571_),
    .A2(net5266),
    .Y(_04615_),
    .B1(net5325));
 sg13g2_nand2_2 _20289_ (.Y(_04616_),
    .A(_04614_),
    .B(_04615_));
 sg13g2_a21oi_1 _20290_ (.A1(_10502_),
    .A2(net5319),
    .Y(_04617_),
    .B1(net5092));
 sg13g2_a221oi_1 _20291_ (.B2(_04617_),
    .C1(net4890),
    .B1(_04616_),
    .A1(net5092),
    .Y(_04618_),
    .A2(_10491_));
 sg13g2_a21o_1 _20292_ (.A2(net4890),
    .A1(net1968),
    .B1(_04618_),
    .X(_01390_));
 sg13g2_nand2_2 _20293_ (.Y(_04619_),
    .A(_04152_),
    .B(net5259));
 sg13g2_a21oi_1 _20294_ (.A1(_02589_),
    .A2(net5264),
    .Y(_04620_),
    .B1(net5326));
 sg13g2_a221oi_1 _20295_ (.B2(_04620_),
    .C1(net5092),
    .B1(_04619_),
    .A1(_10515_),
    .Y(_04621_),
    .A2(net5319));
 sg13g2_nor2_1 _20296_ (.A(net5176),
    .B(_10505_),
    .Y(_04622_));
 sg13g2_nor3_1 _20297_ (.A(net4890),
    .B(_04621_),
    .C(_04622_),
    .Y(_04623_));
 sg13g2_a21o_1 _20298_ (.A2(net4890),
    .A1(net2043),
    .B1(_04623_),
    .X(_01391_));
 sg13g2_nand2_1 _20299_ (.Y(_04624_),
    .A(_04164_),
    .B(net5257));
 sg13g2_a21oi_1 _20300_ (.A1(_02607_),
    .A2(net5262),
    .Y(_04625_),
    .B1(net5322));
 sg13g2_a221oi_1 _20301_ (.B2(_04625_),
    .C1(net4894),
    .B1(_04624_),
    .A1(_09708_),
    .Y(_04626_),
    .A2(net5319));
 sg13g2_nor2_1 _20302_ (.A(net2064),
    .B(net4817),
    .Y(_04627_));
 sg13g2_nor2_1 _20303_ (.A(net5176),
    .B(_09678_),
    .Y(_04628_));
 sg13g2_nor3_1 _20304_ (.A(_04626_),
    .B(_04627_),
    .C(_04628_),
    .Y(_01392_));
 sg13g2_a21oi_1 _20305_ (.A1(_02623_),
    .A2(net5266),
    .Y(_04629_),
    .B1(net5326));
 sg13g2_o21ai_1 _20306_ (.B1(_04629_),
    .Y(_04630_),
    .A1(_04174_),
    .A2(net5267));
 sg13g2_a21oi_1 _20307_ (.A1(_09729_),
    .A2(net5319),
    .Y(_04631_),
    .B1(net5093));
 sg13g2_a22oi_1 _20308_ (.Y(_04632_),
    .B1(_04630_),
    .B2(_04631_),
    .A2(_09712_),
    .A1(net5093));
 sg13g2_mux2_1 _20309_ (.A0(net2552),
    .A1(_04632_),
    .S(net4817),
    .X(_01393_));
 sg13g2_nand2_2 _20310_ (.Y(_04633_),
    .A(_04184_),
    .B(net5260));
 sg13g2_a21oi_1 _20311_ (.A1(_02641_),
    .A2(net5262),
    .Y(_04634_),
    .B1(net5322));
 sg13g2_a221oi_1 _20312_ (.B2(_04634_),
    .C1(net4895),
    .B1(_04633_),
    .A1(_09742_),
    .Y(_04635_),
    .A2(net5323));
 sg13g2_nor2_1 _20313_ (.A(net2185),
    .B(net4817),
    .Y(_04636_));
 sg13g2_nor2_1 _20314_ (.A(net5175),
    .B(_09732_),
    .Y(_04637_));
 sg13g2_nor3_1 _20315_ (.A(_04635_),
    .B(_04636_),
    .C(_04637_),
    .Y(_01394_));
 sg13g2_o21ai_1 _20316_ (.B1(net5318),
    .Y(_04638_),
    .A1(_02659_),
    .A2(net5259));
 sg13g2_a21oi_2 _20317_ (.B1(_04638_),
    .Y(_04639_),
    .A2(net5259),
    .A1(_04195_));
 sg13g2_a21o_1 _20318_ (.A2(net5321),
    .A1(_09754_),
    .B1(net4894),
    .X(_04640_));
 sg13g2_a22oi_1 _20319_ (.Y(_04641_),
    .B1(net4892),
    .B2(net6097),
    .A2(_09746_),
    .A1(net5095));
 sg13g2_o21ai_1 _20320_ (.B1(_04641_),
    .Y(_01395_),
    .A1(_04639_),
    .A2(_04640_));
 sg13g2_nand2_2 _20321_ (.Y(_04642_),
    .A(_04208_),
    .B(net5259));
 sg13g2_a21oi_1 _20322_ (.A1(_02677_),
    .A2(net5262),
    .Y(_04643_),
    .B1(net5320));
 sg13g2_a221oi_1 _20323_ (.B2(_04643_),
    .C1(net4894),
    .B1(_04642_),
    .A1(_09765_),
    .Y(_04644_),
    .A2(net5320));
 sg13g2_nor2_1 _20324_ (.A(net2135),
    .B(net4816),
    .Y(_04645_));
 sg13g2_nor2_1 _20325_ (.A(net5175),
    .B(_09757_),
    .Y(_04646_));
 sg13g2_nor3_1 _20326_ (.A(_04644_),
    .B(_04645_),
    .C(_04646_),
    .Y(_01396_));
 sg13g2_nand2_2 _20327_ (.Y(_04647_),
    .A(_04217_),
    .B(net5260));
 sg13g2_a21oi_1 _20328_ (.A1(_02695_),
    .A2(net5262),
    .Y(_04648_),
    .B1(net5322));
 sg13g2_a221oi_1 _20329_ (.B2(_04648_),
    .C1(net4895),
    .B1(_04647_),
    .A1(_09776_),
    .Y(_04649_),
    .A2(net5322));
 sg13g2_nor2_1 _20330_ (.A(net3771),
    .B(net4816),
    .Y(_04650_));
 sg13g2_nor2_1 _20331_ (.A(net5175),
    .B(_09769_),
    .Y(_04651_));
 sg13g2_nor3_1 _20332_ (.A(_04649_),
    .B(_04650_),
    .C(_04651_),
    .Y(_01397_));
 sg13g2_nand2_1 _20333_ (.Y(_04652_),
    .A(_04229_),
    .B(net5259));
 sg13g2_a21oi_1 _20334_ (.A1(_02713_),
    .A2(net5266),
    .Y(_04653_),
    .B1(net5325));
 sg13g2_nand2_2 _20335_ (.Y(_04654_),
    .A(_04652_),
    .B(_04653_));
 sg13g2_a21oi_1 _20336_ (.A1(_09787_),
    .A2(net5321),
    .Y(_04655_),
    .B1(net5095));
 sg13g2_a221oi_1 _20337_ (.B2(_04655_),
    .C1(net4892),
    .B1(_04654_),
    .A1(net5095),
    .Y(_04656_),
    .A2(_09779_));
 sg13g2_a21o_1 _20338_ (.A2(net4892),
    .A1(net2082),
    .B1(_04656_),
    .X(_01398_));
 sg13g2_a21oi_1 _20339_ (.A1(_02731_),
    .A2(net5267),
    .Y(_04657_),
    .B1(net5326));
 sg13g2_o21ai_1 _20340_ (.B1(_04657_),
    .Y(_04658_),
    .A1(_04243_),
    .A2(net5267));
 sg13g2_a21oi_1 _20341_ (.A1(_09799_),
    .A2(net5319),
    .Y(_04659_),
    .B1(net5092));
 sg13g2_a22oi_1 _20342_ (.Y(_04660_),
    .B1(_04658_),
    .B2(_04659_),
    .A2(_09790_),
    .A1(net5093));
 sg13g2_mux2_1 _20343_ (.A0(net3480),
    .A1(_04660_),
    .S(net4817),
    .X(_01399_));
 sg13g2_nand3_1 _20344_ (.B(net5227),
    .C(_07004_),
    .A(_06954_),
    .Y(_04661_));
 sg13g2_nand3_1 _20345_ (.B(_08826_),
    .C(_04661_),
    .A(net5624),
    .Y(_04662_));
 sg13g2_nand2_1 _20346_ (.Y(_01400_),
    .A(_08714_),
    .B(net6379));
 sg13g2_a22oi_1 _20347_ (.Y(_04663_),
    .B1(_07021_),
    .B2(_07004_),
    .A2(_07014_),
    .A1(_07012_));
 sg13g2_nor2_1 _20348_ (.A(_06546_),
    .B(_04663_),
    .Y(_04664_));
 sg13g2_nand2b_2 _20349_ (.Y(_04665_),
    .B(net5633),
    .A_N(_04663_));
 sg13g2_nor4_1 _20350_ (.A(_08733_),
    .B(_08736_),
    .C(_09556_),
    .D(net4888),
    .Y(_04666_));
 sg13g2_or4_1 _20351_ (.A(_08733_),
    .B(_08736_),
    .C(_09556_),
    .D(net4889),
    .X(_04667_));
 sg13g2_nand2_1 _20352_ (.Y(_04668_),
    .A(net5616),
    .B(net4815));
 sg13g2_nand2_1 _20353_ (.Y(_04669_),
    .A(net6396),
    .B(net4881));
 sg13g2_o21ai_1 _20354_ (.B1(_04669_),
    .Y(_04670_),
    .A1(net5664),
    .A2(net4881));
 sg13g2_o21ai_1 _20355_ (.B1(_04668_),
    .Y(_01401_),
    .A1(net4815),
    .A2(_04670_));
 sg13g2_xnor2_1 _20356_ (.Y(_04671_),
    .A(\fpga_top.bus_gather.u_read_adr[2] ),
    .B(net5615));
 sg13g2_nand2_1 _20357_ (.Y(_04672_),
    .A(_04665_),
    .B(_04671_));
 sg13g2_o21ai_1 _20358_ (.B1(_04672_),
    .Y(_04673_),
    .A1(net5662),
    .A2(_04665_));
 sg13g2_nor2_1 _20359_ (.A(net3851),
    .B(net4811),
    .Y(_04674_));
 sg13g2_a21oi_1 _20360_ (.A1(net4811),
    .A2(_04673_),
    .Y(_01402_),
    .B1(_04674_));
 sg13g2_a21oi_1 _20361_ (.A1(net5616),
    .A2(net5615),
    .Y(_04675_),
    .B1(net6449));
 sg13g2_nand3_1 _20362_ (.B(net5615),
    .C(\fpga_top.bus_gather.u_read_adr[4] ),
    .A(net5616),
    .Y(_04676_));
 sg13g2_nand2_1 _20363_ (.Y(_04677_),
    .A(net4881),
    .B(_04676_));
 sg13g2_or2_1 _20364_ (.X(_04678_),
    .B(_04677_),
    .A(_04675_));
 sg13g2_a21oi_1 _20365_ (.A1(net5660),
    .A2(net4888),
    .Y(_04679_),
    .B1(net4815));
 sg13g2_a22oi_1 _20366_ (.Y(_01403_),
    .B1(_04678_),
    .B2(_04679_),
    .A2(net4815),
    .A1(_06508_));
 sg13g2_a21oi_1 _20367_ (.A1(net4811),
    .A2(_04677_),
    .Y(_04680_),
    .B1(net6303));
 sg13g2_or2_1 _20368_ (.X(_04681_),
    .B(_04676_),
    .A(_06507_));
 sg13g2_a21o_1 _20369_ (.A2(_04681_),
    .A1(net4881),
    .B1(net4815),
    .X(_04682_));
 sg13g2_a21oi_1 _20370_ (.A1(net5658),
    .A2(net4888),
    .Y(_04683_),
    .B1(_04682_));
 sg13g2_nor2_1 _20371_ (.A(net6304),
    .B(_04683_),
    .Y(_01404_));
 sg13g2_nor2_1 _20372_ (.A(_06514_),
    .B(_04681_),
    .Y(_04684_));
 sg13g2_o21ai_1 _20373_ (.B1(net4811),
    .Y(_04685_),
    .A1(net4888),
    .A2(_04684_));
 sg13g2_a21oi_1 _20374_ (.A1(\fpga_top.cpu_start_adr[6] ),
    .A2(net4888),
    .Y(_04686_),
    .B1(_04685_));
 sg13g2_a21oi_1 _20375_ (.A1(_06514_),
    .A2(_04682_),
    .Y(_01405_),
    .B1(_04686_));
 sg13g2_nor3_1 _20376_ (.A(_06513_),
    .B(_06514_),
    .C(_04681_),
    .Y(_04687_));
 sg13g2_o21ai_1 _20377_ (.B1(net4811),
    .Y(_04688_),
    .A1(net4887),
    .A2(_04687_));
 sg13g2_a21oi_1 _20378_ (.A1(net5656),
    .A2(net4888),
    .Y(_04689_),
    .B1(_04688_));
 sg13g2_a21oi_1 _20379_ (.A1(_06513_),
    .A2(_04685_),
    .Y(_01406_),
    .B1(_04689_));
 sg13g2_nand2_1 _20380_ (.Y(_04690_),
    .A(net5654),
    .B(net4887));
 sg13g2_nand2_1 _20381_ (.Y(_04691_),
    .A(net6364),
    .B(_04687_));
 sg13g2_a21oi_1 _20382_ (.A1(net4880),
    .A2(_04691_),
    .Y(_04692_),
    .B1(net4814));
 sg13g2_a22oi_1 _20383_ (.Y(_01407_),
    .B1(_04690_),
    .B2(_04692_),
    .A2(_04688_),
    .A1(_06511_));
 sg13g2_nor2_1 _20384_ (.A(net6119),
    .B(_04692_),
    .Y(_04693_));
 sg13g2_nor2_1 _20385_ (.A(_06509_),
    .B(_04691_),
    .Y(_04694_));
 sg13g2_o21ai_1 _20386_ (.B1(net4810),
    .Y(_04695_),
    .A1(net4887),
    .A2(_04694_));
 sg13g2_a21oi_1 _20387_ (.A1(net5653),
    .A2(net4887),
    .Y(_04696_),
    .B1(_04695_));
 sg13g2_nor2_1 _20388_ (.A(net6120),
    .B(_04696_),
    .Y(_01408_));
 sg13g2_nand2_1 _20389_ (.Y(_04697_),
    .A(net5652),
    .B(net4889));
 sg13g2_a21oi_1 _20390_ (.A1(net6341),
    .A2(_04694_),
    .Y(_04698_),
    .B1(net4887));
 sg13g2_nor2_1 _20391_ (.A(net4814),
    .B(_04698_),
    .Y(_04699_));
 sg13g2_a22oi_1 _20392_ (.Y(_01409_),
    .B1(_04697_),
    .B2(_04699_),
    .A2(_04695_),
    .A1(_06523_));
 sg13g2_nor4_1 _20393_ (.A(_06509_),
    .B(_06522_),
    .C(_06523_),
    .D(_04691_),
    .Y(_04700_));
 sg13g2_o21ai_1 _20394_ (.B1(net4810),
    .Y(_04701_),
    .A1(net4887),
    .A2(_04700_));
 sg13g2_a21oi_1 _20395_ (.A1(net5651),
    .A2(net4887),
    .Y(_04702_),
    .B1(_04701_));
 sg13g2_nor2_1 _20396_ (.A(net6214),
    .B(_04699_),
    .Y(_04703_));
 sg13g2_nor2_1 _20397_ (.A(_04702_),
    .B(net6215),
    .Y(_01410_));
 sg13g2_nor2_1 _20398_ (.A(net5375),
    .B(net4880),
    .Y(_04704_));
 sg13g2_a21oi_1 _20399_ (.A1(net6301),
    .A2(_04700_),
    .Y(_04705_),
    .B1(net4887));
 sg13g2_nor3_1 _20400_ (.A(net4814),
    .B(_04704_),
    .C(_04705_),
    .Y(_04706_));
 sg13g2_a21oi_1 _20401_ (.A1(_06521_),
    .A2(_04701_),
    .Y(_01411_),
    .B1(_04706_));
 sg13g2_nor2b_2 _20402_ (.A(_09565_),
    .B_N(_04700_),
    .Y(_04707_));
 sg13g2_nor2_1 _20403_ (.A(net4882),
    .B(_04707_),
    .Y(_04708_));
 sg13g2_o21ai_1 _20404_ (.B1(net4808),
    .Y(_04709_),
    .A1(net4883),
    .A2(_04707_));
 sg13g2_a21oi_1 _20405_ (.A1(\fpga_top.cpu_start_adr[13] ),
    .A2(net4886),
    .Y(_04710_),
    .B1(_04708_));
 sg13g2_nor3_1 _20406_ (.A(net4814),
    .B(_04705_),
    .C(_04710_),
    .Y(_04711_));
 sg13g2_a21o_1 _20407_ (.A2(_04709_),
    .A1(net6286),
    .B1(_04711_),
    .X(_01412_));
 sg13g2_nand2_1 _20408_ (.Y(_04712_),
    .A(net5650),
    .B(net4883));
 sg13g2_a21oi_1 _20409_ (.A1(_06518_),
    .A2(net4880),
    .Y(_04713_),
    .B1(_04709_));
 sg13g2_a22oi_1 _20410_ (.Y(_01413_),
    .B1(_04712_),
    .B2(_04713_),
    .A2(_04709_),
    .A1(_06518_));
 sg13g2_nor2_1 _20411_ (.A(net6224),
    .B(_04713_),
    .Y(_04714_));
 sg13g2_and3_1 _20412_ (.X(_04715_),
    .A(\fpga_top.bus_gather.u_read_adr[14] ),
    .B(net6224),
    .C(_04707_));
 sg13g2_a21oi_1 _20413_ (.A1(\fpga_top.cpu_start_adr[15] ),
    .A2(net4883),
    .Y(_04716_),
    .B1(net4812));
 sg13g2_o21ai_1 _20414_ (.B1(_04716_),
    .Y(_04717_),
    .A1(net4883),
    .A2(_04715_));
 sg13g2_nor2b_1 _20415_ (.A(net6225),
    .B_N(_04717_),
    .Y(_01414_));
 sg13g2_nand2_1 _20416_ (.Y(_04718_),
    .A(net5649),
    .B(net4884));
 sg13g2_and2_1 _20417_ (.A(\fpga_top.bus_gather.u_read_adr[16] ),
    .B(_04715_),
    .X(_04719_));
 sg13g2_o21ai_1 _20418_ (.B1(net4810),
    .Y(_04720_),
    .A1(net4883),
    .A2(_04719_));
 sg13g2_o21ai_1 _20419_ (.B1(_04720_),
    .Y(_04721_),
    .A1(net6231),
    .A2(_04715_));
 sg13g2_nand4_1 _20420_ (.B(\fpga_top.bus_gather.u_read_adr[14] ),
    .C(\fpga_top.bus_gather.u_read_adr[15] ),
    .A(\fpga_top.bus_gather.u_read_adr[16] ),
    .Y(_04722_),
    .D(_04707_));
 sg13g2_a22oi_1 _20421_ (.Y(_01415_),
    .B1(_04718_),
    .B2(_04721_),
    .A2(net4813),
    .A1(_06517_));
 sg13g2_and2_1 _20422_ (.A(net6255),
    .B(_04719_),
    .X(_04723_));
 sg13g2_o21ai_1 _20423_ (.B1(net4881),
    .Y(_04724_),
    .A1(net6255),
    .A2(_04719_));
 sg13g2_or2_1 _20424_ (.X(_04725_),
    .B(_04724_),
    .A(_04723_));
 sg13g2_a21oi_1 _20425_ (.A1(net5648),
    .A2(net4883),
    .Y(_04726_),
    .B1(net4812));
 sg13g2_a22oi_1 _20426_ (.Y(_01416_),
    .B1(_04725_),
    .B2(_04726_),
    .A2(net4813),
    .A1(_06515_));
 sg13g2_nand2_1 _20427_ (.Y(_04727_),
    .A(net5647),
    .B(net4884));
 sg13g2_and2_1 _20428_ (.A(net6289),
    .B(_04723_),
    .X(_04728_));
 sg13g2_o21ai_1 _20429_ (.B1(net4808),
    .Y(_04729_),
    .A1(net4884),
    .A2(_04728_));
 sg13g2_o21ai_1 _20430_ (.B1(_04729_),
    .Y(_04730_),
    .A1(net6289),
    .A2(_04723_));
 sg13g2_a22oi_1 _20431_ (.Y(_01417_),
    .B1(_04727_),
    .B2(_04730_),
    .A2(net4813),
    .A1(_06529_));
 sg13g2_nor2_1 _20432_ (.A(net6264),
    .B(_04728_),
    .Y(_04731_));
 sg13g2_nor4_1 _20433_ (.A(_06515_),
    .B(_06527_),
    .C(_06529_),
    .D(_04722_),
    .Y(_04732_));
 sg13g2_or3_1 _20434_ (.A(net4884),
    .B(_04731_),
    .C(_04732_),
    .X(_04733_));
 sg13g2_a21oi_1 _20435_ (.A1(\fpga_top.cpu_start_adr[19] ),
    .A2(net4883),
    .Y(_04734_),
    .B1(net4812));
 sg13g2_a22oi_1 _20436_ (.Y(_01418_),
    .B1(_04733_),
    .B2(_04734_),
    .A2(net4813),
    .A1(_06527_));
 sg13g2_nor2_1 _20437_ (.A(net6291),
    .B(net4808),
    .Y(_04735_));
 sg13g2_and3_2 _20438_ (.X(_04736_),
    .A(\fpga_top.bus_gather.u_read_adr[20] ),
    .B(\fpga_top.bus_gather.u_read_adr[19] ),
    .C(_04728_));
 sg13g2_o21ai_1 _20439_ (.B1(net4881),
    .Y(_04737_),
    .A1(net6291),
    .A2(_04732_));
 sg13g2_nor2_1 _20440_ (.A(_04736_),
    .B(_04737_),
    .Y(_04738_));
 sg13g2_a21oi_1 _20441_ (.A1(net5646),
    .A2(net4885),
    .Y(_04739_),
    .B1(_04738_));
 sg13g2_a21oi_1 _20442_ (.A1(net4808),
    .A2(_04739_),
    .Y(_01419_),
    .B1(_04735_));
 sg13g2_o21ai_1 _20443_ (.B1(net4880),
    .Y(_04740_),
    .A1(net5614),
    .A2(_04736_));
 sg13g2_a21o_1 _20444_ (.A2(_04736_),
    .A1(net5614),
    .B1(_04740_),
    .X(_04741_));
 sg13g2_a21oi_1 _20445_ (.A1(net5644),
    .A2(net4883),
    .Y(_04742_),
    .B1(net4813));
 sg13g2_a22oi_1 _20446_ (.Y(_01420_),
    .B1(_04741_),
    .B2(_04742_),
    .A2(net4812),
    .A1(_06525_));
 sg13g2_nor2_1 _20447_ (.A(net6233),
    .B(net4808),
    .Y(_04743_));
 sg13g2_nand3_1 _20448_ (.B(net6233),
    .C(_04736_),
    .A(net5614),
    .Y(_04744_));
 sg13g2_a21oi_1 _20449_ (.A1(net5614),
    .A2(_04736_),
    .Y(_04745_),
    .B1(net6233));
 sg13g2_nor2_1 _20450_ (.A(net4885),
    .B(_04745_),
    .Y(_04746_));
 sg13g2_nand4_1 _20451_ (.B(\fpga_top.bus_gather.u_read_adr[20] ),
    .C(net6494),
    .A(net5614),
    .Y(_04747_),
    .D(_04732_));
 sg13g2_a22oi_1 _20452_ (.Y(_04748_),
    .B1(_04744_),
    .B2(_04746_),
    .A2(net4885),
    .A1(net5643));
 sg13g2_a21oi_1 _20453_ (.A1(net4808),
    .A2(_04748_),
    .Y(_01421_),
    .B1(_04743_));
 sg13g2_nor2_1 _20454_ (.A(net3901),
    .B(net4808),
    .Y(_04749_));
 sg13g2_nor2_2 _20455_ (.A(_06532_),
    .B(_04744_),
    .Y(_04750_));
 sg13g2_a21oi_1 _20456_ (.A1(_06532_),
    .A2(_04747_),
    .Y(_04751_),
    .B1(net4885));
 sg13g2_nor2b_1 _20457_ (.A(_04750_),
    .B_N(_04751_),
    .Y(_04752_));
 sg13g2_a21oi_1 _20458_ (.A1(net5642),
    .A2(net4885),
    .Y(_04753_),
    .B1(_04752_));
 sg13g2_a21oi_1 _20459_ (.A1(net4808),
    .A2(_04753_),
    .Y(_01422_),
    .B1(_04749_));
 sg13g2_o21ai_1 _20460_ (.B1(net4880),
    .Y(_04754_),
    .A1(net6319),
    .A2(_04750_));
 sg13g2_a21o_1 _20461_ (.A2(_04750_),
    .A1(net6319),
    .B1(_04754_),
    .X(_04755_));
 sg13g2_a21oi_1 _20462_ (.A1(\fpga_top.cpu_start_adr[24] ),
    .A2(net4885),
    .Y(_04756_),
    .B1(net4812));
 sg13g2_a22oi_1 _20463_ (.Y(_01423_),
    .B1(_04755_),
    .B2(_04756_),
    .A2(net4812),
    .A1(_06531_));
 sg13g2_a21oi_1 _20464_ (.A1(\fpga_top.bus_gather.u_read_adr[24] ),
    .A2(_04750_),
    .Y(_04757_),
    .B1(net6239));
 sg13g2_nor4_1 _20465_ (.A(_06530_),
    .B(_06531_),
    .C(_06532_),
    .D(_04747_),
    .Y(_04758_));
 sg13g2_or3_1 _20466_ (.A(net4885),
    .B(_04757_),
    .C(_04758_),
    .X(_04759_));
 sg13g2_a21oi_1 _20467_ (.A1(\fpga_top.cpu_start_adr[25] ),
    .A2(net4885),
    .Y(_04760_),
    .B1(net4812));
 sg13g2_a22oi_1 _20468_ (.Y(_01424_),
    .B1(_04759_),
    .B2(_04760_),
    .A2(net4812),
    .A1(_06530_));
 sg13g2_nor2_1 _20469_ (.A(net3954),
    .B(net4809),
    .Y(_04761_));
 sg13g2_and4_1 _20470_ (.A(\fpga_top.bus_gather.u_read_adr[25] ),
    .B(\fpga_top.bus_gather.u_read_adr[24] ),
    .C(\fpga_top.bus_gather.u_read_adr[26] ),
    .D(_04750_),
    .X(_04762_));
 sg13g2_o21ai_1 _20471_ (.B1(net4880),
    .Y(_04763_),
    .A1(net3954),
    .A2(_04758_));
 sg13g2_nor2_1 _20472_ (.A(_04762_),
    .B(_04763_),
    .Y(_04764_));
 sg13g2_a21oi_1 _20473_ (.A1(\fpga_top.cpu_start_adr[26] ),
    .A2(net4882),
    .Y(_04765_),
    .B1(_04764_));
 sg13g2_a21oi_1 _20474_ (.A1(net4809),
    .A2(_04765_),
    .Y(_01425_),
    .B1(_04761_));
 sg13g2_nor2_1 _20475_ (.A(net3945),
    .B(net4809),
    .Y(_04766_));
 sg13g2_and2_1 _20476_ (.A(net3945),
    .B(_04762_),
    .X(_04767_));
 sg13g2_o21ai_1 _20477_ (.B1(net4880),
    .Y(_04768_),
    .A1(net3945),
    .A2(_04762_));
 sg13g2_nor2_1 _20478_ (.A(_04767_),
    .B(_04768_),
    .Y(_04769_));
 sg13g2_a21oi_1 _20479_ (.A1(net5640),
    .A2(net4882),
    .Y(_04770_),
    .B1(_04769_));
 sg13g2_a21oi_1 _20480_ (.A1(net4809),
    .A2(_04770_),
    .Y(_01426_),
    .B1(_04766_));
 sg13g2_nor2_1 _20481_ (.A(net3909),
    .B(net4809),
    .Y(_04771_));
 sg13g2_nor2_1 _20482_ (.A(net3909),
    .B(_04767_),
    .Y(_04772_));
 sg13g2_and4_1 _20483_ (.A(net3909),
    .B(net3945),
    .C(net3954),
    .D(_04758_),
    .X(_04773_));
 sg13g2_nor3_1 _20484_ (.A(net4882),
    .B(_04772_),
    .C(_04773_),
    .Y(_04774_));
 sg13g2_a21oi_1 _20485_ (.A1(net5638),
    .A2(net4882),
    .Y(_04775_),
    .B1(_04774_));
 sg13g2_a21oi_1 _20486_ (.A1(net4809),
    .A2(_04775_),
    .Y(_01427_),
    .B1(_04771_));
 sg13g2_xnor2_1 _20487_ (.Y(_04776_),
    .A(_06534_),
    .B(_04773_));
 sg13g2_nand2_1 _20488_ (.Y(_04777_),
    .A(net4880),
    .B(_04776_));
 sg13g2_a21oi_1 _20489_ (.A1(net5637),
    .A2(net4882),
    .Y(_04778_),
    .B1(net4814));
 sg13g2_a22oi_1 _20490_ (.Y(_01428_),
    .B1(_04777_),
    .B2(_04778_),
    .A2(net4814),
    .A1(_06534_));
 sg13g2_nor2_1 _20491_ (.A(net5613),
    .B(net4809),
    .Y(_04779_));
 sg13g2_nand4_1 _20492_ (.B(net3909),
    .C(net5613),
    .A(net6317),
    .Y(_04780_),
    .D(_04767_));
 sg13g2_a21oi_1 _20493_ (.A1(net6317),
    .A2(_04773_),
    .Y(_04781_),
    .B1(net5613));
 sg13g2_nor2_1 _20494_ (.A(net4882),
    .B(_04781_),
    .Y(_04782_));
 sg13g2_a22oi_1 _20495_ (.Y(_04783_),
    .B1(_04780_),
    .B2(_04782_),
    .A2(net4882),
    .A1(net5635));
 sg13g2_a21oi_1 _20496_ (.A1(net4809),
    .A2(_04783_),
    .Y(_01429_),
    .B1(_04779_));
 sg13g2_xnor2_1 _20497_ (.Y(_04784_),
    .A(net6524),
    .B(_04780_));
 sg13g2_a21oi_1 _20498_ (.A1(_06811_),
    .A2(net4888),
    .Y(_04785_),
    .B1(net4815));
 sg13g2_o21ai_1 _20499_ (.B1(_04785_),
    .Y(_04786_),
    .A1(net4888),
    .A2(_04784_));
 sg13g2_o21ai_1 _20500_ (.B1(_04786_),
    .Y(_01430_),
    .A1(_06540_),
    .A2(net4811));
 sg13g2_nor3_1 _20501_ (.A(_06540_),
    .B(net4815),
    .C(_04780_),
    .Y(_04787_));
 sg13g2_o21ai_1 _20502_ (.B1(net4881),
    .Y(_04788_),
    .A1(net1641),
    .A2(_04787_));
 sg13g2_a21oi_1 _20503_ (.A1(net1641),
    .A2(_04787_),
    .Y(_01431_),
    .B1(_04788_));
 sg13g2_nand2_1 _20504_ (.Y(_04789_),
    .A(net5612),
    .B(net5069));
 sg13g2_nand2_1 _20505_ (.Y(_04790_),
    .A(net5611),
    .B(net5070));
 sg13g2_o21ai_1 _20506_ (.B1(_04789_),
    .Y(_01432_),
    .A1(_09543_),
    .A2(_04790_));
 sg13g2_nand2_1 _20507_ (.Y(_04791_),
    .A(net5611),
    .B(net5069));
 sg13g2_nand2_1 _20508_ (.Y(_04792_),
    .A(net5610),
    .B(net5070));
 sg13g2_o21ai_1 _20509_ (.B1(_04791_),
    .Y(_01433_),
    .A1(_09543_),
    .A2(_04792_));
 sg13g2_nand2_1 _20510_ (.Y(_04793_),
    .A(net5610),
    .B(_09294_));
 sg13g2_nand2_1 _20511_ (.Y(_04794_),
    .A(net5609),
    .B(net5070));
 sg13g2_o21ai_1 _20512_ (.B1(_04793_),
    .Y(_01434_),
    .A1(_09543_),
    .A2(_04794_));
 sg13g2_nand2_1 _20513_ (.Y(_04795_),
    .A(net5609),
    .B(net5069));
 sg13g2_nand2_1 _20514_ (.Y(_04796_),
    .A(net5608),
    .B(net5070));
 sg13g2_o21ai_1 _20515_ (.B1(_04795_),
    .Y(_01435_),
    .A1(_09543_),
    .A2(_04796_));
 sg13g2_nand2_1 _20516_ (.Y(_04797_),
    .A(net5608),
    .B(net5069));
 sg13g2_nand2_1 _20517_ (.Y(_04798_),
    .A(net3659),
    .B(net5070));
 sg13g2_o21ai_1 _20518_ (.B1(_04797_),
    .Y(_01436_),
    .A1(_09543_),
    .A2(_04798_));
 sg13g2_nand2_1 _20519_ (.Y(_04799_),
    .A(net5607),
    .B(net5069));
 sg13g2_nand2_1 _20520_ (.Y(_04800_),
    .A(net3488),
    .B(net5070));
 sg13g2_o21ai_1 _20521_ (.B1(_04799_),
    .Y(_01437_),
    .A1(_09543_),
    .A2(_04800_));
 sg13g2_nand2_1 _20522_ (.Y(_04801_),
    .A(net3488),
    .B(net5069));
 sg13g2_nand2_1 _20523_ (.Y(_04802_),
    .A(net3168),
    .B(net5070));
 sg13g2_o21ai_1 _20524_ (.B1(_04801_),
    .Y(_01438_),
    .A1(_09543_),
    .A2(_04802_));
 sg13g2_nand2_1 _20525_ (.Y(_04803_),
    .A(net3168),
    .B(net5069));
 sg13g2_o21ai_1 _20526_ (.B1(_04803_),
    .Y(_01439_),
    .A1(net5069),
    .A2(_09541_));
 sg13g2_a21oi_1 _20527_ (.A1(_06663_),
    .A2(_09557_),
    .Y(_01440_),
    .B1(_08855_));
 sg13g2_or2_1 _20528_ (.X(_04804_),
    .B(_03656_),
    .A(_06929_));
 sg13g2_mux2_1 _20529_ (.A0(\fpga_top.io_uart_out.rout[0] ),
    .A1(\fpga_top.io_uart_out.uart_io_char[0] ),
    .S(net5711),
    .X(_04805_));
 sg13g2_nand2b_2 _20530_ (.Y(_04806_),
    .B(\fpga_top.uart_top.uart_send_char.send_cntr[2] ),
    .A_N(net5422));
 sg13g2_nor3_2 _20531_ (.A(net5424),
    .B(net5423),
    .C(_04806_),
    .Y(_04807_));
 sg13g2_and2_1 _20532_ (.A(net5422),
    .B(_08744_),
    .X(_04808_));
 sg13g2_and3_2 _20533_ (.X(_04809_),
    .A(net5424),
    .B(net5422),
    .C(_08739_));
 sg13g2_nand3_1 _20534_ (.B(net5422),
    .C(_08739_),
    .A(net5424),
    .Y(_04810_));
 sg13g2_nor3_2 _20535_ (.A(_06501_),
    .B(net5423),
    .C(_04806_),
    .Y(_04811_));
 sg13g2_nand2_1 _20536_ (.Y(_04812_),
    .A(net5425),
    .B(\fpga_top.uart_top.uart_send_char.send_cntr[1] ));
 sg13g2_nor2_2 _20537_ (.A(_04806_),
    .B(_04812_),
    .Y(_04813_));
 sg13g2_nor3_2 _20538_ (.A(net5422),
    .B(\fpga_top.uart_top.uart_send_char.send_cntr[2] ),
    .C(_04812_),
    .Y(_04814_));
 sg13g2_nand2_1 _20539_ (.Y(_04815_),
    .A(_06501_),
    .B(\fpga_top.uart_top.uart_send_char.send_cntr[1] ));
 sg13g2_nor2_2 _20540_ (.A(_04806_),
    .B(_04815_),
    .Y(_04816_));
 sg13g2_a221oi_1 _20541_ (.B2(\fpga_top.bus_gather.i_read_adr[20] ),
    .C1(net5229),
    .B1(_04813_),
    .A1(net5590),
    .Y(_04817_),
    .A2(_04809_));
 sg13g2_a22oi_1 _20542_ (.Y(_04818_),
    .B1(_04816_),
    .B2(net5593),
    .A2(_04807_),
    .A1(net5595));
 sg13g2_a22oi_1 _20543_ (.Y(_04819_),
    .B1(_04814_),
    .B2(net5597),
    .A2(_04808_),
    .A1(\fpga_top.bus_gather.i_read_adr[24] ));
 sg13g2_nand3_1 _20544_ (.B(_04818_),
    .C(_04819_),
    .A(_04817_),
    .Y(_04820_));
 sg13g2_a21oi_1 _20545_ (.A1(\fpga_top.bus_gather.i_read_adr[12] ),
    .A2(_04811_),
    .Y(_04821_),
    .B1(_04820_));
 sg13g2_nand2_1 _20546_ (.Y(_04822_),
    .A(\fpga_top.uart_top.uart_logics.data_0[8] ),
    .B(_04807_));
 sg13g2_nor3_2 _20547_ (.A(\fpga_top.uart_top.uart_send_char.send_cntr[3] ),
    .B(\fpga_top.uart_top.uart_send_char.send_cntr[2] ),
    .C(_04815_),
    .Y(_04823_));
 sg13g2_nand2_1 _20548_ (.Y(_04824_),
    .A(\fpga_top.uart_top.uart_logics.data_0[0] ),
    .B(_04823_));
 sg13g2_a221oi_1 _20549_ (.B2(\fpga_top.uart_top.uart_logics.data_0[12] ),
    .C1(net5234),
    .B1(_04811_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[28] ),
    .Y(_04825_),
    .A2(_04809_));
 sg13g2_a22oi_1 _20550_ (.Y(_04826_),
    .B1(_04816_),
    .B2(\fpga_top.uart_top.uart_logics.data_0[16] ),
    .A2(_04814_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[4] ));
 sg13g2_a22oi_1 _20551_ (.Y(_04827_),
    .B1(_04813_),
    .B2(\fpga_top.uart_top.uart_logics.data_0[20] ),
    .A2(_04808_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[24] ));
 sg13g2_and4_1 _20552_ (.A(_04822_),
    .B(_04824_),
    .C(_04826_),
    .D(_04827_),
    .X(_04828_));
 sg13g2_a21oi_2 _20553_ (.B1(_04821_),
    .Y(_04829_),
    .A2(_04828_),
    .A1(_04825_));
 sg13g2_a21o_1 _20554_ (.A2(_08740_),
    .A1(net5425),
    .B1(_04829_),
    .X(_04830_));
 sg13g2_o21ai_1 _20555_ (.B1(_04807_),
    .Y(_04831_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[11] ),
    .A2(net5231));
 sg13g2_a21oi_1 _20556_ (.A1(_06597_),
    .A2(net5230),
    .Y(_04832_),
    .B1(_04831_));
 sg13g2_o21ai_1 _20557_ (.B1(_04814_),
    .Y(_04833_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[7] ),
    .A2(net5232));
 sg13g2_a21oi_1 _20558_ (.A1(_06590_),
    .A2(net5232),
    .Y(_04834_),
    .B1(_04833_));
 sg13g2_o21ai_1 _20559_ (.B1(_04816_),
    .Y(_04835_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[19] ),
    .A2(net5231));
 sg13g2_a21oi_1 _20560_ (.A1(_06617_),
    .A2(net5231),
    .Y(_04836_),
    .B1(_04835_));
 sg13g2_o21ai_1 _20561_ (.B1(_04823_),
    .Y(_04837_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[3] ),
    .A2(net5233));
 sg13g2_a21oi_1 _20562_ (.A1(_06584_),
    .A2(net5232),
    .Y(_04838_),
    .B1(_04837_));
 sg13g2_o21ai_1 _20563_ (.B1(_04808_),
    .Y(_04839_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[27] ),
    .A2(net5231));
 sg13g2_a21oi_1 _20564_ (.A1(_06636_),
    .A2(net5230),
    .Y(_04840_),
    .B1(_04839_));
 sg13g2_o21ai_1 _20565_ (.B1(_04809_),
    .Y(_04841_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[31] ),
    .A2(net5232));
 sg13g2_a21oi_1 _20566_ (.A1(_06646_),
    .A2(net5232),
    .Y(_04842_),
    .B1(_04841_));
 sg13g2_o21ai_1 _20567_ (.B1(_04811_),
    .Y(_04843_),
    .A1(\fpga_top.bus_gather.i_read_adr[15] ),
    .A2(net5229));
 sg13g2_a21oi_1 _20568_ (.A1(_06857_),
    .A2(net5229),
    .Y(_04844_),
    .B1(_04843_));
 sg13g2_o21ai_1 _20569_ (.B1(_04813_),
    .Y(_04845_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[23] ),
    .A2(net5234));
 sg13g2_a21oi_1 _20570_ (.A1(_06626_),
    .A2(net5232),
    .Y(_04846_),
    .B1(_04845_));
 sg13g2_nor4_1 _20571_ (.A(_04832_),
    .B(_04836_),
    .C(_04840_),
    .D(_04844_),
    .Y(_04847_));
 sg13g2_nor4_1 _20572_ (.A(_04834_),
    .B(_04838_),
    .C(_04842_),
    .D(_04846_),
    .Y(_04848_));
 sg13g2_and2_1 _20573_ (.A(_04847_),
    .B(_04848_),
    .X(_04849_));
 sg13g2_nand2_1 _20574_ (.Y(_04850_),
    .A(\fpga_top.uart_top.uart_logics.data_0[13] ),
    .B(_04811_));
 sg13g2_a22oi_1 _20575_ (.Y(_04851_),
    .B1(_04823_),
    .B2(\fpga_top.uart_top.uart_logics.data_0[1] ),
    .A2(_04814_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[5] ));
 sg13g2_a21oi_1 _20576_ (.A1(\fpga_top.uart_top.uart_logics.data_0[25] ),
    .A2(_04808_),
    .Y(_04852_),
    .B1(net5234));
 sg13g2_a22oi_1 _20577_ (.Y(_04853_),
    .B1(_04813_),
    .B2(\fpga_top.uart_top.uart_logics.data_0[21] ),
    .A2(_04807_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[9] ));
 sg13g2_nand4_1 _20578_ (.B(_04851_),
    .C(_04852_),
    .A(_04850_),
    .Y(_04854_),
    .D(_04853_));
 sg13g2_a21oi_1 _20579_ (.A1(\fpga_top.bus_gather.i_read_adr[5] ),
    .A2(_04814_),
    .Y(_04855_),
    .B1(net5229));
 sg13g2_a22oi_1 _20580_ (.Y(_04856_),
    .B1(_04813_),
    .B2(\fpga_top.bus_gather.i_read_adr[21] ),
    .A2(_04808_),
    .A1(\fpga_top.bus_gather.i_read_adr[25] ));
 sg13g2_a22oi_1 _20581_ (.Y(_04857_),
    .B1(_04811_),
    .B2(\fpga_top.bus_gather.i_read_adr[13] ),
    .A2(_04807_),
    .A1(\fpga_top.bus_gather.i_read_adr[9] ));
 sg13g2_nand3_1 _20582_ (.B(_04856_),
    .C(_04857_),
    .A(_04855_),
    .Y(_04858_));
 sg13g2_a21oi_1 _20583_ (.A1(_06641_),
    .A2(net5234),
    .Y(_04859_),
    .B1(_04810_));
 sg13g2_o21ai_1 _20584_ (.B1(_04859_),
    .Y(_04860_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[29] ),
    .A2(net5234));
 sg13g2_o21ai_1 _20585_ (.B1(_04816_),
    .Y(_04861_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[17] ),
    .A2(net5235));
 sg13g2_a21o_1 _20586_ (.A2(net5234),
    .A1(_06611_),
    .B1(_04861_),
    .X(_04862_));
 sg13g2_nand3_1 _20587_ (.B(_04860_),
    .C(_04862_),
    .A(_08745_),
    .Y(_04863_));
 sg13g2_a21oi_2 _20588_ (.B1(_04863_),
    .Y(_04864_),
    .A2(_04858_),
    .A1(_04854_));
 sg13g2_o21ai_1 _20589_ (.B1(_04813_),
    .Y(_04865_),
    .A1(net5591),
    .A2(net5229));
 sg13g2_a21oi_1 _20590_ (.A1(_06861_),
    .A2(net5229),
    .Y(_04866_),
    .B1(_04865_));
 sg13g2_o21ai_1 _20591_ (.B1(_04809_),
    .Y(_04867_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[30] ),
    .A2(net5231));
 sg13g2_a21oi_1 _20592_ (.A1(_06643_),
    .A2(net5230),
    .Y(_04868_),
    .B1(_04867_));
 sg13g2_o21ai_1 _20593_ (.B1(_04808_),
    .Y(_04869_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[26] ),
    .A2(net5233));
 sg13g2_a21oi_1 _20594_ (.A1(_06634_),
    .A2(net5230),
    .Y(_04870_),
    .B1(_04869_));
 sg13g2_o21ai_1 _20595_ (.B1(_04811_),
    .Y(_04871_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[14] ),
    .A2(net5230));
 sg13g2_a21oi_1 _20596_ (.A1(_06603_),
    .A2(net5230),
    .Y(_04872_),
    .B1(_04871_));
 sg13g2_o21ai_1 _20597_ (.B1(_04814_),
    .Y(_04873_),
    .A1(net5596),
    .A2(net5229));
 sg13g2_a21oi_1 _20598_ (.A1(_06860_),
    .A2(_06992_),
    .Y(_04874_),
    .B1(_04873_));
 sg13g2_o21ai_1 _20599_ (.B1(_04807_),
    .Y(_04875_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[10] ),
    .A2(net5231));
 sg13g2_a21oi_1 _20600_ (.A1(_06594_),
    .A2(net5230),
    .Y(_04876_),
    .B1(_04875_));
 sg13g2_o21ai_1 _20601_ (.B1(_04816_),
    .Y(_04877_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[18] ),
    .A2(net5232));
 sg13g2_a21oi_1 _20602_ (.A1(_06614_),
    .A2(net5230),
    .Y(_04878_),
    .B1(_04877_));
 sg13g2_o21ai_1 _20603_ (.B1(_04823_),
    .Y(_04879_),
    .A1(\fpga_top.uart_top.uart_logics.data_0[2] ),
    .A2(net5234));
 sg13g2_a21oi_1 _20604_ (.A1(net5386),
    .A2(net5232),
    .Y(_04880_),
    .B1(_04879_));
 sg13g2_nor4_1 _20605_ (.A(_04866_),
    .B(_04870_),
    .C(_04874_),
    .D(_04878_),
    .Y(_04881_));
 sg13g2_nor4_1 _20606_ (.A(_04868_),
    .B(_04872_),
    .C(_04876_),
    .D(_04880_),
    .Y(_04882_));
 sg13g2_and2_1 _20607_ (.A(_04881_),
    .B(_04882_),
    .X(_04883_));
 sg13g2_nand2_1 _20608_ (.Y(_04884_),
    .A(_04864_),
    .B(_04883_));
 sg13g2_a21oi_1 _20609_ (.A1(_04864_),
    .A2(_04883_),
    .Y(_04885_),
    .B1(_04849_));
 sg13g2_o21ai_1 _20610_ (.B1(net5341),
    .Y(_04886_),
    .A1(_04830_),
    .A2(_04885_));
 sg13g2_a21oi_1 _20611_ (.A1(_04830_),
    .A2(_04885_),
    .Y(_04887_),
    .B1(_04886_));
 sg13g2_a21oi_2 _20612_ (.B1(_04887_),
    .Y(_04888_),
    .A2(_04805_),
    .A1(net5340));
 sg13g2_nand2_1 _20613_ (.Y(_04889_),
    .A(net1431),
    .B(net4879));
 sg13g2_o21ai_1 _20614_ (.B1(_04889_),
    .Y(_01441_),
    .A1(net4879),
    .A2(_04888_));
 sg13g2_nand2b_1 _20615_ (.Y(_04890_),
    .B(net5711),
    .A_N(\fpga_top.io_uart_out.uart_io_char[1] ));
 sg13g2_o21ai_1 _20616_ (.B1(_04890_),
    .Y(_04891_),
    .A1(net5711),
    .A2(\fpga_top.io_uart_out.rout[1] ));
 sg13g2_or2_1 _20617_ (.X(_04892_),
    .B(_04849_),
    .A(_04830_));
 sg13g2_inv_1 _20618_ (.Y(_04893_),
    .A(_04892_));
 sg13g2_xor2_1 _20619_ (.B(_04892_),
    .A(_04864_),
    .X(_04894_));
 sg13g2_nand3_1 _20620_ (.B(_04884_),
    .C(_04894_),
    .A(net5341),
    .Y(_04895_));
 sg13g2_o21ai_1 _20621_ (.B1(_04895_),
    .Y(_04896_),
    .A1(net5341),
    .A2(_04891_));
 sg13g2_mux2_1 _20622_ (.A0(_04896_),
    .A1(net2533),
    .S(net4879),
    .X(_01442_));
 sg13g2_a21o_1 _20623_ (.A2(_04893_),
    .A1(_04864_),
    .B1(_04883_),
    .X(_04897_));
 sg13g2_a21oi_1 _20624_ (.A1(net5425),
    .A2(_08740_),
    .Y(_04898_),
    .B1(net5340));
 sg13g2_nor2b_1 _20625_ (.A(net5711),
    .B_N(\fpga_top.io_uart_out.rout[2] ),
    .Y(_04899_));
 sg13g2_a21oi_1 _20626_ (.A1(net5712),
    .A2(\fpga_top.io_uart_out.uart_io_char[2] ),
    .Y(_04900_),
    .B1(_04899_));
 sg13g2_a22oi_1 _20627_ (.Y(_04901_),
    .B1(_04900_),
    .B2(net5340),
    .A2(_04898_),
    .A1(_04897_));
 sg13g2_mux2_1 _20628_ (.A0(_04901_),
    .A1(net3679),
    .S(net4879),
    .X(_01443_));
 sg13g2_or2_1 _20629_ (.X(_04902_),
    .B(_04884_),
    .A(_04849_));
 sg13g2_nor2_1 _20630_ (.A(_08740_),
    .B(net5340),
    .Y(_04903_));
 sg13g2_nor2b_1 _20631_ (.A(net5711),
    .B_N(\fpga_top.io_uart_out.rout[3] ),
    .Y(_04904_));
 sg13g2_a21oi_1 _20632_ (.A1(net5712),
    .A2(\fpga_top.io_uart_out.uart_io_char[3] ),
    .Y(_04905_),
    .B1(_04904_));
 sg13g2_a22oi_1 _20633_ (.Y(_04906_),
    .B1(_04905_),
    .B2(net5340),
    .A2(_04903_),
    .A1(_04902_));
 sg13g2_mux2_1 _20634_ (.A0(_04906_),
    .A1(net2881),
    .S(net4879),
    .X(_01444_));
 sg13g2_o21ai_1 _20635_ (.B1(net5422),
    .Y(_04907_),
    .A1(net5423),
    .A2(\fpga_top.uart_top.uart_send_char.send_cntr[2] ));
 sg13g2_nand3b_1 _20636_ (.B(_04903_),
    .C(_04907_),
    .Y(_04908_),
    .A_N(_04885_));
 sg13g2_nand2b_1 _20637_ (.Y(_04909_),
    .B(net5713),
    .A_N(\fpga_top.io_uart_out.uart_io_char[4] ));
 sg13g2_o21ai_1 _20638_ (.B1(_04909_),
    .Y(_04910_),
    .A1(net5711),
    .A2(\fpga_top.io_uart_out.rout[4] ));
 sg13g2_o21ai_1 _20639_ (.B1(_04908_),
    .Y(_04911_),
    .A1(net5341),
    .A2(_04910_));
 sg13g2_mux2_1 _20640_ (.A0(_04911_),
    .A1(net2177),
    .S(_04804_),
    .X(_01445_));
 sg13g2_mux2_1 _20641_ (.A0(\fpga_top.io_uart_out.rout[5] ),
    .A1(\fpga_top.io_uart_out.uart_io_char[5] ),
    .S(net5711),
    .X(_04912_));
 sg13g2_a21o_2 _20642_ (.A2(_04912_),
    .A1(net5340),
    .B1(_04903_),
    .X(_04913_));
 sg13g2_mux2_1 _20643_ (.A0(_04913_),
    .A1(net2886),
    .S(net4879),
    .X(_01446_));
 sg13g2_nand2b_1 _20644_ (.Y(_04914_),
    .B(net5713),
    .A_N(\fpga_top.io_uart_out.uart_io_char[6] ));
 sg13g2_o21ai_1 _20645_ (.B1(_04914_),
    .Y(_04915_),
    .A1(net5711),
    .A2(\fpga_top.io_uart_out.rout[6] ));
 sg13g2_nand2_1 _20646_ (.Y(_04916_),
    .A(net5341),
    .B(_04885_));
 sg13g2_o21ai_1 _20647_ (.B1(_04916_),
    .Y(_04917_),
    .A1(net5341),
    .A2(_04915_));
 sg13g2_mux2_1 _20648_ (.A0(_04917_),
    .A1(net3240),
    .S(net4879),
    .X(_01447_));
 sg13g2_o21ai_1 _20649_ (.B1(net5340),
    .Y(_04918_),
    .A1(net5713),
    .A2(\fpga_top.io_uart_out.rout[7] ));
 sg13g2_a21oi_2 _20650_ (.B1(_04918_),
    .Y(_04919_),
    .A2(_06862_),
    .A1(net5713));
 sg13g2_mux2_1 _20651_ (.A0(_04919_),
    .A1(net2809),
    .S(net4879),
    .X(_01448_));
 sg13g2_nand3_1 _20652_ (.B(_07575_),
    .C(_03921_),
    .A(_06557_),
    .Y(_04920_));
 sg13g2_nor3_2 _20653_ (.A(_07290_),
    .B(_03915_),
    .C(_04920_),
    .Y(_04921_));
 sg13g2_nand2_2 _20654_ (.Y(_04922_),
    .A(\fpga_top.cpu_top.csr_rmie ),
    .B(_04921_));
 sg13g2_nand2_2 _20655_ (.Y(_04923_),
    .A(_03929_),
    .B(_04922_));
 sg13g2_nand2_2 _20656_ (.Y(_04924_),
    .A(_06773_),
    .B(_08916_));
 sg13g2_and2_1 _20657_ (.A(net4777),
    .B(net5255),
    .X(_04925_));
 sg13g2_nand2_1 _20658_ (.Y(_04926_),
    .A(net4777),
    .B(net5256));
 sg13g2_nor2_1 _20659_ (.A(net1810),
    .B(net4741),
    .Y(_04927_));
 sg13g2_a21oi_1 _20660_ (.A1(net5386),
    .A2(net4741),
    .Y(_01449_),
    .B1(_04927_));
 sg13g2_nand2_1 _20661_ (.Y(_04928_),
    .A(net1699),
    .B(net4727));
 sg13g2_o21ai_1 _20662_ (.B1(_04928_),
    .Y(_01450_),
    .A1(_06584_),
    .A2(net4727));
 sg13g2_mux2_1 _20663_ (.A0(net5598),
    .A1(net3367),
    .S(net4727),
    .X(_01451_));
 sg13g2_nand2_1 _20664_ (.Y(_04929_),
    .A(net1520),
    .B(net4728));
 sg13g2_o21ai_1 _20665_ (.B1(_04929_),
    .Y(_01452_),
    .A1(_06587_),
    .A2(net4728));
 sg13g2_nand2_1 _20666_ (.Y(_04930_),
    .A(net1475),
    .B(net4728));
 sg13g2_o21ai_1 _20667_ (.B1(_04930_),
    .Y(_01453_),
    .A1(_06588_),
    .A2(net4728));
 sg13g2_nand2_1 _20668_ (.Y(_04931_),
    .A(net1541),
    .B(net4729));
 sg13g2_o21ai_1 _20669_ (.B1(_04931_),
    .Y(_01454_),
    .A1(_06590_),
    .A2(net4729));
 sg13g2_mux2_1 _20670_ (.A0(net2541),
    .A1(net3312),
    .S(net4727),
    .X(_01455_));
 sg13g2_nand2_1 _20671_ (.Y(_04932_),
    .A(net1477),
    .B(net4731));
 sg13g2_o21ai_1 _20672_ (.B1(_04932_),
    .Y(_01456_),
    .A1(_06592_),
    .A2(net4731));
 sg13g2_nand2_1 _20673_ (.Y(_04933_),
    .A(net1417),
    .B(net4731));
 sg13g2_o21ai_1 _20674_ (.B1(_04933_),
    .Y(_01457_),
    .A1(_06594_),
    .A2(net4731));
 sg13g2_nand2_1 _20675_ (.Y(_04934_),
    .A(net1509),
    .B(net4729));
 sg13g2_o21ai_1 _20676_ (.B1(_04934_),
    .Y(_01458_),
    .A1(_06597_),
    .A2(net4729));
 sg13g2_nand2_1 _20677_ (.Y(_04935_),
    .A(net1531),
    .B(net4731));
 sg13g2_o21ai_1 _20678_ (.B1(_04935_),
    .Y(_01459_),
    .A1(_06599_),
    .A2(net4730));
 sg13g2_nand2_1 _20679_ (.Y(_04936_),
    .A(net1495),
    .B(net4730));
 sg13g2_o21ai_1 _20680_ (.B1(_04936_),
    .Y(_01460_),
    .A1(_06601_),
    .A2(net4730));
 sg13g2_nand2_1 _20681_ (.Y(_04937_),
    .A(net1550),
    .B(net4730));
 sg13g2_o21ai_1 _20682_ (.B1(_04937_),
    .Y(_01461_),
    .A1(_06603_),
    .A2(net4730));
 sg13g2_nand2_1 _20683_ (.Y(_04938_),
    .A(net1446),
    .B(net4732));
 sg13g2_o21ai_1 _20684_ (.B1(_04938_),
    .Y(_01462_),
    .A1(_06605_),
    .A2(net4730));
 sg13g2_mux2_1 _20685_ (.A0(net5594),
    .A1(net3753),
    .S(net4734),
    .X(_01463_));
 sg13g2_nand2_1 _20686_ (.Y(_04939_),
    .A(net1440),
    .B(net4735));
 sg13g2_o21ai_1 _20687_ (.B1(_04939_),
    .Y(_01464_),
    .A1(_06611_),
    .A2(net4735));
 sg13g2_nand2_1 _20688_ (.Y(_04940_),
    .A(net1524),
    .B(net4733));
 sg13g2_o21ai_1 _20689_ (.B1(_04940_),
    .Y(_01465_),
    .A1(_06614_),
    .A2(net4733));
 sg13g2_nand2_1 _20690_ (.Y(_04941_),
    .A(net1582),
    .B(net4736));
 sg13g2_o21ai_1 _20691_ (.B1(_04941_),
    .Y(_01466_),
    .A1(_06617_),
    .A2(net4736));
 sg13g2_nand2_1 _20692_ (.Y(_04942_),
    .A(net1512),
    .B(net4734));
 sg13g2_o21ai_1 _20693_ (.B1(_04942_),
    .Y(_01467_),
    .A1(_06620_),
    .A2(net4734));
 sg13g2_nand2_1 _20694_ (.Y(_04943_),
    .A(net1506),
    .B(net4735));
 sg13g2_o21ai_1 _20695_ (.B1(_04943_),
    .Y(_01468_),
    .A1(_06623_),
    .A2(net4737));
 sg13g2_mux2_1 _20696_ (.A0(net5592),
    .A1(net3779),
    .S(net4735),
    .X(_01469_));
 sg13g2_nand2_1 _20697_ (.Y(_04944_),
    .A(net1555),
    .B(net4735));
 sg13g2_o21ai_1 _20698_ (.B1(_04944_),
    .Y(_01470_),
    .A1(_06626_),
    .A2(net4735));
 sg13g2_nand2_1 _20699_ (.Y(_04945_),
    .A(net1546),
    .B(net4738));
 sg13g2_o21ai_1 _20700_ (.B1(_04945_),
    .Y(_01471_),
    .A1(_06629_),
    .A2(net4735));
 sg13g2_nor2_1 _20701_ (.A(net1944),
    .B(net4742),
    .Y(_04946_));
 sg13g2_a21oi_1 _20702_ (.A1(_06631_),
    .A2(net4742),
    .Y(_01472_),
    .B1(_04946_));
 sg13g2_nand2_1 _20703_ (.Y(_04947_),
    .A(net1600),
    .B(net4737));
 sg13g2_o21ai_1 _20704_ (.B1(_04947_),
    .Y(_01473_),
    .A1(_06634_),
    .A2(net4737));
 sg13g2_nand2_1 _20705_ (.Y(_04948_),
    .A(net1591),
    .B(net4736));
 sg13g2_o21ai_1 _20706_ (.B1(_04948_),
    .Y(_01474_),
    .A1(_06636_),
    .A2(net4736));
 sg13g2_mux2_1 _20707_ (.A0(\fpga_top.bus_gather.i_read_adr[28] ),
    .A1(net3647),
    .S(net4738),
    .X(_01475_));
 sg13g2_nor2_1 _20708_ (.A(net2027),
    .B(net4743),
    .Y(_04949_));
 sg13g2_a21oi_1 _20709_ (.A1(_06641_),
    .A2(net4742),
    .Y(_01476_),
    .B1(_04949_));
 sg13g2_nand2_1 _20710_ (.Y(_04950_),
    .A(net1676),
    .B(net4736));
 sg13g2_o21ai_1 _20711_ (.B1(_04950_),
    .Y(_01477_),
    .A1(_06643_),
    .A2(net4735));
 sg13g2_nand2_1 _20712_ (.Y(_04951_),
    .A(net1438),
    .B(net4733));
 sg13g2_o21ai_1 _20713_ (.B1(_04951_),
    .Y(_01478_),
    .A1(_06646_),
    .A2(net4733));
 sg13g2_and4_1 _20714_ (.A(\fpga_top.cpu_top.br_ofs[8] ),
    .B(\fpga_top.cpu_top.br_ofs[9] ),
    .C(_07288_),
    .D(_03914_),
    .X(_04952_));
 sg13g2_nand4_1 _20715_ (.B(_06563_),
    .C(_06575_),
    .A(\fpga_top.cpu_top.alui_shamt[1] ),
    .Y(_04953_),
    .D(_04952_));
 sg13g2_nor2_1 _20716_ (.A(_04920_),
    .B(_04953_),
    .Y(_04954_));
 sg13g2_nor3_2 _20717_ (.A(net5273),
    .B(_04920_),
    .C(_04953_),
    .Y(_04955_));
 sg13g2_nand3b_1 _20718_ (.B(_06557_),
    .C(_03913_),
    .Y(_04956_),
    .A_N(_04953_));
 sg13g2_o21ai_1 _20719_ (.B1(net4727),
    .Y(_01479_),
    .A1(_06772_),
    .A2(_04955_));
 sg13g2_nand3_1 _20720_ (.B(_07036_),
    .C(_09892_),
    .A(net5574),
    .Y(_04957_));
 sg13g2_nand4_1 _20721_ (.B(_09853_),
    .C(_09857_),
    .A(_07706_),
    .Y(_04958_),
    .D(_09870_));
 sg13g2_o21ai_1 _20722_ (.B1(_04958_),
    .Y(_04959_),
    .A1(net5574),
    .A2(_07303_));
 sg13g2_o21ai_1 _20723_ (.B1(_04959_),
    .Y(_04960_),
    .A1(_07037_),
    .A2(_04958_));
 sg13g2_or2_1 _20724_ (.X(_04961_),
    .B(_09892_),
    .A(_07602_));
 sg13g2_mux2_1 _20725_ (.A0(_07607_),
    .A1(_07609_),
    .S(_09893_),
    .X(_04962_));
 sg13g2_nand4_1 _20726_ (.B(_04960_),
    .C(_04961_),
    .A(_04957_),
    .Y(_04963_),
    .D(_04962_));
 sg13g2_a21oi_2 _20727_ (.B1(net5213),
    .Y(_04964_),
    .A2(_04963_),
    .A1(_03905_));
 sg13g2_inv_1 _20728_ (.Y(_04965_),
    .A(net4578));
 sg13g2_o21ai_1 _20729_ (.B1(\fpga_top.cpu_top.csr_rmie ),
    .Y(_04966_),
    .A1(\fpga_top.cpu_top.pc_stage.frc_cntr_val_leq_latch ),
    .A2(\fpga_top.cpu_top.pc_stage.g_interrupt_latch ));
 sg13g2_nand3_1 _20730_ (.B(_04922_),
    .C(_04966_),
    .A(_03929_),
    .Y(_04967_));
 sg13g2_nor2_2 _20731_ (.A(net4875),
    .B(_04967_),
    .Y(_04968_));
 sg13g2_nand2b_2 _20732_ (.Y(_04969_),
    .B(net5043),
    .A_N(_04967_));
 sg13g2_nor2_2 _20733_ (.A(net4562),
    .B(net4723),
    .Y(_04970_));
 sg13g2_nor2_1 _20734_ (.A(net5275),
    .B(_04970_),
    .Y(_04971_));
 sg13g2_o21ai_1 _20735_ (.B1(net5278),
    .Y(_04972_),
    .A1(net4561),
    .A2(net4724));
 sg13g2_nor2_1 _20736_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[0] ),
    .B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[1] ),
    .Y(_04973_));
 sg13g2_or2_1 _20737_ (.X(_04974_),
    .B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[1] ),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[0] ));
 sg13g2_nor4_2 _20738_ (.A(\fpga_top.cpu_top.pc_stage.frc_cntr_val_leq_latch ),
    .B(\fpga_top.cpu_top.pc_stage.g_interrupt_latch ),
    .C(_06771_),
    .Y(_04975_),
    .D(net5272));
 sg13g2_nand2_1 _20739_ (.Y(_04976_),
    .A(\fpga_top.cpu_top.pc_stage.cmd_ecall_pc_pre ),
    .B(_04975_));
 sg13g2_and2_1 _20740_ (.A(\fpga_top.cpu_top.pc_stage.cmd_ebreak_pc_pre ),
    .B(_04975_),
    .X(_04977_));
 sg13g2_nand2_2 _20741_ (.Y(_04978_),
    .A(\fpga_top.cpu_top.pc_stage.cmd_ebreak_pc_pre ),
    .B(_04975_));
 sg13g2_nor2_1 _20742_ (.A(net5253),
    .B(net5042),
    .Y(_04979_));
 sg13g2_nand4_1 _20743_ (.B(_03928_),
    .C(_04976_),
    .A(_03927_),
    .Y(_04980_),
    .D(_04979_));
 sg13g2_a21oi_1 _20744_ (.A1(_04974_),
    .A2(_04980_),
    .Y(_04981_),
    .B1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[2] ));
 sg13g2_and2_1 _20745_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[2] ),
    .B(_04980_),
    .X(_04982_));
 sg13g2_and2_1 _20746_ (.A(net5043),
    .B(_04967_),
    .X(_04983_));
 sg13g2_nand2_2 _20747_ (.Y(_04984_),
    .A(net5043),
    .B(_04967_));
 sg13g2_a21oi_1 _20748_ (.A1(net5315),
    .A2(_04982_),
    .Y(_04985_),
    .B1(_04981_));
 sg13g2_nor2_1 _20749_ (.A(_08155_),
    .B(net4724),
    .Y(_04986_));
 sg13g2_a221oi_1 _20750_ (.B2(_04985_),
    .C1(_04986_),
    .B1(net4719),
    .A1(net1964),
    .Y(_04987_),
    .A2(net4875));
 sg13g2_nand2b_1 _20751_ (.Y(_04988_),
    .B(net4497),
    .A_N(_04987_));
 sg13g2_nor2_2 _20752_ (.A(net5588),
    .B(net5273),
    .Y(_04989_));
 sg13g2_nand2_2 _20753_ (.Y(_04990_),
    .A(_06775_),
    .B(net5279));
 sg13g2_a21oi_1 _20754_ (.A1(net5386),
    .A2(_04970_),
    .Y(_04991_),
    .B1(_04990_));
 sg13g2_nor2_1 _20755_ (.A(net6410),
    .B(net5278),
    .Y(_04992_));
 sg13g2_nor2_1 _20756_ (.A(_06775_),
    .B(net5273),
    .Y(_04993_));
 sg13g2_nand2_2 _20757_ (.Y(_04994_),
    .A(net5588),
    .B(net5279));
 sg13g2_a221oi_1 _20758_ (.B2(_06684_),
    .C1(_04992_),
    .B1(net5117),
    .A1(_04988_),
    .Y(_01480_),
    .A2(_04991_));
 sg13g2_nor2_1 _20759_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[3] ),
    .B(_04982_),
    .Y(_04995_));
 sg13g2_a21o_1 _20760_ (.A2(_04980_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[2] ),
    .B1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[3] ),
    .X(_04996_));
 sg13g2_o21ai_1 _20761_ (.B1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[3] ),
    .Y(_04997_),
    .A1(_04973_),
    .A2(_04982_));
 sg13g2_a21oi_1 _20762_ (.A1(net5315),
    .A2(_04995_),
    .Y(_04998_),
    .B1(_04984_));
 sg13g2_or2_1 _20763_ (.X(_04999_),
    .B(net5043),
    .A(\fpga_top.cpu_top.csr_mepc_ex[3] ));
 sg13g2_o21ai_1 _20764_ (.B1(_04999_),
    .Y(_05000_),
    .A1(_08186_),
    .A2(net4724));
 sg13g2_a21oi_1 _20765_ (.A1(_04997_),
    .A2(_04998_),
    .Y(_05001_),
    .B1(_05000_));
 sg13g2_a21oi_1 _20766_ (.A1(_08189_),
    .A2(net4540),
    .Y(_05002_),
    .B1(net5117));
 sg13g2_o21ai_1 _20767_ (.B1(_05002_),
    .Y(_05003_),
    .A1(net4540),
    .A2(_05001_));
 sg13g2_a21oi_1 _20768_ (.A1(net5587),
    .A2(net5662),
    .Y(_05004_),
    .B1(net5271));
 sg13g2_a22oi_1 _20769_ (.Y(_01481_),
    .B1(_05003_),
    .B2(_05004_),
    .A2(net5271),
    .A1(_06584_));
 sg13g2_a221oi_1 _20770_ (.B2(\fpga_top.cpu_top.pc_stage.cmd_ecall_pc_pre ),
    .C1(net5042),
    .B1(_04975_),
    .A1(_03927_),
    .Y(_05005_),
    .A2(_03928_));
 sg13g2_nand3_1 _20771_ (.B(_04976_),
    .C(net5033),
    .A(_03929_),
    .Y(_05006_));
 sg13g2_a21oi_1 _20772_ (.A1(_06773_),
    .A2(_05006_),
    .Y(_05007_),
    .B1(\fpga_top.cpu_top.execution.csr_array.g_interrupt ));
 sg13g2_o21ai_1 _20773_ (.B1(_08916_),
    .Y(_05008_),
    .A1(\fpga_top.cpu_top.execution.csr_array.frc_cntr_val_leq ),
    .A2(_05005_));
 sg13g2_nor2_1 _20774_ (.A(_06887_),
    .B(_05008_),
    .Y(_05009_));
 sg13g2_nand2_1 _20775_ (.Y(_05010_),
    .A(_06887_),
    .B(_05008_));
 sg13g2_nor2b_1 _20776_ (.A(_05009_),
    .B_N(_05010_),
    .Y(_05011_));
 sg13g2_xnor2_1 _20777_ (.Y(_05012_),
    .A(_04996_),
    .B(_05011_));
 sg13g2_o21ai_1 _20778_ (.B1(net4719),
    .Y(_05013_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[4] ),
    .A2(_04974_));
 sg13g2_a21oi_1 _20779_ (.A1(_04974_),
    .A2(_05012_),
    .Y(_05014_),
    .B1(_05013_));
 sg13g2_a221oi_1 _20780_ (.B2(_08218_),
    .C1(_05014_),
    .B1(net4726),
    .A1(net1878),
    .Y(_05015_),
    .A2(net4875));
 sg13g2_inv_1 _20781_ (.Y(_05016_),
    .A(_05015_));
 sg13g2_o21ai_1 _20782_ (.B1(_04989_),
    .Y(_05017_),
    .A1(_08221_),
    .A2(net4497));
 sg13g2_a21oi_1 _20783_ (.A1(net4499),
    .A2(_05016_),
    .Y(_05018_),
    .B1(_05017_));
 sg13g2_nor2_1 _20784_ (.A(net5597),
    .B(net5278),
    .Y(_05019_));
 sg13g2_nor2_1 _20785_ (.A(net5660),
    .B(_04994_),
    .Y(_05020_));
 sg13g2_nor3_1 _20786_ (.A(_05018_),
    .B(_05019_),
    .C(_05020_),
    .Y(_01482_));
 sg13g2_a21oi_1 _20787_ (.A1(_04996_),
    .A2(_05010_),
    .Y(_05021_),
    .B1(_05009_));
 sg13g2_a22oi_1 _20788_ (.Y(_05022_),
    .B1(net5033),
    .B2(_03929_),
    .A2(_04975_),
    .A1(\fpga_top.cpu_top.pc_stage.cmd_ecall_pc_pre ));
 sg13g2_o21ai_1 _20789_ (.B1(_08916_),
    .Y(_05023_),
    .A1(\fpga_top.cpu_top.execution.csr_array.frc_cntr_val_leq ),
    .A2(_05022_));
 sg13g2_nand2_1 _20790_ (.Y(_05024_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[5] ),
    .B(_05023_));
 sg13g2_xnor2_1 _20791_ (.Y(_05025_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[5] ),
    .B(_05023_));
 sg13g2_xnor2_1 _20792_ (.Y(_05026_),
    .A(_05021_),
    .B(_05025_));
 sg13g2_o21ai_1 _20793_ (.B1(net4719),
    .Y(_05027_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[5] ),
    .A2(net5315));
 sg13g2_a21oi_1 _20794_ (.A1(net5315),
    .A2(_05026_),
    .Y(_05028_),
    .B1(_05027_));
 sg13g2_a221oi_1 _20795_ (.B2(_08097_),
    .C1(_05028_),
    .B1(net4726),
    .A1(net1923),
    .Y(_05029_),
    .A2(net4875));
 sg13g2_nand2_1 _20796_ (.Y(_05030_),
    .A(_08099_),
    .B(net4540));
 sg13g2_nand2_1 _20797_ (.Y(_05031_),
    .A(net4497),
    .B(_05029_));
 sg13g2_nand3_1 _20798_ (.B(_05030_),
    .C(_05031_),
    .A(_04994_),
    .Y(_05032_));
 sg13g2_a21oi_1 _20799_ (.A1(net5587),
    .A2(net5659),
    .Y(_05033_),
    .B1(net5271));
 sg13g2_a22oi_1 _20800_ (.Y(_01483_),
    .B1(_05032_),
    .B2(_05033_),
    .A2(net5271),
    .A1(_06587_));
 sg13g2_nor2_2 _20801_ (.A(net5253),
    .B(_05006_),
    .Y(_05034_));
 sg13g2_and2_1 _20802_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[6] ),
    .B(_05034_),
    .X(_05035_));
 sg13g2_or2_1 _20803_ (.X(_05036_),
    .B(_05034_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[6] ));
 sg13g2_nand2b_1 _20804_ (.Y(_05037_),
    .B(_05036_),
    .A_N(_05035_));
 sg13g2_o21ai_1 _20805_ (.B1(_05024_),
    .Y(_05038_),
    .A1(_05021_),
    .A2(_05025_));
 sg13g2_xnor2_1 _20806_ (.Y(_05039_),
    .A(_05037_),
    .B(_05038_));
 sg13g2_mux2_1 _20807_ (.A0(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[6] ),
    .A1(_05039_),
    .S(net5315),
    .X(_05040_));
 sg13g2_and2_1 _20808_ (.A(_08243_),
    .B(net4726),
    .X(_05041_));
 sg13g2_a221oi_1 _20809_ (.B2(_05040_),
    .C1(_05041_),
    .B1(net4719),
    .A1(net2311),
    .Y(_05042_),
    .A2(net4875));
 sg13g2_inv_1 _20810_ (.Y(_05043_),
    .A(_05042_));
 sg13g2_o21ai_1 _20811_ (.B1(_04989_),
    .Y(_05044_),
    .A1(_08245_),
    .A2(net4497));
 sg13g2_a21oi_1 _20812_ (.A1(net4497),
    .A2(_05043_),
    .Y(_05045_),
    .B1(_05044_));
 sg13g2_a221oi_1 _20813_ (.B2(_06790_),
    .C1(_05045_),
    .B1(net5117),
    .A1(_06588_),
    .Y(_01484_),
    .A2(net5272));
 sg13g2_a21o_1 _20814_ (.A2(_05038_),
    .A1(_05036_),
    .B1(_05035_),
    .X(_05046_));
 sg13g2_xnor2_1 _20815_ (.Y(_05047_),
    .A(_06894_),
    .B(_05034_));
 sg13g2_a21oi_1 _20816_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[7] ),
    .A2(_05034_),
    .Y(_05048_),
    .B1(_05046_));
 sg13g2_xnor2_1 _20817_ (.Y(_05049_),
    .A(_05046_),
    .B(_05047_));
 sg13g2_o21ai_1 _20818_ (.B1(net4719),
    .Y(_05050_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[7] ),
    .A2(net5315));
 sg13g2_a21oi_1 _20819_ (.A1(net5315),
    .A2(_05049_),
    .Y(_05051_),
    .B1(_05050_));
 sg13g2_nand2_1 _20820_ (.Y(_05052_),
    .A(net2104),
    .B(net4875));
 sg13g2_a21oi_1 _20821_ (.A1(_08068_),
    .A2(net4726),
    .Y(_05053_),
    .B1(_05051_));
 sg13g2_nand3_1 _20822_ (.B(_05052_),
    .C(_05053_),
    .A(net4497),
    .Y(_05054_));
 sg13g2_a21oi_1 _20823_ (.A1(_08071_),
    .A2(net4540),
    .Y(_05055_),
    .B1(net5117));
 sg13g2_a221oi_1 _20824_ (.B2(_05055_),
    .C1(net5273),
    .B1(_05054_),
    .A1(net5587),
    .Y(_05056_),
    .A2(net5656));
 sg13g2_a21oi_1 _20825_ (.A1(_06590_),
    .A2(net5272),
    .Y(_01485_),
    .B1(_05056_));
 sg13g2_nand2_1 _20826_ (.Y(_05057_),
    .A(net2541),
    .B(net5273));
 sg13g2_o21ai_1 _20827_ (.B1(net5315),
    .Y(_05058_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[7] ),
    .A2(_05034_));
 sg13g2_or3_1 _20828_ (.A(_06900_),
    .B(_05048_),
    .C(_05058_),
    .X(_05059_));
 sg13g2_o21ai_1 _20829_ (.B1(_06900_),
    .Y(_05060_),
    .A1(_05048_),
    .A2(_05058_));
 sg13g2_and2_1 _20830_ (.A(net4719),
    .B(_05060_),
    .X(_05061_));
 sg13g2_and2_1 _20831_ (.A(_08124_),
    .B(net4726),
    .X(_05062_));
 sg13g2_a221oi_1 _20832_ (.B2(_05061_),
    .C1(_05062_),
    .B1(_05059_),
    .A1(\fpga_top.cpu_top.csr_mepc_ex[8] ),
    .Y(_05063_),
    .A2(net4875));
 sg13g2_nor2_1 _20833_ (.A(_08126_),
    .B(net4497),
    .Y(_05064_));
 sg13g2_o21ai_1 _20834_ (.B1(_06775_),
    .Y(_05065_),
    .A1(net4540),
    .A2(_05063_));
 sg13g2_nor2_1 _20835_ (.A(_05064_),
    .B(_05065_),
    .Y(_05066_));
 sg13g2_o21ai_1 _20836_ (.B1(net5278),
    .Y(_05067_),
    .A1(_06775_),
    .A2(net5655));
 sg13g2_o21ai_1 _20837_ (.B1(_05057_),
    .Y(_01486_),
    .A1(_05066_),
    .A2(_05067_));
 sg13g2_nor2_2 _20838_ (.A(_06902_),
    .B(_05059_),
    .Y(_05068_));
 sg13g2_xnor2_1 _20839_ (.Y(_05069_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[9] ),
    .B(_05059_));
 sg13g2_a22oi_1 _20840_ (.Y(_05070_),
    .B1(net4719),
    .B2(_05069_),
    .A2(net4878),
    .A1(net2122));
 sg13g2_o21ai_1 _20841_ (.B1(_05070_),
    .Y(_05071_),
    .A1(_08309_),
    .A2(net4724));
 sg13g2_o21ai_1 _20842_ (.B1(_04989_),
    .Y(_05072_),
    .A1(_08311_),
    .A2(net4498));
 sg13g2_a21oi_1 _20843_ (.A1(net4498),
    .A2(_05071_),
    .Y(_05073_),
    .B1(_05072_));
 sg13g2_a221oi_1 _20844_ (.B2(_06792_),
    .C1(_05073_),
    .B1(net5117),
    .A1(_06592_),
    .Y(_01487_),
    .A2(net5274));
 sg13g2_o21ai_1 _20845_ (.B1(_04989_),
    .Y(_05074_),
    .A1(_08010_),
    .A2(net4498));
 sg13g2_xnor2_1 _20846_ (.Y(_05075_),
    .A(net6229),
    .B(_05068_));
 sg13g2_or2_1 _20847_ (.X(_05076_),
    .B(net5043),
    .A(net2284));
 sg13g2_o21ai_1 _20848_ (.B1(_05076_),
    .Y(_05077_),
    .A1(_08008_),
    .A2(net4724));
 sg13g2_a21oi_1 _20849_ (.A1(net4720),
    .A2(_05075_),
    .Y(_05078_),
    .B1(_05077_));
 sg13g2_a21oi_1 _20850_ (.A1(net4498),
    .A2(_05078_),
    .Y(_05079_),
    .B1(_05074_));
 sg13g2_a221oi_1 _20851_ (.B2(_06679_),
    .C1(_05079_),
    .B1(net5117),
    .A1(_06594_),
    .Y(_01488_),
    .A2(net5273));
 sg13g2_nand3_1 _20852_ (.B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[11] ),
    .C(_05068_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[10] ),
    .Y(_05080_));
 sg13g2_a21o_1 _20853_ (.A2(_05068_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[10] ),
    .B1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[11] ),
    .X(_05081_));
 sg13g2_nand2_1 _20854_ (.Y(_05082_),
    .A(_05080_),
    .B(_05081_));
 sg13g2_nor3_1 _20855_ (.A(\fpga_top.cpu_top.csr_mepc_ex[11] ),
    .B(_04920_),
    .C(_04953_),
    .Y(_05083_));
 sg13g2_a221oi_1 _20856_ (.B2(_05082_),
    .C1(_05083_),
    .B1(net4719),
    .A1(_08251_),
    .Y(_05084_),
    .A2(net4726));
 sg13g2_a21oi_1 _20857_ (.A1(net4497),
    .A2(_05084_),
    .Y(_05085_),
    .B1(net5588));
 sg13g2_o21ai_1 _20858_ (.B1(_05085_),
    .Y(_05086_),
    .A1(_08275_),
    .A2(net4499));
 sg13g2_a21oi_1 _20859_ (.A1(net5587),
    .A2(_06793_),
    .Y(_05087_),
    .B1(net5271));
 sg13g2_a22oi_1 _20860_ (.Y(_05088_),
    .B1(_05086_),
    .B2(_05087_),
    .A2(net5274),
    .A1(net6510));
 sg13g2_inv_1 _20861_ (.Y(_01489_),
    .A(_05088_));
 sg13g2_nor2_1 _20862_ (.A(_08343_),
    .B(net4498),
    .Y(_05089_));
 sg13g2_nand4_1 _20863_ (.B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[11] ),
    .C(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[12] ),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[10] ),
    .Y(_05090_),
    .D(_05068_));
 sg13g2_xnor2_1 _20864_ (.Y(_05091_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[12] ),
    .B(_05080_));
 sg13g2_nor2_1 _20865_ (.A(_08339_),
    .B(net4724),
    .Y(_05092_));
 sg13g2_a221oi_1 _20866_ (.B2(_05091_),
    .C1(_05092_),
    .B1(net4720),
    .A1(\fpga_top.cpu_top.csr_mepc_ex[12] ),
    .Y(_05093_),
    .A2(net4878));
 sg13g2_o21ai_1 _20867_ (.B1(_04994_),
    .Y(_05094_),
    .A1(net4540),
    .A2(_05093_));
 sg13g2_o21ai_1 _20868_ (.B1(net5279),
    .Y(_05095_),
    .A1(_05089_),
    .A2(_05094_));
 sg13g2_a21oi_1 _20869_ (.A1(net5587),
    .A2(net5375),
    .Y(_05096_),
    .B1(_05095_));
 sg13g2_a21o_1 _20870_ (.A2(net5274),
    .A1(net6488),
    .B1(_05096_),
    .X(_01490_));
 sg13g2_o21ai_1 _20871_ (.B1(_04989_),
    .Y(_05097_),
    .A1(_07968_),
    .A2(net4499));
 sg13g2_nor2_2 _20872_ (.A(_06907_),
    .B(_05090_),
    .Y(_05098_));
 sg13g2_xnor2_1 _20873_ (.Y(_05099_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[13] ),
    .B(_05090_));
 sg13g2_nor2_1 _20874_ (.A(_07965_),
    .B(net4724),
    .Y(_05100_));
 sg13g2_a221oi_1 _20875_ (.B2(_05099_),
    .C1(_05100_),
    .B1(net4720),
    .A1(net2103),
    .Y(_05101_),
    .A2(net4875));
 sg13g2_inv_1 _20876_ (.Y(_05102_),
    .A(_05101_));
 sg13g2_a21oi_1 _20877_ (.A1(net4499),
    .A2(_05102_),
    .Y(_05103_),
    .B1(_05097_));
 sg13g2_a221oi_1 _20878_ (.B2(net5374),
    .C1(_05103_),
    .B1(net5120),
    .A1(_06601_),
    .Y(_01491_),
    .A2(net5277));
 sg13g2_xnor2_1 _20879_ (.Y(_05104_),
    .A(net6199),
    .B(_05098_));
 sg13g2_nor2_1 _20880_ (.A(net1979),
    .B(net5043),
    .Y(_05105_));
 sg13g2_a221oi_1 _20881_ (.B2(_05104_),
    .C1(_05105_),
    .B1(net4720),
    .A1(_07939_),
    .Y(_05106_),
    .A2(net4726));
 sg13g2_o21ai_1 _20882_ (.B1(_04989_),
    .Y(_05107_),
    .A1(_07941_),
    .A2(net4498));
 sg13g2_a21oi_1 _20883_ (.A1(net4498),
    .A2(_05106_),
    .Y(_05108_),
    .B1(_05107_));
 sg13g2_a221oi_1 _20884_ (.B2(_06796_),
    .C1(_05108_),
    .B1(net5120),
    .A1(_06603_),
    .Y(_01492_),
    .A2(net5277));
 sg13g2_nand3_1 _20885_ (.B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[15] ),
    .C(_05098_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[14] ),
    .Y(_05109_));
 sg13g2_a21oi_1 _20886_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[14] ),
    .A2(_05098_),
    .Y(_05110_),
    .B1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[15] ));
 sg13g2_nor2_1 _20887_ (.A(_04984_),
    .B(_05110_),
    .Y(_05111_));
 sg13g2_nand2_1 _20888_ (.Y(_05112_),
    .A(net1817),
    .B(net4876));
 sg13g2_a22oi_1 _20889_ (.Y(_05113_),
    .B1(_05109_),
    .B2(_05111_),
    .A2(net4725),
    .A1(_08530_));
 sg13g2_a21oi_1 _20890_ (.A1(_05112_),
    .A2(_05113_),
    .Y(_05114_),
    .B1(net4539));
 sg13g2_o21ai_1 _20891_ (.B1(_06775_),
    .Y(_05115_),
    .A1(_08546_),
    .A2(net4498));
 sg13g2_a21oi_1 _20892_ (.A1(net5589),
    .A2(net5373),
    .Y(_05116_),
    .B1(net5277));
 sg13g2_o21ai_1 _20893_ (.B1(_05116_),
    .Y(_05117_),
    .A1(_05114_),
    .A2(_05115_));
 sg13g2_o21ai_1 _20894_ (.B1(_05117_),
    .Y(_01493_),
    .A1(_06605_),
    .A2(net5279));
 sg13g2_and4_1 _20895_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[14] ),
    .B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[15] ),
    .C(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[16] ),
    .D(_05098_),
    .X(_05118_));
 sg13g2_xnor2_1 _20896_ (.Y(_05119_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[16] ),
    .B(_05109_));
 sg13g2_nor2_1 _20897_ (.A(_08032_),
    .B(net4723),
    .Y(_05120_));
 sg13g2_a221oi_1 _20898_ (.B2(_05119_),
    .C1(_05120_),
    .B1(net4721),
    .A1(\fpga_top.cpu_top.csr_mepc_ex[16] ),
    .Y(_05121_),
    .A2(net4876));
 sg13g2_nand2b_1 _20899_ (.Y(_05122_),
    .B(net4500),
    .A_N(_05121_));
 sg13g2_a21oi_1 _20900_ (.A1(_08036_),
    .A2(net4539),
    .Y(_05123_),
    .B1(net5119));
 sg13g2_a221oi_1 _20901_ (.B2(_05123_),
    .C1(net5277),
    .B1(_05122_),
    .A1(net5589),
    .Y(_05124_),
    .A2(_06798_));
 sg13g2_a21o_1 _20902_ (.A2(net5277),
    .A1(net5594),
    .B1(_05124_),
    .X(_01494_));
 sg13g2_xnor2_1 _20903_ (.Y(_05125_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[17] ),
    .B(_05118_));
 sg13g2_nand2_1 _20904_ (.Y(_05126_),
    .A(net4721),
    .B(_05125_));
 sg13g2_a221oi_1 _20905_ (.B2(_08371_),
    .C1(net4539),
    .B1(net4725),
    .A1(_06910_),
    .Y(_05127_),
    .A2(net4876));
 sg13g2_a221oi_1 _20906_ (.B2(_05127_),
    .C1(net5121),
    .B1(_05126_),
    .A1(_08375_),
    .Y(_05128_),
    .A2(net4539));
 sg13g2_a221oi_1 _20907_ (.B2(_06799_),
    .C1(_05128_),
    .B1(net5117),
    .A1(_06611_),
    .Y(_01495_),
    .A2(net5274));
 sg13g2_nor4_1 _20908_ (.A(_06909_),
    .B(_06911_),
    .C(_06912_),
    .D(_05109_),
    .Y(_05129_));
 sg13g2_a21oi_1 _20909_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[17] ),
    .A2(_05118_),
    .Y(_05130_),
    .B1(net3948));
 sg13g2_or2_1 _20910_ (.X(_05131_),
    .B(_05130_),
    .A(_05129_));
 sg13g2_nor2_1 _20911_ (.A(net2489),
    .B(_04956_),
    .Y(_05132_));
 sg13g2_a221oi_1 _20912_ (.B2(_05131_),
    .C1(_05132_),
    .B1(net4721),
    .A1(_08520_),
    .Y(_05133_),
    .A2(_04968_));
 sg13g2_a21oi_1 _20913_ (.A1(_08523_),
    .A2(net4539),
    .Y(_05134_),
    .B1(net5121));
 sg13g2_o21ai_1 _20914_ (.B1(_05134_),
    .Y(_05135_),
    .A1(net4539),
    .A2(_05133_));
 sg13g2_a22oi_1 _20915_ (.Y(_05136_),
    .B1(net5119),
    .B2(net5647),
    .A2(net5277),
    .A1(net6547));
 sg13g2_nand2_1 _20916_ (.Y(_01496_),
    .A(_05135_),
    .B(net6548));
 sg13g2_and4_1 _20917_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[17] ),
    .B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[18] ),
    .C(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[19] ),
    .D(_05118_),
    .X(_05137_));
 sg13g2_nor2_1 _20918_ (.A(_04984_),
    .B(_05137_),
    .Y(_05138_));
 sg13g2_o21ai_1 _20919_ (.B1(_05138_),
    .Y(_05139_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[19] ),
    .A2(_05129_));
 sg13g2_a221oi_1 _20920_ (.B2(_08381_),
    .C1(net4537),
    .B1(net4725),
    .A1(\fpga_top.cpu_top.csr_mepc_ex[19] ),
    .Y(_05140_),
    .A2(net4876));
 sg13g2_a22oi_1 _20921_ (.Y(_05141_),
    .B1(_05139_),
    .B2(_05140_),
    .A2(net4538),
    .A1(_08402_));
 sg13g2_nor2_2 _20922_ (.A(net5121),
    .B(_05141_),
    .Y(_05142_));
 sg13g2_a221oi_1 _20923_ (.B2(_06801_),
    .C1(_05142_),
    .B1(net5117),
    .A1(_06617_),
    .Y(_01497_),
    .A2(net5271));
 sg13g2_and2_1 _20924_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[20] ),
    .B(_05137_),
    .X(_05143_));
 sg13g2_o21ai_1 _20925_ (.B1(net4721),
    .Y(_05144_),
    .A1(net3886),
    .A2(_05137_));
 sg13g2_nand2_1 _20926_ (.Y(_05145_),
    .A(_08424_),
    .B(net4538));
 sg13g2_o21ai_1 _20927_ (.B1(net4500),
    .Y(_05146_),
    .A1(_08421_),
    .A2(net4723));
 sg13g2_a21oi_1 _20928_ (.A1(net2210),
    .A2(net4877),
    .Y(_05147_),
    .B1(_05146_));
 sg13g2_o21ai_1 _20929_ (.B1(_05147_),
    .Y(_05148_),
    .A1(_05143_),
    .A2(_05144_));
 sg13g2_a21oi_1 _20930_ (.A1(_05145_),
    .A2(_05148_),
    .Y(_05149_),
    .B1(net5121));
 sg13g2_a221oi_1 _20931_ (.B2(_06802_),
    .C1(_05149_),
    .B1(net5118),
    .A1(_06620_),
    .Y(_01498_),
    .A2(net5276));
 sg13g2_nand2_1 _20932_ (.Y(_05150_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ),
    .B(_05143_));
 sg13g2_o21ai_1 _20933_ (.B1(net4721),
    .Y(_05151_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ),
    .A2(_05143_));
 sg13g2_nand2b_1 _20934_ (.Y(_05152_),
    .B(_05150_),
    .A_N(_05151_));
 sg13g2_nor2_1 _20935_ (.A(_07861_),
    .B(net4723),
    .Y(_05153_));
 sg13g2_a21oi_1 _20936_ (.A1(net3749),
    .A2(net4877),
    .Y(_05154_),
    .B1(_05153_));
 sg13g2_nand3_1 _20937_ (.B(_05152_),
    .C(_05154_),
    .A(net4500),
    .Y(_05155_));
 sg13g2_a21oi_1 _20938_ (.A1(_07864_),
    .A2(net4537),
    .Y(_05156_),
    .B1(net5118));
 sg13g2_a221oi_1 _20939_ (.B2(_05156_),
    .C1(net5275),
    .B1(_05155_),
    .A1(net5589),
    .Y(_05157_),
    .A2(net5645));
 sg13g2_a21oi_1 _20940_ (.A1(_06623_),
    .A2(net5276),
    .Y(_01499_),
    .B1(_05157_));
 sg13g2_nand3_1 _20941_ (.B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[22] ),
    .C(_05143_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ),
    .Y(_05158_));
 sg13g2_xor2_1 _20942_ (.B(_05150_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[22] ),
    .X(_05159_));
 sg13g2_or2_1 _20943_ (.X(_05160_),
    .B(net5043),
    .A(\fpga_top.cpu_top.csr_mepc_ex[22] ));
 sg13g2_o21ai_1 _20944_ (.B1(_05160_),
    .Y(_05161_),
    .A1(_07832_),
    .A2(net4723));
 sg13g2_a21oi_1 _20945_ (.A1(net4721),
    .A2(_05159_),
    .Y(_05162_),
    .B1(_05161_));
 sg13g2_a21oi_1 _20946_ (.A1(_07835_),
    .A2(_04970_),
    .Y(_05163_),
    .B1(net5121));
 sg13g2_o21ai_1 _20947_ (.B1(_05163_),
    .Y(_05164_),
    .A1(net4536),
    .A2(_05162_));
 sg13g2_a22oi_1 _20948_ (.Y(_05165_),
    .B1(net5118),
    .B2(net5643),
    .A2(net5275),
    .A1(net5592));
 sg13g2_nand2_1 _20949_ (.Y(_01500_),
    .A(_05164_),
    .B(_05165_));
 sg13g2_nand4_1 _20950_ (.B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[22] ),
    .C(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[23] ),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ),
    .Y(_05166_),
    .D(_05143_));
 sg13g2_xor2_1 _20951_ (.B(_05158_),
    .A(net6201),
    .X(_05167_));
 sg13g2_a221oi_1 _20952_ (.B2(_08455_),
    .C1(net4536),
    .B1(net4725),
    .A1(net2789),
    .Y(_05168_),
    .A2(net4877));
 sg13g2_o21ai_1 _20953_ (.B1(_05168_),
    .Y(_05169_),
    .A1(_04984_),
    .A2(_05167_));
 sg13g2_a21oi_1 _20954_ (.A1(_08472_),
    .A2(net4537),
    .Y(_05170_),
    .B1(net5118));
 sg13g2_a221oi_1 _20955_ (.B2(_05170_),
    .C1(net5275),
    .B1(_05169_),
    .A1(net6475),
    .Y(_05171_),
    .A2(net5642));
 sg13g2_a21oi_1 _20956_ (.A1(_06626_),
    .A2(net5275),
    .Y(_01501_),
    .B1(_05171_));
 sg13g2_or2_1 _20957_ (.X(_05172_),
    .B(_05166_),
    .A(_06917_));
 sg13g2_a21oi_1 _20958_ (.A1(_06917_),
    .A2(_05166_),
    .Y(_05173_),
    .B1(_04984_));
 sg13g2_o21ai_1 _20959_ (.B1(net4500),
    .Y(_05174_),
    .A1(_07901_),
    .A2(net4723));
 sg13g2_a221oi_1 _20960_ (.B2(_05173_),
    .C1(_05174_),
    .B1(_05172_),
    .A1(net2329),
    .Y(_05175_),
    .A2(net4877));
 sg13g2_a21oi_1 _20961_ (.A1(_07903_),
    .A2(net4538),
    .Y(_05176_),
    .B1(_05175_));
 sg13g2_nor2_1 _20962_ (.A(_04990_),
    .B(_05176_),
    .Y(_05177_));
 sg13g2_a221oi_1 _20963_ (.B2(_06805_),
    .C1(_05177_),
    .B1(net5118),
    .A1(_06629_),
    .Y(_01502_),
    .A2(net5276));
 sg13g2_nor2_2 _20964_ (.A(_06918_),
    .B(_05172_),
    .Y(_05178_));
 sg13g2_a21oi_1 _20965_ (.A1(_06918_),
    .A2(_05172_),
    .Y(_05179_),
    .B1(_04984_));
 sg13g2_nand2b_1 _20966_ (.Y(_05180_),
    .B(_05179_),
    .A_N(_05178_));
 sg13g2_nand2_1 _20967_ (.Y(_05181_),
    .A(_08495_),
    .B(net4561));
 sg13g2_a221oi_1 _20968_ (.B2(_05181_),
    .C1(net5276),
    .B1(net4725),
    .A1(net1996),
    .Y(_05182_),
    .A2(net4876));
 sg13g2_a22oi_1 _20969_ (.Y(_05183_),
    .B1(_05180_),
    .B2(_05182_),
    .A2(net4538),
    .A1(_08497_));
 sg13g2_nor2_1 _20970_ (.A(net5121),
    .B(_05183_),
    .Y(_05184_));
 sg13g2_a221oi_1 _20971_ (.B2(_06806_),
    .C1(_05184_),
    .B1(net5118),
    .A1(_06631_),
    .Y(_01503_),
    .A2(net5276));
 sg13g2_xnor2_1 _20972_ (.Y(_05185_),
    .A(net3916),
    .B(_05178_));
 sg13g2_a221oi_1 _20973_ (.B2(_08593_),
    .C1(net4536),
    .B1(net4725),
    .A1(net2312),
    .Y(_05186_),
    .A2(net4876));
 sg13g2_o21ai_1 _20974_ (.B1(_05186_),
    .Y(_05187_),
    .A1(_04984_),
    .A2(_05185_));
 sg13g2_a21oi_1 _20975_ (.A1(_08596_),
    .A2(net4536),
    .Y(_05188_),
    .B1(net5118));
 sg13g2_a221oi_1 _20976_ (.B2(_05188_),
    .C1(net5275),
    .B1(_05187_),
    .A1(net5589),
    .Y(_05189_),
    .A2(\fpga_top.cpu_start_adr[26] ));
 sg13g2_a21oi_1 _20977_ (.A1(_06634_),
    .A2(net5276),
    .Y(_01504_),
    .B1(_05189_));
 sg13g2_a21oi_1 _20978_ (.A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[26] ),
    .A2(_05178_),
    .Y(_05190_),
    .B1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[27] ));
 sg13g2_and3_1 _20979_ (.X(_05191_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[26] ),
    .B(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[27] ),
    .C(_05178_));
 sg13g2_o21ai_1 _20980_ (.B1(net4722),
    .Y(_05192_),
    .A1(_05190_),
    .A2(_05191_));
 sg13g2_or2_1 _20981_ (.X(_05193_),
    .B(net5043),
    .A(\fpga_top.cpu_top.csr_mepc_ex[27] ));
 sg13g2_o21ai_1 _20982_ (.B1(_05193_),
    .Y(_05194_),
    .A1(_08432_),
    .A2(net4723));
 sg13g2_nor2b_1 _20983_ (.A(_05194_),
    .B_N(_05192_),
    .Y(_05195_));
 sg13g2_a21oi_1 _20984_ (.A1(_08450_),
    .A2(_04970_),
    .Y(_05196_),
    .B1(net5121));
 sg13g2_o21ai_1 _20985_ (.B1(_05196_),
    .Y(_05197_),
    .A1(net4536),
    .A2(_05195_));
 sg13g2_a22oi_1 _20986_ (.Y(_05198_),
    .B1(net5118),
    .B2(net5641),
    .A2(net5276),
    .A1(net6569));
 sg13g2_nand2_1 _20987_ (.Y(_01505_),
    .A(_05197_),
    .B(_05198_));
 sg13g2_nand2_1 _20988_ (.Y(_05199_),
    .A(net5590),
    .B(net5275));
 sg13g2_nor2_1 _20989_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[28] ),
    .B(_05191_),
    .Y(_05200_));
 sg13g2_and2_1 _20990_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[28] ),
    .B(_05191_),
    .X(_05201_));
 sg13g2_o21ai_1 _20991_ (.B1(net4722),
    .Y(_05202_),
    .A1(_05200_),
    .A2(_05201_));
 sg13g2_nor2_1 _20992_ (.A(_08569_),
    .B(net4723),
    .Y(_05203_));
 sg13g2_nor2_1 _20993_ (.A(net2048),
    .B(_04956_),
    .Y(_05204_));
 sg13g2_nor3_1 _20994_ (.A(net4536),
    .B(_05203_),
    .C(_05204_),
    .Y(_05205_));
 sg13g2_a221oi_1 _20995_ (.B2(_05205_),
    .C1(net5589),
    .B1(_05202_),
    .A1(_08571_),
    .Y(_05206_),
    .A2(net4536));
 sg13g2_a21oi_2 _20996_ (.B1(_04989_),
    .Y(_05207_),
    .A2(net5278),
    .A1(net5638));
 sg13g2_o21ai_1 _20997_ (.B1(_05199_),
    .Y(_01506_),
    .A1(_05206_),
    .A2(_05207_));
 sg13g2_and2_1 _20998_ (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[29] ),
    .B(_05201_),
    .X(_05208_));
 sg13g2_xnor2_1 _20999_ (.Y(_05209_),
    .A(net6132),
    .B(_05201_));
 sg13g2_or2_1 _21000_ (.X(_05210_),
    .B(_04956_),
    .A(net1792));
 sg13g2_o21ai_1 _21001_ (.B1(_05210_),
    .Y(_05211_),
    .A1(_07752_),
    .A2(_04969_));
 sg13g2_a21oi_1 _21002_ (.A1(net4721),
    .A2(_05209_),
    .Y(_05212_),
    .B1(_05211_));
 sg13g2_a21oi_1 _21003_ (.A1(_07796_),
    .A2(_04970_),
    .Y(_05213_),
    .B1(net5121));
 sg13g2_o21ai_1 _21004_ (.B1(_05213_),
    .Y(_05214_),
    .A1(net4536),
    .A2(_05212_));
 sg13g2_a22oi_1 _21005_ (.Y(_05215_),
    .B1(net5119),
    .B2(net5637),
    .A2(net5275),
    .A1(net6565));
 sg13g2_nand2_1 _21006_ (.Y(_01507_),
    .A(_05214_),
    .B(_05215_));
 sg13g2_or2_1 _21007_ (.X(_05216_),
    .B(_05208_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[30] ));
 sg13g2_nand2_2 _21008_ (.Y(_05217_),
    .A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[30] ),
    .B(_05208_));
 sg13g2_a21o_1 _21009_ (.A2(_05217_),
    .A1(_05216_),
    .B1(_04984_),
    .X(_05218_));
 sg13g2_a221oi_1 _21010_ (.B2(_07676_),
    .C1(net4537),
    .B1(net4725),
    .A1(_06920_),
    .Y(_05219_),
    .A2(net4876));
 sg13g2_a21oi_1 _21011_ (.A1(_05218_),
    .A2(_05219_),
    .Y(_05220_),
    .B1(net5589));
 sg13g2_o21ai_1 _21012_ (.B1(_05220_),
    .Y(_05221_),
    .A1(_07746_),
    .A2(net4500));
 sg13g2_a21oi_1 _21013_ (.A1(net5587),
    .A2(_06810_),
    .Y(_05222_),
    .B1(net5272));
 sg13g2_a22oi_1 _21014_ (.Y(_05223_),
    .B1(_05221_),
    .B2(_05222_),
    .A2(net5271),
    .A1(net6479));
 sg13g2_inv_1 _21015_ (.Y(_01508_),
    .A(_05223_));
 sg13g2_nor2_1 _21016_ (.A(_06646_),
    .B(net5278),
    .Y(_05224_));
 sg13g2_xnor2_1 _21017_ (.Y(_05225_),
    .A(_06923_),
    .B(_05217_));
 sg13g2_nand2_1 _21018_ (.Y(_05226_),
    .A(net4721),
    .B(_05225_));
 sg13g2_a221oi_1 _21019_ (.B2(_07287_),
    .C1(net4539),
    .B1(net4725),
    .A1(_06922_),
    .Y(_05227_),
    .A2(net4876));
 sg13g2_a21oi_1 _21020_ (.A1(_05226_),
    .A2(_05227_),
    .Y(_05228_),
    .B1(net5119));
 sg13g2_o21ai_1 _21021_ (.B1(_05228_),
    .Y(_05229_),
    .A1(_07671_),
    .A2(net4500));
 sg13g2_a21oi_1 _21022_ (.A1(net5587),
    .A2(_06811_),
    .Y(_05230_),
    .B1(net5272));
 sg13g2_a21o_1 _21023_ (.A2(_05230_),
    .A1(_05229_),
    .B1(_05224_),
    .X(_01509_));
 sg13g2_nand2_1 _21024_ (.Y(_05231_),
    .A(\fpga_top.cpu_top.pc_stage.g_interrupt_latch ),
    .B(net5272));
 sg13g2_o21ai_1 _21025_ (.B1(_05231_),
    .Y(_01510_),
    .A1(net1376),
    .A2(_08916_));
 sg13g2_o21ai_1 _21026_ (.B1(net5272),
    .Y(_05232_),
    .A1(net6544),
    .A2(net5587));
 sg13g2_inv_1 _21027_ (.Y(_01511_),
    .A(_05232_));
 sg13g2_a22oi_1 _21028_ (.Y(_05233_),
    .B1(net5272),
    .B2(net3414),
    .A2(_06774_),
    .A1(\fpga_top.cpu_top.execution.csr_array.frc_cntr_val_leq ));
 sg13g2_inv_1 _21029_ (.Y(_01512_),
    .A(net3415));
 sg13g2_o21ai_1 _21030_ (.B1(net5427),
    .Y(_05234_),
    .A1(net1380),
    .A2(net6401));
 sg13g2_nor2_1 _21031_ (.A(net5097),
    .B(_05234_),
    .Y(_01513_));
 sg13g2_a21oi_1 _21032_ (.A1(net5572),
    .A2(_04921_),
    .Y(_05235_),
    .B1(net1843));
 sg13g2_nor2_1 _21033_ (.A(net5278),
    .B(net1844),
    .Y(_01514_));
 sg13g2_nand3_1 _21034_ (.B(_09663_),
    .C(_09666_),
    .A(_09661_),
    .Y(_05236_));
 sg13g2_or2_1 _21035_ (.X(_05237_),
    .B(_05236_),
    .A(_09659_));
 sg13g2_mux2_1 _21036_ (.A0(net4366),
    .A1(net2687),
    .S(net4125),
    .X(_01515_));
 sg13g2_mux2_1 _21037_ (.A0(net4358),
    .A1(net2261),
    .S(net4127),
    .X(_01516_));
 sg13g2_mux2_1 _21038_ (.A0(net4352),
    .A1(net2310),
    .S(net4126),
    .X(_01517_));
 sg13g2_mux2_1 _21039_ (.A0(net4347),
    .A1(net2940),
    .S(net4126),
    .X(_01518_));
 sg13g2_mux2_1 _21040_ (.A0(net4342),
    .A1(net2226),
    .S(net4127),
    .X(_01519_));
 sg13g2_mux2_1 _21041_ (.A0(net4197),
    .A1(net3592),
    .S(net4129),
    .X(_01520_));
 sg13g2_mux2_1 _21042_ (.A0(net4336),
    .A1(net3275),
    .S(net4126),
    .X(_01521_));
 sg13g2_mux2_1 _21043_ (.A0(net4333),
    .A1(net2692),
    .S(net4128),
    .X(_01522_));
 sg13g2_mux2_1 _21044_ (.A0(net4326),
    .A1(net3130),
    .S(net4127),
    .X(_01523_));
 sg13g2_mux2_1 _21045_ (.A0(net4323),
    .A1(net3332),
    .S(net4125),
    .X(_01524_));
 sg13g2_mux2_1 _21046_ (.A0(net4192),
    .A1(net3118),
    .S(net4128),
    .X(_01525_));
 sg13g2_mux2_1 _21047_ (.A0(net4188),
    .A1(net2375),
    .S(net4125),
    .X(_01526_));
 sg13g2_mux2_1 _21048_ (.A0(net4316),
    .A1(net2842),
    .S(net4128),
    .X(_01527_));
 sg13g2_mux2_1 _21049_ (.A0(net4310),
    .A1(net2435),
    .S(net4125),
    .X(_01528_));
 sg13g2_mux2_1 _21050_ (.A0(net4305),
    .A1(net3280),
    .S(net4125),
    .X(_01529_));
 sg13g2_mux2_1 _21051_ (.A0(net4298),
    .A1(net3154),
    .S(net4127),
    .X(_01530_));
 sg13g2_mux2_1 _21052_ (.A0(net4294),
    .A1(net3345),
    .S(net4129),
    .X(_01531_));
 sg13g2_mux2_1 _21053_ (.A0(net4289),
    .A1(net3050),
    .S(net4125),
    .X(_01532_));
 sg13g2_mux2_1 _21054_ (.A0(net4281),
    .A1(net3285),
    .S(net4128),
    .X(_01533_));
 sg13g2_mux2_1 _21055_ (.A0(net4278),
    .A1(net2694),
    .S(net4126),
    .X(_01534_));
 sg13g2_mux2_1 _21056_ (.A0(net4272),
    .A1(net3108),
    .S(net4127),
    .X(_01535_));
 sg13g2_mux2_1 _21057_ (.A0(net4266),
    .A1(net3131),
    .S(net4125),
    .X(_01536_));
 sg13g2_mux2_1 _21058_ (.A0(net4263),
    .A1(net2561),
    .S(net4127),
    .X(_01537_));
 sg13g2_mux2_1 _21059_ (.A0(net4257),
    .A1(net2712),
    .S(net4129),
    .X(_01538_));
 sg13g2_mux2_1 _21060_ (.A0(net4405),
    .A1(net2455),
    .S(net4128),
    .X(_01539_));
 sg13g2_mux2_1 _21061_ (.A0(net4402),
    .A1(net2370),
    .S(net4127),
    .X(_01540_));
 sg13g2_mux2_1 _21062_ (.A0(net4395),
    .A1(net2584),
    .S(net4126),
    .X(_01541_));
 sg13g2_mux2_1 _21063_ (.A0(net4391),
    .A1(net2470),
    .S(net4126),
    .X(_01542_));
 sg13g2_mux2_1 _21064_ (.A0(net4383),
    .A1(net3400),
    .S(net4125),
    .X(_01543_));
 sg13g2_mux2_1 _21065_ (.A0(net4379),
    .A1(net3341),
    .S(net4128),
    .X(_01544_));
 sg13g2_mux2_1 _21066_ (.A0(net4375),
    .A1(net3042),
    .S(net4127),
    .X(_01545_));
 sg13g2_mux2_1 _21067_ (.A0(net4369),
    .A1(net3313),
    .S(net4128),
    .X(_01546_));
 sg13g2_or2_1 _21068_ (.X(_05238_),
    .B(_05236_),
    .A(_09805_));
 sg13g2_mux2_1 _21069_ (.A0(net4366),
    .A1(net3579),
    .S(net4120),
    .X(_01547_));
 sg13g2_mux2_1 _21070_ (.A0(net4359),
    .A1(net3476),
    .S(net4122),
    .X(_01548_));
 sg13g2_mux2_1 _21071_ (.A0(net4352),
    .A1(net2987),
    .S(net4121),
    .X(_01549_));
 sg13g2_mux2_1 _21072_ (.A0(net4348),
    .A1(net2372),
    .S(net4121),
    .X(_01550_));
 sg13g2_mux2_1 _21073_ (.A0(net4342),
    .A1(net2713),
    .S(net4122),
    .X(_01551_));
 sg13g2_mux2_1 _21074_ (.A0(net4197),
    .A1(net2884),
    .S(net4124),
    .X(_01552_));
 sg13g2_mux2_1 _21075_ (.A0(net4336),
    .A1(net3024),
    .S(net4121),
    .X(_01553_));
 sg13g2_mux2_1 _21076_ (.A0(net4333),
    .A1(net2671),
    .S(net4123),
    .X(_01554_));
 sg13g2_mux2_1 _21077_ (.A0(net4326),
    .A1(net3106),
    .S(net4122),
    .X(_01555_));
 sg13g2_mux2_1 _21078_ (.A0(net4323),
    .A1(net2992),
    .S(net4120),
    .X(_01556_));
 sg13g2_mux2_1 _21079_ (.A0(net4192),
    .A1(net3084),
    .S(net4123),
    .X(_01557_));
 sg13g2_mux2_1 _21080_ (.A0(net4188),
    .A1(net2276),
    .S(net4120),
    .X(_01558_));
 sg13g2_mux2_1 _21081_ (.A0(net4316),
    .A1(net3064),
    .S(net4123),
    .X(_01559_));
 sg13g2_mux2_1 _21082_ (.A0(net4310),
    .A1(net3256),
    .S(net4120),
    .X(_01560_));
 sg13g2_mux2_1 _21083_ (.A0(net4305),
    .A1(net2603),
    .S(net4120),
    .X(_01561_));
 sg13g2_mux2_1 _21084_ (.A0(net4298),
    .A1(net3330),
    .S(net4122),
    .X(_01562_));
 sg13g2_mux2_1 _21085_ (.A0(net4294),
    .A1(net3626),
    .S(net4124),
    .X(_01563_));
 sg13g2_mux2_1 _21086_ (.A0(net4289),
    .A1(net3514),
    .S(net4120),
    .X(_01564_));
 sg13g2_mux2_1 _21087_ (.A0(net4281),
    .A1(net2469),
    .S(net4123),
    .X(_01565_));
 sg13g2_mux2_1 _21088_ (.A0(net4278),
    .A1(net3274),
    .S(net4121),
    .X(_01566_));
 sg13g2_mux2_1 _21089_ (.A0(net4272),
    .A1(net3208),
    .S(net4122),
    .X(_01567_));
 sg13g2_mux2_1 _21090_ (.A0(net4267),
    .A1(net3543),
    .S(net4120),
    .X(_01568_));
 sg13g2_mux2_1 _21091_ (.A0(net4263),
    .A1(net3314),
    .S(net4122),
    .X(_01569_));
 sg13g2_mux2_1 _21092_ (.A0(net4257),
    .A1(net2487),
    .S(net4124),
    .X(_01570_));
 sg13g2_mux2_1 _21093_ (.A0(net4405),
    .A1(net2386),
    .S(net4123),
    .X(_01571_));
 sg13g2_mux2_1 _21094_ (.A0(net4402),
    .A1(net3608),
    .S(net4122),
    .X(_01572_));
 sg13g2_mux2_1 _21095_ (.A0(net4395),
    .A1(net2283),
    .S(net4121),
    .X(_01573_));
 sg13g2_mux2_1 _21096_ (.A0(net4391),
    .A1(net2855),
    .S(net4121),
    .X(_01574_));
 sg13g2_mux2_1 _21097_ (.A0(net4383),
    .A1(net3317),
    .S(net4120),
    .X(_01575_));
 sg13g2_mux2_1 _21098_ (.A0(net4379),
    .A1(net3184),
    .S(net4123),
    .X(_01576_));
 sg13g2_mux2_1 _21099_ (.A0(net4375),
    .A1(net3381),
    .S(net4122),
    .X(_01577_));
 sg13g2_mux2_1 _21100_ (.A0(net4369),
    .A1(net3384),
    .S(net4123),
    .X(_01578_));
 sg13g2_mux2_1 _21101_ (.A0(net3583),
    .A1(_03861_),
    .S(net5054),
    .X(_01579_));
 sg13g2_mux2_1 _21102_ (.A0(net3723),
    .A1(_03879_),
    .S(net5051),
    .X(_01580_));
 sg13g2_nor2_1 _21103_ (.A(net5138),
    .B(_03895_),
    .Y(_05239_));
 sg13g2_a21oi_1 _21104_ (.A1(_06583_),
    .A2(net5138),
    .Y(_01581_),
    .B1(_05239_));
 sg13g2_nand2_1 _21105_ (.Y(_05240_),
    .A(net1455),
    .B(net5138));
 sg13g2_o21ai_1 _21106_ (.B1(_05240_),
    .Y(_01582_),
    .A1(net5138),
    .A2(_03943_));
 sg13g2_mux2_1 _21107_ (.A0(net3155),
    .A1(_04528_),
    .S(net5051),
    .X(_01583_));
 sg13g2_nor2_1 _21108_ (.A(net5138),
    .B(_04540_),
    .Y(_05241_));
 sg13g2_a21oi_1 _21109_ (.A1(_06585_),
    .A2(net5138),
    .Y(_01584_),
    .B1(_05241_));
 sg13g2_nor2_1 _21110_ (.A(net1937),
    .B(net5051),
    .Y(_05242_));
 sg13g2_a21oi_1 _21111_ (.A1(net5051),
    .A2(_03956_),
    .Y(_01585_),
    .B1(_05242_));
 sg13g2_mux2_1 _21112_ (.A0(net2752),
    .A1(_03969_),
    .S(net5051),
    .X(_01586_));
 sg13g2_mux2_1 _21113_ (.A0(net2793),
    .A1(_03981_),
    .S(net5051),
    .X(_01587_));
 sg13g2_nor2_1 _21114_ (.A(net1716),
    .B(net5053),
    .Y(_05243_));
 sg13g2_a21oi_1 _21115_ (.A1(net5053),
    .A2(_03995_),
    .Y(_01588_),
    .B1(_05243_));
 sg13g2_nor2_1 _21116_ (.A(net1859),
    .B(net5052),
    .Y(_05244_));
 sg13g2_a21oi_1 _21117_ (.A1(net5052),
    .A2(_04005_),
    .Y(_01589_),
    .B1(_05244_));
 sg13g2_nor2_1 _21118_ (.A(net1639),
    .B(net5051),
    .Y(_05245_));
 sg13g2_a21oi_1 _21119_ (.A1(net5051),
    .A2(_04019_),
    .Y(_01590_),
    .B1(_05245_));
 sg13g2_nor2_1 _21120_ (.A(net1794),
    .B(net5054),
    .Y(_05246_));
 sg13g2_a21oi_1 _21121_ (.A1(net5054),
    .A2(_04033_),
    .Y(_01591_),
    .B1(_05246_));
 sg13g2_nor2_1 _21122_ (.A(net1661),
    .B(net5052),
    .Y(_05247_));
 sg13g2_a21oi_1 _21123_ (.A1(net5052),
    .A2(_04044_),
    .Y(_01592_),
    .B1(_05247_));
 sg13g2_nor2_1 _21124_ (.A(net1646),
    .B(net5052),
    .Y(_05248_));
 sg13g2_a21oi_1 _21125_ (.A1(net5052),
    .A2(_04058_),
    .Y(_01593_),
    .B1(_05248_));
 sg13g2_nor2_1 _21126_ (.A(net1651),
    .B(net5052),
    .Y(_05249_));
 sg13g2_a21oi_1 _21127_ (.A1(net5052),
    .A2(_04067_),
    .Y(_01594_),
    .B1(_05249_));
 sg13g2_nor2_1 _21128_ (.A(net5145),
    .B(_04079_),
    .Y(_05250_));
 sg13g2_a21oi_1 _21129_ (.A1(_06607_),
    .A2(net5145),
    .Y(_01595_),
    .B1(_05250_));
 sg13g2_mux2_1 _21130_ (.A0(net3438),
    .A1(_04089_),
    .S(net5063),
    .X(_01596_));
 sg13g2_nor2_1 _21131_ (.A(net5145),
    .B(_04097_),
    .Y(_05251_));
 sg13g2_a21oi_1 _21132_ (.A1(_06613_),
    .A2(net5145),
    .Y(_01597_),
    .B1(_05251_));
 sg13g2_nor2_1 _21133_ (.A(net1914),
    .B(net5062),
    .Y(_05252_));
 sg13g2_a21oi_1 _21134_ (.A1(net5062),
    .A2(_04107_),
    .Y(_01598_),
    .B1(_05252_));
 sg13g2_nor2_1 _21135_ (.A(net1832),
    .B(net5061),
    .Y(_05253_));
 sg13g2_a21oi_1 _21136_ (.A1(net5062),
    .A2(_04120_),
    .Y(_01599_),
    .B1(_05253_));
 sg13g2_nor2_1 _21137_ (.A(net2040),
    .B(net5062),
    .Y(_05254_));
 sg13g2_a21oi_1 _21138_ (.A1(net5062),
    .A2(_04130_),
    .Y(_01600_),
    .B1(_05254_));
 sg13g2_nor2_1 _21139_ (.A(net1742),
    .B(net5061),
    .Y(_05255_));
 sg13g2_a21oi_1 _21140_ (.A1(net5062),
    .A2(_04142_),
    .Y(_01601_),
    .B1(_05255_));
 sg13g2_nor2_1 _21141_ (.A(net1768),
    .B(net5061),
    .Y(_05256_));
 sg13g2_a21oi_1 _21142_ (.A1(net5061),
    .A2(_04152_),
    .Y(_01602_),
    .B1(_05256_));
 sg13g2_nor2_1 _21143_ (.A(net1867),
    .B(net5063),
    .Y(_05257_));
 sg13g2_a21oi_1 _21144_ (.A1(net5063),
    .A2(_04164_),
    .Y(_01603_),
    .B1(_05257_));
 sg13g2_mux2_1 _21145_ (.A0(net2705),
    .A1(_04174_),
    .S(net5063),
    .X(_01604_));
 sg13g2_nor2_1 _21146_ (.A(net1717),
    .B(net5061),
    .Y(_05258_));
 sg13g2_a21oi_1 _21147_ (.A1(net5061),
    .A2(_04184_),
    .Y(_01605_),
    .B1(_05258_));
 sg13g2_mux2_1 _21148_ (.A0(net2970),
    .A1(_04195_),
    .S(net5061),
    .X(_01606_));
 sg13g2_nor2_1 _21149_ (.A(net1941),
    .B(net5062),
    .Y(_05259_));
 sg13g2_a21oi_1 _21150_ (.A1(net5062),
    .A2(_04208_),
    .Y(_01607_),
    .B1(_05259_));
 sg13g2_nor2_1 _21151_ (.A(net1680),
    .B(net5064),
    .Y(_05260_));
 sg13g2_a21oi_1 _21152_ (.A1(net5061),
    .A2(_04217_),
    .Y(_01608_),
    .B1(_05260_));
 sg13g2_nor2_1 _21153_ (.A(net2032),
    .B(net5063),
    .Y(_05261_));
 sg13g2_a21oi_1 _21154_ (.A1(net5063),
    .A2(_04229_),
    .Y(_01609_),
    .B1(_05261_));
 sg13g2_mux2_1 _21155_ (.A0(net3385),
    .A1(_04243_),
    .S(net5053),
    .X(_01610_));
 sg13g2_nand2_2 _21156_ (.Y(_05262_),
    .A(net1380),
    .B(net5097));
 sg13g2_nand2_1 _21157_ (.Y(_05263_),
    .A(net3864),
    .B(net4872));
 sg13g2_o21ai_1 _21158_ (.B1(_05263_),
    .Y(_01611_),
    .A1(_09808_),
    .A2(net4867));
 sg13g2_nand2_1 _21159_ (.Y(_05264_),
    .A(net3922),
    .B(net4872));
 sg13g2_o21ai_1 _21160_ (.B1(_05264_),
    .Y(_01612_),
    .A1(_09963_),
    .A2(net4868));
 sg13g2_nand2_1 _21161_ (.Y(_05265_),
    .A(net3572),
    .B(net4867));
 sg13g2_o21ai_1 _21162_ (.B1(_05265_),
    .Y(_01613_),
    .A1(_10028_),
    .A2(net4867));
 sg13g2_nand2_1 _21163_ (.Y(_05266_),
    .A(net6282),
    .B(net4871));
 sg13g2_o21ai_1 _21164_ (.B1(_05266_),
    .Y(_01614_),
    .A1(_10082_),
    .A2(net4870));
 sg13g2_mux2_1 _21165_ (.A0(_10126_),
    .A1(net6439),
    .S(net4871),
    .X(_01615_));
 sg13g2_nand2_1 _21166_ (.Y(_05267_),
    .A(net6314),
    .B(net4868));
 sg13g2_o21ai_1 _21167_ (.B1(_05267_),
    .Y(_01616_),
    .A1(net6392),
    .A2(net4868));
 sg13g2_nand2_1 _21168_ (.Y(_05268_),
    .A(net3806),
    .B(net4871));
 sg13g2_o21ai_1 _21169_ (.B1(_05268_),
    .Y(_01617_),
    .A1(_10202_),
    .A2(net4870));
 sg13g2_nand2_1 _21170_ (.Y(_05269_),
    .A(net4042),
    .B(net4869));
 sg13g2_o21ai_1 _21171_ (.B1(_05269_),
    .Y(_01618_),
    .A1(_09671_),
    .A2(net4874));
 sg13g2_nand2_1 _21172_ (.Y(_05270_),
    .A(net3395),
    .B(net4867));
 sg13g2_o21ai_1 _21173_ (.B1(_05270_),
    .Y(_01619_),
    .A1(_10272_),
    .A2(net4867));
 sg13g2_nand2_1 _21174_ (.Y(_05271_),
    .A(net6090),
    .B(net4872));
 sg13g2_o21ai_1 _21175_ (.B1(_05271_),
    .Y(_01620_),
    .A1(_10301_),
    .A2(net4868));
 sg13g2_nand2_1 _21176_ (.Y(_05272_),
    .A(net3938),
    .B(net4867));
 sg13g2_o21ai_1 _21177_ (.B1(_05272_),
    .Y(_01621_),
    .A1(_10324_),
    .A2(net4869));
 sg13g2_nand2_1 _21178_ (.Y(_05273_),
    .A(net3939),
    .B(net4867));
 sg13g2_o21ai_1 _21179_ (.B1(_05273_),
    .Y(_01622_),
    .A1(_10340_),
    .A2(net4869));
 sg13g2_nand2_1 _21180_ (.Y(_05274_),
    .A(net5584),
    .B(net4872));
 sg13g2_o21ai_1 _21181_ (.B1(_05274_),
    .Y(_01623_),
    .A1(_10354_),
    .A2(net4872));
 sg13g2_nand2_1 _21182_ (.Y(_05275_),
    .A(net5581),
    .B(net4872));
 sg13g2_o21ai_1 _21183_ (.B1(_05275_),
    .Y(_01624_),
    .A1(_10367_),
    .A2(net4872));
 sg13g2_nand2_1 _21184_ (.Y(_05276_),
    .A(net5577),
    .B(net4873));
 sg13g2_o21ai_1 _21185_ (.B1(_05276_),
    .Y(_01625_),
    .A1(_10381_),
    .A2(net4872));
 sg13g2_nand2_1 _21186_ (.Y(_05277_),
    .A(net6217),
    .B(net4871));
 sg13g2_o21ai_1 _21187_ (.B1(_05277_),
    .Y(_01626_),
    .A1(_09675_),
    .A2(net4871));
 sg13g2_nand2_1 _21188_ (.Y(_05278_),
    .A(net6093),
    .B(net4871));
 sg13g2_o21ai_1 _21189_ (.B1(_05278_),
    .Y(_01627_),
    .A1(_10405_),
    .A2(net4871));
 sg13g2_nand2_1 _21190_ (.Y(_05279_),
    .A(net6211),
    .B(net4873));
 sg13g2_o21ai_1 _21191_ (.B1(_05279_),
    .Y(_01628_),
    .A1(_10421_),
    .A2(net4873));
 sg13g2_mux2_1 _21192_ (.A0(_10436_),
    .A1(net6455),
    .S(net4873),
    .X(_01629_));
 sg13g2_mux2_1 _21193_ (.A0(_10450_),
    .A1(net6375),
    .S(net4871),
    .X(_01630_));
 sg13g2_nand2_1 _21194_ (.Y(_05280_),
    .A(net5573),
    .B(net4874));
 sg13g2_o21ai_1 _21195_ (.B1(_05280_),
    .Y(_01631_),
    .A1(_10463_),
    .A2(net4874));
 sg13g2_mux2_1 _21196_ (.A0(_10477_),
    .A1(net6520),
    .S(net4869),
    .X(_01632_));
 sg13g2_nand2_1 _21197_ (.Y(_05281_),
    .A(net6390),
    .B(net4874));
 sg13g2_o21ai_1 _21198_ (.B1(_05281_),
    .Y(_01633_),
    .A1(_10491_),
    .A2(net4874));
 sg13g2_mux2_1 _21199_ (.A0(_10505_),
    .A1(net6522),
    .S(net4874),
    .X(_01634_));
 sg13g2_mux2_1 _21200_ (.A0(_09678_),
    .A1(net6517),
    .S(net4874),
    .X(_01635_));
 sg13g2_mux2_1 _21201_ (.A0(_09711_),
    .A1(net6445),
    .S(net4870),
    .X(_01636_));
 sg13g2_mux2_1 _21202_ (.A0(_09732_),
    .A1(net5571),
    .S(net4874),
    .X(_01637_));
 sg13g2_mux2_1 _21203_ (.A0(_09746_),
    .A1(net6425),
    .S(net4873),
    .X(_01638_));
 sg13g2_mux2_1 _21204_ (.A0(_09757_),
    .A1(net6470),
    .S(net4867),
    .X(_01639_));
 sg13g2_mux2_1 _21205_ (.A0(_09769_),
    .A1(net5570),
    .S(net4868),
    .X(_01640_));
 sg13g2_nand2_1 _21206_ (.Y(_05282_),
    .A(net6406),
    .B(net4870));
 sg13g2_o21ai_1 _21207_ (.B1(_05282_),
    .Y(_01641_),
    .A1(_09779_),
    .A2(net4870));
 sg13g2_nand2_1 _21208_ (.Y(_05283_),
    .A(net5569),
    .B(net4870));
 sg13g2_o21ai_1 _21209_ (.B1(_05283_),
    .Y(_01642_),
    .A1(_09790_),
    .A2(net4870));
 sg13g2_a21oi_2 _21210_ (.B1(_03917_),
    .Y(_05284_),
    .A2(_09436_),
    .A1(net3894));
 sg13g2_nand2_1 _21211_ (.Y(_05285_),
    .A(net3695),
    .B(net5032));
 sg13g2_or2_1 _21212_ (.X(_05286_),
    .B(_03917_),
    .A(_09444_));
 sg13g2_o21ai_1 _21213_ (.B1(net3696),
    .Y(_01643_),
    .A1(_10642_),
    .A2(net5025));
 sg13g2_nand2_1 _21214_ (.Y(_05287_),
    .A(net3303),
    .B(net5027));
 sg13g2_o21ai_1 _21215_ (.B1(_05287_),
    .Y(_01644_),
    .A1(_10660_),
    .A2(net5022));
 sg13g2_nand2_1 _21216_ (.Y(_05288_),
    .A(net6218),
    .B(net5027));
 sg13g2_o21ai_1 _21217_ (.B1(_05288_),
    .Y(_01645_),
    .A1(_10678_),
    .A2(net5021));
 sg13g2_nand2_1 _21218_ (.Y(_05289_),
    .A(net3571),
    .B(net5027));
 sg13g2_o21ai_1 _21219_ (.B1(_05289_),
    .Y(_01646_),
    .A1(_10696_),
    .A2(net5022));
 sg13g2_nand2_1 _21220_ (.Y(_05290_),
    .A(net3633),
    .B(net5027));
 sg13g2_o21ai_1 _21221_ (.B1(_05290_),
    .Y(_01647_),
    .A1(_10714_),
    .A2(net5021));
 sg13g2_nand2_1 _21222_ (.Y(_05291_),
    .A(net2160),
    .B(net5028));
 sg13g2_o21ai_1 _21223_ (.B1(_05291_),
    .Y(_01648_),
    .A1(_10732_),
    .A2(net5021));
 sg13g2_nand2_1 _21224_ (.Y(_05292_),
    .A(net6336),
    .B(net5028));
 sg13g2_o21ai_1 _21225_ (.B1(_05292_),
    .Y(_01649_),
    .A1(_10750_),
    .A2(net5021));
 sg13g2_nand2_1 _21226_ (.Y(_05293_),
    .A(net6242),
    .B(net5027));
 sg13g2_o21ai_1 _21227_ (.B1(_05293_),
    .Y(_01650_),
    .A1(_10768_),
    .A2(net5021));
 sg13g2_nand2_1 _21228_ (.Y(_05294_),
    .A(net6285),
    .B(net5028));
 sg13g2_o21ai_1 _21229_ (.B1(_05294_),
    .Y(_01651_),
    .A1(_10784_),
    .A2(net5022));
 sg13g2_nand2_1 _21230_ (.Y(_05295_),
    .A(net6124),
    .B(net5027));
 sg13g2_o21ai_1 _21231_ (.B1(_05295_),
    .Y(_01652_),
    .A1(_10802_),
    .A2(net5021));
 sg13g2_nand2_1 _21232_ (.Y(_05296_),
    .A(net2938),
    .B(net5027));
 sg13g2_o21ai_1 _21233_ (.B1(_05296_),
    .Y(_01653_),
    .A1(_10820_),
    .A2(net5021));
 sg13g2_nand2_1 _21234_ (.Y(_05297_),
    .A(net6293),
    .B(net5029));
 sg13g2_o21ai_1 _21235_ (.B1(_05297_),
    .Y(_01654_),
    .A1(_10838_),
    .A2(net5022));
 sg13g2_nand2_1 _21236_ (.Y(_05298_),
    .A(net6363),
    .B(net5029));
 sg13g2_o21ai_1 _21237_ (.B1(_05298_),
    .Y(_01655_),
    .A1(_10856_),
    .A2(net5026));
 sg13g2_nand2_1 _21238_ (.Y(_05299_),
    .A(net6345),
    .B(net5029));
 sg13g2_o21ai_1 _21239_ (.B1(_05299_),
    .Y(_01656_),
    .A1(_10874_),
    .A2(net5026));
 sg13g2_nand2_1 _21240_ (.Y(_05300_),
    .A(net6423),
    .B(net5030));
 sg13g2_o21ai_1 _21241_ (.B1(_05300_),
    .Y(_01657_),
    .A1(_10892_),
    .A2(net5023));
 sg13g2_nand2_1 _21242_ (.Y(_05301_),
    .A(net3505),
    .B(net5029));
 sg13g2_o21ai_1 _21243_ (.B1(_05301_),
    .Y(_01658_),
    .A1(_10910_),
    .A2(net5022));
 sg13g2_nand2_1 _21244_ (.Y(_05302_),
    .A(net6125),
    .B(net5029));
 sg13g2_o21ai_1 _21245_ (.B1(_05302_),
    .Y(_01659_),
    .A1(_10928_),
    .A2(net5022));
 sg13g2_nand2_1 _21246_ (.Y(_05303_),
    .A(net6276),
    .B(net5031));
 sg13g2_o21ai_1 _21247_ (.B1(_05303_),
    .Y(_01660_),
    .A1(_10944_),
    .A2(net5024));
 sg13g2_nand2_1 _21248_ (.Y(_05304_),
    .A(net6337),
    .B(net5032));
 sg13g2_o21ai_1 _21249_ (.B1(_05304_),
    .Y(_01661_),
    .A1(_10962_),
    .A2(net5025));
 sg13g2_nand2_1 _21250_ (.Y(_05305_),
    .A(net6156),
    .B(net5030));
 sg13g2_o21ai_1 _21251_ (.B1(_05305_),
    .Y(_01662_),
    .A1(_10980_),
    .A2(net5023));
 sg13g2_nand2_1 _21252_ (.Y(_05306_),
    .A(net4038),
    .B(net5030));
 sg13g2_o21ai_1 _21253_ (.B1(_05306_),
    .Y(_01663_),
    .A1(_10998_),
    .A2(net5023));
 sg13g2_nand2_1 _21254_ (.Y(_05307_),
    .A(net6431),
    .B(net5030));
 sg13g2_o21ai_1 _21255_ (.B1(_05307_),
    .Y(_01664_),
    .A1(_02553_),
    .A2(net5023));
 sg13g2_nand2_1 _21256_ (.Y(_05308_),
    .A(net6204),
    .B(net5030));
 sg13g2_o21ai_1 _21257_ (.B1(_05308_),
    .Y(_01665_),
    .A1(_02571_),
    .A2(net5023));
 sg13g2_nand2_1 _21258_ (.Y(_05309_),
    .A(net6352),
    .B(net5031));
 sg13g2_o21ai_1 _21259_ (.B1(_05309_),
    .Y(_01666_),
    .A1(_02589_),
    .A2(net5024));
 sg13g2_nand2_1 _21260_ (.Y(_05310_),
    .A(net6393),
    .B(net5031));
 sg13g2_o21ai_1 _21261_ (.B1(_05310_),
    .Y(_01667_),
    .A1(_02607_),
    .A2(net5024));
 sg13g2_nand2_1 _21262_ (.Y(_05311_),
    .A(net6376),
    .B(net5031));
 sg13g2_o21ai_1 _21263_ (.B1(_05311_),
    .Y(_01668_),
    .A1(_02623_),
    .A2(net5024));
 sg13g2_nand2_1 _21264_ (.Y(_05312_),
    .A(net6270),
    .B(net5027));
 sg13g2_o21ai_1 _21265_ (.B1(_05312_),
    .Y(_01669_),
    .A1(_02641_),
    .A2(net5021));
 sg13g2_nand2_1 _21266_ (.Y(_05313_),
    .A(net6422),
    .B(net5030));
 sg13g2_o21ai_1 _21267_ (.B1(_05313_),
    .Y(_01670_),
    .A1(_02659_),
    .A2(net5023));
 sg13g2_nand2_1 _21268_ (.Y(_05314_),
    .A(net4073),
    .B(net5030));
 sg13g2_o21ai_1 _21269_ (.B1(_05314_),
    .Y(_01671_),
    .A1(_02677_),
    .A2(net5023));
 sg13g2_nand2_1 _21270_ (.Y(_05315_),
    .A(net6326),
    .B(net5032));
 sg13g2_o21ai_1 _21271_ (.B1(_05315_),
    .Y(_01672_),
    .A1(_02695_),
    .A2(net5025));
 sg13g2_nand2_1 _21272_ (.Y(_05316_),
    .A(net6457),
    .B(net5030));
 sg13g2_o21ai_1 _21273_ (.B1(_05316_),
    .Y(_01673_),
    .A1(_02713_),
    .A2(net5023));
 sg13g2_nand2_1 _21274_ (.Y(_05317_),
    .A(net6269),
    .B(net5029));
 sg13g2_o21ai_1 _21275_ (.B1(_05317_),
    .Y(_01674_),
    .A1(_02731_),
    .A2(net5022));
 sg13g2_a21oi_1 _21276_ (.A1(_06563_),
    .A2(_04921_),
    .Y(_05318_),
    .B1(net1938));
 sg13g2_nor2_1 _21277_ (.A(net5278),
    .B(net1939),
    .Y(_01675_));
 sg13g2_nand2_1 _21278_ (.Y(_05319_),
    .A(_09667_),
    .B(_09802_));
 sg13g2_or2_1 _21279_ (.X(_05320_),
    .B(_05319_),
    .A(_09805_));
 sg13g2_mux2_1 _21280_ (.A0(net4365),
    .A1(net2407),
    .S(net4115),
    .X(_01676_));
 sg13g2_mux2_1 _21281_ (.A0(net4359),
    .A1(net2982),
    .S(net4117),
    .X(_01677_));
 sg13g2_mux2_1 _21282_ (.A0(net4353),
    .A1(net3128),
    .S(net4116),
    .X(_01678_));
 sg13g2_mux2_1 _21283_ (.A0(net4345),
    .A1(net2613),
    .S(net4115),
    .X(_01679_));
 sg13g2_mux2_1 _21284_ (.A0(net4341),
    .A1(net2481),
    .S(net4117),
    .X(_01680_));
 sg13g2_mux2_1 _21285_ (.A0(net4198),
    .A1(net3418),
    .S(net4117),
    .X(_01681_));
 sg13g2_mux2_1 _21286_ (.A0(net4338),
    .A1(net3392),
    .S(net4115),
    .X(_01682_));
 sg13g2_mux2_1 _21287_ (.A0(net4333),
    .A1(net2927),
    .S(net4118),
    .X(_01683_));
 sg13g2_mux2_1 _21288_ (.A0(net4327),
    .A1(net2688),
    .S(net4119),
    .X(_01684_));
 sg13g2_mux2_1 _21289_ (.A0(net4319),
    .A1(net3200),
    .S(net4116),
    .X(_01685_));
 sg13g2_mux2_1 _21290_ (.A0(net4192),
    .A1(net3613),
    .S(net4118),
    .X(_01686_));
 sg13g2_mux2_1 _21291_ (.A0(net4187),
    .A1(net2498),
    .S(net4116),
    .X(_01687_));
 sg13g2_mux2_1 _21292_ (.A0(net4315),
    .A1(net2539),
    .S(net4118),
    .X(_01688_));
 sg13g2_mux2_1 _21293_ (.A0(net4310),
    .A1(net2747),
    .S(net4116),
    .X(_01689_));
 sg13g2_mux2_1 _21294_ (.A0(net4301),
    .A1(net3559),
    .S(net4115),
    .X(_01690_));
 sg13g2_mux2_1 _21295_ (.A0(net4298),
    .A1(net3464),
    .S(net4119),
    .X(_01691_));
 sg13g2_mux2_1 _21296_ (.A0(net4295),
    .A1(net3565),
    .S(net4118),
    .X(_01692_));
 sg13g2_mux2_1 _21297_ (.A0(net4287),
    .A1(net2511),
    .S(net4115),
    .X(_01693_));
 sg13g2_mux2_1 _21298_ (.A0(net4282),
    .A1(net3515),
    .S(net4118),
    .X(_01694_));
 sg13g2_mux2_1 _21299_ (.A0(net4277),
    .A1(net3428),
    .S(net4115),
    .X(_01695_));
 sg13g2_mux2_1 _21300_ (.A0(net4271),
    .A1(net3110),
    .S(net4117),
    .X(_01696_));
 sg13g2_mux2_1 _21301_ (.A0(net4266),
    .A1(net2517),
    .S(net4115),
    .X(_01697_));
 sg13g2_mux2_1 _21302_ (.A0(net4262),
    .A1(net2837),
    .S(net4117),
    .X(_01698_));
 sg13g2_mux2_1 _21303_ (.A0(net4258),
    .A1(net2371),
    .S(net4118),
    .X(_01699_));
 sg13g2_mux2_1 _21304_ (.A0(net4406),
    .A1(net2624),
    .S(net4118),
    .X(_01700_));
 sg13g2_mux2_1 _21305_ (.A0(net4401),
    .A1(net3248),
    .S(net4117),
    .X(_01701_));
 sg13g2_mux2_1 _21306_ (.A0(net4396),
    .A1(net2997),
    .S(net4116),
    .X(_01702_));
 sg13g2_mux2_1 _21307_ (.A0(net4390),
    .A1(net2277),
    .S(net4115),
    .X(_01703_));
 sg13g2_mux2_1 _21308_ (.A0(net4382),
    .A1(net2786),
    .S(net4116),
    .X(_01704_));
 sg13g2_mux2_1 _21309_ (.A0(net4380),
    .A1(net3539),
    .S(net4118),
    .X(_01705_));
 sg13g2_mux2_1 _21310_ (.A0(net4375),
    .A1(net2867),
    .S(net4117),
    .X(_01706_));
 sg13g2_mux2_1 _21311_ (.A0(net4369),
    .A1(net2693),
    .S(net4117),
    .X(_01707_));
 sg13g2_or2_1 _21312_ (.X(_05321_),
    .B(_05319_),
    .A(_03169_));
 sg13g2_mux2_1 _21313_ (.A0(net4364),
    .A1(net2543),
    .S(net4110),
    .X(_01708_));
 sg13g2_mux2_1 _21314_ (.A0(net4359),
    .A1(net3410),
    .S(net4112),
    .X(_01709_));
 sg13g2_mux2_1 _21315_ (.A0(net4353),
    .A1(net3051),
    .S(net4111),
    .X(_01710_));
 sg13g2_mux2_1 _21316_ (.A0(net4345),
    .A1(net3101),
    .S(net4110),
    .X(_01711_));
 sg13g2_mux2_1 _21317_ (.A0(net4341),
    .A1(net3191),
    .S(net4112),
    .X(_01712_));
 sg13g2_mux2_1 _21318_ (.A0(net4198),
    .A1(net2964),
    .S(net4112),
    .X(_01713_));
 sg13g2_mux2_1 _21319_ (.A0(net4338),
    .A1(net2814),
    .S(net4110),
    .X(_01714_));
 sg13g2_mux2_1 _21320_ (.A0(net4333),
    .A1(net3566),
    .S(net4113),
    .X(_01715_));
 sg13g2_mux2_1 _21321_ (.A0(net4327),
    .A1(net3518),
    .S(net4114),
    .X(_01716_));
 sg13g2_mux2_1 _21322_ (.A0(net4319),
    .A1(net3662),
    .S(net4111),
    .X(_01717_));
 sg13g2_mux2_1 _21323_ (.A0(net4192),
    .A1(net2499),
    .S(net4113),
    .X(_01718_));
 sg13g2_mux2_1 _21324_ (.A0(net4187),
    .A1(net2265),
    .S(net4111),
    .X(_01719_));
 sg13g2_mux2_1 _21325_ (.A0(net4316),
    .A1(net2766),
    .S(net4113),
    .X(_01720_));
 sg13g2_mux2_1 _21326_ (.A0(_10379_),
    .A1(net2392),
    .S(net4111),
    .X(_01721_));
 sg13g2_mux2_1 _21327_ (.A0(net4301),
    .A1(net3637),
    .S(net4110),
    .X(_01722_));
 sg13g2_mux2_1 _21328_ (.A0(net4300),
    .A1(net3393),
    .S(net4114),
    .X(_01723_));
 sg13g2_mux2_1 _21329_ (.A0(net4295),
    .A1(net3140),
    .S(net4113),
    .X(_01724_));
 sg13g2_mux2_1 _21330_ (.A0(net4287),
    .A1(net3259),
    .S(net4110),
    .X(_01725_));
 sg13g2_mux2_1 _21331_ (.A0(net4282),
    .A1(net3533),
    .S(net4113),
    .X(_01726_));
 sg13g2_mux2_1 _21332_ (.A0(net4277),
    .A1(net2652),
    .S(net4110),
    .X(_01727_));
 sg13g2_mux2_1 _21333_ (.A0(net4271),
    .A1(net2751),
    .S(net4112),
    .X(_01728_));
 sg13g2_mux2_1 _21334_ (.A0(net4266),
    .A1(net3137),
    .S(net4110),
    .X(_01729_));
 sg13g2_mux2_1 _21335_ (.A0(net4262),
    .A1(net2390),
    .S(net4112),
    .X(_01730_));
 sg13g2_mux2_1 _21336_ (.A0(net4258),
    .A1(net2659),
    .S(net4113),
    .X(_01731_));
 sg13g2_mux2_1 _21337_ (.A0(net4406),
    .A1(net2641),
    .S(net4113),
    .X(_01732_));
 sg13g2_mux2_1 _21338_ (.A0(net4401),
    .A1(net3422),
    .S(net4112),
    .X(_01733_));
 sg13g2_mux2_1 _21339_ (.A0(net4396),
    .A1(net2462),
    .S(net4111),
    .X(_01734_));
 sg13g2_mux2_1 _21340_ (.A0(net4390),
    .A1(net2529),
    .S(net4110),
    .X(_01735_));
 sg13g2_mux2_1 _21341_ (.A0(net4382),
    .A1(net3504),
    .S(net4111),
    .X(_01736_));
 sg13g2_mux2_1 _21342_ (.A0(net4380),
    .A1(net2784),
    .S(net4113),
    .X(_01737_));
 sg13g2_mux2_1 _21343_ (.A0(net4375),
    .A1(net2289),
    .S(net4112),
    .X(_01738_));
 sg13g2_mux2_1 _21344_ (.A0(net4370),
    .A1(net2589),
    .S(net4112),
    .X(_01739_));
 sg13g2_or2_1 _21345_ (.X(_05322_),
    .B(_05236_),
    .A(_02993_));
 sg13g2_mux2_1 _21346_ (.A0(net4366),
    .A1(net2437),
    .S(net4105),
    .X(_01740_));
 sg13g2_mux2_1 _21347_ (.A0(net4359),
    .A1(net2480),
    .S(net4107),
    .X(_01741_));
 sg13g2_mux2_1 _21348_ (.A0(net4352),
    .A1(net3020),
    .S(net4106),
    .X(_01742_));
 sg13g2_mux2_1 _21349_ (.A0(net4348),
    .A1(net2628),
    .S(net4106),
    .X(_01743_));
 sg13g2_mux2_1 _21350_ (.A0(net4342),
    .A1(net2684),
    .S(net4107),
    .X(_01744_));
 sg13g2_mux2_1 _21351_ (.A0(net4197),
    .A1(net2935),
    .S(net4109),
    .X(_01745_));
 sg13g2_mux2_1 _21352_ (.A0(net4336),
    .A1(net2263),
    .S(net4106),
    .X(_01746_));
 sg13g2_mux2_1 _21353_ (.A0(_10269_),
    .A1(net2660),
    .S(net4108),
    .X(_01747_));
 sg13g2_mux2_1 _21354_ (.A0(net4326),
    .A1(net2527),
    .S(net4107),
    .X(_01748_));
 sg13g2_mux2_1 _21355_ (.A0(net4323),
    .A1(net2990),
    .S(net4105),
    .X(_01749_));
 sg13g2_mux2_1 _21356_ (.A0(net4194),
    .A1(net3115),
    .S(net4108),
    .X(_01750_));
 sg13g2_mux2_1 _21357_ (.A0(net4188),
    .A1(net2290),
    .S(net4105),
    .X(_01751_));
 sg13g2_mux2_1 _21358_ (.A0(net4316),
    .A1(net2169),
    .S(net4108),
    .X(_01752_));
 sg13g2_mux2_1 _21359_ (.A0(net4310),
    .A1(net2807),
    .S(net4105),
    .X(_01753_));
 sg13g2_mux2_1 _21360_ (.A0(net4305),
    .A1(net3374),
    .S(net4105),
    .X(_01754_));
 sg13g2_mux2_1 _21361_ (.A0(net4298),
    .A1(net2439),
    .S(net4107),
    .X(_01755_));
 sg13g2_mux2_1 _21362_ (.A0(net4294),
    .A1(net2902),
    .S(net4109),
    .X(_01756_));
 sg13g2_mux2_1 _21363_ (.A0(net4289),
    .A1(net2909),
    .S(net4105),
    .X(_01757_));
 sg13g2_mux2_1 _21364_ (.A0(net4281),
    .A1(net2980),
    .S(net4108),
    .X(_01758_));
 sg13g2_mux2_1 _21365_ (.A0(net4278),
    .A1(net2330),
    .S(net4106),
    .X(_01759_));
 sg13g2_mux2_1 _21366_ (.A0(net4272),
    .A1(net2883),
    .S(net4107),
    .X(_01760_));
 sg13g2_mux2_1 _21367_ (.A0(net4267),
    .A1(net2932),
    .S(net4105),
    .X(_01761_));
 sg13g2_mux2_1 _21368_ (.A0(net4263),
    .A1(net2708),
    .S(net4107),
    .X(_01762_));
 sg13g2_mux2_1 _21369_ (.A0(net4257),
    .A1(net3263),
    .S(net4109),
    .X(_01763_));
 sg13g2_mux2_1 _21370_ (.A0(net4405),
    .A1(net2831),
    .S(net4108),
    .X(_01764_));
 sg13g2_mux2_1 _21371_ (.A0(net4402),
    .A1(net2846),
    .S(net4107),
    .X(_01765_));
 sg13g2_mux2_1 _21372_ (.A0(net4395),
    .A1(net2449),
    .S(net4106),
    .X(_01766_));
 sg13g2_mux2_1 _21373_ (.A0(net4391),
    .A1(net2532),
    .S(net4106),
    .X(_01767_));
 sg13g2_mux2_1 _21374_ (.A0(net4383),
    .A1(net2898),
    .S(net4105),
    .X(_01768_));
 sg13g2_mux2_1 _21375_ (.A0(net4379),
    .A1(net2316),
    .S(net4108),
    .X(_01769_));
 sg13g2_mux2_1 _21376_ (.A0(net4375),
    .A1(net2367),
    .S(net4107),
    .X(_01770_));
 sg13g2_mux2_1 _21377_ (.A0(net4369),
    .A1(net2685),
    .S(net4108),
    .X(_01771_));
 sg13g2_or2_1 _21378_ (.X(_05323_),
    .B(_03191_),
    .A(_02993_));
 sg13g2_mux2_1 _21379_ (.A0(net4365),
    .A1(net2841),
    .S(net4100),
    .X(_01772_));
 sg13g2_mux2_1 _21380_ (.A0(net4358),
    .A1(net2364),
    .S(net4102),
    .X(_01773_));
 sg13g2_mux2_1 _21381_ (.A0(net4352),
    .A1(net2978),
    .S(net4101),
    .X(_01774_));
 sg13g2_mux2_1 _21382_ (.A0(net4347),
    .A1(net3359),
    .S(net4101),
    .X(_01775_));
 sg13g2_mux2_1 _21383_ (.A0(net4342),
    .A1(net2860),
    .S(net4102),
    .X(_01776_));
 sg13g2_mux2_1 _21384_ (.A0(net4197),
    .A1(net2155),
    .S(net4104),
    .X(_01777_));
 sg13g2_mux2_1 _21385_ (.A0(net4337),
    .A1(net3630),
    .S(net4104),
    .X(_01778_));
 sg13g2_mux2_1 _21386_ (.A0(net4332),
    .A1(net2191),
    .S(net4103),
    .X(_01779_));
 sg13g2_mux2_1 _21387_ (.A0(net4327),
    .A1(net3023),
    .S(net4102),
    .X(_01780_));
 sg13g2_mux2_1 _21388_ (.A0(net4318),
    .A1(net2753),
    .S(net4100),
    .X(_01781_));
 sg13g2_mux2_1 _21389_ (.A0(net4192),
    .A1(net3228),
    .S(net4103),
    .X(_01782_));
 sg13g2_mux2_1 _21390_ (.A0(net4188),
    .A1(net3547),
    .S(net4100),
    .X(_01783_));
 sg13g2_mux2_1 _21391_ (.A0(net4315),
    .A1(net2680),
    .S(net4103),
    .X(_01784_));
 sg13g2_mux2_1 _21392_ (.A0(net4311),
    .A1(net2655),
    .S(net4100),
    .X(_01785_));
 sg13g2_mux2_1 _21393_ (.A0(net4305),
    .A1(net2691),
    .S(net4100),
    .X(_01786_));
 sg13g2_mux2_1 _21394_ (.A0(net4299),
    .A1(net2468),
    .S(net4102),
    .X(_01787_));
 sg13g2_mux2_1 _21395_ (.A0(net4293),
    .A1(net2506),
    .S(net4103),
    .X(_01788_));
 sg13g2_mux2_1 _21396_ (.A0(net4289),
    .A1(net2501),
    .S(net4100),
    .X(_01789_));
 sg13g2_mux2_1 _21397_ (.A0(net4281),
    .A1(net2348),
    .S(net4103),
    .X(_01790_));
 sg13g2_mux2_1 _21398_ (.A0(_10462_),
    .A1(net3059),
    .S(net4101),
    .X(_01791_));
 sg13g2_mux2_1 _21399_ (.A0(net4272),
    .A1(net3019),
    .S(net4102),
    .X(_01792_));
 sg13g2_mux2_1 _21400_ (.A0(net4267),
    .A1(net2207),
    .S(net4100),
    .X(_01793_));
 sg13g2_mux2_1 _21401_ (.A0(net4263),
    .A1(net3230),
    .S(net4102),
    .X(_01794_));
 sg13g2_mux2_1 _21402_ (.A0(net4257),
    .A1(net2764),
    .S(net4104),
    .X(_01795_));
 sg13g2_mux2_1 _21403_ (.A0(net4405),
    .A1(net3074),
    .S(net4103),
    .X(_01796_));
 sg13g2_mux2_1 _21404_ (.A0(net4402),
    .A1(net3167),
    .S(net4102),
    .X(_01797_));
 sg13g2_mux2_1 _21405_ (.A0(net4395),
    .A1(net2929),
    .S(net4101),
    .X(_01798_));
 sg13g2_mux2_1 _21406_ (.A0(net4391),
    .A1(net2545),
    .S(net4101),
    .X(_01799_));
 sg13g2_mux2_1 _21407_ (.A0(net4386),
    .A1(net3209),
    .S(net4100),
    .X(_01800_));
 sg13g2_mux2_1 _21408_ (.A0(net4379),
    .A1(net3037),
    .S(net4103),
    .X(_01801_));
 sg13g2_mux2_1 _21409_ (.A0(net4374),
    .A1(net2314),
    .S(net4102),
    .X(_01802_));
 sg13g2_mux2_1 _21410_ (.A0(net4369),
    .A1(net3235),
    .S(net4103),
    .X(_01803_));
 sg13g2_or2_1 _21411_ (.X(_05324_),
    .B(_03191_),
    .A(_09805_));
 sg13g2_mux2_1 _21412_ (.A0(net4365),
    .A1(net2595),
    .S(net4095),
    .X(_01804_));
 sg13g2_mux2_1 _21413_ (.A0(net4358),
    .A1(net3617),
    .S(net4097),
    .X(_01805_));
 sg13g2_mux2_1 _21414_ (.A0(net4352),
    .A1(net3523),
    .S(net4096),
    .X(_01806_));
 sg13g2_mux2_1 _21415_ (.A0(net4347),
    .A1(net3166),
    .S(net4096),
    .X(_01807_));
 sg13g2_mux2_1 _21416_ (.A0(net4342),
    .A1(net2924),
    .S(net4097),
    .X(_01808_));
 sg13g2_mux2_1 _21417_ (.A0(net4197),
    .A1(net3082),
    .S(net4099),
    .X(_01809_));
 sg13g2_mux2_1 _21418_ (.A0(net4337),
    .A1(net3324),
    .S(net4096),
    .X(_01810_));
 sg13g2_mux2_1 _21419_ (.A0(net4332),
    .A1(net2781),
    .S(net4098),
    .X(_01811_));
 sg13g2_mux2_1 _21420_ (.A0(net4327),
    .A1(net3654),
    .S(net4097),
    .X(_01812_));
 sg13g2_mux2_1 _21421_ (.A0(net4318),
    .A1(net3542),
    .S(net4095),
    .X(_01813_));
 sg13g2_mux2_1 _21422_ (.A0(net4193),
    .A1(net2711),
    .S(net4098),
    .X(_01814_));
 sg13g2_mux2_1 _21423_ (.A0(net4188),
    .A1(net3503),
    .S(net4095),
    .X(_01815_));
 sg13g2_mux2_1 _21424_ (.A0(net4315),
    .A1(net2714),
    .S(net4098),
    .X(_01816_));
 sg13g2_mux2_1 _21425_ (.A0(net4310),
    .A1(net3224),
    .S(net4095),
    .X(_01817_));
 sg13g2_mux2_1 _21426_ (.A0(net4306),
    .A1(net3245),
    .S(net4095),
    .X(_01818_));
 sg13g2_mux2_1 _21427_ (.A0(net4298),
    .A1(net2732),
    .S(net4097),
    .X(_01819_));
 sg13g2_mux2_1 _21428_ (.A0(net4294),
    .A1(net2486),
    .S(net4098),
    .X(_01820_));
 sg13g2_mux2_1 _21429_ (.A0(net4287),
    .A1(net2803),
    .S(net4095),
    .X(_01821_));
 sg13g2_mux2_1 _21430_ (.A0(net4281),
    .A1(net2981),
    .S(net4098),
    .X(_01822_));
 sg13g2_mux2_1 _21431_ (.A0(net4277),
    .A1(net3283),
    .S(net4096),
    .X(_01823_));
 sg13g2_mux2_1 _21432_ (.A0(net4272),
    .A1(net2700),
    .S(net4097),
    .X(_01824_));
 sg13g2_mux2_1 _21433_ (.A0(net4267),
    .A1(net3591),
    .S(net4095),
    .X(_01825_));
 sg13g2_mux2_1 _21434_ (.A0(net4263),
    .A1(net3205),
    .S(net4097),
    .X(_01826_));
 sg13g2_mux2_1 _21435_ (.A0(net4257),
    .A1(net2857),
    .S(net4099),
    .X(_01827_));
 sg13g2_mux2_1 _21436_ (.A0(net4405),
    .A1(net2385),
    .S(net4098),
    .X(_01828_));
 sg13g2_mux2_1 _21437_ (.A0(net4402),
    .A1(net3398),
    .S(net4097),
    .X(_01829_));
 sg13g2_mux2_1 _21438_ (.A0(net4395),
    .A1(net3304),
    .S(net4096),
    .X(_01830_));
 sg13g2_mux2_1 _21439_ (.A0(net4391),
    .A1(net3276),
    .S(net4096),
    .X(_01831_));
 sg13g2_mux2_1 _21440_ (.A0(net4386),
    .A1(net3519),
    .S(net4095),
    .X(_01832_));
 sg13g2_mux2_1 _21441_ (.A0(net4379),
    .A1(net3472),
    .S(net4098),
    .X(_01833_));
 sg13g2_mux2_1 _21442_ (.A0(net4374),
    .A1(net2476),
    .S(net4097),
    .X(_01834_));
 sg13g2_mux2_1 _21443_ (.A0(net4370),
    .A1(net2979),
    .S(net4098),
    .X(_01835_));
 sg13g2_or2_1 _21444_ (.X(_05325_),
    .B(_05236_),
    .A(_03169_));
 sg13g2_mux2_1 _21445_ (.A0(net4364),
    .A1(net2931),
    .S(net4090),
    .X(_01836_));
 sg13g2_mux2_1 _21446_ (.A0(net4359),
    .A1(net2648),
    .S(net4092),
    .X(_01837_));
 sg13g2_mux2_1 _21447_ (.A0(net4352),
    .A1(net2934),
    .S(net4091),
    .X(_01838_));
 sg13g2_mux2_1 _21448_ (.A0(net4348),
    .A1(net3002),
    .S(net4091),
    .X(_01839_));
 sg13g2_mux2_1 _21449_ (.A0(net4342),
    .A1(net3604),
    .S(net4092),
    .X(_01840_));
 sg13g2_mux2_1 _21450_ (.A0(net4197),
    .A1(net3484),
    .S(net4094),
    .X(_01841_));
 sg13g2_mux2_1 _21451_ (.A0(net4336),
    .A1(net3148),
    .S(net4091),
    .X(_01842_));
 sg13g2_mux2_1 _21452_ (.A0(net4333),
    .A1(net3573),
    .S(net4093),
    .X(_01843_));
 sg13g2_mux2_1 _21453_ (.A0(net4326),
    .A1(net3473),
    .S(net4092),
    .X(_01844_));
 sg13g2_mux2_1 _21454_ (.A0(net4323),
    .A1(net3146),
    .S(net4090),
    .X(_01845_));
 sg13g2_mux2_1 _21455_ (.A0(net4192),
    .A1(net2408),
    .S(net4093),
    .X(_01846_));
 sg13g2_mux2_1 _21456_ (.A0(net4188),
    .A1(net2785),
    .S(net4090),
    .X(_01847_));
 sg13g2_mux2_1 _21457_ (.A0(net4316),
    .A1(net3025),
    .S(net4093),
    .X(_01848_));
 sg13g2_mux2_1 _21458_ (.A0(net4310),
    .A1(net2484),
    .S(net4090),
    .X(_01849_));
 sg13g2_mux2_1 _21459_ (.A0(net4306),
    .A1(net2411),
    .S(net4090),
    .X(_01850_));
 sg13g2_mux2_1 _21460_ (.A0(net4298),
    .A1(net2307),
    .S(net4092),
    .X(_01851_));
 sg13g2_mux2_1 _21461_ (.A0(net4293),
    .A1(net2707),
    .S(net4094),
    .X(_01852_));
 sg13g2_mux2_1 _21462_ (.A0(net4289),
    .A1(net2380),
    .S(net4090),
    .X(_01853_));
 sg13g2_mux2_1 _21463_ (.A0(net4281),
    .A1(net3562),
    .S(net4093),
    .X(_01854_));
 sg13g2_mux2_1 _21464_ (.A0(net4278),
    .A1(net3218),
    .S(net4091),
    .X(_01855_));
 sg13g2_mux2_1 _21465_ (.A0(net4272),
    .A1(net3417),
    .S(net4092),
    .X(_01856_));
 sg13g2_mux2_1 _21466_ (.A0(net4267),
    .A1(net2535),
    .S(net4090),
    .X(_01857_));
 sg13g2_mux2_1 _21467_ (.A0(net4263),
    .A1(net3529),
    .S(net4092),
    .X(_01858_));
 sg13g2_mux2_1 _21468_ (.A0(net4257),
    .A1(net2636),
    .S(net4094),
    .X(_01859_));
 sg13g2_mux2_1 _21469_ (.A0(net4405),
    .A1(net2704),
    .S(net4093),
    .X(_01860_));
 sg13g2_mux2_1 _21470_ (.A0(net4402),
    .A1(net2977),
    .S(net4092),
    .X(_01861_));
 sg13g2_mux2_1 _21471_ (.A0(net4395),
    .A1(net2223),
    .S(net4091),
    .X(_01862_));
 sg13g2_mux2_1 _21472_ (.A0(net4391),
    .A1(net3495),
    .S(net4091),
    .X(_01863_));
 sg13g2_mux2_1 _21473_ (.A0(net4383),
    .A1(net3250),
    .S(net4090),
    .X(_01864_));
 sg13g2_mux2_1 _21474_ (.A0(net4379),
    .A1(net3169),
    .S(net4093),
    .X(_01865_));
 sg13g2_mux2_1 _21475_ (.A0(net4375),
    .A1(net3322),
    .S(net4092),
    .X(_01866_));
 sg13g2_mux2_1 _21476_ (.A0(net4370),
    .A1(net2637),
    .S(net4093),
    .X(_01867_));
 sg13g2_or2_1 _21477_ (.X(_05326_),
    .B(_09805_),
    .A(_09668_));
 sg13g2_mux2_1 _21478_ (.A0(net4363),
    .A1(net3394),
    .S(net4085),
    .X(_01868_));
 sg13g2_mux2_1 _21479_ (.A0(net4355),
    .A1(net2640),
    .S(net4087),
    .X(_01869_));
 sg13g2_mux2_1 _21480_ (.A0(net4351),
    .A1(net2795),
    .S(net4086),
    .X(_01870_));
 sg13g2_mux2_1 _21481_ (.A0(net4344),
    .A1(net2596),
    .S(net4085),
    .X(_01871_));
 sg13g2_mux2_1 _21482_ (.A0(net4340),
    .A1(net3293),
    .S(net4087),
    .X(_01872_));
 sg13g2_mux2_1 _21483_ (.A0(net4195),
    .A1(net2950),
    .S(net4087),
    .X(_01873_));
 sg13g2_mux2_1 _21484_ (.A0(net4335),
    .A1(net3170),
    .S(net4086),
    .X(_01874_));
 sg13g2_mux2_1 _21485_ (.A0(net4330),
    .A1(net2683),
    .S(net4089),
    .X(_01875_));
 sg13g2_mux2_1 _21486_ (.A0(net4325),
    .A1(net2397),
    .S(net4087),
    .X(_01876_));
 sg13g2_mux2_1 _21487_ (.A0(net4320),
    .A1(net2890),
    .S(net4086),
    .X(_01877_));
 sg13g2_mux2_1 _21488_ (.A0(net4191),
    .A1(net2736),
    .S(net4088),
    .X(_01878_));
 sg13g2_mux2_1 _21489_ (.A0(net4187),
    .A1(net2910),
    .S(net4085),
    .X(_01879_));
 sg13g2_mux2_1 _21490_ (.A0(net4312),
    .A1(net3391),
    .S(net4088),
    .X(_01880_));
 sg13g2_mux2_1 _21491_ (.A0(net4309),
    .A1(net3211),
    .S(net4085),
    .X(_01881_));
 sg13g2_mux2_1 _21492_ (.A0(net4303),
    .A1(net3277),
    .S(net4085),
    .X(_01882_));
 sg13g2_mux2_1 _21493_ (.A0(net4297),
    .A1(net3067),
    .S(net4088),
    .X(_01883_));
 sg13g2_mux2_1 _21494_ (.A0(net4292),
    .A1(net3094),
    .S(net4088),
    .X(_01884_));
 sg13g2_mux2_1 _21495_ (.A0(net4285),
    .A1(net3261),
    .S(net4085),
    .X(_01885_));
 sg13g2_mux2_1 _21496_ (.A0(net4280),
    .A1(net3487),
    .S(net4088),
    .X(_01886_));
 sg13g2_mux2_1 _21497_ (.A0(net4274),
    .A1(net3182),
    .S(net4087),
    .X(_01887_));
 sg13g2_mux2_1 _21498_ (.A0(net4270),
    .A1(net3511),
    .S(net4087),
    .X(_01888_));
 sg13g2_mux2_1 _21499_ (.A0(net4266),
    .A1(net3054),
    .S(net4085),
    .X(_01889_));
 sg13g2_mux2_1 _21500_ (.A0(net4259),
    .A1(net3227),
    .S(net4089),
    .X(_01890_));
 sg13g2_mux2_1 _21501_ (.A0(net4255),
    .A1(net3550),
    .S(net4088),
    .X(_01891_));
 sg13g2_mux2_1 _21502_ (.A0(net4403),
    .A1(net3270),
    .S(net4088),
    .X(_01892_));
 sg13g2_mux2_1 _21503_ (.A0(net4400),
    .A1(net2445),
    .S(net4087),
    .X(_01893_));
 sg13g2_mux2_1 _21504_ (.A0(net4397),
    .A1(net3213),
    .S(net4086),
    .X(_01894_));
 sg13g2_mux2_1 _21505_ (.A0(net4388),
    .A1(net3047),
    .S(net4085),
    .X(_01895_));
 sg13g2_mux2_1 _21506_ (.A0(net4385),
    .A1(net3133),
    .S(net4086),
    .X(_01896_));
 sg13g2_mux2_1 _21507_ (.A0(net4378),
    .A1(net2516),
    .S(net4089),
    .X(_01897_));
 sg13g2_mux2_1 _21508_ (.A0(net4372),
    .A1(net2806),
    .S(net4087),
    .X(_01898_));
 sg13g2_mux2_1 _21509_ (.A0(net4368),
    .A1(net2733),
    .S(net4088),
    .X(_01899_));
 sg13g2_nor2_1 _21510_ (.A(net5271),
    .B(_04966_),
    .Y(_05327_));
 sg13g2_nor2_1 _21511_ (.A(_05006_),
    .B(_05327_),
    .Y(_05328_));
 sg13g2_nand2b_2 _21512_ (.Y(_05329_),
    .B(_05005_),
    .A_N(_05327_));
 sg13g2_nor2_2 _21513_ (.A(_04955_),
    .B(net4803),
    .Y(_05330_));
 sg13g2_nand2_2 _21514_ (.Y(_05331_),
    .A(net4828),
    .B(net4658));
 sg13g2_nor2_2 _21515_ (.A(_03832_),
    .B(_03873_),
    .Y(_05332_));
 sg13g2_nand2_1 _21516_ (.Y(_05333_),
    .A(_05330_),
    .B(_05331_));
 sg13g2_nand2_2 _21517_ (.Y(_05334_),
    .A(net5047),
    .B(net4658));
 sg13g2_nor2_1 _21518_ (.A(_03945_),
    .B(_05334_),
    .Y(_05335_));
 sg13g2_nor2_1 _21519_ (.A(net5135),
    .B(_03873_),
    .Y(_05336_));
 sg13g2_o21ai_1 _21520_ (.B1(_05330_),
    .Y(_05337_),
    .A1(net5662),
    .A2(_05336_));
 sg13g2_nand3_1 _21521_ (.B(net2066),
    .C(_04955_),
    .A(_06772_),
    .Y(_05338_));
 sg13g2_o21ai_1 _21522_ (.B1(_05338_),
    .Y(_05339_),
    .A1(_05335_),
    .A2(_05337_));
 sg13g2_nand2_1 _21523_ (.Y(_05340_),
    .A(_05333_),
    .B(_05339_));
 sg13g2_o21ai_1 _21524_ (.B1(_05340_),
    .Y(_01900_),
    .A1(_06771_),
    .A2(_05333_));
 sg13g2_nand2_1 _21525_ (.Y(_05341_),
    .A(net1467),
    .B(net4570));
 sg13g2_o21ai_1 _21526_ (.B1(net1468),
    .Y(_01901_),
    .A1(net5379),
    .A2(net4570));
 sg13g2_and2_1 _21527_ (.A(net4828),
    .B(_03936_),
    .X(_05342_));
 sg13g2_nor3_1 _21528_ (.A(net5134),
    .B(_03853_),
    .C(_03902_),
    .Y(_05343_));
 sg13g2_nand3_1 _21529_ (.B(_03936_),
    .C(_03946_),
    .A(net5050),
    .Y(_05344_));
 sg13g2_nand3_1 _21530_ (.B(_05342_),
    .C(_05344_),
    .A(_03947_),
    .Y(_05345_));
 sg13g2_o21ai_1 _21531_ (.B1(_05345_),
    .Y(_01902_),
    .A1(_06883_),
    .A2(_05342_));
 sg13g2_a22oi_1 _21532_ (.Y(_05346_),
    .B1(_03971_),
    .B2(_05343_),
    .A2(net5135),
    .A1(net5657));
 sg13g2_nor2_1 _21533_ (.A(net6212),
    .B(_05342_),
    .Y(_05347_));
 sg13g2_a21oi_1 _21534_ (.A1(_05342_),
    .A2(_05346_),
    .Y(_01903_),
    .B1(_05347_));
 sg13g2_a22oi_1 _21535_ (.Y(_05348_),
    .B1(_04021_),
    .B2(_05343_),
    .A2(net5135),
    .A1(net2190));
 sg13g2_nor2_1 _21536_ (.A(net6407),
    .B(_05342_),
    .Y(_05349_));
 sg13g2_a21oi_1 _21537_ (.A1(_05342_),
    .A2(_05348_),
    .Y(_01904_),
    .B1(_05349_));
 sg13g2_and2_1 _21538_ (.A(\fpga_top.cpu_top.pc_stage.pc_int_ecall_syn_state ),
    .B(_04955_),
    .X(_05350_));
 sg13g2_nand2_2 _21539_ (.Y(_05351_),
    .A(\fpga_top.cpu_top.pc_stage.pc_int_ecall_syn_state ),
    .B(_04955_));
 sg13g2_a21oi_2 _21540_ (.B1(net4798),
    .Y(_05352_),
    .A2(_05331_),
    .A1(_05330_));
 sg13g2_nand2b_1 _21541_ (.Y(_05353_),
    .B(net2066),
    .A_N(_05352_));
 sg13g2_nand2_1 _21542_ (.Y(_05354_),
    .A(_03971_),
    .B(_05336_));
 sg13g2_nand2_1 _21543_ (.Y(_05355_),
    .A(_05330_),
    .B(_05354_));
 sg13g2_a21oi_1 _21544_ (.A1(net5656),
    .A2(_05334_),
    .Y(_05356_),
    .B1(_05355_));
 sg13g2_o21ai_1 _21545_ (.B1(_05352_),
    .Y(_05357_),
    .A1(\fpga_top.cpu_top.csr_rmie ),
    .A2(_03929_));
 sg13g2_o21ai_1 _21546_ (.B1(_05353_),
    .Y(_01905_),
    .A1(_05356_),
    .A2(_05357_));
 sg13g2_a21oi_2 _21547_ (.B1(net4803),
    .Y(_05358_),
    .A2(net4671),
    .A1(net4828));
 sg13g2_nor3_2 _21548_ (.A(_03800_),
    .B(net5134),
    .C(_03844_),
    .Y(_05359_));
 sg13g2_o21ai_1 _21549_ (.B1(net4764),
    .Y(_05360_),
    .A1(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .A2(net4650));
 sg13g2_a21o_1 _21550_ (.A2(net4650),
    .A1(_03866_),
    .B1(_05360_),
    .X(_05361_));
 sg13g2_nand4_1 _21551_ (.B(_03927_),
    .C(_03928_),
    .A(\fpga_top.cpu_top.decoder.illegal_ops_inst[0] ),
    .Y(_05362_),
    .D(_04979_));
 sg13g2_a21oi_1 _21552_ (.A1(_05361_),
    .A2(_05362_),
    .Y(_05363_),
    .B1(net4620));
 sg13g2_a21o_1 _21553_ (.A2(net4620),
    .A1(net2080),
    .B1(_05363_),
    .X(_01906_));
 sg13g2_o21ai_1 _21554_ (.B1(net4762),
    .Y(_05364_),
    .A1(\fpga_top.cpu_top.csr_wdata_mon[1] ),
    .A2(net4649));
 sg13g2_a21oi_1 _21555_ (.A1(_03880_),
    .A2(net4649),
    .Y(_05365_),
    .B1(_05364_));
 sg13g2_and4_1 _21556_ (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[1] ),
    .B(_03927_),
    .C(_03928_),
    .D(_04979_),
    .X(_05366_));
 sg13g2_nor3_1 _21557_ (.A(net4619),
    .B(_05365_),
    .C(_05366_),
    .Y(_05367_));
 sg13g2_a21oi_1 _21558_ (.A1(_06877_),
    .A2(net4618),
    .Y(_01907_),
    .B1(_05367_));
 sg13g2_nor2_1 _21559_ (.A(\fpga_top.cpu_start_adr[2] ),
    .B(net4651),
    .Y(_05368_));
 sg13g2_a21oi_1 _21560_ (.A1(_03897_),
    .A2(_05359_),
    .Y(_05369_),
    .B1(_05368_));
 sg13g2_a21oi_2 _21561_ (.B1(net5253),
    .Y(_05370_),
    .A2(net5033),
    .A1(_03929_));
 sg13g2_nor2_1 _21562_ (.A(net5585),
    .B(_04977_),
    .Y(_05371_));
 sg13g2_a21oi_1 _21563_ (.A1(_06547_),
    .A2(net5041),
    .Y(_05372_),
    .B1(_05371_));
 sg13g2_a221oi_1 _21564_ (.B2(_05372_),
    .C1(net4620),
    .B1(net4788),
    .A1(net4774),
    .Y(_05373_),
    .A2(_05369_));
 sg13g2_a21oi_1 _21565_ (.A1(_06881_),
    .A2(net4621),
    .Y(_01908_),
    .B1(_05373_));
 sg13g2_o21ai_1 _21566_ (.B1(net4762),
    .Y(_05374_),
    .A1(net5662),
    .A2(net4648));
 sg13g2_a21oi_1 _21567_ (.A1(_03946_),
    .A2(net4648),
    .Y(_05375_),
    .B1(_05374_));
 sg13g2_nor2_1 _21568_ (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[3] ),
    .B(net5042),
    .Y(_05376_));
 sg13g2_a21oi_1 _21569_ (.A1(_06584_),
    .A2(net5042),
    .Y(_05377_),
    .B1(_05376_));
 sg13g2_a21oi_1 _21570_ (.A1(net4787),
    .A2(_05377_),
    .Y(_05378_),
    .B1(_05375_));
 sg13g2_nand2_1 _21571_ (.Y(_05379_),
    .A(net1574),
    .B(net4619));
 sg13g2_o21ai_1 _21572_ (.B1(_05379_),
    .Y(_01909_),
    .A1(net4618),
    .A2(_05378_));
 sg13g2_nor2_1 _21573_ (.A(net5577),
    .B(net5815),
    .Y(_05380_));
 sg13g2_a21oi_1 _21574_ (.A1(net5576),
    .A2(_06618_),
    .Y(_05381_),
    .B1(_05380_));
 sg13g2_nor2_1 _21575_ (.A(net5381),
    .B(_05381_),
    .Y(_05382_));
 sg13g2_a22oi_1 _21576_ (.Y(_05383_),
    .B1(_05382_),
    .B2(_04528_),
    .A2(_05381_),
    .A1(net5129));
 sg13g2_nor2_1 _21577_ (.A(net5661),
    .B(net4650),
    .Y(_05384_));
 sg13g2_a21oi_1 _21578_ (.A1(net4650),
    .A2(_05383_),
    .Y(_05385_),
    .B1(_05384_));
 sg13g2_mux2_1 _21579_ (.A0(\fpga_top.cpu_top.decoder.illegal_ops_inst[4] ),
    .A1(net5598),
    .S(net5042),
    .X(_05386_));
 sg13g2_a221oi_1 _21580_ (.B2(net4787),
    .C1(net4620),
    .B1(_05386_),
    .A1(net4764),
    .Y(_05387_),
    .A2(_05385_));
 sg13g2_a21oi_1 _21581_ (.A1(_06885_),
    .A2(net4620),
    .Y(_01910_),
    .B1(_05387_));
 sg13g2_nand2_1 _21582_ (.Y(_05388_),
    .A(net5379),
    .B(net5812));
 sg13g2_nand3_1 _21583_ (.B(_04540_),
    .C(_05388_),
    .A(net5581),
    .Y(_05389_));
 sg13g2_o21ai_1 _21584_ (.B1(_05389_),
    .Y(_05390_),
    .A1(_03838_),
    .A2(_05388_));
 sg13g2_inv_2 _21585_ (.Y(_05391_),
    .A(_05390_));
 sg13g2_nor2_1 _21586_ (.A(net5659),
    .B(net4650),
    .Y(_05392_));
 sg13g2_a21oi_1 _21587_ (.A1(net4650),
    .A2(_05391_),
    .Y(_05393_),
    .B1(_05392_));
 sg13g2_nor2_1 _21588_ (.A(\fpga_top.bus_gather.i_read_adr[5] ),
    .B(net5034),
    .Y(_05394_));
 sg13g2_a21oi_1 _21589_ (.A1(_06550_),
    .A2(net5034),
    .Y(_05395_),
    .B1(_05394_));
 sg13g2_a221oi_1 _21590_ (.B2(net4787),
    .C1(net4620),
    .B1(_05395_),
    .A1(net4764),
    .Y(_05396_),
    .A2(_05393_));
 sg13g2_a21oi_1 _21591_ (.A1(_06888_),
    .A2(net4620),
    .Y(_01911_),
    .B1(_05396_));
 sg13g2_nor2_1 _21592_ (.A(\fpga_top.cpu_start_adr[6] ),
    .B(net4648),
    .Y(_05397_));
 sg13g2_a21oi_1 _21593_ (.A1(_03958_),
    .A2(net4648),
    .Y(_05398_),
    .B1(_05397_));
 sg13g2_nor2_1 _21594_ (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[6] ),
    .B(net5042),
    .Y(_05399_));
 sg13g2_a21oi_1 _21595_ (.A1(_06588_),
    .A2(net5042),
    .Y(_05400_),
    .B1(_05399_));
 sg13g2_a221oi_1 _21596_ (.B2(net4787),
    .C1(net4619),
    .B1(_05400_),
    .A1(net4763),
    .Y(_05401_),
    .A2(_05398_));
 sg13g2_a21oi_1 _21597_ (.A1(_06892_),
    .A2(net4618),
    .Y(_01912_),
    .B1(_05401_));
 sg13g2_o21ai_1 _21598_ (.B1(net4763),
    .Y(_05402_),
    .A1(net5657),
    .A2(net4648));
 sg13g2_a21oi_1 _21599_ (.A1(_03972_),
    .A2(net4648),
    .Y(_05403_),
    .B1(_05402_));
 sg13g2_nor2_1 _21600_ (.A(\fpga_top.bus_gather.i_read_adr[7] ),
    .B(net5034),
    .Y(_05404_));
 sg13g2_a21oi_1 _21601_ (.A1(_06564_),
    .A2(net5033),
    .Y(_05405_),
    .B1(_05404_));
 sg13g2_a21oi_1 _21602_ (.A1(net4787),
    .A2(_05405_),
    .Y(_05406_),
    .B1(_05403_));
 sg13g2_nand2_1 _21603_ (.Y(_05407_),
    .A(net1415),
    .B(net4618));
 sg13g2_o21ai_1 _21604_ (.B1(_05407_),
    .Y(_01913_),
    .A1(net4618),
    .A2(_05406_));
 sg13g2_nor2_1 _21605_ (.A(net5655),
    .B(net4649),
    .Y(_05408_));
 sg13g2_a21oi_1 _21606_ (.A1(_03982_),
    .A2(net4649),
    .Y(_05409_),
    .B1(_05408_));
 sg13g2_nor2_1 _21607_ (.A(net5595),
    .B(net5033),
    .Y(_05410_));
 sg13g2_a21oi_1 _21608_ (.A1(_06560_),
    .A2(net5033),
    .Y(_05411_),
    .B1(_05410_));
 sg13g2_a221oi_1 _21609_ (.B2(net4787),
    .C1(net4619),
    .B1(_05411_),
    .A1(net4762),
    .Y(_05412_),
    .A2(_05409_));
 sg13g2_a21oi_1 _21610_ (.A1(_06899_),
    .A2(net4618),
    .Y(_01914_),
    .B1(_05412_));
 sg13g2_nor2_1 _21611_ (.A(net5653),
    .B(net4651),
    .Y(_05413_));
 sg13g2_a21oi_1 _21612_ (.A1(_03997_),
    .A2(net4651),
    .Y(_05414_),
    .B1(_05413_));
 sg13g2_nor2_1 _21613_ (.A(\fpga_top.cpu_top.br_ofs[2] ),
    .B(_04977_),
    .Y(_05415_));
 sg13g2_a21oi_1 _21614_ (.A1(_06592_),
    .A2(net5041),
    .Y(_05416_),
    .B1(_05415_));
 sg13g2_a22oi_1 _21615_ (.Y(_05417_),
    .B1(_05416_),
    .B2(net4788),
    .A2(_05414_),
    .A1(net4774));
 sg13g2_nand2_1 _21616_ (.Y(_05418_),
    .A(net1465),
    .B(net4621));
 sg13g2_o21ai_1 _21617_ (.B1(_05418_),
    .Y(_01915_),
    .A1(net4621),
    .A2(_05417_));
 sg13g2_nor2_1 _21618_ (.A(net5652),
    .B(net4653),
    .Y(_05419_));
 sg13g2_a21oi_1 _21619_ (.A1(_04007_),
    .A2(net4653),
    .Y(_05420_),
    .B1(_05419_));
 sg13g2_nor2_1 _21620_ (.A(\fpga_top.bus_gather.i_read_adr[10] ),
    .B(net5035),
    .Y(_05421_));
 sg13g2_a21oi_2 _21621_ (.B1(_05421_),
    .Y(_05422_),
    .A2(net5035),
    .A1(_06569_));
 sg13g2_a22oi_1 _21622_ (.Y(_05423_),
    .B1(_05422_),
    .B2(net4790),
    .A2(_05420_),
    .A1(net4769));
 sg13g2_nand2_1 _21623_ (.Y(_05424_),
    .A(net1533),
    .B(net4623));
 sg13g2_o21ai_1 _21624_ (.B1(_05424_),
    .Y(_01916_),
    .A1(net4623),
    .A2(_05423_));
 sg13g2_o21ai_1 _21625_ (.B1(net4762),
    .Y(_05425_),
    .A1(net5651),
    .A2(net4648));
 sg13g2_a21oi_1 _21626_ (.A1(_04022_),
    .A2(net4648),
    .Y(_05426_),
    .B1(_05425_));
 sg13g2_nor2_1 _21627_ (.A(\fpga_top.bus_gather.i_read_adr[11] ),
    .B(net5033),
    .Y(_05427_));
 sg13g2_a21oi_1 _21628_ (.A1(_06576_),
    .A2(net5033),
    .Y(_05428_),
    .B1(_05427_));
 sg13g2_a21oi_1 _21629_ (.A1(net4787),
    .A2(_05428_),
    .Y(_05429_),
    .B1(_05426_));
 sg13g2_nand2_1 _21630_ (.Y(_05430_),
    .A(net1500),
    .B(net4618));
 sg13g2_o21ai_1 _21631_ (.B1(_05430_),
    .Y(_01917_),
    .A1(net4618),
    .A2(_05429_));
 sg13g2_nor2_1 _21632_ (.A(\fpga_top.cpu_start_adr[12] ),
    .B(net4649),
    .Y(_05431_));
 sg13g2_a21oi_1 _21633_ (.A1(_04035_),
    .A2(net4649),
    .Y(_05432_),
    .B1(_05431_));
 sg13g2_nor2_1 _21634_ (.A(\fpga_top.bus_gather.i_read_adr[12] ),
    .B(net5034),
    .Y(_05433_));
 sg13g2_a21oi_1 _21635_ (.A1(_06552_),
    .A2(net5034),
    .Y(_05434_),
    .B1(_05433_));
 sg13g2_a22oi_1 _21636_ (.Y(_05435_),
    .B1(_05434_),
    .B2(net4787),
    .A2(_05432_),
    .A1(net4762));
 sg13g2_nand2_1 _21637_ (.Y(_05436_),
    .A(net1432),
    .B(net4619));
 sg13g2_o21ai_1 _21638_ (.B1(_05436_),
    .Y(_01918_),
    .A1(net4619),
    .A2(_05435_));
 sg13g2_nor2_1 _21639_ (.A(\fpga_top.cpu_start_adr[13] ),
    .B(net4652),
    .Y(_05437_));
 sg13g2_a21oi_1 _21640_ (.A1(_04046_),
    .A2(net4652),
    .Y(_05438_),
    .B1(_05437_));
 sg13g2_nor2_1 _21641_ (.A(\fpga_top.bus_gather.i_read_adr[13] ),
    .B(net5040),
    .Y(_05439_));
 sg13g2_a21oi_1 _21642_ (.A1(net5381),
    .A2(net5040),
    .Y(_05440_),
    .B1(_05439_));
 sg13g2_a22oi_1 _21643_ (.Y(_05441_),
    .B1(_05440_),
    .B2(net4791),
    .A2(_05438_),
    .A1(net4767));
 sg13g2_nand2_1 _21644_ (.Y(_05442_),
    .A(net1503),
    .B(net4622));
 sg13g2_o21ai_1 _21645_ (.B1(_05442_),
    .Y(_01919_),
    .A1(net4622),
    .A2(_05441_));
 sg13g2_o21ai_1 _21646_ (.B1(net4766),
    .Y(_05443_),
    .A1(net5650),
    .A2(net4651));
 sg13g2_a21oi_1 _21647_ (.A1(_04060_),
    .A2(net4651),
    .Y(_05444_),
    .B1(_05443_));
 sg13g2_o21ai_1 _21648_ (.B1(net4788),
    .Y(_05445_),
    .A1(\fpga_top.bus_gather.i_read_adr[14] ),
    .A2(net5035));
 sg13g2_a21oi_1 _21649_ (.A1(net5380),
    .A2(net5035),
    .Y(_05446_),
    .B1(_05445_));
 sg13g2_nor3_1 _21650_ (.A(net4621),
    .B(_05444_),
    .C(_05446_),
    .Y(_05447_));
 sg13g2_a21oi_1 _21651_ (.A1(_06908_),
    .A2(net4621),
    .Y(_01920_),
    .B1(_05447_));
 sg13g2_nor2_1 _21652_ (.A(\fpga_top.cpu_start_adr[15] ),
    .B(net4652),
    .Y(_05448_));
 sg13g2_a21oi_1 _21653_ (.A1(_04069_),
    .A2(net4652),
    .Y(_05449_),
    .B1(_05448_));
 sg13g2_nor2_1 _21654_ (.A(\fpga_top.cpu_top.csr_uimm[0] ),
    .B(net5041),
    .Y(_05450_));
 sg13g2_a21oi_1 _21655_ (.A1(_06605_),
    .A2(net5041),
    .Y(_05451_),
    .B1(_05450_));
 sg13g2_a22oi_1 _21656_ (.Y(_05452_),
    .B1(_05451_),
    .B2(net4791),
    .A2(_05449_),
    .A1(net4767));
 sg13g2_nand2_1 _21657_ (.Y(_05453_),
    .A(net1474),
    .B(net4622));
 sg13g2_o21ai_1 _21658_ (.B1(_05453_),
    .Y(_01921_),
    .A1(net4622),
    .A2(_05452_));
 sg13g2_mux2_1 _21659_ (.A0(net5649),
    .A1(_04081_),
    .S(net4652),
    .X(_05454_));
 sg13g2_nor2_1 _21660_ (.A(net5594),
    .B(net5040),
    .Y(_05455_));
 sg13g2_a21oi_1 _21661_ (.A1(_06608_),
    .A2(net5040),
    .Y(_05456_),
    .B1(_05455_));
 sg13g2_a22oi_1 _21662_ (.Y(_05457_),
    .B1(_05456_),
    .B2(net4791),
    .A2(_05454_),
    .A1(net4767));
 sg13g2_nand2_1 _21663_ (.Y(_05458_),
    .A(net1416),
    .B(net4622));
 sg13g2_o21ai_1 _21664_ (.B1(_05458_),
    .Y(_01922_),
    .A1(net4627),
    .A2(_05457_));
 sg13g2_nor2_1 _21665_ (.A(net5648),
    .B(net4653),
    .Y(_05459_));
 sg13g2_a21oi_1 _21666_ (.A1(_04091_),
    .A2(net4653),
    .Y(_05460_),
    .B1(_05459_));
 sg13g2_nor2_1 _21667_ (.A(net6614),
    .B(net5041),
    .Y(_05461_));
 sg13g2_a21oi_2 _21668_ (.B1(_05461_),
    .Y(_05462_),
    .A2(net5041),
    .A1(_06611_));
 sg13g2_a22oi_1 _21669_ (.Y(_05463_),
    .B1(_05462_),
    .B2(net4790),
    .A2(_05460_),
    .A1(net4769));
 sg13g2_nand2_1 _21670_ (.Y(_05464_),
    .A(net1462),
    .B(net4626));
 sg13g2_o21ai_1 _21671_ (.B1(_05464_),
    .Y(_01923_),
    .A1(net4623),
    .A2(_05463_));
 sg13g2_nor2_1 _21672_ (.A(net5647),
    .B(net4652),
    .Y(_05465_));
 sg13g2_a21oi_1 _21673_ (.A1(_04099_),
    .A2(net4657),
    .Y(_05466_),
    .B1(_05465_));
 sg13g2_nand2_1 _21674_ (.Y(_05467_),
    .A(\fpga_top.cpu_top.csr_uimm[3] ),
    .B(net5040));
 sg13g2_o21ai_1 _21675_ (.B1(_05467_),
    .Y(_05468_),
    .A1(_06614_),
    .A2(net5040));
 sg13g2_a22oi_1 _21676_ (.Y(_05469_),
    .B1(_05468_),
    .B2(net4791),
    .A2(_05466_),
    .A1(net4768));
 sg13g2_nand2_1 _21677_ (.Y(_05470_),
    .A(net1544),
    .B(net4623));
 sg13g2_o21ai_1 _21678_ (.B1(_05470_),
    .Y(_01924_),
    .A1(net4627),
    .A2(_05469_));
 sg13g2_nor2_1 _21679_ (.A(\fpga_top.cpu_start_adr[19] ),
    .B(net4654),
    .Y(_05471_));
 sg13g2_a21oi_1 _21680_ (.A1(_04109_),
    .A2(net4654),
    .Y(_05472_),
    .B1(_05471_));
 sg13g2_nor2_1 _21681_ (.A(\fpga_top.bus_gather.i_read_adr[19] ),
    .B(net5037),
    .Y(_05473_));
 sg13g2_a21oi_1 _21682_ (.A1(_06618_),
    .A2(net5037),
    .Y(_05474_),
    .B1(_05473_));
 sg13g2_a221oi_1 _21683_ (.B2(net4790),
    .C1(net4624),
    .B1(_05474_),
    .A1(net4770),
    .Y(_05475_),
    .A2(_05472_));
 sg13g2_a21oi_1 _21684_ (.A1(_06914_),
    .A2(net4624),
    .Y(_01925_),
    .B1(_05475_));
 sg13g2_nor2_1 _21685_ (.A(net5646),
    .B(net4653),
    .Y(_05476_));
 sg13g2_a21oi_1 _21686_ (.A1(_04122_),
    .A2(net4656),
    .Y(_05477_),
    .B1(_05476_));
 sg13g2_nor2_1 _21687_ (.A(\fpga_top.bus_gather.i_read_adr[20] ),
    .B(net5037),
    .Y(_05478_));
 sg13g2_a21oi_1 _21688_ (.A1(_06563_),
    .A2(net5037),
    .Y(_05479_),
    .B1(_05478_));
 sg13g2_a22oi_1 _21689_ (.Y(_05480_),
    .B1(_05479_),
    .B2(net4789),
    .A2(_05477_),
    .A1(net4769));
 sg13g2_nand2_1 _21690_ (.Y(_05481_),
    .A(net1593),
    .B(net4623));
 sg13g2_o21ai_1 _21691_ (.B1(_05481_),
    .Y(_01926_),
    .A1(net4623),
    .A2(_05480_));
 sg13g2_nor2_1 _21692_ (.A(net5645),
    .B(net4655),
    .Y(_05482_));
 sg13g2_a21oi_1 _21693_ (.A1(_04132_),
    .A2(net4655),
    .Y(_05483_),
    .B1(_05482_));
 sg13g2_nor2_1 _21694_ (.A(\fpga_top.bus_gather.i_read_adr[21] ),
    .B(net5036),
    .Y(_05484_));
 sg13g2_a21oi_1 _21695_ (.A1(_06559_),
    .A2(net5038),
    .Y(_05485_),
    .B1(_05484_));
 sg13g2_a221oi_1 _21696_ (.B2(net4789),
    .C1(net4625),
    .B1(_05485_),
    .A1(net4770),
    .Y(_05486_),
    .A2(_05483_));
 sg13g2_a21oi_1 _21697_ (.A1(_06915_),
    .A2(net4625),
    .Y(_01927_),
    .B1(_05486_));
 sg13g2_nor2_1 _21698_ (.A(net5643),
    .B(net4657),
    .Y(_05487_));
 sg13g2_a21oi_1 _21699_ (.A1(_04144_),
    .A2(net4653),
    .Y(_05488_),
    .B1(_05487_));
 sg13g2_nor2_1 _21700_ (.A(net5592),
    .B(net5037),
    .Y(_05489_));
 sg13g2_a21oi_1 _21701_ (.A1(_06548_),
    .A2(net5037),
    .Y(_05490_),
    .B1(_05489_));
 sg13g2_a22oi_1 _21702_ (.Y(_05491_),
    .B1(_05490_),
    .B2(net4789),
    .A2(_05488_),
    .A1(net4769));
 sg13g2_nand2_1 _21703_ (.Y(_05492_),
    .A(net1424),
    .B(net4625));
 sg13g2_o21ai_1 _21704_ (.B1(_05492_),
    .Y(_01928_),
    .A1(net4623),
    .A2(_05491_));
 sg13g2_nor2_1 _21705_ (.A(net5642),
    .B(net4654),
    .Y(_05493_));
 sg13g2_a21oi_1 _21706_ (.A1(_04154_),
    .A2(net4654),
    .Y(_05494_),
    .B1(_05493_));
 sg13g2_nor2_1 _21707_ (.A(\fpga_top.bus_gather.i_read_adr[23] ),
    .B(net5037),
    .Y(_05495_));
 sg13g2_a21oi_1 _21708_ (.A1(_06568_),
    .A2(net5036),
    .Y(_05496_),
    .B1(_05495_));
 sg13g2_a221oi_1 _21709_ (.B2(net4789),
    .C1(net4625),
    .B1(_05496_),
    .A1(net4770),
    .Y(_05497_),
    .A2(_05494_));
 sg13g2_a21oi_1 _21710_ (.A1(_06916_),
    .A2(net4624),
    .Y(_01929_),
    .B1(_05497_));
 sg13g2_nor2_1 _21711_ (.A(\fpga_top.cpu_start_adr[24] ),
    .B(net4652),
    .Y(_05498_));
 sg13g2_a21oi_1 _21712_ (.A1(_04166_),
    .A2(net4657),
    .Y(_05499_),
    .B1(_05498_));
 sg13g2_nor2_1 _21713_ (.A(\fpga_top.bus_gather.i_read_adr[24] ),
    .B(net5039),
    .Y(_05500_));
 sg13g2_a21oi_1 _21714_ (.A1(_06575_),
    .A2(net5039),
    .Y(_05501_),
    .B1(_05500_));
 sg13g2_a22oi_1 _21715_ (.Y(_05502_),
    .B1(_05501_),
    .B2(net4791),
    .A2(_05499_),
    .A1(net4768));
 sg13g2_nand2_1 _21716_ (.Y(_05503_),
    .A(net1508),
    .B(net4622));
 sg13g2_o21ai_1 _21717_ (.B1(_05503_),
    .Y(_01930_),
    .A1(net4622),
    .A2(_05502_));
 sg13g2_o21ai_1 _21718_ (.B1(net4768),
    .Y(_05504_),
    .A1(\fpga_top.cpu_start_adr[25] ),
    .A2(net4652));
 sg13g2_a21oi_1 _21719_ (.A1(_04176_),
    .A2(net4657),
    .Y(_05505_),
    .B1(_05504_));
 sg13g2_o21ai_1 _21720_ (.B1(net4791),
    .Y(_05506_),
    .A1(\fpga_top.bus_gather.i_read_adr[25] ),
    .A2(net5040));
 sg13g2_a21oi_1 _21721_ (.A1(_06558_),
    .A2(net5039),
    .Y(_05507_),
    .B1(_05506_));
 sg13g2_nor2_1 _21722_ (.A(_05505_),
    .B(_05507_),
    .Y(_05508_));
 sg13g2_nand2_1 _21723_ (.Y(_05509_),
    .A(net1444),
    .B(net4627));
 sg13g2_o21ai_1 _21724_ (.B1(_05509_),
    .Y(_01931_),
    .A1(net4622),
    .A2(_05508_));
 sg13g2_nor2_1 _21725_ (.A(\fpga_top.cpu_start_adr[26] ),
    .B(net4655),
    .Y(_05510_));
 sg13g2_a21oi_1 _21726_ (.A1(_04186_),
    .A2(net4655),
    .Y(_05511_),
    .B1(_05510_));
 sg13g2_nor2_1 _21727_ (.A(\fpga_top.bus_gather.i_read_adr[26] ),
    .B(net5036),
    .Y(_05512_));
 sg13g2_a21oi_1 _21728_ (.A1(_06549_),
    .A2(net5036),
    .Y(_05513_),
    .B1(_05512_));
 sg13g2_a22oi_1 _21729_ (.Y(_05514_),
    .B1(_05513_),
    .B2(net4789),
    .A2(_05511_),
    .A1(net4770));
 sg13g2_nand2_1 _21730_ (.Y(_05515_),
    .A(net1430),
    .B(net4624));
 sg13g2_o21ai_1 _21731_ (.B1(_05515_),
    .Y(_01932_),
    .A1(net4624),
    .A2(_05514_));
 sg13g2_nor2_1 _21732_ (.A(net5641),
    .B(net4654),
    .Y(_05516_));
 sg13g2_a21oi_1 _21733_ (.A1(_04197_),
    .A2(net4654),
    .Y(_05517_),
    .B1(_05516_));
 sg13g2_nor2_1 _21734_ (.A(\fpga_top.bus_gather.i_read_adr[27] ),
    .B(net5036),
    .Y(_05518_));
 sg13g2_a21oi_1 _21735_ (.A1(_06554_),
    .A2(net5036),
    .Y(_05519_),
    .B1(_05518_));
 sg13g2_a22oi_1 _21736_ (.Y(_05520_),
    .B1(_05519_),
    .B2(net4789),
    .A2(_05517_),
    .A1(net4773));
 sg13g2_nand2_1 _21737_ (.Y(_05521_),
    .A(net1473),
    .B(net4624));
 sg13g2_o21ai_1 _21738_ (.B1(_05521_),
    .Y(_01933_),
    .A1(net4624),
    .A2(_05520_));
 sg13g2_o21ai_1 _21739_ (.B1(net4773),
    .Y(_05522_),
    .A1(net5638),
    .A2(net4656));
 sg13g2_a21oi_1 _21740_ (.A1(_04210_),
    .A2(net4656),
    .Y(_05523_),
    .B1(_05522_));
 sg13g2_o21ai_1 _21741_ (.B1(net4789),
    .Y(_05524_),
    .A1(net5590),
    .A2(net5038));
 sg13g2_a21oi_1 _21742_ (.A1(_06555_),
    .A2(net5038),
    .Y(_05525_),
    .B1(_05524_));
 sg13g2_nor2_1 _21743_ (.A(_05523_),
    .B(_05525_),
    .Y(_05526_));
 sg13g2_nand2_1 _21744_ (.Y(_05527_),
    .A(net1463),
    .B(net4626));
 sg13g2_o21ai_1 _21745_ (.B1(_05527_),
    .Y(_01934_),
    .A1(net4626),
    .A2(_05526_));
 sg13g2_nor2_1 _21746_ (.A(net5637),
    .B(net4654),
    .Y(_05528_));
 sg13g2_a21oi_1 _21747_ (.A1(_04219_),
    .A2(net4654),
    .Y(_05529_),
    .B1(_05528_));
 sg13g2_nor2_1 _21748_ (.A(\fpga_top.bus_gather.i_read_adr[29] ),
    .B(net5036),
    .Y(_05530_));
 sg13g2_a21oi_1 _21749_ (.A1(_06556_),
    .A2(net5036),
    .Y(_05531_),
    .B1(_05530_));
 sg13g2_a22oi_1 _21750_ (.Y(_05532_),
    .B1(_05531_),
    .B2(net4789),
    .A2(_05529_),
    .A1(net4772));
 sg13g2_nand2_1 _21751_ (.Y(_05533_),
    .A(net1594),
    .B(net4624));
 sg13g2_o21ai_1 _21752_ (.B1(_05533_),
    .Y(_01935_),
    .A1(net4625),
    .A2(_05532_));
 sg13g2_nor2_1 _21753_ (.A(net5635),
    .B(net4653),
    .Y(_05534_));
 sg13g2_a21oi_1 _21754_ (.A1(_04231_),
    .A2(net4653),
    .Y(_05535_),
    .B1(_05534_));
 sg13g2_nor2_1 _21755_ (.A(\fpga_top.bus_gather.i_read_adr[30] ),
    .B(net5039),
    .Y(_05536_));
 sg13g2_a21oi_1 _21756_ (.A1(_06557_),
    .A2(net5039),
    .Y(_05537_),
    .B1(_05536_));
 sg13g2_a22oi_1 _21757_ (.Y(_05538_),
    .B1(_05537_),
    .B2(net4790),
    .A2(_05535_),
    .A1(net4773));
 sg13g2_nand2_1 _21758_ (.Y(_05539_),
    .A(net1410),
    .B(net4626));
 sg13g2_o21ai_1 _21759_ (.B1(_05539_),
    .Y(_01936_),
    .A1(net4623),
    .A2(_05538_));
 sg13g2_nor2_1 _21760_ (.A(\fpga_top.cpu_start_adr[31] ),
    .B(net4651),
    .Y(_05540_));
 sg13g2_a21oi_1 _21761_ (.A1(_04244_),
    .A2(net4651),
    .Y(_05541_),
    .B1(_05540_));
 sg13g2_nor2_1 _21762_ (.A(\fpga_top.cpu_top.br_ofs[12] ),
    .B(net5041),
    .Y(_05542_));
 sg13g2_a21oi_1 _21763_ (.A1(_06646_),
    .A2(net5041),
    .Y(_05543_),
    .B1(_05542_));
 sg13g2_a221oi_1 _21764_ (.B2(net4788),
    .C1(net4620),
    .B1(_05543_),
    .A1(net4766),
    .Y(_05544_),
    .A2(_05541_));
 sg13g2_a21oi_1 _21765_ (.A1(_06921_),
    .A2(net4621),
    .Y(_01937_),
    .B1(_05544_));
 sg13g2_and2_1 _21766_ (.A(net5048),
    .B(_03866_),
    .X(_05545_));
 sg13g2_nor2_2 _21767_ (.A(net5137),
    .B(_03847_),
    .Y(_05546_));
 sg13g2_nand2_1 _21768_ (.Y(_05547_),
    .A(net5047),
    .B(net4670));
 sg13g2_nor3_2 _21769_ (.A(_03832_),
    .B(_03847_),
    .C(net4803),
    .Y(_05548_));
 sg13g2_o21ai_1 _21770_ (.B1(_05548_),
    .Y(_05549_),
    .A1(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .A2(net4580));
 sg13g2_a21oi_2 _21771_ (.B1(net4803),
    .Y(_05550_),
    .A2(net4670),
    .A1(net4829));
 sg13g2_a22oi_1 _21772_ (.Y(_05551_),
    .B1(_05550_),
    .B2(net3493),
    .A2(net4804),
    .A1(_04980_));
 sg13g2_o21ai_1 _21773_ (.B1(_05551_),
    .Y(_01938_),
    .A1(_05545_),
    .A2(_05549_));
 sg13g2_nor2_1 _21774_ (.A(_03880_),
    .B(_05547_),
    .Y(_05552_));
 sg13g2_a21oi_1 _21775_ (.A1(\fpga_top.cpu_top.csr_wdata_mon[1] ),
    .A2(_05547_),
    .Y(_05553_),
    .B1(_05552_));
 sg13g2_a22oi_1 _21776_ (.Y(_01939_),
    .B1(_05553_),
    .B2(_05548_),
    .A2(_05550_),
    .A1(_06876_));
 sg13g2_a22oi_1 _21777_ (.Y(_05554_),
    .B1(_05550_),
    .B2(net3781),
    .A2(net4803),
    .A1(_05007_));
 sg13g2_o21ai_1 _21778_ (.B1(_05548_),
    .Y(_05555_),
    .A1(\fpga_top.cpu_start_adr[2] ),
    .A2(_05546_));
 sg13g2_a21oi_1 _21779_ (.A1(_03897_),
    .A2(_05546_),
    .Y(_05556_),
    .B1(_05555_));
 sg13g2_nand2b_1 _21780_ (.Y(_01940_),
    .B(_05554_),
    .A_N(_05556_));
 sg13g2_a22oi_1 _21781_ (.Y(_05557_),
    .B1(_05550_),
    .B2(net3489),
    .A2(net4803),
    .A1(_05023_));
 sg13g2_nor2_1 _21782_ (.A(_03945_),
    .B(_05547_),
    .Y(_05558_));
 sg13g2_o21ai_1 _21783_ (.B1(_05548_),
    .Y(_05559_),
    .A1(net5663),
    .A2(net4580));
 sg13g2_o21ai_1 _21784_ (.B1(_05557_),
    .Y(_01941_),
    .A1(_05558_),
    .A2(_05559_));
 sg13g2_a21oi_1 _21785_ (.A1(_05034_),
    .A2(_05327_),
    .Y(_05560_),
    .B1(_05550_));
 sg13g2_o21ai_1 _21786_ (.B1(net4765),
    .Y(_05561_),
    .A1(net5661),
    .A2(net4580));
 sg13g2_a21o_1 _21787_ (.A2(net4580),
    .A1(_05383_),
    .B1(_05561_),
    .X(_05562_));
 sg13g2_a22oi_1 _21788_ (.Y(_01942_),
    .B1(_05560_),
    .B2(_05562_),
    .A2(_05550_),
    .A1(_06886_));
 sg13g2_o21ai_1 _21789_ (.B1(net4764),
    .Y(_05563_),
    .A1(net5659),
    .A2(net4580));
 sg13g2_a21o_1 _21790_ (.A2(net4580),
    .A1(_05391_),
    .B1(_05563_),
    .X(_05564_));
 sg13g2_a22oi_1 _21791_ (.Y(_01943_),
    .B1(_05560_),
    .B2(_05564_),
    .A2(_05550_),
    .A1(_06889_));
 sg13g2_a22oi_1 _21792_ (.Y(_05565_),
    .B1(_05550_),
    .B2(net3598),
    .A2(net4804),
    .A1(net5254));
 sg13g2_o21ai_1 _21793_ (.B1(_05548_),
    .Y(_05566_),
    .A1(\fpga_top.cpu_start_adr[31] ),
    .A2(net4580));
 sg13g2_a21oi_1 _21794_ (.A1(_04244_),
    .A2(net4580),
    .Y(_05567_),
    .B1(_05566_));
 sg13g2_nand2b_1 _21795_ (.Y(_01944_),
    .B(_05565_),
    .A_N(_05567_));
 sg13g2_nand2_1 _21796_ (.Y(_05568_),
    .A(net4828),
    .B(net4686));
 sg13g2_and3_1 _21797_ (.X(_05569_),
    .A(net4764),
    .B(net4792),
    .C(_05568_));
 sg13g2_nand3_1 _21798_ (.B(net4792),
    .C(_05568_),
    .A(net4765),
    .Y(_05570_));
 sg13g2_nand2_1 _21799_ (.Y(_05571_),
    .A(net1964),
    .B(net4611));
 sg13g2_a21oi_1 _21800_ (.A1(net5386),
    .A2(net4573),
    .Y(_05572_),
    .B1(net4775));
 sg13g2_o21ai_1 _21801_ (.B1(_05572_),
    .Y(_05573_),
    .A1(_08155_),
    .A2(net4573));
 sg13g2_a21oi_2 _21802_ (.B1(net5253),
    .Y(_05574_),
    .A2(_04922_),
    .A1(_03929_));
 sg13g2_a22oi_1 _21803_ (.Y(_05575_),
    .B1(net4757),
    .B2(_06547_),
    .A2(net4741),
    .A1(_06882_));
 sg13g2_nand3_1 _21804_ (.B(_05573_),
    .C(_05575_),
    .A(net4804),
    .Y(_05576_));
 sg13g2_and2_1 _21805_ (.A(net5057),
    .B(net4687),
    .X(_05577_));
 sg13g2_a21oi_1 _21806_ (.A1(_03897_),
    .A2(net4641),
    .Y(_05578_),
    .B1(net4804));
 sg13g2_o21ai_1 _21807_ (.B1(_05578_),
    .Y(_05579_),
    .A1(\fpga_top.cpu_start_adr[2] ),
    .A2(net4639));
 sg13g2_nand3_1 _21808_ (.B(_05576_),
    .C(_05579_),
    .A(net4792),
    .Y(_05580_));
 sg13g2_o21ai_1 _21809_ (.B1(_05580_),
    .Y(_05581_),
    .A1(net1810),
    .A2(net4792));
 sg13g2_o21ai_1 _21810_ (.B1(_05571_),
    .Y(_01945_),
    .A1(net4611),
    .A2(_05581_));
 sg13g2_nand2_1 _21811_ (.Y(_05582_),
    .A(net1752),
    .B(net4611));
 sg13g2_nand2_1 _21812_ (.Y(_05583_),
    .A(_08189_),
    .B(net4571));
 sg13g2_o21ai_1 _21813_ (.B1(_05583_),
    .Y(_05584_),
    .A1(_08186_),
    .A2(net4571));
 sg13g2_o21ai_1 _21814_ (.B1(net4775),
    .Y(_05585_),
    .A1(\fpga_top.bus_gather.i_read_adr[3] ),
    .A2(net5253));
 sg13g2_o21ai_1 _21815_ (.B1(_05585_),
    .Y(_05586_),
    .A1(net4757),
    .A2(_05584_));
 sg13g2_o21ai_1 _21816_ (.B1(_05586_),
    .Y(_05587_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[3] ),
    .A2(net4727));
 sg13g2_o21ai_1 _21817_ (.B1(net4762),
    .Y(_05588_),
    .A1(net5663),
    .A2(net4638));
 sg13g2_a21oi_1 _21818_ (.A1(_03946_),
    .A2(net4638),
    .Y(_05589_),
    .B1(_05588_));
 sg13g2_nor2_1 _21819_ (.A(net4798),
    .B(_05589_),
    .Y(_05590_));
 sg13g2_o21ai_1 _21820_ (.B1(_05590_),
    .Y(_05591_),
    .A1(net4765),
    .A2(_05587_));
 sg13g2_o21ai_1 _21821_ (.B1(_05591_),
    .Y(_05592_),
    .A1(net1699),
    .A2(net4792));
 sg13g2_o21ai_1 _21822_ (.B1(_05582_),
    .Y(_01946_),
    .A1(net4611),
    .A2(_05592_));
 sg13g2_nand2_1 _21823_ (.Y(_05593_),
    .A(net1878),
    .B(net4612));
 sg13g2_a21oi_1 _21824_ (.A1(_08221_),
    .A2(net4572),
    .Y(_05594_),
    .B1(net4757));
 sg13g2_o21ai_1 _21825_ (.B1(_05594_),
    .Y(_05595_),
    .A1(_08218_),
    .A2(net4572));
 sg13g2_o21ai_1 _21826_ (.B1(net4775),
    .Y(_05596_),
    .A1(net5598),
    .A2(net5254));
 sg13g2_a221oi_1 _21827_ (.B2(_05596_),
    .C1(net4765),
    .B1(_05595_),
    .A1(_06887_),
    .Y(_05597_),
    .A2(net4741));
 sg13g2_o21ai_1 _21828_ (.B1(net4765),
    .Y(_05598_),
    .A1(net5661),
    .A2(net4639));
 sg13g2_a21oi_1 _21829_ (.A1(_05383_),
    .A2(net4641),
    .Y(_05599_),
    .B1(_05598_));
 sg13g2_nor3_1 _21830_ (.A(net4798),
    .B(_05597_),
    .C(_05599_),
    .Y(_05600_));
 sg13g2_o21ai_1 _21831_ (.B1(net4608),
    .Y(_05601_),
    .A1(\fpga_top.cpu_top.execution.csr_array.pc_excep2[4] ),
    .A2(net4792));
 sg13g2_o21ai_1 _21832_ (.B1(_05593_),
    .Y(_01947_),
    .A1(_05600_),
    .A2(_05601_));
 sg13g2_nand2_1 _21833_ (.Y(_05602_),
    .A(net1923),
    .B(net4611));
 sg13g2_a21oi_1 _21834_ (.A1(_08099_),
    .A2(net4571),
    .Y(_05603_),
    .B1(net4757));
 sg13g2_o21ai_1 _21835_ (.B1(_05603_),
    .Y(_05604_),
    .A1(_08097_),
    .A2(net4571));
 sg13g2_o21ai_1 _21836_ (.B1(net4775),
    .Y(_05605_),
    .A1(\fpga_top.bus_gather.i_read_adr[5] ),
    .A2(net5253));
 sg13g2_o21ai_1 _21837_ (.B1(net4803),
    .Y(_05606_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[5] ),
    .A2(net4727));
 sg13g2_a21oi_1 _21838_ (.A1(_05604_),
    .A2(_05605_),
    .Y(_05607_),
    .B1(_05606_));
 sg13g2_o21ai_1 _21839_ (.B1(net4764),
    .Y(_05608_),
    .A1(net5659),
    .A2(net4639));
 sg13g2_a21oi_1 _21840_ (.A1(_05391_),
    .A2(net4641),
    .Y(_05609_),
    .B1(_05608_));
 sg13g2_nor3_1 _21841_ (.A(net4798),
    .B(_05607_),
    .C(_05609_),
    .Y(_05610_));
 sg13g2_o21ai_1 _21842_ (.B1(net4608),
    .Y(_05611_),
    .A1(net1520),
    .A2(net4793));
 sg13g2_o21ai_1 _21843_ (.B1(_05602_),
    .Y(_01948_),
    .A1(_05610_),
    .A2(_05611_));
 sg13g2_nand2_1 _21844_ (.Y(_05612_),
    .A(net2311),
    .B(net4611));
 sg13g2_a21oi_1 _21845_ (.A1(_08245_),
    .A2(net4571),
    .Y(_05613_),
    .B1(net4757));
 sg13g2_o21ai_1 _21846_ (.B1(_05613_),
    .Y(_05614_),
    .A1(_08243_),
    .A2(net4571));
 sg13g2_o21ai_1 _21847_ (.B1(net4775),
    .Y(_05615_),
    .A1(net6604),
    .A2(net5253));
 sg13g2_o21ai_1 _21848_ (.B1(net4803),
    .Y(_05616_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[6] ),
    .A2(net4727));
 sg13g2_a21oi_1 _21849_ (.A1(_05614_),
    .A2(_05615_),
    .Y(_05617_),
    .B1(_05616_));
 sg13g2_o21ai_1 _21850_ (.B1(net4763),
    .Y(_05618_),
    .A1(\fpga_top.cpu_start_adr[6] ),
    .A2(net4638));
 sg13g2_a21oi_1 _21851_ (.A1(_03958_),
    .A2(net4638),
    .Y(_05619_),
    .B1(_05618_));
 sg13g2_nor3_1 _21852_ (.A(net4798),
    .B(net6605),
    .C(_05619_),
    .Y(_05620_));
 sg13g2_o21ai_1 _21853_ (.B1(net4608),
    .Y(_05621_),
    .A1(net1475),
    .A2(net4793));
 sg13g2_o21ai_1 _21854_ (.B1(_05612_),
    .Y(_01949_),
    .A1(_05620_),
    .A2(_05621_));
 sg13g2_nand2_1 _21855_ (.Y(_05622_),
    .A(net2104),
    .B(net4611));
 sg13g2_a21oi_1 _21856_ (.A1(_08071_),
    .A2(net4571),
    .Y(_05623_),
    .B1(net4757));
 sg13g2_o21ai_1 _21857_ (.B1(_05623_),
    .Y(_05624_),
    .A1(_08068_),
    .A2(net4571));
 sg13g2_o21ai_1 _21858_ (.B1(net4775),
    .Y(_05625_),
    .A1(\fpga_top.bus_gather.i_read_adr[7] ),
    .A2(net5253));
 sg13g2_a221oi_1 _21859_ (.B2(_05625_),
    .C1(net4762),
    .B1(_05624_),
    .A1(_06894_),
    .Y(_05626_),
    .A2(net4741));
 sg13g2_o21ai_1 _21860_ (.B1(net4763),
    .Y(_05627_),
    .A1(net5657),
    .A2(net4638));
 sg13g2_a21oi_1 _21861_ (.A1(_03972_),
    .A2(net4638),
    .Y(_05628_),
    .B1(_05627_));
 sg13g2_nor3_1 _21862_ (.A(net4798),
    .B(_05626_),
    .C(_05628_),
    .Y(_05629_));
 sg13g2_o21ai_1 _21863_ (.B1(net4608),
    .Y(_05630_),
    .A1(net1541),
    .A2(net4793));
 sg13g2_o21ai_1 _21864_ (.B1(_05622_),
    .Y(_01950_),
    .A1(_05629_),
    .A2(_05630_));
 sg13g2_nand2_1 _21865_ (.Y(_05631_),
    .A(net2127),
    .B(net4611));
 sg13g2_a21oi_1 _21866_ (.A1(_08126_),
    .A2(net4572),
    .Y(_05632_),
    .B1(net4757));
 sg13g2_o21ai_1 _21867_ (.B1(_05632_),
    .Y(_05633_),
    .A1(_08124_),
    .A2(net4572));
 sg13g2_o21ai_1 _21868_ (.B1(net4775),
    .Y(_05634_),
    .A1(\fpga_top.bus_gather.i_read_adr[8] ),
    .A2(net5254));
 sg13g2_a221oi_1 _21869_ (.B2(_05634_),
    .C1(net4765),
    .B1(_05633_),
    .A1(_06900_),
    .Y(_05635_),
    .A2(net4741));
 sg13g2_o21ai_1 _21870_ (.B1(net4764),
    .Y(_05636_),
    .A1(net5655),
    .A2(net4639));
 sg13g2_a21oi_1 _21871_ (.A1(_03982_),
    .A2(net4639),
    .Y(_05637_),
    .B1(_05636_));
 sg13g2_nor3_1 _21872_ (.A(net4798),
    .B(_05635_),
    .C(_05637_),
    .Y(_05638_));
 sg13g2_o21ai_1 _21873_ (.B1(net4608),
    .Y(_05639_),
    .A1(\fpga_top.cpu_top.execution.csr_array.pc_excep2[8] ),
    .A2(net4792));
 sg13g2_o21ai_1 _21874_ (.B1(_05631_),
    .Y(_01951_),
    .A1(_05638_),
    .A2(_05639_));
 sg13g2_nand2_1 _21875_ (.Y(_05640_),
    .A(net2122),
    .B(net4613));
 sg13g2_nand2_1 _21876_ (.Y(_05641_),
    .A(_08311_),
    .B(net4574));
 sg13g2_a21oi_1 _21877_ (.A1(_08309_),
    .A2(net4561),
    .Y(_05642_),
    .B1(net4758));
 sg13g2_a221oi_1 _21878_ (.B2(_05642_),
    .C1(net4741),
    .B1(_05641_),
    .A1(\fpga_top.bus_gather.i_read_adr[9] ),
    .Y(_05643_),
    .A2(net4776));
 sg13g2_o21ai_1 _21879_ (.B1(net4805),
    .Y(_05644_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[9] ),
    .A2(net4730));
 sg13g2_nor2_1 _21880_ (.A(_05643_),
    .B(_05644_),
    .Y(_05645_));
 sg13g2_o21ai_1 _21881_ (.B1(net4774),
    .Y(_05646_),
    .A1(net5653),
    .A2(net4640));
 sg13g2_a21oi_1 _21882_ (.A1(_03997_),
    .A2(net4640),
    .Y(_05647_),
    .B1(_05646_));
 sg13g2_nor3_1 _21883_ (.A(net4799),
    .B(_05645_),
    .C(_05647_),
    .Y(_05648_));
 sg13g2_o21ai_1 _21884_ (.B1(net4608),
    .Y(_05649_),
    .A1(net1477),
    .A2(net4794));
 sg13g2_o21ai_1 _21885_ (.B1(_05640_),
    .Y(_01952_),
    .A1(_05648_),
    .A2(_05649_));
 sg13g2_nand2_1 _21886_ (.Y(_05650_),
    .A(net2284),
    .B(net4616));
 sg13g2_nand2_1 _21887_ (.Y(_05651_),
    .A(_08010_),
    .B(net4574));
 sg13g2_o21ai_1 _21888_ (.B1(_05651_),
    .Y(_05652_),
    .A1(_08008_),
    .A2(net4574));
 sg13g2_o21ai_1 _21889_ (.B1(net4776),
    .Y(_05653_),
    .A1(\fpga_top.bus_gather.i_read_adr[10] ),
    .A2(net5254));
 sg13g2_o21ai_1 _21890_ (.B1(_05653_),
    .Y(_05654_),
    .A1(net4758),
    .A2(_05652_));
 sg13g2_o21ai_1 _21891_ (.B1(_05654_),
    .Y(_05655_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[10] ),
    .A2(net4731));
 sg13g2_o21ai_1 _21892_ (.B1(net4767),
    .Y(_05656_),
    .A1(\fpga_top.cpu_start_adr[10] ),
    .A2(net4640));
 sg13g2_a21oi_1 _21893_ (.A1(_04007_),
    .A2(net4640),
    .Y(_05657_),
    .B1(_05656_));
 sg13g2_nor2_1 _21894_ (.A(net4799),
    .B(_05657_),
    .Y(_05658_));
 sg13g2_o21ai_1 _21895_ (.B1(_05658_),
    .Y(_05659_),
    .A1(net4766),
    .A2(_05655_));
 sg13g2_o21ai_1 _21896_ (.B1(_05659_),
    .Y(_05660_),
    .A1(net1417),
    .A2(net4794));
 sg13g2_o21ai_1 _21897_ (.B1(_05650_),
    .Y(_01953_),
    .A1(net4613),
    .A2(_05660_));
 sg13g2_nand2_1 _21898_ (.Y(_05661_),
    .A(net1819),
    .B(net4612));
 sg13g2_nor2_1 _21899_ (.A(_08275_),
    .B(net4561),
    .Y(_05662_));
 sg13g2_nor2_1 _21900_ (.A(_08251_),
    .B(net4573),
    .Y(_05663_));
 sg13g2_nor3_1 _21901_ (.A(net4775),
    .B(_05662_),
    .C(_05663_),
    .Y(_05664_));
 sg13g2_a21oi_1 _21902_ (.A1(_06597_),
    .A2(net4757),
    .Y(_05665_),
    .B1(net4765));
 sg13g2_o21ai_1 _21903_ (.B1(_05665_),
    .Y(_05666_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[11] ),
    .A2(net4729));
 sg13g2_o21ai_1 _21904_ (.B1(net4762),
    .Y(_05667_),
    .A1(net5651),
    .A2(net4638));
 sg13g2_a21oi_1 _21905_ (.A1(_04022_),
    .A2(net4638),
    .Y(_05668_),
    .B1(_05667_));
 sg13g2_nor2_1 _21906_ (.A(net4798),
    .B(_05668_),
    .Y(_05669_));
 sg13g2_o21ai_1 _21907_ (.B1(_05669_),
    .Y(_05670_),
    .A1(_05664_),
    .A2(_05666_));
 sg13g2_o21ai_1 _21908_ (.B1(_05670_),
    .Y(_05671_),
    .A1(net1509),
    .A2(net4792));
 sg13g2_o21ai_1 _21909_ (.B1(_05661_),
    .Y(_01954_),
    .A1(net4612),
    .A2(_05671_));
 sg13g2_nand2_1 _21910_ (.Y(_05672_),
    .A(net2084),
    .B(net4613));
 sg13g2_nand2_1 _21911_ (.Y(_05673_),
    .A(_08343_),
    .B(net4574));
 sg13g2_a21oi_1 _21912_ (.A1(_08339_),
    .A2(net4561),
    .Y(_05674_),
    .B1(net4758));
 sg13g2_a221oi_1 _21913_ (.B2(_05674_),
    .C1(net4741),
    .B1(_05673_),
    .A1(\fpga_top.bus_gather.i_read_adr[12] ),
    .Y(_05675_),
    .A2(net4776));
 sg13g2_o21ai_1 _21914_ (.B1(net4805),
    .Y(_05676_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[12] ),
    .A2(net4730));
 sg13g2_nor2_1 _21915_ (.A(_05675_),
    .B(_05676_),
    .Y(_05677_));
 sg13g2_o21ai_1 _21916_ (.B1(net4764),
    .Y(_05678_),
    .A1(\fpga_top.cpu_start_adr[12] ),
    .A2(net4639));
 sg13g2_a21oi_1 _21917_ (.A1(_04035_),
    .A2(net4639),
    .Y(_05679_),
    .B1(_05678_));
 sg13g2_nor3_1 _21918_ (.A(net4799),
    .B(_05677_),
    .C(_05679_),
    .Y(_05680_));
 sg13g2_o21ai_1 _21919_ (.B1(net4608),
    .Y(_05681_),
    .A1(net1531),
    .A2(net4794));
 sg13g2_o21ai_1 _21920_ (.B1(_05672_),
    .Y(_01955_),
    .A1(_05680_),
    .A2(_05681_));
 sg13g2_nand2_1 _21921_ (.Y(_05682_),
    .A(net2103),
    .B(net4613));
 sg13g2_nand2_1 _21922_ (.Y(_05683_),
    .A(_07968_),
    .B(net4574));
 sg13g2_a21oi_1 _21923_ (.A1(_07965_),
    .A2(net4561),
    .Y(_05684_),
    .B1(net4758));
 sg13g2_a221oi_1 _21924_ (.B2(_05684_),
    .C1(net4744),
    .B1(_05683_),
    .A1(\fpga_top.bus_gather.i_read_adr[13] ),
    .Y(_05685_),
    .A2(net4776));
 sg13g2_o21ai_1 _21925_ (.B1(net4807),
    .Y(_05686_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[13] ),
    .A2(net4732));
 sg13g2_nor2_1 _21926_ (.A(_05685_),
    .B(_05686_),
    .Y(_05687_));
 sg13g2_o21ai_1 _21927_ (.B1(net4767),
    .Y(_05688_),
    .A1(\fpga_top.cpu_start_adr[13] ),
    .A2(net4640));
 sg13g2_a21oi_1 _21928_ (.A1(_04046_),
    .A2(net4641),
    .Y(_05689_),
    .B1(_05688_));
 sg13g2_nor3_1 _21929_ (.A(net4799),
    .B(_05687_),
    .C(_05689_),
    .Y(_05690_));
 sg13g2_o21ai_1 _21930_ (.B1(net4608),
    .Y(_05691_),
    .A1(net1495),
    .A2(net4794));
 sg13g2_o21ai_1 _21931_ (.B1(_05682_),
    .Y(_01956_),
    .A1(_05690_),
    .A2(_05691_));
 sg13g2_nand2_1 _21932_ (.Y(_05692_),
    .A(net1979),
    .B(net4613));
 sg13g2_mux2_1 _21933_ (.A0(_07939_),
    .A1(_07941_),
    .S(net4574),
    .X(_05693_));
 sg13g2_o21ai_1 _21934_ (.B1(net4776),
    .Y(_05694_),
    .A1(\fpga_top.bus_gather.i_read_adr[14] ),
    .A2(net5254));
 sg13g2_o21ai_1 _21935_ (.B1(_05694_),
    .Y(_05695_),
    .A1(net4758),
    .A2(_05693_));
 sg13g2_o21ai_1 _21936_ (.B1(_05695_),
    .Y(_05696_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[14] ),
    .A2(net4731));
 sg13g2_o21ai_1 _21937_ (.B1(net4766),
    .Y(_05697_),
    .A1(net5650),
    .A2(net4640));
 sg13g2_a21oi_1 _21938_ (.A1(_04060_),
    .A2(net4640),
    .Y(_05698_),
    .B1(_05697_));
 sg13g2_nor2_1 _21939_ (.A(net4799),
    .B(_05698_),
    .Y(_05699_));
 sg13g2_o21ai_1 _21940_ (.B1(_05699_),
    .Y(_05700_),
    .A1(net4766),
    .A2(_05696_));
 sg13g2_o21ai_1 _21941_ (.B1(_05700_),
    .Y(_05701_),
    .A1(net1550),
    .A2(net4794));
 sg13g2_o21ai_1 _21942_ (.B1(_05692_),
    .Y(_01957_),
    .A1(net4613),
    .A2(_05701_));
 sg13g2_nand2_1 _21943_ (.Y(_05702_),
    .A(net1817),
    .B(net4617));
 sg13g2_a21oi_1 _21944_ (.A1(_08546_),
    .A2(net4574),
    .Y(_05703_),
    .B1(net4758));
 sg13g2_o21ai_1 _21945_ (.B1(_05703_),
    .Y(_05704_),
    .A1(_08530_),
    .A2(_04964_));
 sg13g2_o21ai_1 _21946_ (.B1(net4776),
    .Y(_05705_),
    .A1(\fpga_top.bus_gather.i_read_adr[15] ),
    .A2(net5254));
 sg13g2_o21ai_1 _21947_ (.B1(net4807),
    .Y(_05706_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[15] ),
    .A2(net4732));
 sg13g2_a21oi_1 _21948_ (.A1(_05704_),
    .A2(_05705_),
    .Y(_05707_),
    .B1(_05706_));
 sg13g2_o21ai_1 _21949_ (.B1(net4767),
    .Y(_05708_),
    .A1(\fpga_top.cpu_start_adr[15] ),
    .A2(net4642));
 sg13g2_a21oi_1 _21950_ (.A1(_04069_),
    .A2(net4642),
    .Y(_05709_),
    .B1(_05708_));
 sg13g2_nor3_1 _21951_ (.A(net4799),
    .B(_05707_),
    .C(_05709_),
    .Y(_05710_));
 sg13g2_o21ai_1 _21952_ (.B1(_05570_),
    .Y(_05711_),
    .A1(net1446),
    .A2(net4794));
 sg13g2_o21ai_1 _21953_ (.B1(_05702_),
    .Y(_01958_),
    .A1(_05710_),
    .A2(_05711_));
 sg13g2_nand2_1 _21954_ (.Y(_05712_),
    .A(net3348),
    .B(net4616));
 sg13g2_nand2_1 _21955_ (.Y(_05713_),
    .A(_08035_),
    .B(net4579));
 sg13g2_a21oi_1 _21956_ (.A1(_08032_),
    .A2(net4562),
    .Y(_05714_),
    .B1(net4761));
 sg13g2_a221oi_1 _21957_ (.B2(_05714_),
    .C1(net4742),
    .B1(_05713_),
    .A1(net5593),
    .Y(_05715_),
    .A2(net4779));
 sg13g2_o21ai_1 _21958_ (.B1(net4807),
    .Y(_05716_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[16] ),
    .A2(net4733));
 sg13g2_nor2_1 _21959_ (.A(_05715_),
    .B(_05716_),
    .Y(_05717_));
 sg13g2_nor2b_1 _21960_ (.A(_04081_),
    .B_N(net4647),
    .Y(_05718_));
 sg13g2_o21ai_1 _21961_ (.B1(net4768),
    .Y(_05719_),
    .A1(net5649),
    .A2(net4642));
 sg13g2_o21ai_1 _21962_ (.B1(net4797),
    .Y(_05720_),
    .A1(_05718_),
    .A2(_05719_));
 sg13g2_nor2_1 _21963_ (.A(_05717_),
    .B(_05720_),
    .Y(_05721_));
 sg13g2_o21ai_1 _21964_ (.B1(net4610),
    .Y(_05722_),
    .A1(\fpga_top.cpu_top.execution.csr_array.pc_excep2[16] ),
    .A2(net4797));
 sg13g2_o21ai_1 _21965_ (.B1(_05712_),
    .Y(_01959_),
    .A1(_05721_),
    .A2(_05722_));
 sg13g2_nand2_1 _21966_ (.Y(_05723_),
    .A(net3706),
    .B(net4614));
 sg13g2_a21oi_1 _21967_ (.A1(_08375_),
    .A2(net4579),
    .Y(_05724_),
    .B1(net4779));
 sg13g2_o21ai_1 _21968_ (.B1(_05724_),
    .Y(_05725_),
    .A1(_08371_),
    .A2(net4579));
 sg13g2_a221oi_1 _21969_ (.B2(_06611_),
    .C1(net4769),
    .B1(net4760),
    .A1(_06911_),
    .Y(_05726_),
    .A2(net4743));
 sg13g2_o21ai_1 _21970_ (.B1(net4773),
    .Y(_05727_),
    .A1(net5648),
    .A2(net4646));
 sg13g2_a21oi_1 _21971_ (.A1(_04091_),
    .A2(net4646),
    .Y(_05728_),
    .B1(_05727_));
 sg13g2_or2_1 _21972_ (.X(_05729_),
    .B(_05728_),
    .A(net4801));
 sg13g2_a21o_1 _21973_ (.A2(_05726_),
    .A1(_05725_),
    .B1(_05729_),
    .X(_05730_));
 sg13g2_o21ai_1 _21974_ (.B1(_05730_),
    .Y(_05731_),
    .A1(net1440),
    .A2(net4795));
 sg13g2_o21ai_1 _21975_ (.B1(_05723_),
    .Y(_01960_),
    .A1(net4614),
    .A2(_05731_));
 sg13g2_nand2_1 _21976_ (.Y(_05732_),
    .A(net2489),
    .B(net4616));
 sg13g2_nand2_1 _21977_ (.Y(_05733_),
    .A(_08523_),
    .B(net4579));
 sg13g2_a21oi_1 _21978_ (.A1(_08520_),
    .A2(net4562),
    .Y(_05734_),
    .B1(net4761));
 sg13g2_a221oi_1 _21979_ (.B2(_05734_),
    .C1(net4742),
    .B1(_05733_),
    .A1(\fpga_top.bus_gather.i_read_adr[18] ),
    .Y(_05735_),
    .A2(net4779));
 sg13g2_o21ai_1 _21980_ (.B1(net4806),
    .Y(_05736_),
    .A1(net6611),
    .A2(net4734));
 sg13g2_nor2_1 _21981_ (.A(_05735_),
    .B(_05736_),
    .Y(_05737_));
 sg13g2_o21ai_1 _21982_ (.B1(net4768),
    .Y(_05738_),
    .A1(\fpga_top.cpu_start_adr[18] ),
    .A2(net4642));
 sg13g2_a21oi_1 _21983_ (.A1(_04099_),
    .A2(net4647),
    .Y(_05739_),
    .B1(_05738_));
 sg13g2_nor3_1 _21984_ (.A(net4802),
    .B(_05737_),
    .C(_05739_),
    .Y(_05740_));
 sg13g2_o21ai_1 _21985_ (.B1(net4610),
    .Y(_05741_),
    .A1(net1524),
    .A2(net4797));
 sg13g2_o21ai_1 _21986_ (.B1(_05732_),
    .Y(_01961_),
    .A1(_05740_),
    .A2(_05741_));
 sg13g2_nand2_1 _21987_ (.Y(_05742_),
    .A(net3558),
    .B(net4614));
 sg13g2_a21oi_1 _21988_ (.A1(_08402_),
    .A2(net4577),
    .Y(_05743_),
    .B1(net4759));
 sg13g2_o21ai_1 _21989_ (.B1(_05743_),
    .Y(_05744_),
    .A1(_08381_),
    .A2(net4577));
 sg13g2_o21ai_1 _21990_ (.B1(net4778),
    .Y(_05745_),
    .A1(\fpga_top.bus_gather.i_read_adr[19] ),
    .A2(net5255));
 sg13g2_o21ai_1 _21991_ (.B1(net4806),
    .Y(_05746_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[19] ),
    .A2(net4739));
 sg13g2_a21oi_1 _21992_ (.A1(_05744_),
    .A2(_05745_),
    .Y(_05747_),
    .B1(_05746_));
 sg13g2_o21ai_1 _21993_ (.B1(net4771),
    .Y(_05748_),
    .A1(\fpga_top.cpu_start_adr[19] ),
    .A2(net4644));
 sg13g2_a21oi_1 _21994_ (.A1(_04109_),
    .A2(net4643),
    .Y(_05749_),
    .B1(_05748_));
 sg13g2_nor3_1 _21995_ (.A(net4800),
    .B(_05747_),
    .C(_05749_),
    .Y(_05750_));
 sg13g2_o21ai_1 _21996_ (.B1(net4609),
    .Y(_05751_),
    .A1(net1582),
    .A2(net4795));
 sg13g2_o21ai_1 _21997_ (.B1(_05742_),
    .Y(_01962_),
    .A1(_05750_),
    .A2(_05751_));
 sg13g2_nand2_1 _21998_ (.Y(_05752_),
    .A(net2210),
    .B(net4616));
 sg13g2_nand2_1 _21999_ (.Y(_05753_),
    .A(_08424_),
    .B(net4577));
 sg13g2_a21oi_1 _22000_ (.A1(_08421_),
    .A2(net4561),
    .Y(_05754_),
    .B1(net4759));
 sg13g2_a221oi_1 _22001_ (.B2(_05754_),
    .C1(net4743),
    .B1(_05753_),
    .A1(\fpga_top.bus_gather.i_read_adr[20] ),
    .Y(_05755_),
    .A2(net4778));
 sg13g2_o21ai_1 _22002_ (.B1(net4807),
    .Y(_05756_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[20] ),
    .A2(net4739));
 sg13g2_nor2_1 _22003_ (.A(_05755_),
    .B(_05756_),
    .Y(_05757_));
 sg13g2_o21ai_1 _22004_ (.B1(net4773),
    .Y(_05758_),
    .A1(\fpga_top.cpu_start_adr[20] ),
    .A2(net4646));
 sg13g2_a21oi_1 _22005_ (.A1(_04122_),
    .A2(net4646),
    .Y(_05759_),
    .B1(_05758_));
 sg13g2_nor3_1 _22006_ (.A(net4801),
    .B(_05757_),
    .C(_05759_),
    .Y(_05760_));
 sg13g2_o21ai_1 _22007_ (.B1(net4610),
    .Y(_05761_),
    .A1(net1512),
    .A2(net4797));
 sg13g2_o21ai_1 _22008_ (.B1(_05752_),
    .Y(_01963_),
    .A1(_05760_),
    .A2(_05761_));
 sg13g2_nand2_1 _22009_ (.Y(_05762_),
    .A(net3749),
    .B(net4615));
 sg13g2_nand2_1 _22010_ (.Y(_05763_),
    .A(_07864_),
    .B(net4576));
 sg13g2_a21oi_1 _22011_ (.A1(_07861_),
    .A2(net4561),
    .Y(_05764_),
    .B1(net4759));
 sg13g2_a221oi_1 _22012_ (.B2(_05764_),
    .C1(net4742),
    .B1(_05763_),
    .A1(\fpga_top.bus_gather.i_read_adr[21] ),
    .Y(_05765_),
    .A2(net4777));
 sg13g2_o21ai_1 _22013_ (.B1(net4806),
    .Y(_05766_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ),
    .A2(net4738));
 sg13g2_nor2_1 _22014_ (.A(_05765_),
    .B(_05766_),
    .Y(_05767_));
 sg13g2_o21ai_1 _22015_ (.B1(net4770),
    .Y(_05768_),
    .A1(net5645),
    .A2(net4644));
 sg13g2_a21oi_1 _22016_ (.A1(_04132_),
    .A2(net4644),
    .Y(_05769_),
    .B1(_05768_));
 sg13g2_nor3_1 _22017_ (.A(net4800),
    .B(_05767_),
    .C(_05769_),
    .Y(_05770_));
 sg13g2_o21ai_1 _22018_ (.B1(net4610),
    .Y(_05771_),
    .A1(net1506),
    .A2(net4796));
 sg13g2_o21ai_1 _22019_ (.B1(_05762_),
    .Y(_01964_),
    .A1(_05770_),
    .A2(_05771_));
 sg13g2_nand2_1 _22020_ (.Y(_05772_),
    .A(net3337),
    .B(net4614));
 sg13g2_a21oi_1 _22021_ (.A1(_07835_),
    .A2(net4575),
    .Y(_05773_),
    .B1(net4759));
 sg13g2_o21ai_1 _22022_ (.B1(_05773_),
    .Y(_05774_),
    .A1(_07832_),
    .A2(net4576));
 sg13g2_o21ai_1 _22023_ (.B1(net4777),
    .Y(_05775_),
    .A1(net5592),
    .A2(net5255));
 sg13g2_o21ai_1 _22024_ (.B1(net4807),
    .Y(_05776_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[22] ),
    .A2(net4739));
 sg13g2_a21oi_1 _22025_ (.A1(_05774_),
    .A2(_05775_),
    .Y(_05777_),
    .B1(_05776_));
 sg13g2_o21ai_1 _22026_ (.B1(net4772),
    .Y(_05778_),
    .A1(net5643),
    .A2(net4646));
 sg13g2_a21oi_1 _22027_ (.A1(_04144_),
    .A2(net4645),
    .Y(_05779_),
    .B1(_05778_));
 sg13g2_nor3_1 _22028_ (.A(net4800),
    .B(_05777_),
    .C(_05779_),
    .Y(_05780_));
 sg13g2_o21ai_1 _22029_ (.B1(net4610),
    .Y(_05781_),
    .A1(\fpga_top.cpu_top.execution.csr_array.pc_excep2[22] ),
    .A2(net4796));
 sg13g2_o21ai_1 _22030_ (.B1(_05772_),
    .Y(_01965_),
    .A1(_05780_),
    .A2(_05781_));
 sg13g2_nand2_1 _22031_ (.Y(_05782_),
    .A(net2789),
    .B(net4615));
 sg13g2_a21oi_1 _22032_ (.A1(_08472_),
    .A2(net4576),
    .Y(_05783_),
    .B1(net4759));
 sg13g2_o21ai_1 _22033_ (.B1(_05783_),
    .Y(_05784_),
    .A1(_08455_),
    .A2(net4576));
 sg13g2_o21ai_1 _22034_ (.B1(net4777),
    .Y(_05785_),
    .A1(\fpga_top.bus_gather.i_read_adr[23] ),
    .A2(net5255));
 sg13g2_o21ai_1 _22035_ (.B1(net4806),
    .Y(_05786_),
    .A1(net6613),
    .A2(net4739));
 sg13g2_a21oi_1 _22036_ (.A1(_05784_),
    .A2(_05785_),
    .Y(_05787_),
    .B1(_05786_));
 sg13g2_o21ai_1 _22037_ (.B1(net4771),
    .Y(_05788_),
    .A1(net5642),
    .A2(net4643));
 sg13g2_a21oi_1 _22038_ (.A1(_04154_),
    .A2(net4644),
    .Y(_05789_),
    .B1(_05788_));
 sg13g2_nor3_1 _22039_ (.A(net4801),
    .B(_05787_),
    .C(_05789_),
    .Y(_05790_));
 sg13g2_o21ai_1 _22040_ (.B1(net4609),
    .Y(_05791_),
    .A1(net1555),
    .A2(net4795));
 sg13g2_o21ai_1 _22041_ (.B1(_05782_),
    .Y(_01966_),
    .A1(_05790_),
    .A2(_05791_));
 sg13g2_nand2_1 _22042_ (.Y(_05792_),
    .A(net2329),
    .B(net4615));
 sg13g2_nand2_1 _22043_ (.Y(_05793_),
    .A(_07903_),
    .B(net4578));
 sg13g2_a21oi_1 _22044_ (.A1(_07901_),
    .A2(net4562),
    .Y(_05794_),
    .B1(net4760));
 sg13g2_a221oi_1 _22045_ (.B2(_05794_),
    .C1(net4742),
    .B1(_05793_),
    .A1(\fpga_top.bus_gather.i_read_adr[24] ),
    .Y(_05795_),
    .A2(net4778));
 sg13g2_o21ai_1 _22046_ (.B1(net4806),
    .Y(_05796_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[24] ),
    .A2(net4733));
 sg13g2_nor2_1 _22047_ (.A(_05795_),
    .B(_05796_),
    .Y(_05797_));
 sg13g2_o21ai_1 _22048_ (.B1(net4769),
    .Y(_05798_),
    .A1(\fpga_top.cpu_start_adr[24] ),
    .A2(net4642));
 sg13g2_a21oi_1 _22049_ (.A1(_04166_),
    .A2(net4646),
    .Y(_05799_),
    .B1(_05798_));
 sg13g2_nor3_1 _22050_ (.A(net4801),
    .B(_05797_),
    .C(_05799_),
    .Y(_05800_));
 sg13g2_o21ai_1 _22051_ (.B1(net4609),
    .Y(_05801_),
    .A1(net1546),
    .A2(net4796));
 sg13g2_o21ai_1 _22052_ (.B1(_05792_),
    .Y(_01967_),
    .A1(_05800_),
    .A2(_05801_));
 sg13g2_nand2_1 _22053_ (.Y(_05802_),
    .A(net1996),
    .B(net4616));
 sg13g2_o21ai_1 _22054_ (.B1(net4806),
    .Y(_05803_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[25] ),
    .A2(net4733));
 sg13g2_a21oi_1 _22055_ (.A1(_08497_),
    .A2(net4578),
    .Y(_05804_),
    .B1(net4760));
 sg13g2_a221oi_1 _22056_ (.B2(_05804_),
    .C1(net4742),
    .B1(_05181_),
    .A1(\fpga_top.bus_gather.i_read_adr[25] ),
    .Y(_05805_),
    .A2(net4778));
 sg13g2_o21ai_1 _22057_ (.B1(net4768),
    .Y(_05806_),
    .A1(\fpga_top.cpu_start_adr[25] ),
    .A2(net4642));
 sg13g2_a21oi_1 _22058_ (.A1(_04176_),
    .A2(net4642),
    .Y(_05807_),
    .B1(_05806_));
 sg13g2_nor2_1 _22059_ (.A(net4802),
    .B(_05807_),
    .Y(_05808_));
 sg13g2_o21ai_1 _22060_ (.B1(_05808_),
    .Y(_05809_),
    .A1(_05803_),
    .A2(_05805_));
 sg13g2_o21ai_1 _22061_ (.B1(_05809_),
    .Y(_05810_),
    .A1(net1944),
    .A2(net4797));
 sg13g2_o21ai_1 _22062_ (.B1(_05802_),
    .Y(_01968_),
    .A1(net4616),
    .A2(_05810_));
 sg13g2_nand2_1 _22063_ (.Y(_05811_),
    .A(net2312),
    .B(net4614));
 sg13g2_a21oi_1 _22064_ (.A1(_08596_),
    .A2(net4575),
    .Y(_05812_),
    .B1(net4759));
 sg13g2_o21ai_1 _22065_ (.B1(_05812_),
    .Y(_05813_),
    .A1(_08593_),
    .A2(net4575));
 sg13g2_o21ai_1 _22066_ (.B1(net4778),
    .Y(_05814_),
    .A1(\fpga_top.bus_gather.i_read_adr[26] ),
    .A2(net5255));
 sg13g2_o21ai_1 _22067_ (.B1(net4806),
    .Y(_05815_),
    .A1(net6596),
    .A2(net4738));
 sg13g2_a21oi_1 _22068_ (.A1(_05813_),
    .A2(_05814_),
    .Y(_05816_),
    .B1(_05815_));
 sg13g2_o21ai_1 _22069_ (.B1(net4770),
    .Y(_05817_),
    .A1(\fpga_top.cpu_start_adr[26] ),
    .A2(net4643));
 sg13g2_a21oi_1 _22070_ (.A1(_04186_),
    .A2(net4643),
    .Y(_05818_),
    .B1(_05817_));
 sg13g2_nor3_1 _22071_ (.A(net4800),
    .B(_05816_),
    .C(_05818_),
    .Y(_05819_));
 sg13g2_o21ai_1 _22072_ (.B1(net4609),
    .Y(_05820_),
    .A1(net1600),
    .A2(net4795));
 sg13g2_o21ai_1 _22073_ (.B1(_05811_),
    .Y(_01969_),
    .A1(_05819_),
    .A2(_05820_));
 sg13g2_nand2_1 _22074_ (.Y(_05821_),
    .A(net2154),
    .B(net4614));
 sg13g2_a21oi_1 _22075_ (.A1(_08450_),
    .A2(net4575),
    .Y(_05822_),
    .B1(net4759));
 sg13g2_o21ai_1 _22076_ (.B1(_05822_),
    .Y(_05823_),
    .A1(_08432_),
    .A2(net4575));
 sg13g2_o21ai_1 _22077_ (.B1(net4777),
    .Y(_05824_),
    .A1(\fpga_top.bus_gather.i_read_adr[27] ),
    .A2(net5255));
 sg13g2_a221oi_1 _22078_ (.B2(_05824_),
    .C1(net4772),
    .B1(_05823_),
    .A1(_06919_),
    .Y(_05825_),
    .A2(net4743));
 sg13g2_o21ai_1 _22079_ (.B1(net4771),
    .Y(_05826_),
    .A1(net5641),
    .A2(net4643));
 sg13g2_a21oi_1 _22080_ (.A1(_04197_),
    .A2(net4643),
    .Y(_05827_),
    .B1(_05826_));
 sg13g2_nor3_1 _22081_ (.A(net4800),
    .B(_05825_),
    .C(_05827_),
    .Y(_05828_));
 sg13g2_o21ai_1 _22082_ (.B1(net4609),
    .Y(_05829_),
    .A1(net1591),
    .A2(net4795));
 sg13g2_o21ai_1 _22083_ (.B1(_05821_),
    .Y(_01970_),
    .A1(_05828_),
    .A2(_05829_));
 sg13g2_nand2_1 _22084_ (.Y(_05830_),
    .A(net2048),
    .B(net4615));
 sg13g2_a21oi_1 _22085_ (.A1(_08572_),
    .A2(net4575),
    .Y(_05831_),
    .B1(net4760));
 sg13g2_o21ai_1 _22086_ (.B1(_05831_),
    .Y(_05832_),
    .A1(_08569_),
    .A2(net4576));
 sg13g2_o21ai_1 _22087_ (.B1(net4777),
    .Y(_05833_),
    .A1(\fpga_top.bus_gather.i_read_adr[28] ),
    .A2(net5255));
 sg13g2_o21ai_1 _22088_ (.B1(net4806),
    .Y(_05834_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[28] ),
    .A2(net4738));
 sg13g2_a21oi_1 _22089_ (.A1(_05832_),
    .A2(_05833_),
    .Y(_05835_),
    .B1(_05834_));
 sg13g2_o21ai_1 _22090_ (.B1(net4770),
    .Y(_05836_),
    .A1(net5639),
    .A2(net4645));
 sg13g2_a21oi_1 _22091_ (.A1(_04210_),
    .A2(net4645),
    .Y(_05837_),
    .B1(_05836_));
 sg13g2_nor3_1 _22092_ (.A(net4800),
    .B(_05835_),
    .C(_05837_),
    .Y(_05838_));
 sg13g2_o21ai_1 _22093_ (.B1(net4609),
    .Y(_05839_),
    .A1(\fpga_top.cpu_top.execution.csr_array.pc_excep2[28] ),
    .A2(net4795));
 sg13g2_o21ai_1 _22094_ (.B1(_05830_),
    .Y(_01971_),
    .A1(_05838_),
    .A2(_05839_));
 sg13g2_nand2_1 _22095_ (.Y(_05840_),
    .A(net1792),
    .B(net4614));
 sg13g2_a21oi_1 _22096_ (.A1(_07796_),
    .A2(net4575),
    .Y(_05841_),
    .B1(net4759));
 sg13g2_o21ai_1 _22097_ (.B1(_05841_),
    .Y(_05842_),
    .A1(_07752_),
    .A2(net4575));
 sg13g2_o21ai_1 _22098_ (.B1(net4777),
    .Y(_05843_),
    .A1(\fpga_top.bus_gather.i_read_adr[29] ),
    .A2(net5255));
 sg13g2_o21ai_1 _22099_ (.B1(net4807),
    .Y(_05844_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[29] ),
    .A2(net4739));
 sg13g2_a21oi_1 _22100_ (.A1(_05842_),
    .A2(_05843_),
    .Y(_05845_),
    .B1(_05844_));
 sg13g2_o21ai_1 _22101_ (.B1(net4770),
    .Y(_05846_),
    .A1(\fpga_top.cpu_start_adr[29] ),
    .A2(net4643));
 sg13g2_a21oi_1 _22102_ (.A1(_04219_),
    .A2(net4643),
    .Y(_05847_),
    .B1(_05846_));
 sg13g2_nor3_1 _22103_ (.A(net4800),
    .B(_05845_),
    .C(_05847_),
    .Y(_05848_));
 sg13g2_o21ai_1 _22104_ (.B1(net4609),
    .Y(_05849_),
    .A1(\fpga_top.cpu_top.execution.csr_array.pc_excep2[29] ),
    .A2(net4795));
 sg13g2_o21ai_1 _22105_ (.B1(_05840_),
    .Y(_01972_),
    .A1(_05848_),
    .A2(_05849_));
 sg13g2_nand2_1 _22106_ (.Y(_05850_),
    .A(net2936),
    .B(net4614));
 sg13g2_mux2_1 _22107_ (.A0(_07676_),
    .A1(_07746_),
    .S(net4578),
    .X(_05851_));
 sg13g2_o21ai_1 _22108_ (.B1(net4778),
    .Y(_05852_),
    .A1(\fpga_top.bus_gather.i_read_adr[30] ),
    .A2(net5256));
 sg13g2_o21ai_1 _22109_ (.B1(_05852_),
    .Y(_05853_),
    .A1(net4760),
    .A2(_05851_));
 sg13g2_o21ai_1 _22110_ (.B1(_05853_),
    .Y(_05854_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[30] ),
    .A2(net4739));
 sg13g2_nor2_1 _22111_ (.A(net4769),
    .B(_05854_),
    .Y(_05855_));
 sg13g2_o21ai_1 _22112_ (.B1(net4769),
    .Y(_05856_),
    .A1(net5636),
    .A2(net4646));
 sg13g2_a21oi_1 _22113_ (.A1(_04231_),
    .A2(net4646),
    .Y(_05857_),
    .B1(_05856_));
 sg13g2_nor3_1 _22114_ (.A(net4800),
    .B(_05855_),
    .C(_05857_),
    .Y(_05858_));
 sg13g2_o21ai_1 _22115_ (.B1(net4609),
    .Y(_05859_),
    .A1(net1676),
    .A2(net4795));
 sg13g2_o21ai_1 _22116_ (.B1(_05850_),
    .Y(_01973_),
    .A1(_05858_),
    .A2(_05859_));
 sg13g2_nand2_1 _22117_ (.Y(_05860_),
    .A(net2010),
    .B(net4613));
 sg13g2_nor2_1 _22118_ (.A(_07287_),
    .B(net4579),
    .Y(_05861_));
 sg13g2_nor2_1 _22119_ (.A(_07671_),
    .B(net4562),
    .Y(_05862_));
 sg13g2_nor3_1 _22120_ (.A(net4779),
    .B(_05861_),
    .C(_05862_),
    .Y(_05863_));
 sg13g2_a21oi_1 _22121_ (.A1(_06646_),
    .A2(net4761),
    .Y(_05864_),
    .B1(net4767));
 sg13g2_o21ai_1 _22122_ (.B1(_05864_),
    .Y(_05865_),
    .A1(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[31] ),
    .A2(net4733));
 sg13g2_o21ai_1 _22123_ (.B1(net4767),
    .Y(_05866_),
    .A1(\fpga_top.cpu_start_adr[31] ),
    .A2(net4640));
 sg13g2_a21oi_1 _22124_ (.A1(_04244_),
    .A2(net4642),
    .Y(_05867_),
    .B1(_05866_));
 sg13g2_nor2_1 _22125_ (.A(net4802),
    .B(_05867_),
    .Y(_05868_));
 sg13g2_o21ai_1 _22126_ (.B1(_05868_),
    .Y(_05869_),
    .A1(_05863_),
    .A2(_05865_));
 sg13g2_o21ai_1 _22127_ (.B1(_05869_),
    .Y(_05870_),
    .A1(net1438),
    .A2(net4794));
 sg13g2_o21ai_1 _22128_ (.B1(_05860_),
    .Y(_01974_),
    .A1(net4613),
    .A2(_05870_));
 sg13g2_nor2_1 _22129_ (.A(net3770),
    .B(_05352_),
    .Y(_05871_));
 sg13g2_nand2b_1 _22130_ (.Y(_05872_),
    .B(_04021_),
    .A_N(_05334_));
 sg13g2_nand3_1 _22131_ (.B(net4658),
    .C(_05330_),
    .A(net4828),
    .Y(_05873_));
 sg13g2_a21oi_1 _22132_ (.A1(net5651),
    .A2(_05334_),
    .Y(_05874_),
    .B1(_05873_));
 sg13g2_a21oi_1 _22133_ (.A1(_05872_),
    .A2(_05874_),
    .Y(_01975_),
    .B1(_05871_));
 sg13g2_a21oi_1 _22134_ (.A1(\fpga_top.cpu_start_adr[12] ),
    .A2(_05334_),
    .Y(_05875_),
    .B1(_05873_));
 sg13g2_o21ai_1 _22135_ (.B1(_05875_),
    .Y(_05876_),
    .A1(_04035_),
    .A2(_05334_));
 sg13g2_o21ai_1 _22136_ (.B1(_05876_),
    .Y(_05877_),
    .A1(net6259),
    .A2(_05352_));
 sg13g2_inv_1 _22137_ (.Y(_01976_),
    .A(net6260));
 sg13g2_nor3_2 _22138_ (.A(_03819_),
    .B(_03832_),
    .C(_03849_),
    .Y(_05878_));
 sg13g2_nand2_1 _22139_ (.Y(_05879_),
    .A(net4828),
    .B(net4665));
 sg13g2_nor3_1 _22140_ (.A(_03867_),
    .B(_05545_),
    .C(net4601),
    .Y(_05880_));
 sg13g2_a21o_1 _22141_ (.A2(net4601),
    .A1(net2147),
    .B1(_05880_),
    .X(_01977_));
 sg13g2_nand2_1 _22142_ (.Y(_05881_),
    .A(net1554),
    .B(net4599));
 sg13g2_o21ai_1 _22143_ (.B1(_05881_),
    .Y(_01978_),
    .A1(_03882_),
    .A2(net4599));
 sg13g2_nor2_1 _22144_ (.A(net1990),
    .B(net4636),
    .Y(_05882_));
 sg13g2_nor3_2 _22145_ (.A(_03819_),
    .B(net5135),
    .C(_03849_),
    .Y(_05883_));
 sg13g2_nand2_2 _22146_ (.Y(_05884_),
    .A(net5047),
    .B(net4665));
 sg13g2_a21oi_1 _22147_ (.A1(_03899_),
    .A2(net4636),
    .Y(_01979_),
    .B1(_05882_));
 sg13g2_nand2_1 _22148_ (.Y(_05885_),
    .A(net1505),
    .B(net4599));
 sg13g2_o21ai_1 _22149_ (.B1(_03947_),
    .Y(_05886_),
    .A1(_03945_),
    .A2(_05884_));
 sg13g2_o21ai_1 _22150_ (.B1(_05885_),
    .Y(_01980_),
    .A1(net4600),
    .A2(_05886_));
 sg13g2_nand2_1 _22151_ (.Y(_05887_),
    .A(net5048),
    .B(_05383_));
 sg13g2_nor2_1 _22152_ (.A(net5661),
    .B(net5048),
    .Y(_05888_));
 sg13g2_nor2_1 _22153_ (.A(net4601),
    .B(_05888_),
    .Y(_05889_));
 sg13g2_a22oi_1 _22154_ (.Y(_05890_),
    .B1(_05887_),
    .B2(_05889_),
    .A2(net4601),
    .A1(net2893));
 sg13g2_inv_1 _22155_ (.Y(_01981_),
    .A(_05890_));
 sg13g2_nor2_2 _22156_ (.A(net5659),
    .B(net5047),
    .Y(_05891_));
 sg13g2_nor2_2 _22157_ (.A(net5137),
    .B(_05390_),
    .Y(_05892_));
 sg13g2_nor3_1 _22158_ (.A(net4600),
    .B(_05891_),
    .C(_05892_),
    .Y(_05893_));
 sg13g2_a21o_1 _22159_ (.A2(net4600),
    .A1(net2076),
    .B1(_05893_),
    .X(_01982_));
 sg13g2_o21ai_1 _22160_ (.B1(_03959_),
    .Y(_05894_),
    .A1(_03957_),
    .A2(_05884_));
 sg13g2_nor2_1 _22161_ (.A(net1643),
    .B(net4636),
    .Y(_05895_));
 sg13g2_a21oi_1 _22162_ (.A1(net4636),
    .A2(_05894_),
    .Y(_01983_),
    .B1(_05895_));
 sg13g2_nand2_1 _22163_ (.Y(_05896_),
    .A(net1584),
    .B(net4599));
 sg13g2_nand2_1 _22164_ (.Y(_05897_),
    .A(_06791_),
    .B(net5134));
 sg13g2_o21ai_1 _22165_ (.B1(_05897_),
    .Y(_05898_),
    .A1(_03971_),
    .A2(_05884_));
 sg13g2_o21ai_1 _22166_ (.B1(_05896_),
    .Y(_01984_),
    .A1(net4600),
    .A2(_05898_));
 sg13g2_nand3_1 _22167_ (.B(_03984_),
    .C(net4636),
    .A(_03983_),
    .Y(_05899_));
 sg13g2_o21ai_1 _22168_ (.B1(_05899_),
    .Y(_01985_),
    .A1(_06896_),
    .A2(net4636));
 sg13g2_nand2_1 _22169_ (.Y(_05900_),
    .A(net1552),
    .B(net4602));
 sg13g2_o21ai_1 _22170_ (.B1(net4637),
    .Y(_05901_),
    .A1(\fpga_top.cpu_start_adr[9] ),
    .A2(net5055));
 sg13g2_o21ai_1 _22171_ (.B1(_05900_),
    .Y(_01986_),
    .A1(_03999_),
    .A2(_05901_));
 sg13g2_nor3_1 _22172_ (.A(_04008_),
    .B(_04009_),
    .C(net4605),
    .Y(_05902_));
 sg13g2_a21o_1 _22173_ (.A2(net4603),
    .A1(net1988),
    .B1(_05902_),
    .X(_01987_));
 sg13g2_nand2_1 _22174_ (.Y(_05903_),
    .A(net1741),
    .B(net4599));
 sg13g2_nand2_1 _22175_ (.Y(_05904_),
    .A(_06793_),
    .B(net5135));
 sg13g2_o21ai_1 _22176_ (.B1(_05904_),
    .Y(_05905_),
    .A1(_04021_),
    .A2(_05884_));
 sg13g2_o21ai_1 _22177_ (.B1(_05903_),
    .Y(_01988_),
    .A1(net4599),
    .A2(_05905_));
 sg13g2_a221oi_1 _22178_ (.B2(net4635),
    .C1(net4599),
    .B1(_04035_),
    .A1(net5376),
    .Y(_05906_),
    .A2(net5136));
 sg13g2_a21o_1 _22179_ (.A2(net4599),
    .A1(net2068),
    .B1(_05906_),
    .X(_01989_));
 sg13g2_a221oi_1 _22180_ (.B2(net4635),
    .C1(net4601),
    .B1(_04046_),
    .A1(net5374),
    .Y(_05907_),
    .A2(net5140));
 sg13g2_a21o_1 _22181_ (.A2(net4607),
    .A1(net2050),
    .B1(_05907_),
    .X(_01990_));
 sg13g2_nand2_1 _22182_ (.Y(_05908_),
    .A(net1540),
    .B(net4601));
 sg13g2_o21ai_1 _22183_ (.B1(net4637),
    .Y(_05909_),
    .A1(net5650),
    .A2(net5049));
 sg13g2_o21ai_1 _22184_ (.B1(_05908_),
    .Y(_01991_),
    .A1(_04061_),
    .A2(_05909_));
 sg13g2_a221oi_1 _22185_ (.B2(net4635),
    .C1(net4602),
    .B1(_04069_),
    .A1(net5373),
    .Y(_05910_),
    .A2(net5140));
 sg13g2_a21o_1 _22186_ (.A2(net4602),
    .A1(net1930),
    .B1(_05910_),
    .X(_01992_));
 sg13g2_nand2_1 _22187_ (.Y(_05911_),
    .A(net1612),
    .B(net4602));
 sg13g2_o21ai_1 _22188_ (.B1(net4637),
    .Y(_05912_),
    .A1(\fpga_top.cpu_start_adr[16] ),
    .A2(net5055));
 sg13g2_o21ai_1 _22189_ (.B1(_05911_),
    .Y(_01993_),
    .A1(_04082_),
    .A2(_05912_));
 sg13g2_nand2_1 _22190_ (.Y(_05913_),
    .A(net2111),
    .B(net4605));
 sg13g2_o21ai_1 _22191_ (.B1(net4636),
    .Y(_05914_),
    .A1(\fpga_top.cpu_start_adr[17] ),
    .A2(net5058));
 sg13g2_o21ai_1 _22192_ (.B1(_05913_),
    .Y(_01994_),
    .A1(_04092_),
    .A2(_05914_));
 sg13g2_a221oi_1 _22193_ (.B2(net4635),
    .C1(net4602),
    .B1(_04099_),
    .A1(_06800_),
    .Y(_05915_),
    .A2(net5143));
 sg13g2_a21o_1 _22194_ (.A2(net4606),
    .A1(net2026),
    .B1(_05915_),
    .X(_01995_));
 sg13g2_nor2_1 _22195_ (.A(_04111_),
    .B(net4603),
    .Y(_05916_));
 sg13g2_a22oi_1 _22196_ (.Y(_05917_),
    .B1(_05916_),
    .B2(_04110_),
    .A2(net4603),
    .A1(net3056));
 sg13g2_inv_1 _22197_ (.Y(_01996_),
    .A(_05917_));
 sg13g2_a221oi_1 _22198_ (.B2(net4635),
    .C1(net4605),
    .B1(_04122_),
    .A1(_06802_),
    .Y(_05918_),
    .A2(net5143));
 sg13g2_a21o_1 _22199_ (.A2(net4605),
    .A1(net3497),
    .B1(_05918_),
    .X(_01997_));
 sg13g2_nor3_1 _22200_ (.A(_04133_),
    .B(_04134_),
    .C(net4603),
    .Y(_05919_));
 sg13g2_a21o_1 _22201_ (.A2(net4604),
    .A1(net2092),
    .B1(_05919_),
    .X(_01998_));
 sg13g2_a221oi_1 _22202_ (.B2(net4635),
    .C1(net4605),
    .B1(_04144_),
    .A1(_06803_),
    .Y(_05920_),
    .A2(net5142));
 sg13g2_a21o_1 _22203_ (.A2(net4605),
    .A1(net1989),
    .B1(_05920_),
    .X(_01999_));
 sg13g2_nor3_1 _22204_ (.A(_04155_),
    .B(_04156_),
    .C(net4604),
    .Y(_05921_));
 sg13g2_a21o_1 _22205_ (.A2(net4604),
    .A1(net2038),
    .B1(_05921_),
    .X(_02000_));
 sg13g2_a221oi_1 _22206_ (.B2(net4635),
    .C1(net4602),
    .B1(_04166_),
    .A1(_06805_),
    .Y(_05922_),
    .A2(net5141));
 sg13g2_a21o_1 _22207_ (.A2(net4606),
    .A1(net2098),
    .B1(_05922_),
    .X(_02001_));
 sg13g2_a221oi_1 _22208_ (.B2(_05883_),
    .C1(net4602),
    .B1(_04176_),
    .A1(_06806_),
    .Y(_05923_),
    .A2(net5141));
 sg13g2_a21o_1 _22209_ (.A2(net4602),
    .A1(net3085),
    .B1(_05923_),
    .X(_02002_));
 sg13g2_nor3_1 _22210_ (.A(_04187_),
    .B(_04188_),
    .C(net4603),
    .Y(_05924_));
 sg13g2_a21o_1 _22211_ (.A2(net4603),
    .A1(net2625),
    .B1(_05924_),
    .X(_02003_));
 sg13g2_o21ai_1 _22212_ (.B1(net4637),
    .Y(_05925_),
    .A1(net5641),
    .A2(net5057));
 sg13g2_a21oi_1 _22213_ (.A1(_04197_),
    .A2(net4635),
    .Y(_05926_),
    .B1(_05925_));
 sg13g2_a21o_1 _22214_ (.A2(net4603),
    .A1(net1995),
    .B1(_05926_),
    .X(_02004_));
 sg13g2_nand2_1 _22215_ (.Y(_05927_),
    .A(net1466),
    .B(net4605));
 sg13g2_o21ai_1 _22216_ (.B1(net4636),
    .Y(_05928_),
    .A1(net5639),
    .A2(net5058));
 sg13g2_o21ai_1 _22217_ (.B1(_05927_),
    .Y(_02005_),
    .A1(_04211_),
    .A2(_05928_));
 sg13g2_nor3_1 _22218_ (.A(_04220_),
    .B(_04221_),
    .C(net4603),
    .Y(_05929_));
 sg13g2_a21o_1 _22219_ (.A2(net4604),
    .A1(net2125),
    .B1(_05929_),
    .X(_02006_));
 sg13g2_nand2_1 _22220_ (.Y(_05930_),
    .A(net1482),
    .B(net4605));
 sg13g2_o21ai_1 _22221_ (.B1(net4637),
    .Y(_05931_),
    .A1(net5636),
    .A2(net5059));
 sg13g2_nor2_1 _22222_ (.A(net5142),
    .B(_04232_),
    .Y(_05932_));
 sg13g2_o21ai_1 _22223_ (.B1(_05930_),
    .Y(_02007_),
    .A1(_05931_),
    .A2(_05932_));
 sg13g2_nor2_1 _22224_ (.A(_04246_),
    .B(net4601),
    .Y(_05933_));
 sg13g2_a22oi_1 _22225_ (.Y(_05934_),
    .B1(_05933_),
    .B2(_04245_),
    .A2(net4601),
    .A1(net3674));
 sg13g2_inv_1 _22226_ (.Y(_02008_),
    .A(_05934_));
 sg13g2_or3_1 _22227_ (.A(_05331_),
    .B(_05891_),
    .C(_05892_),
    .X(_05935_));
 sg13g2_o21ai_1 _22228_ (.B1(_05935_),
    .Y(_02009_),
    .A1(_06890_),
    .A2(_05332_));
 sg13g2_nor3_2 _22229_ (.A(_03818_),
    .B(_03832_),
    .C(_03849_),
    .Y(_05936_));
 sg13g2_nand2_2 _22230_ (.Y(_05937_),
    .A(net4829),
    .B(net4664));
 sg13g2_nand2_2 _22231_ (.Y(_05938_),
    .A(net4828),
    .B(net4660));
 sg13g2_nor3_1 _22232_ (.A(_03867_),
    .B(_05545_),
    .C(net4593),
    .Y(_05939_));
 sg13g2_a21o_1 _22233_ (.A2(net4593),
    .A1(net2594),
    .B1(_05939_),
    .X(_02010_));
 sg13g2_nand2_1 _22234_ (.Y(_05940_),
    .A(net1543),
    .B(net4594));
 sg13g2_o21ai_1 _22235_ (.B1(_05940_),
    .Y(_02011_),
    .A1(_03882_),
    .A2(net4594));
 sg13g2_nand2_1 _22236_ (.Y(_05941_),
    .A(net1530),
    .B(net4593));
 sg13g2_o21ai_1 _22237_ (.B1(_05941_),
    .Y(_02012_),
    .A1(_03899_),
    .A2(net4593));
 sg13g2_nand2_1 _22238_ (.Y(_05942_),
    .A(net1504),
    .B(net4594));
 sg13g2_and2_1 _22239_ (.A(net5049),
    .B(net4661),
    .X(_05943_));
 sg13g2_nand2_2 _22240_ (.Y(_05944_),
    .A(net5047),
    .B(net4660));
 sg13g2_o21ai_1 _22241_ (.B1(_03947_),
    .Y(_05945_),
    .A1(_03945_),
    .A2(_05944_));
 sg13g2_o21ai_1 _22242_ (.B1(_05942_),
    .Y(_02013_),
    .A1(net4591),
    .A2(_05945_));
 sg13g2_nand2_1 _22243_ (.Y(_05946_),
    .A(net1538),
    .B(net4593));
 sg13g2_nand2_1 _22244_ (.Y(_05947_),
    .A(_05887_),
    .B(net4633));
 sg13g2_o21ai_1 _22245_ (.B1(_05946_),
    .Y(_02014_),
    .A1(_05888_),
    .A2(_05947_));
 sg13g2_nand2_1 _22246_ (.Y(_05948_),
    .A(net1486),
    .B(net4594));
 sg13g2_nand2b_1 _22247_ (.Y(_05949_),
    .B(net4633),
    .A_N(_05891_));
 sg13g2_o21ai_1 _22248_ (.B1(_05948_),
    .Y(_02015_),
    .A1(_05892_),
    .A2(_05949_));
 sg13g2_o21ai_1 _22249_ (.B1(_03959_),
    .Y(_05950_),
    .A1(_03957_),
    .A2(_05944_));
 sg13g2_nor2_1 _22250_ (.A(net1918),
    .B(net4633),
    .Y(_05951_));
 sg13g2_a21oi_1 _22251_ (.A1(net4633),
    .A2(_05950_),
    .Y(_02016_),
    .B1(_05951_));
 sg13g2_nand2_1 _22252_ (.Y(_05952_),
    .A(net1433),
    .B(net4594));
 sg13g2_o21ai_1 _22253_ (.B1(_05897_),
    .Y(_05953_),
    .A1(_03971_),
    .A2(_05944_));
 sg13g2_o21ai_1 _22254_ (.B1(_05952_),
    .Y(_02017_),
    .A1(net4591),
    .A2(_05953_));
 sg13g2_nand3_1 _22255_ (.B(_03984_),
    .C(net4633),
    .A(_03983_),
    .Y(_05954_));
 sg13g2_o21ai_1 _22256_ (.B1(_05954_),
    .Y(_02018_),
    .A1(_06897_),
    .A2(net4633));
 sg13g2_nand2_1 _22257_ (.Y(_05955_),
    .A(net1585),
    .B(_05937_));
 sg13g2_o21ai_1 _22258_ (.B1(net4633),
    .Y(_05956_),
    .A1(\fpga_top.cpu_start_adr[9] ),
    .A2(net5055));
 sg13g2_o21ai_1 _22259_ (.B1(_05955_),
    .Y(_02019_),
    .A1(_03999_),
    .A2(_05956_));
 sg13g2_nor3_1 _22260_ (.A(_04008_),
    .B(_04009_),
    .C(net4597),
    .Y(_05957_));
 sg13g2_a21o_1 _22261_ (.A2(net4596),
    .A1(net2110),
    .B1(_05957_),
    .X(_02020_));
 sg13g2_nand2_1 _22262_ (.Y(_05958_),
    .A(net1561),
    .B(net4594));
 sg13g2_o21ai_1 _22263_ (.B1(_05904_),
    .Y(_05959_),
    .A1(_04021_),
    .A2(_05944_));
 sg13g2_o21ai_1 _22264_ (.B1(_05958_),
    .Y(_02021_),
    .A1(net4591),
    .A2(_05959_));
 sg13g2_a221oi_1 _22265_ (.B2(net4590),
    .C1(net4591),
    .B1(_04035_),
    .A1(net5376),
    .Y(_05960_),
    .A2(net5137));
 sg13g2_a21o_1 _22266_ (.A2(net4593),
    .A1(net2091),
    .B1(_05960_),
    .X(_02022_));
 sg13g2_a221oi_1 _22267_ (.B2(net4590),
    .C1(net4591),
    .B1(_04046_),
    .A1(_06795_),
    .Y(_05961_),
    .A2(net5139));
 sg13g2_a21o_1 _22268_ (.A2(net4593),
    .A1(net2023),
    .B1(_05961_),
    .X(_02023_));
 sg13g2_a221oi_1 _22269_ (.B2(net4590),
    .C1(net4591),
    .B1(_04060_),
    .A1(_06796_),
    .Y(_05962_),
    .A2(net5139));
 sg13g2_a21o_1 _22270_ (.A2(net4593),
    .A1(net2089),
    .B1(_05962_),
    .X(_02024_));
 sg13g2_a221oi_1 _22271_ (.B2(net4590),
    .C1(net4592),
    .B1(_04069_),
    .A1(net5373),
    .Y(_05963_),
    .A2(net5140));
 sg13g2_a21o_1 _22272_ (.A2(net4598),
    .A1(net2019),
    .B1(_05963_),
    .X(_02025_));
 sg13g2_nand2_1 _22273_ (.Y(_05964_),
    .A(net1517),
    .B(net4598));
 sg13g2_o21ai_1 _22274_ (.B1(net4634),
    .Y(_05965_),
    .A1(\fpga_top.cpu_start_adr[16] ),
    .A2(net5064));
 sg13g2_o21ai_1 _22275_ (.B1(_05964_),
    .Y(_02026_),
    .A1(_04082_),
    .A2(_05965_));
 sg13g2_nand2_1 _22276_ (.Y(_05966_),
    .A(net1589),
    .B(net4597));
 sg13g2_o21ai_1 _22277_ (.B1(net4634),
    .Y(_05967_),
    .A1(\fpga_top.cpu_start_adr[17] ),
    .A2(net5058));
 sg13g2_o21ai_1 _22278_ (.B1(_05966_),
    .Y(_02027_),
    .A1(_04092_),
    .A2(_05967_));
 sg13g2_a221oi_1 _22279_ (.B2(net4590),
    .C1(net4591),
    .B1(_04099_),
    .A1(_06800_),
    .Y(_05968_),
    .A2(net5143));
 sg13g2_a21o_1 _22280_ (.A2(net4598),
    .A1(net2944),
    .B1(_05968_),
    .X(_02028_));
 sg13g2_nand2_1 _22281_ (.Y(_05969_),
    .A(net1464),
    .B(net4595));
 sg13g2_nand2_1 _22282_ (.Y(_05970_),
    .A(_04110_),
    .B(net4634));
 sg13g2_o21ai_1 _22283_ (.B1(_05969_),
    .Y(_02029_),
    .A1(_04111_),
    .A2(_05970_));
 sg13g2_a221oi_1 _22284_ (.B2(net4590),
    .C1(net4592),
    .B1(_04122_),
    .A1(_06802_),
    .Y(_05971_),
    .A2(net5142));
 sg13g2_a21o_1 _22285_ (.A2(net4597),
    .A1(net2041),
    .B1(_05971_),
    .X(_02030_));
 sg13g2_nor3_1 _22286_ (.A(_04133_),
    .B(_04134_),
    .C(net4595),
    .Y(_05972_));
 sg13g2_a21o_1 _22287_ (.A2(net4595),
    .A1(net2097),
    .B1(_05972_),
    .X(_02031_));
 sg13g2_a221oi_1 _22288_ (.B2(net4590),
    .C1(net4592),
    .B1(_04144_),
    .A1(_06803_),
    .Y(_05973_),
    .A2(net5142));
 sg13g2_a21o_1 _22289_ (.A2(net4597),
    .A1(net2090),
    .B1(_05973_),
    .X(_02032_));
 sg13g2_nor3_1 _22290_ (.A(_04155_),
    .B(_04156_),
    .C(net4595),
    .Y(_05974_));
 sg13g2_a21o_1 _22291_ (.A2(net4596),
    .A1(net1942),
    .B1(_05974_),
    .X(_02033_));
 sg13g2_a221oi_1 _22292_ (.B2(_05943_),
    .C1(net4592),
    .B1(_04166_),
    .A1(_06805_),
    .Y(_05975_),
    .A2(net5141));
 sg13g2_a21o_1 _22293_ (.A2(net4598),
    .A1(net1998),
    .B1(_05975_),
    .X(_02034_));
 sg13g2_a221oi_1 _22294_ (.B2(net4590),
    .C1(net4591),
    .B1(_04176_),
    .A1(_06806_),
    .Y(_05976_),
    .A2(net5141));
 sg13g2_a21o_1 _22295_ (.A2(net4598),
    .A1(net2055),
    .B1(_05976_),
    .X(_02035_));
 sg13g2_nor3_1 _22296_ (.A(_04187_),
    .B(_04188_),
    .C(net4595),
    .Y(_05977_));
 sg13g2_a21o_1 _22297_ (.A2(net4595),
    .A1(net2132),
    .B1(_05977_),
    .X(_02036_));
 sg13g2_nand2_1 _22298_ (.Y(_05978_),
    .A(net1501),
    .B(net4596));
 sg13g2_o21ai_1 _22299_ (.B1(net4634),
    .Y(_05979_),
    .A1(net5641),
    .A2(net5056));
 sg13g2_o21ai_1 _22300_ (.B1(_05978_),
    .Y(_02037_),
    .A1(_04198_),
    .A2(_05979_));
 sg13g2_nand2_1 _22301_ (.Y(_05980_),
    .A(net1924),
    .B(net4597));
 sg13g2_o21ai_1 _22302_ (.B1(net4634),
    .Y(_05981_),
    .A1(net5639),
    .A2(net5058));
 sg13g2_o21ai_1 _22303_ (.B1(_05980_),
    .Y(_02038_),
    .A1(_04211_),
    .A2(_05981_));
 sg13g2_nor3_1 _22304_ (.A(_04220_),
    .B(_04221_),
    .C(net4595),
    .Y(_05982_));
 sg13g2_a21o_1 _22305_ (.A2(net4595),
    .A1(net1972),
    .B1(_05982_),
    .X(_02039_));
 sg13g2_nand2_1 _22306_ (.Y(_05983_),
    .A(net1595),
    .B(net4597));
 sg13g2_o21ai_1 _22307_ (.B1(net4634),
    .Y(_05984_),
    .A1(net5636),
    .A2(net5059));
 sg13g2_o21ai_1 _22308_ (.B1(_05983_),
    .Y(_02040_),
    .A1(_05932_),
    .A2(_05984_));
 sg13g2_nand2_1 _22309_ (.Y(_05985_),
    .A(net1452),
    .B(net4594));
 sg13g2_nand2_1 _22310_ (.Y(_05986_),
    .A(_04245_),
    .B(net4633));
 sg13g2_o21ai_1 _22311_ (.B1(_05985_),
    .Y(_02041_),
    .A1(_04246_),
    .A2(_05986_));
 sg13g2_nor2_1 _22312_ (.A(_03832_),
    .B(net4695),
    .Y(_05987_));
 sg13g2_nor2_2 _22313_ (.A(_03832_),
    .B(_03864_),
    .Y(_05988_));
 sg13g2_nand2_1 _22314_ (.Y(_05989_),
    .A(net4829),
    .B(net4692));
 sg13g2_nor3_1 _22315_ (.A(_03867_),
    .B(_05545_),
    .C(net4678),
    .Y(_05990_));
 sg13g2_a21o_1 _22316_ (.A2(net4678),
    .A1(net3897),
    .B1(_05990_),
    .X(_02042_));
 sg13g2_nand2_1 _22317_ (.Y(_05991_),
    .A(net2201),
    .B(net4677));
 sg13g2_o21ai_1 _22318_ (.B1(_05991_),
    .Y(_02043_),
    .A1(_03882_),
    .A2(net4677));
 sg13g2_nand2_1 _22319_ (.Y(_05992_),
    .A(net3135),
    .B(net4679));
 sg13g2_o21ai_1 _22320_ (.B1(_05992_),
    .Y(_02044_),
    .A1(_03899_),
    .A2(net4683));
 sg13g2_nor2_1 _22321_ (.A(net6080),
    .B(net4685),
    .Y(_05993_));
 sg13g2_nor2_2 _22322_ (.A(net5137),
    .B(_03864_),
    .Y(_05994_));
 sg13g2_nand2_2 _22323_ (.Y(_05995_),
    .A(net5048),
    .B(net4694));
 sg13g2_a22oi_1 _22324_ (.Y(_05996_),
    .B1(_03945_),
    .B2(_05994_),
    .A2(net5135),
    .A1(net5663));
 sg13g2_a21oi_1 _22325_ (.A1(_05988_),
    .A2(_05996_),
    .Y(_02045_),
    .B1(_05993_));
 sg13g2_nor2_1 _22326_ (.A(_05888_),
    .B(net4678),
    .Y(_05997_));
 sg13g2_a22oi_1 _22327_ (.Y(_05998_),
    .B1(_05997_),
    .B2(_05887_),
    .A2(net4678),
    .A1(net3993));
 sg13g2_inv_1 _22328_ (.Y(_02046_),
    .A(_05998_));
 sg13g2_nand2_1 _22329_ (.Y(_05999_),
    .A(net3786),
    .B(net4677));
 sg13g2_a21o_1 _22330_ (.A2(_05994_),
    .A1(_05391_),
    .B1(_05891_),
    .X(_06000_));
 sg13g2_o21ai_1 _22331_ (.B1(_05999_),
    .Y(_02047_),
    .A1(net4677),
    .A2(_06000_));
 sg13g2_nand2_1 _22332_ (.Y(_06001_),
    .A(net3675),
    .B(net4677));
 sg13g2_o21ai_1 _22333_ (.B1(_03959_),
    .Y(_06002_),
    .A1(net5134),
    .A2(_03957_));
 sg13g2_o21ai_1 _22334_ (.B1(_06001_),
    .Y(_02048_),
    .A1(net4677),
    .A2(_06002_));
 sg13g2_nand2_1 _22335_ (.Y(_06003_),
    .A(net3846),
    .B(net4677));
 sg13g2_o21ai_1 _22336_ (.B1(_05897_),
    .Y(_06004_),
    .A1(_03971_),
    .A2(_05995_));
 sg13g2_o21ai_1 _22337_ (.B1(_06003_),
    .Y(_02049_),
    .A1(net4677),
    .A2(_06004_));
 sg13g2_nand3_1 _22338_ (.B(_03984_),
    .C(net4685),
    .A(_03983_),
    .Y(_06005_));
 sg13g2_o21ai_1 _22339_ (.B1(_06005_),
    .Y(_02050_),
    .A1(_06900_),
    .A2(_05988_));
 sg13g2_a221oi_1 _22340_ (.B2(_05994_),
    .C1(net4679),
    .B1(_03998_),
    .A1(\fpga_top.cpu_start_adr[9] ),
    .Y(_06006_),
    .A2(net5139));
 sg13g2_a21oi_1 _22341_ (.A1(_06902_),
    .A2(net4679),
    .Y(_02051_),
    .B1(_06006_));
 sg13g2_nand2_1 _22342_ (.Y(_06007_),
    .A(net6229),
    .B(net4681));
 sg13g2_nand2b_1 _22343_ (.Y(_06008_),
    .B(net4684),
    .A_N(_04009_));
 sg13g2_o21ai_1 _22344_ (.B1(_06007_),
    .Y(_02052_),
    .A1(_04008_),
    .A2(_06008_));
 sg13g2_nand2_1 _22345_ (.Y(_06009_),
    .A(net3869),
    .B(net4678));
 sg13g2_o21ai_1 _22346_ (.B1(_05904_),
    .Y(_06010_),
    .A1(_04021_),
    .A2(_05995_));
 sg13g2_o21ai_1 _22347_ (.B1(_06009_),
    .Y(_02053_),
    .A1(net4678),
    .A2(_06010_));
 sg13g2_a221oi_1 _22348_ (.B2(_05994_),
    .C1(net4679),
    .B1(_04035_),
    .A1(net5376),
    .Y(_06011_),
    .A2(net5137));
 sg13g2_a21o_1 _22349_ (.A2(net4679),
    .A1(net6100),
    .B1(_06011_),
    .X(_02054_));
 sg13g2_nor2_1 _22350_ (.A(net3950),
    .B(net4685),
    .Y(_06012_));
 sg13g2_nor2_1 _22351_ (.A(_04046_),
    .B(_05995_),
    .Y(_06013_));
 sg13g2_a21oi_1 _22352_ (.A1(\fpga_top.cpu_start_adr[13] ),
    .A2(net5139),
    .Y(_06014_),
    .B1(_06013_));
 sg13g2_a21oi_1 _22353_ (.A1(_05988_),
    .A2(_06014_),
    .Y(_02055_),
    .B1(_06012_));
 sg13g2_nor2_1 _22354_ (.A(net6199),
    .B(net4685),
    .Y(_06015_));
 sg13g2_nor2_1 _22355_ (.A(_04060_),
    .B(_05995_),
    .Y(_06016_));
 sg13g2_a21oi_1 _22356_ (.A1(\fpga_top.cpu_start_adr[14] ),
    .A2(net5139),
    .Y(_06017_),
    .B1(_06016_));
 sg13g2_a21oi_1 _22357_ (.A1(_05988_),
    .A2(_06017_),
    .Y(_02056_),
    .B1(_06015_));
 sg13g2_a221oi_1 _22358_ (.B2(_05994_),
    .C1(net4682),
    .B1(_04069_),
    .A1(_06797_),
    .Y(_06018_),
    .A2(net5139));
 sg13g2_a21o_1 _22359_ (.A2(net4682),
    .A1(net6088),
    .B1(_06018_),
    .X(_02057_));
 sg13g2_a221oi_1 _22360_ (.B2(_05994_),
    .C1(net4682),
    .B1(_04081_),
    .A1(\fpga_top.cpu_start_adr[16] ),
    .Y(_06019_),
    .A2(net5144));
 sg13g2_a21oi_1 _22361_ (.A1(_06909_),
    .A2(net4682),
    .Y(_02058_),
    .B1(_06019_));
 sg13g2_nand2_1 _22362_ (.Y(_06020_),
    .A(net3941),
    .B(net4681));
 sg13g2_o21ai_1 _22363_ (.B1(net4685),
    .Y(_06021_),
    .A1(\fpga_top.cpu_start_adr[17] ),
    .A2(net5057));
 sg13g2_o21ai_1 _22364_ (.B1(_06020_),
    .Y(_02059_),
    .A1(_04092_),
    .A2(_06021_));
 sg13g2_a221oi_1 _22365_ (.B2(_05994_),
    .C1(net4682),
    .B1(_04099_),
    .A1(_06800_),
    .Y(_06022_),
    .A2(net5144));
 sg13g2_a21o_1 _22366_ (.A2(net4682),
    .A1(net3948),
    .B1(_06022_),
    .X(_02060_));
 sg13g2_nor2_1 _22367_ (.A(_04111_),
    .B(net4680),
    .Y(_06023_));
 sg13g2_a22oi_1 _22368_ (.Y(_06024_),
    .B1(_06023_),
    .B2(_04110_),
    .A2(net4680),
    .A1(net6329));
 sg13g2_inv_1 _22369_ (.Y(_02061_),
    .A(_06024_));
 sg13g2_nor2_1 _22370_ (.A(net3886),
    .B(net4684),
    .Y(_06025_));
 sg13g2_nor2_1 _22371_ (.A(_04122_),
    .B(_05995_),
    .Y(_06026_));
 sg13g2_a21oi_1 _22372_ (.A1(\fpga_top.cpu_start_adr[20] ),
    .A2(net5143),
    .Y(_06027_),
    .B1(_06026_));
 sg13g2_a21oi_1 _22373_ (.A1(_05988_),
    .A2(_06027_),
    .Y(_02062_),
    .B1(_06025_));
 sg13g2_nor3_1 _22374_ (.A(_04133_),
    .B(_04134_),
    .C(net4680),
    .Y(_06028_));
 sg13g2_a21o_1 _22375_ (.A2(net4680),
    .A1(net6294),
    .B1(_06028_),
    .X(_02063_));
 sg13g2_nor2_1 _22376_ (.A(net6106),
    .B(net4684),
    .Y(_06029_));
 sg13g2_nor2_1 _22377_ (.A(_04144_),
    .B(_05995_),
    .Y(_06030_));
 sg13g2_a21oi_1 _22378_ (.A1(\fpga_top.cpu_start_adr[22] ),
    .A2(net5143),
    .Y(_06031_),
    .B1(_06030_));
 sg13g2_a21oi_1 _22379_ (.A1(_05988_),
    .A2(_06031_),
    .Y(_02064_),
    .B1(_06029_));
 sg13g2_nor3_1 _22380_ (.A(_04155_),
    .B(_04156_),
    .C(net4680),
    .Y(_06032_));
 sg13g2_a21o_1 _22381_ (.A2(net4681),
    .A1(net6201),
    .B1(_06032_),
    .X(_02065_));
 sg13g2_nand2b_1 _22382_ (.Y(_06033_),
    .B(_05994_),
    .A_N(_04166_));
 sg13g2_a21oi_1 _22383_ (.A1(\fpga_top.cpu_start_adr[24] ),
    .A2(net5144),
    .Y(_06034_),
    .B1(net4682));
 sg13g2_a22oi_1 _22384_ (.Y(_02066_),
    .B1(_06033_),
    .B2(_06034_),
    .A2(net4682),
    .A1(_06917_));
 sg13g2_nor2_1 _22385_ (.A(net3612),
    .B(net4684),
    .Y(_06035_));
 sg13g2_nor2_1 _22386_ (.A(_04176_),
    .B(_05995_),
    .Y(_06036_));
 sg13g2_a21oi_1 _22387_ (.A1(net6587),
    .A2(net5141),
    .Y(_06037_),
    .B1(_06036_));
 sg13g2_a21oi_1 _22388_ (.A1(_05988_),
    .A2(_06037_),
    .Y(_02067_),
    .B1(_06035_));
 sg13g2_nand2_1 _22389_ (.Y(_06038_),
    .A(net3916),
    .B(net4680));
 sg13g2_nand2b_1 _22390_ (.Y(_06039_),
    .B(net4684),
    .A_N(_04188_));
 sg13g2_o21ai_1 _22391_ (.B1(_06038_),
    .Y(_02068_),
    .A1(_04187_),
    .A2(_06039_));
 sg13g2_nand2_1 _22392_ (.Y(_06040_),
    .A(net2001),
    .B(net4681));
 sg13g2_o21ai_1 _22393_ (.B1(net4684),
    .Y(_06041_),
    .A1(net5641),
    .A2(net5057));
 sg13g2_o21ai_1 _22394_ (.B1(_06040_),
    .Y(_02069_),
    .A1(_04198_),
    .A2(_06041_));
 sg13g2_nand2_1 _22395_ (.Y(_06042_),
    .A(net3649),
    .B(net4681));
 sg13g2_o21ai_1 _22396_ (.B1(net4684),
    .Y(_06043_),
    .A1(net5639),
    .A2(net5057));
 sg13g2_o21ai_1 _22397_ (.B1(_06042_),
    .Y(_02070_),
    .A1(_04211_),
    .A2(_06043_));
 sg13g2_nor3_1 _22398_ (.A(_04220_),
    .B(_04221_),
    .C(net4680),
    .Y(_06044_));
 sg13g2_a21o_1 _22399_ (.A2(net4680),
    .A1(net6132),
    .B1(_06044_),
    .X(_02071_));
 sg13g2_nand2_1 _22400_ (.Y(_06045_),
    .A(net3739),
    .B(net4681));
 sg13g2_o21ai_1 _22401_ (.B1(net4684),
    .Y(_06046_),
    .A1(net5636),
    .A2(net5059));
 sg13g2_o21ai_1 _22402_ (.B1(_06045_),
    .Y(_02072_),
    .A1(_05932_),
    .A2(_06046_));
 sg13g2_nor2_1 _22403_ (.A(_04246_),
    .B(net4683),
    .Y(_06047_));
 sg13g2_a22oi_1 _22404_ (.Y(_06048_),
    .B1(_06047_),
    .B2(_04245_),
    .A2(net4679),
    .A1(net6155));
 sg13g2_inv_1 _22405_ (.Y(_02073_),
    .A(_06048_));
 sg13g2_nand2_1 _22406_ (.Y(_06049_),
    .A(net1445),
    .B(_05331_));
 sg13g2_o21ai_1 _22407_ (.B1(_06049_),
    .Y(_02074_),
    .A1(_03882_),
    .A2(_05331_));
 sg13g2_nand3_1 _22408_ (.B(_03984_),
    .C(_05332_),
    .A(_03983_),
    .Y(_06050_));
 sg13g2_o21ai_1 _22409_ (.B1(_06050_),
    .Y(_02075_),
    .A1(_06901_),
    .A2(_05332_));
 sg13g2_nand2_1 _22410_ (.Y(_06051_),
    .A(net2301),
    .B(_08849_));
 sg13g2_o21ai_1 _22411_ (.B1(net2302),
    .Y(_02076_),
    .A1(_07303_),
    .A2(net4570));
 sg13g2_mux2_1 _22412_ (.A0(_07606_),
    .A1(net5440),
    .S(net4570),
    .X(_02077_));
 sg13g2_or2_1 _22413_ (.X(_06052_),
    .B(\fpga_top.cpu_start ),
    .A(net5426));
 sg13g2_nand3_1 _22414_ (.B(_08684_),
    .C(_06052_),
    .A(net5604),
    .Y(_06053_));
 sg13g2_o21ai_1 _22415_ (.B1(net6281),
    .Y(_02078_),
    .A1(_06924_),
    .A2(net5604));
 sg13g2_nor2_1 _22416_ (.A(\fpga_top.qspi_if.qspi_state[2] ),
    .B(net5350),
    .Y(_06054_));
 sg13g2_a21oi_1 _22417_ (.A1(_06660_),
    .A2(net5351),
    .Y(_02079_),
    .B1(_06054_));
 sg13g2_nor2_2 _22418_ (.A(net4560),
    .B(_02995_),
    .Y(_06055_));
 sg13g2_nor2_1 _22419_ (.A(net3454),
    .B(net4487),
    .Y(_06056_));
 sg13g2_a21oi_1 _22420_ (.A1(net4919),
    .A2(net4487),
    .Y(_02080_),
    .B1(_06056_));
 sg13g2_nor2_1 _22421_ (.A(net3758),
    .B(net4485),
    .Y(_06057_));
 sg13g2_a21oi_1 _22422_ (.A1(net4917),
    .A2(net4485),
    .Y(_02081_),
    .B1(_06057_));
 sg13g2_nor2_1 _22423_ (.A(net3716),
    .B(net4485),
    .Y(_06058_));
 sg13g2_a21oi_1 _22424_ (.A1(net4852),
    .A2(net4485),
    .Y(_02082_),
    .B1(_06058_));
 sg13g2_nand2_1 _22425_ (.Y(_06059_),
    .A(net4843),
    .B(net4485));
 sg13g2_o21ai_1 _22426_ (.B1(_06059_),
    .Y(_02083_),
    .A1(_06688_),
    .A2(net4485));
 sg13g2_nand2_1 _22427_ (.Y(_06060_),
    .A(net4838),
    .B(net4485));
 sg13g2_o21ai_1 _22428_ (.B1(_06060_),
    .Y(_02084_),
    .A1(_06696_),
    .A2(net4485));
 sg13g2_nor2_1 _22429_ (.A(net3646),
    .B(net4486),
    .Y(_06061_));
 sg13g2_a21oi_1 _22430_ (.A1(net4836),
    .A2(net4486),
    .Y(_02085_),
    .B1(_06061_));
 sg13g2_nor2_1 _22431_ (.A(net3634),
    .B(net4486),
    .Y(_06062_));
 sg13g2_a21oi_1 _22432_ (.A1(net4833),
    .A2(net4486),
    .Y(_02086_),
    .B1(_06062_));
 sg13g2_nor2_1 _22433_ (.A(net2077),
    .B(net4488),
    .Y(_06063_));
 sg13g2_a21oi_1 _22434_ (.A1(net4831),
    .A2(net4488),
    .Y(_02087_),
    .B1(_06063_));
 sg13g2_nor2_1 _22435_ (.A(net3362),
    .B(net4488),
    .Y(_06064_));
 sg13g2_a21oi_1 _22436_ (.A1(_02763_),
    .A2(net4488),
    .Y(_02088_),
    .B1(_06064_));
 sg13g2_nor2_1 _22437_ (.A(net3672),
    .B(net4490),
    .Y(_06065_));
 sg13g2_a21oi_1 _22438_ (.A1(_02767_),
    .A2(net4490),
    .Y(_02089_),
    .B1(_06065_));
 sg13g2_nand2_1 _22439_ (.Y(_06066_),
    .A(_08981_),
    .B(net4490));
 sg13g2_o21ai_1 _22440_ (.B1(_06066_),
    .Y(_02090_),
    .A1(_06707_),
    .A2(net4490));
 sg13g2_nor2_1 _22441_ (.A(net1994),
    .B(net4492),
    .Y(_06067_));
 sg13g2_a21oi_1 _22442_ (.A1(_02771_),
    .A2(net4492),
    .Y(_02091_),
    .B1(_06067_));
 sg13g2_nor2_1 _22443_ (.A(net3506),
    .B(net4494),
    .Y(_06068_));
 sg13g2_a21oi_1 _22444_ (.A1(_02775_),
    .A2(net4494),
    .Y(_02092_),
    .B1(_06068_));
 sg13g2_nor2_1 _22445_ (.A(net3817),
    .B(net4494),
    .Y(_06069_));
 sg13g2_a21oi_1 _22446_ (.A1(_02778_),
    .A2(net4494),
    .Y(_02093_),
    .B1(_06069_));
 sg13g2_nor2_1 _22447_ (.A(net3512),
    .B(net4494),
    .Y(_06070_));
 sg13g2_a21oi_1 _22448_ (.A1(_02781_),
    .A2(net4494),
    .Y(_02094_),
    .B1(_06070_));
 sg13g2_nor2_1 _22449_ (.A(net2106),
    .B(net4495),
    .Y(_06071_));
 sg13g2_a21oi_1 _22450_ (.A1(_02784_),
    .A2(net4495),
    .Y(_02095_),
    .B1(_06071_));
 sg13g2_nor2_1 _22451_ (.A(net3769),
    .B(net4491),
    .Y(_06072_));
 sg13g2_a21oi_1 _22452_ (.A1(_10595_),
    .A2(net4491),
    .Y(_02096_),
    .B1(_06072_));
 sg13g2_nor2_1 _22453_ (.A(net3800),
    .B(net4491),
    .Y(_06073_));
 sg13g2_a21oi_1 _22454_ (.A1(_10600_),
    .A2(net4491),
    .Y(_02097_),
    .B1(_06073_));
 sg13g2_nor2_1 _22455_ (.A(net3176),
    .B(net4491),
    .Y(_06074_));
 sg13g2_a21oi_1 _22456_ (.A1(_10603_),
    .A2(net4491),
    .Y(_02098_),
    .B1(_06074_));
 sg13g2_nor2_1 _22457_ (.A(net3814),
    .B(net4490),
    .Y(_06075_));
 sg13g2_a21oi_1 _22458_ (.A1(_02789_),
    .A2(net4490),
    .Y(_02099_),
    .B1(_06075_));
 sg13g2_nor2_1 _22459_ (.A(net3468),
    .B(net4491),
    .Y(_06076_));
 sg13g2_a21oi_1 _22460_ (.A1(_10605_),
    .A2(net4491),
    .Y(_02100_),
    .B1(_06076_));
 sg13g2_nor2_1 _22461_ (.A(net3882),
    .B(net4492),
    .Y(_06077_));
 sg13g2_a21oi_1 _22462_ (.A1(_10609_),
    .A2(net4492),
    .Y(_02101_),
    .B1(_06077_));
 sg13g2_nor2_1 _22463_ (.A(net3540),
    .B(net4492),
    .Y(_06078_));
 sg13g2_a21oi_1 _22464_ (.A1(_10611_),
    .A2(net4493),
    .Y(_02102_),
    .B1(_06078_));
 sg13g2_nor2_1 _22465_ (.A(net3269),
    .B(net4490),
    .Y(_06079_));
 sg13g2_a21oi_1 _22466_ (.A1(_02795_),
    .A2(net4490),
    .Y(_02103_),
    .B1(_06079_));
 sg13g2_nor2_1 _22467_ (.A(net2347),
    .B(net4489),
    .Y(_06080_));
 sg13g2_a21oi_1 _22468_ (.A1(_10615_),
    .A2(net4489),
    .Y(_02104_),
    .B1(_06080_));
 sg13g2_nor2_1 _22469_ (.A(net3364),
    .B(net4496),
    .Y(_06081_));
 sg13g2_a21oi_1 _22470_ (.A1(_10618_),
    .A2(net4496),
    .Y(_02105_),
    .B1(_06081_));
 sg13g2_nor2_1 _22471_ (.A(net3787),
    .B(net4489),
    .Y(_06082_));
 sg13g2_a21oi_1 _22472_ (.A1(_10622_),
    .A2(net4489),
    .Y(_02106_),
    .B1(_06082_));
 sg13g2_nor2_1 _22473_ (.A(net3836),
    .B(net4495),
    .Y(_06083_));
 sg13g2_a21oi_1 _22474_ (.A1(_02803_),
    .A2(net4495),
    .Y(_02107_),
    .B1(_06083_));
 sg13g2_nor2_1 _22475_ (.A(net3759),
    .B(net4496),
    .Y(_06084_));
 sg13g2_a21oi_1 _22476_ (.A1(_02805_),
    .A2(net4496),
    .Y(_02108_),
    .B1(_06084_));
 sg13g2_nor2_1 _22477_ (.A(net3850),
    .B(net4496),
    .Y(_06085_));
 sg13g2_a21oi_1 _22478_ (.A1(_02809_),
    .A2(net4496),
    .Y(_02109_),
    .B1(_06085_));
 sg13g2_nor2_1 _22479_ (.A(net3943),
    .B(net4494),
    .Y(_06086_));
 sg13g2_a21oi_1 _22480_ (.A1(_02814_),
    .A2(net4494),
    .Y(_02110_),
    .B1(_06086_));
 sg13g2_nor2_1 _22481_ (.A(net3642),
    .B(net4489),
    .Y(_06087_));
 sg13g2_a21oi_1 _22482_ (.A1(_02817_),
    .A2(net4489),
    .Y(_02111_),
    .B1(_06087_));
 sg13g2_o21ai_1 _22483_ (.B1(net4468),
    .Y(_06088_),
    .A1(\fpga_top.io_frc.frc_cntrl_val ),
    .A2(_03054_));
 sg13g2_nand2_1 _22484_ (.Y(_06089_),
    .A(net3747),
    .B(net4418));
 sg13g2_a21oi_2 _22485_ (.B1(net4417),
    .Y(_06090_),
    .A2(net4846),
    .A1(_08912_));
 sg13g2_a21o_1 _22486_ (.A2(net4846),
    .A1(_08912_),
    .B1(net4417),
    .X(_06091_));
 sg13g2_xnor2_1 _22487_ (.Y(_06092_),
    .A(net3747),
    .B(_03159_));
 sg13g2_nor2_1 _22488_ (.A(net4510),
    .B(_06092_),
    .Y(_06093_));
 sg13g2_a21oi_1 _22489_ (.A1(_10526_),
    .A2(net4510),
    .Y(_06094_),
    .B1(_06093_));
 sg13g2_o21ai_1 _22490_ (.B1(_06089_),
    .Y(_02112_),
    .A1(net4216),
    .A2(_06094_));
 sg13g2_nand2_1 _22491_ (.Y(_06095_),
    .A(net2182),
    .B(net4418));
 sg13g2_nor4_2 _22492_ (.A(_06712_),
    .B(_06765_),
    .C(_06767_),
    .Y(_06096_),
    .D(_03155_));
 sg13g2_a21oi_1 _22493_ (.A1(\fpga_top.io_frc.frc_cntr_val[32] ),
    .A2(_03159_),
    .Y(_06097_),
    .B1(net2182));
 sg13g2_nor3_1 _22494_ (.A(net4510),
    .B(_06096_),
    .C(_06097_),
    .Y(_06098_));
 sg13g2_a21oi_1 _22495_ (.A1(net4846),
    .A2(net4510),
    .Y(_06099_),
    .B1(_06098_));
 sg13g2_o21ai_1 _22496_ (.B1(_06095_),
    .Y(_02113_),
    .A1(net4216),
    .A2(_06099_));
 sg13g2_nand2_1 _22497_ (.Y(_06100_),
    .A(net3125),
    .B(net4418));
 sg13g2_and2_1 _22498_ (.A(\fpga_top.io_frc.frc_cntr_val[34] ),
    .B(_06096_),
    .X(_06101_));
 sg13g2_xnor2_1 _22499_ (.Y(_06102_),
    .A(net3125),
    .B(_06096_));
 sg13g2_nor2_1 _22500_ (.A(net4510),
    .B(_06102_),
    .Y(_06103_));
 sg13g2_a21oi_1 _22501_ (.A1(_08915_),
    .A2(net4510),
    .Y(_06104_),
    .B1(_06103_));
 sg13g2_o21ai_1 _22502_ (.B1(_06100_),
    .Y(_02114_),
    .A1(net4216),
    .A2(_06104_));
 sg13g2_nand2_1 _22503_ (.Y(_06105_),
    .A(net3971),
    .B(net4418));
 sg13g2_nand2_1 _22504_ (.Y(_06106_),
    .A(\fpga_top.io_frc.frc_cntr_val[35] ),
    .B(_06101_));
 sg13g2_xnor2_1 _22505_ (.Y(_06107_),
    .A(net3971),
    .B(_06101_));
 sg13g2_nor2_1 _22506_ (.A(net4510),
    .B(_06107_),
    .Y(_06108_));
 sg13g2_a21oi_1 _22507_ (.A1(net4843),
    .A2(net4510),
    .Y(_06109_),
    .B1(_06108_));
 sg13g2_o21ai_1 _22508_ (.B1(_06105_),
    .Y(_02115_),
    .A1(net4216),
    .A2(_06109_));
 sg13g2_nand2_1 _22509_ (.Y(_06110_),
    .A(net2212),
    .B(net4418));
 sg13g2_and4_1 _22510_ (.A(\fpga_top.io_frc.frc_cntr_val[36] ),
    .B(\fpga_top.io_frc.frc_cntr_val[35] ),
    .C(\fpga_top.io_frc.frc_cntr_val[34] ),
    .D(_06096_),
    .X(_06111_));
 sg13g2_a21oi_1 _22511_ (.A1(\fpga_top.io_frc.frc_cntr_val[35] ),
    .A2(_06101_),
    .Y(_06112_),
    .B1(net2212));
 sg13g2_nor3_1 _22512_ (.A(net4511),
    .B(_06111_),
    .C(_06112_),
    .Y(_06113_));
 sg13g2_a21oi_1 _22513_ (.A1(net4839),
    .A2(net4511),
    .Y(_06114_),
    .B1(_06113_));
 sg13g2_o21ai_1 _22514_ (.B1(_06110_),
    .Y(_02116_),
    .A1(net4216),
    .A2(_06114_));
 sg13g2_xnor2_1 _22515_ (.Y(_06115_),
    .A(_06760_),
    .B(_06111_));
 sg13g2_nor2_1 _22516_ (.A(net4505),
    .B(_06115_),
    .Y(_06116_));
 sg13g2_a21oi_1 _22517_ (.A1(net4836),
    .A2(net4505),
    .Y(_06117_),
    .B1(_06116_));
 sg13g2_a22oi_1 _22518_ (.Y(_06118_),
    .B1(_06090_),
    .B2(_06117_),
    .A2(net4414),
    .A1(net4004));
 sg13g2_inv_1 _22519_ (.Y(_02117_),
    .A(_06118_));
 sg13g2_nand2_1 _22520_ (.Y(_06119_),
    .A(net3449),
    .B(net4414));
 sg13g2_nor4_1 _22521_ (.A(_06758_),
    .B(_06760_),
    .C(_06761_),
    .D(_06106_),
    .Y(_06120_));
 sg13g2_a21oi_1 _22522_ (.A1(\fpga_top.io_frc.frc_cntr_val[37] ),
    .A2(_06111_),
    .Y(_06121_),
    .B1(net3449));
 sg13g2_nor3_1 _22523_ (.A(net4505),
    .B(_06120_),
    .C(_06121_),
    .Y(_06122_));
 sg13g2_a21oi_1 _22524_ (.A1(_02756_),
    .A2(net4505),
    .Y(_06123_),
    .B1(_06122_));
 sg13g2_o21ai_1 _22525_ (.B1(_06119_),
    .Y(_02118_),
    .A1(net4215),
    .A2(_06123_));
 sg13g2_nand2_1 _22526_ (.Y(_06124_),
    .A(net3904),
    .B(net4414));
 sg13g2_and4_1 _22527_ (.A(\fpga_top.io_frc.frc_cntr_val[39] ),
    .B(\fpga_top.io_frc.frc_cntr_val[38] ),
    .C(\fpga_top.io_frc.frc_cntr_val[37] ),
    .D(_06111_),
    .X(_06125_));
 sg13g2_xnor2_1 _22528_ (.Y(_06126_),
    .A(net3904),
    .B(_06120_));
 sg13g2_nor2_1 _22529_ (.A(net4505),
    .B(_06126_),
    .Y(_06127_));
 sg13g2_a21oi_1 _22530_ (.A1(_02760_),
    .A2(net4505),
    .Y(_06128_),
    .B1(_06127_));
 sg13g2_o21ai_1 _22531_ (.B1(_06124_),
    .Y(_02119_),
    .A1(net4215),
    .A2(_06128_));
 sg13g2_nand2_1 _22532_ (.Y(_06129_),
    .A(net3821),
    .B(net4414));
 sg13g2_xnor2_1 _22533_ (.Y(_06130_),
    .A(net3821),
    .B(_06125_));
 sg13g2_nor2_1 _22534_ (.A(net4506),
    .B(_06130_),
    .Y(_06131_));
 sg13g2_a21oi_1 _22535_ (.A1(_02764_),
    .A2(net4506),
    .Y(_06132_),
    .B1(_06131_));
 sg13g2_o21ai_1 _22536_ (.B1(_06129_),
    .Y(_02120_),
    .A1(net4215),
    .A2(_06132_));
 sg13g2_nand2_1 _22537_ (.Y(_06133_),
    .A(net2074),
    .B(net4414));
 sg13g2_and3_2 _22538_ (.X(_06134_),
    .A(\fpga_top.io_frc.frc_cntr_val[41] ),
    .B(\fpga_top.io_frc.frc_cntr_val[40] ),
    .C(_06125_));
 sg13g2_a21oi_1 _22539_ (.A1(\fpga_top.io_frc.frc_cntr_val[40] ),
    .A2(_06125_),
    .Y(_06135_),
    .B1(net2074));
 sg13g2_nor3_1 _22540_ (.A(net4506),
    .B(_06134_),
    .C(_06135_),
    .Y(_06136_));
 sg13g2_a21oi_1 _22541_ (.A1(_02768_),
    .A2(net4506),
    .Y(_06137_),
    .B1(_06136_));
 sg13g2_o21ai_1 _22542_ (.B1(_06133_),
    .Y(_02121_),
    .A1(net4215),
    .A2(_06137_));
 sg13g2_nand2_1 _22543_ (.Y(_06138_),
    .A(net3709),
    .B(net4414));
 sg13g2_xnor2_1 _22544_ (.Y(_06139_),
    .A(net3709),
    .B(_06134_));
 sg13g2_nor2_1 _22545_ (.A(net4506),
    .B(_06139_),
    .Y(_06140_));
 sg13g2_a21oi_1 _22546_ (.A1(_08981_),
    .A2(net4506),
    .Y(_06141_),
    .B1(_06140_));
 sg13g2_o21ai_1 _22547_ (.B1(_06138_),
    .Y(_02122_),
    .A1(net4215),
    .A2(_06141_));
 sg13g2_nand2_1 _22548_ (.Y(_06142_),
    .A(net3113),
    .B(net4414));
 sg13g2_nand2_1 _22549_ (.Y(_06143_),
    .A(_02771_),
    .B(net4505));
 sg13g2_and3_2 _22550_ (.X(_06144_),
    .A(\fpga_top.io_frc.frc_cntr_val[43] ),
    .B(\fpga_top.io_frc.frc_cntr_val[42] ),
    .C(_06134_));
 sg13g2_a21oi_1 _22551_ (.A1(\fpga_top.io_frc.frc_cntr_val[42] ),
    .A2(_06134_),
    .Y(_06145_),
    .B1(net3113));
 sg13g2_nor2_1 _22552_ (.A(_06144_),
    .B(_06145_),
    .Y(_06146_));
 sg13g2_o21ai_1 _22553_ (.B1(_06143_),
    .Y(_06147_),
    .A1(net4505),
    .A2(_06146_));
 sg13g2_o21ai_1 _22554_ (.B1(_06142_),
    .Y(_02123_),
    .A1(net4215),
    .A2(_06147_));
 sg13g2_or2_1 _22555_ (.X(_06148_),
    .B(_06144_),
    .A(net3618));
 sg13g2_and2_1 _22556_ (.A(\fpga_top.io_frc.frc_cntr_val[44] ),
    .B(_06144_),
    .X(_06149_));
 sg13g2_nor2_1 _22557_ (.A(net4512),
    .B(_06149_),
    .Y(_06150_));
 sg13g2_a22oi_1 _22558_ (.Y(_06151_),
    .B1(_06148_),
    .B2(_06150_),
    .A2(net4512),
    .A1(_02774_));
 sg13g2_nand2_1 _22559_ (.Y(_06152_),
    .A(net3618),
    .B(net4417));
 sg13g2_o21ai_1 _22560_ (.B1(_06152_),
    .Y(_02124_),
    .A1(net4216),
    .A2(_06151_));
 sg13g2_nor2_1 _22561_ (.A(net4417),
    .B(_06150_),
    .Y(_06153_));
 sg13g2_nor2_1 _22562_ (.A(net4009),
    .B(_06153_),
    .Y(_06154_));
 sg13g2_nand2_1 _22563_ (.Y(_06155_),
    .A(net4009),
    .B(_06149_));
 sg13g2_nor2_1 _22564_ (.A(net4515),
    .B(_06155_),
    .Y(_06156_));
 sg13g2_a21oi_1 _22565_ (.A1(_02778_),
    .A2(net4512),
    .Y(_06157_),
    .B1(_06156_));
 sg13g2_a21oi_1 _22566_ (.A1(_03050_),
    .A2(_06157_),
    .Y(_06158_),
    .B1(net4417));
 sg13g2_nor2_1 _22567_ (.A(_06154_),
    .B(_06158_),
    .Y(_02125_));
 sg13g2_nand2_1 _22568_ (.Y(_06159_),
    .A(net2078),
    .B(net4417));
 sg13g2_nor2_1 _22569_ (.A(_06756_),
    .B(_06155_),
    .Y(_06160_));
 sg13g2_a21oi_1 _22570_ (.A1(\fpga_top.io_frc.frc_cntr_val[45] ),
    .A2(_06149_),
    .Y(_06161_),
    .B1(net2078));
 sg13g2_nor3_1 _22571_ (.A(net4512),
    .B(_06160_),
    .C(_06161_),
    .Y(_06162_));
 sg13g2_a21oi_1 _22572_ (.A1(_02782_),
    .A2(net4515),
    .Y(_06163_),
    .B1(_06162_));
 sg13g2_o21ai_1 _22573_ (.B1(_06159_),
    .Y(_02126_),
    .A1(net4217),
    .A2(_06163_));
 sg13g2_nand2_1 _22574_ (.Y(_06164_),
    .A(net1958),
    .B(net4416));
 sg13g2_nor3_2 _22575_ (.A(_06755_),
    .B(_06756_),
    .C(_06155_),
    .Y(_06165_));
 sg13g2_xnor2_1 _22576_ (.Y(_06166_),
    .A(_06755_),
    .B(_06160_));
 sg13g2_nand2_1 _22577_ (.Y(_06167_),
    .A(_02784_),
    .B(net4514));
 sg13g2_o21ai_1 _22578_ (.B1(_06167_),
    .Y(_06168_),
    .A1(net4514),
    .A2(_06166_));
 sg13g2_o21ai_1 _22579_ (.B1(_06164_),
    .Y(_02127_),
    .A1(net4217),
    .A2(_06168_));
 sg13g2_nand2_1 _22580_ (.Y(_06169_),
    .A(net4047),
    .B(net4415));
 sg13g2_xnor2_1 _22581_ (.Y(_06170_),
    .A(net4047),
    .B(_06165_));
 sg13g2_nor2_1 _22582_ (.A(net4508),
    .B(_06170_),
    .Y(_06171_));
 sg13g2_a21oi_1 _22583_ (.A1(_10594_),
    .A2(net4508),
    .Y(_06172_),
    .B1(_06171_));
 sg13g2_o21ai_1 _22584_ (.B1(_06169_),
    .Y(_02128_),
    .A1(net4218),
    .A2(_06172_));
 sg13g2_nand2_1 _22585_ (.Y(_06173_),
    .A(net3774),
    .B(net4414));
 sg13g2_and3_2 _22586_ (.X(_06174_),
    .A(\fpga_top.io_frc.frc_cntr_val[49] ),
    .B(\fpga_top.io_frc.frc_cntr_val[48] ),
    .C(_06165_));
 sg13g2_a21oi_1 _22587_ (.A1(\fpga_top.io_frc.frc_cntr_val[48] ),
    .A2(_06165_),
    .Y(_06175_),
    .B1(net3774));
 sg13g2_nor3_1 _22588_ (.A(net4508),
    .B(_06174_),
    .C(_06175_),
    .Y(_06176_));
 sg13g2_a21oi_1 _22589_ (.A1(_10599_),
    .A2(net4508),
    .Y(_06177_),
    .B1(_06176_));
 sg13g2_o21ai_1 _22590_ (.B1(_06173_),
    .Y(_02129_),
    .A1(net4218),
    .A2(_06177_));
 sg13g2_nand2_1 _22591_ (.Y(_06178_),
    .A(net3645),
    .B(net4415));
 sg13g2_xnor2_1 _22592_ (.Y(_06179_),
    .A(_06746_),
    .B(_06174_));
 sg13g2_nand2_1 _22593_ (.Y(_06180_),
    .A(_10603_),
    .B(net4507));
 sg13g2_o21ai_1 _22594_ (.B1(_06180_),
    .Y(_06181_),
    .A1(net4507),
    .A2(_06179_));
 sg13g2_o21ai_1 _22595_ (.B1(_06178_),
    .Y(_02130_),
    .A1(net4215),
    .A2(_06181_));
 sg13g2_nand3_1 _22596_ (.B(\fpga_top.io_frc.frc_cntr_val[50] ),
    .C(_06174_),
    .A(net6606),
    .Y(_06182_));
 sg13g2_a21o_1 _22597_ (.A2(_06174_),
    .A1(\fpga_top.io_frc.frc_cntr_val[50] ),
    .B1(net4065),
    .X(_06183_));
 sg13g2_a21oi_1 _22598_ (.A1(_06182_),
    .A2(_06183_),
    .Y(_06184_),
    .B1(net4507));
 sg13g2_a21oi_1 _22599_ (.A1(_02789_),
    .A2(net4507),
    .Y(_06185_),
    .B1(_06184_));
 sg13g2_a22oi_1 _22600_ (.Y(_06186_),
    .B1(_06090_),
    .B2(_06185_),
    .A2(net4415),
    .A1(net4065));
 sg13g2_inv_1 _22601_ (.Y(_02131_),
    .A(net4066));
 sg13g2_nand2_1 _22602_ (.Y(_06187_),
    .A(net2138),
    .B(net4415));
 sg13g2_or2_1 _22603_ (.X(_06188_),
    .B(_06182_),
    .A(_06752_));
 sg13g2_xnor2_1 _22604_ (.Y(_06189_),
    .A(_06752_),
    .B(net6607));
 sg13g2_nor2_1 _22605_ (.A(net4507),
    .B(_06189_),
    .Y(_06190_));
 sg13g2_a21oi_1 _22606_ (.A1(_10606_),
    .A2(net4507),
    .Y(_06191_),
    .B1(_06190_));
 sg13g2_o21ai_1 _22607_ (.B1(_06187_),
    .Y(_02132_),
    .A1(net4215),
    .A2(_06191_));
 sg13g2_nor3_2 _22608_ (.A(_06751_),
    .B(_06752_),
    .C(_06182_),
    .Y(_06192_));
 sg13g2_a21oi_1 _22609_ (.A1(_06751_),
    .A2(_06188_),
    .Y(_06193_),
    .B1(_06192_));
 sg13g2_nor2_1 _22610_ (.A(net4507),
    .B(_06193_),
    .Y(_06194_));
 sg13g2_a21oi_1 _22611_ (.A1(_10609_),
    .A2(net4507),
    .Y(_06195_),
    .B1(_06194_));
 sg13g2_a22oi_1 _22612_ (.Y(_06196_),
    .B1(_06090_),
    .B2(_06195_),
    .A2(net4415),
    .A1(net3721));
 sg13g2_inv_1 _22613_ (.Y(_02133_),
    .A(net3722));
 sg13g2_nand2_1 _22614_ (.Y(_06197_),
    .A(net3835),
    .B(net4415));
 sg13g2_nand2_1 _22615_ (.Y(_06198_),
    .A(\fpga_top.io_frc.frc_cntr_val[54] ),
    .B(_06192_));
 sg13g2_xnor2_1 _22616_ (.Y(_06199_),
    .A(net3835),
    .B(_06192_));
 sg13g2_nor2_1 _22617_ (.A(net4509),
    .B(_06199_),
    .Y(_06200_));
 sg13g2_a21oi_1 _22618_ (.A1(_10612_),
    .A2(net4509),
    .Y(_06201_),
    .B1(_06200_));
 sg13g2_o21ai_1 _22619_ (.B1(_06197_),
    .Y(_02134_),
    .A1(net4218),
    .A2(_06201_));
 sg13g2_nor2_1 _22620_ (.A(_06748_),
    .B(_06198_),
    .Y(_06202_));
 sg13g2_xnor2_1 _22621_ (.Y(_06203_),
    .A(net6133),
    .B(_06198_));
 sg13g2_nor2_1 _22622_ (.A(net4512),
    .B(_06203_),
    .Y(_06204_));
 sg13g2_a21oi_1 _22623_ (.A1(_02795_),
    .A2(net4512),
    .Y(_06205_),
    .B1(_06204_));
 sg13g2_a22oi_1 _22624_ (.Y(_06206_),
    .B1(_06090_),
    .B2(_06205_),
    .A2(net4417),
    .A1(net6133));
 sg13g2_inv_1 _22625_ (.Y(_02135_),
    .A(_06206_));
 sg13g2_and4_1 _22626_ (.A(\fpga_top.io_frc.frc_cntr_val[56] ),
    .B(\fpga_top.io_frc.frc_cntr_val[55] ),
    .C(\fpga_top.io_frc.frc_cntr_val[54] ),
    .D(_06192_),
    .X(_06207_));
 sg13g2_xnor2_1 _22627_ (.Y(_06208_),
    .A(_06740_),
    .B(_06202_));
 sg13g2_nor2_1 _22628_ (.A(net4513),
    .B(_06208_),
    .Y(_06209_));
 sg13g2_a21oi_1 _22629_ (.A1(_10615_),
    .A2(net4514),
    .Y(_06210_),
    .B1(_06209_));
 sg13g2_a22oi_1 _22630_ (.Y(_06211_),
    .B1(_06090_),
    .B2(_06210_),
    .A2(net4418),
    .A1(net6102));
 sg13g2_inv_1 _22631_ (.Y(_02136_),
    .A(_06211_));
 sg13g2_nor2_1 _22632_ (.A(net4048),
    .B(_06207_),
    .Y(_06212_));
 sg13g2_and2_1 _22633_ (.A(\fpga_top.io_frc.frc_cntr_val[57] ),
    .B(_06207_),
    .X(_06213_));
 sg13g2_nor3_1 _22634_ (.A(net4513),
    .B(_06212_),
    .C(_06213_),
    .Y(_06214_));
 sg13g2_a21o_1 _22635_ (.A2(net4513),
    .A1(_10619_),
    .B1(_06214_),
    .X(_06215_));
 sg13g2_a22oi_1 _22636_ (.Y(_06216_),
    .B1(_06090_),
    .B2(_06215_),
    .A2(net4416),
    .A1(net4048));
 sg13g2_inv_1 _22637_ (.Y(_02137_),
    .A(_06216_));
 sg13g2_nand2_1 _22638_ (.Y(_06217_),
    .A(net2208),
    .B(net4416));
 sg13g2_xnor2_1 _22639_ (.Y(_06218_),
    .A(_06738_),
    .B(_06213_));
 sg13g2_nand2_1 _22640_ (.Y(_06219_),
    .A(_10622_),
    .B(net4513));
 sg13g2_o21ai_1 _22641_ (.B1(_06219_),
    .Y(_06220_),
    .A1(net4513),
    .A2(_06218_));
 sg13g2_o21ai_1 _22642_ (.B1(_06217_),
    .Y(_02138_),
    .A1(net4216),
    .A2(_06220_));
 sg13g2_nand2_1 _22643_ (.Y(_06221_),
    .A(net3388),
    .B(net4416));
 sg13g2_a21oi_1 _22644_ (.A1(net2208),
    .A2(_06213_),
    .Y(_06222_),
    .B1(net3388));
 sg13g2_and3_2 _22645_ (.X(_06223_),
    .A(net3388),
    .B(\fpga_top.io_frc.frc_cntr_val[58] ),
    .C(_06213_));
 sg13g2_nor3_1 _22646_ (.A(net4514),
    .B(_06222_),
    .C(_06223_),
    .Y(_06224_));
 sg13g2_a21oi_1 _22647_ (.A1(_02802_),
    .A2(net4513),
    .Y(_06225_),
    .B1(_06224_));
 sg13g2_o21ai_1 _22648_ (.B1(_06221_),
    .Y(_02139_),
    .A1(net4216),
    .A2(_06225_));
 sg13g2_nand2_1 _22649_ (.Y(_06226_),
    .A(net3923),
    .B(net4416));
 sg13g2_xor2_1 _22650_ (.B(_06223_),
    .A(net3923),
    .X(_06227_));
 sg13g2_nor2_1 _22651_ (.A(net4513),
    .B(_06227_),
    .Y(_06228_));
 sg13g2_a21o_1 _22652_ (.A2(net4514),
    .A1(_02805_),
    .B1(net4217),
    .X(_06229_));
 sg13g2_o21ai_1 _22653_ (.B1(_06226_),
    .Y(_02140_),
    .A1(_06228_),
    .A2(_06229_));
 sg13g2_nand3_1 _22654_ (.B(\fpga_top.io_frc.frc_cntr_val[60] ),
    .C(_06223_),
    .A(\fpga_top.io_frc.frc_cntr_val[61] ),
    .Y(_06230_));
 sg13g2_a21o_1 _22655_ (.A2(_06223_),
    .A1(\fpga_top.io_frc.frc_cntr_val[60] ),
    .B1(\fpga_top.io_frc.frc_cntr_val[61] ),
    .X(_06231_));
 sg13g2_and2_1 _22656_ (.A(_06230_),
    .B(_06231_),
    .X(_06232_));
 sg13g2_nor3_1 _22657_ (.A(_08893_),
    .B(_02808_),
    .C(_03045_),
    .Y(_06233_));
 sg13g2_o21ai_1 _22658_ (.B1(_06090_),
    .Y(_06234_),
    .A1(net4513),
    .A2(_06232_));
 sg13g2_nand2_1 _22659_ (.Y(_06235_),
    .A(net3615),
    .B(net4416));
 sg13g2_o21ai_1 _22660_ (.B1(_06235_),
    .Y(_02141_),
    .A1(_06233_),
    .A2(_06234_));
 sg13g2_nand4_1 _22661_ (.B(\fpga_top.io_frc.frc_cntr_val[61] ),
    .C(\fpga_top.io_frc.frc_cntr_val[60] ),
    .A(\fpga_top.io_frc.frc_cntr_val[62] ),
    .Y(_06236_),
    .D(_06223_));
 sg13g2_xnor2_1 _22662_ (.Y(_06237_),
    .A(net3407),
    .B(_06230_));
 sg13g2_nor3_1 _22663_ (.A(net4560),
    .B(_02813_),
    .C(_03045_),
    .Y(_06238_));
 sg13g2_o21ai_1 _22664_ (.B1(_06090_),
    .Y(_06239_),
    .A1(net4511),
    .A2(_06237_));
 sg13g2_nand2_1 _22665_ (.Y(_06240_),
    .A(net3407),
    .B(net4416));
 sg13g2_o21ai_1 _22666_ (.B1(_06240_),
    .Y(_02142_),
    .A1(_06238_),
    .A2(_06239_));
 sg13g2_nand2_1 _22667_ (.Y(_06241_),
    .A(net2130),
    .B(net4416));
 sg13g2_xnor2_1 _22668_ (.Y(_06242_),
    .A(net2130),
    .B(_06236_));
 sg13g2_nor2_1 _22669_ (.A(net4514),
    .B(_06242_),
    .Y(_06243_));
 sg13g2_a21o_1 _22670_ (.A2(net4514),
    .A1(_02817_),
    .B1(net4217),
    .X(_06244_));
 sg13g2_o21ai_1 _22671_ (.B1(_06241_),
    .Y(_02143_),
    .A1(_06243_),
    .A2(_06244_));
 sg13g2_nor2b_1 _22672_ (.A(net3998),
    .B_N(net1852),
    .Y(_06245_));
 sg13g2_nor2_1 _22673_ (.A(_08753_),
    .B(_06245_),
    .Y(_06246_));
 sg13g2_nor2b_1 _22674_ (.A(\fpga_top.uart_top.uart_rec_char.next_cmd_status[4] ),
    .B_N(_04356_),
    .Y(_06247_));
 sg13g2_nor3_1 _22675_ (.A(net5426),
    .B(_06958_),
    .C(_06973_),
    .Y(_06248_));
 sg13g2_a21oi_1 _22676_ (.A1(_06966_),
    .A2(_08699_),
    .Y(_06249_),
    .B1(_06994_));
 sg13g2_mux4_1 _22677_ (.S0(\fpga_top.uart_top.uart_rec_char.next_cmd_status[3] ),
    .A0(_06247_),
    .A1(_08688_),
    .A2(_07003_),
    .A3(_07006_),
    .S1(\fpga_top.uart_top.uart_rec_char.next_cmd_status[2] ),
    .X(_06250_));
 sg13g2_or3_1 _22678_ (.A(_06248_),
    .B(_06249_),
    .C(_06250_),
    .X(_06251_));
 sg13g2_nor2_1 _22679_ (.A(_07015_),
    .B(_08836_),
    .Y(_06252_));
 sg13g2_nor4_1 _22680_ (.A(_06986_),
    .B(_07022_),
    .C(_08698_),
    .D(_08751_),
    .Y(_06253_));
 sg13g2_or4_1 _22681_ (.A(\fpga_top.uart_top.uart_rec_char.g_crlf ),
    .B(_06251_),
    .C(_06252_),
    .D(_06253_),
    .X(_06254_));
 sg13g2_or3_1 _22682_ (.A(_08753_),
    .B(_06245_),
    .C(_06254_),
    .X(_06255_));
 sg13g2_xnor2_1 _22683_ (.Y(_06256_),
    .A(net5424),
    .B(net5341));
 sg13g2_nand2b_1 _22684_ (.Y(_02144_),
    .B(_06256_),
    .A_N(_06255_));
 sg13g2_o21ai_1 _22685_ (.B1(net5423),
    .Y(_06257_),
    .A1(net5424),
    .A2(_08742_));
 sg13g2_a21oi_1 _22686_ (.A1(_08743_),
    .A2(net6508),
    .Y(_02145_),
    .B1(_06255_));
 sg13g2_nand2_1 _22687_ (.Y(_06258_),
    .A(_08741_),
    .B(_08744_));
 sg13g2_nand2_1 _22688_ (.Y(_06259_),
    .A(net6297),
    .B(_08743_));
 sg13g2_a21oi_1 _22689_ (.A1(_06258_),
    .A2(_06259_),
    .Y(_02146_),
    .B1(_06255_));
 sg13g2_a21oi_1 _22690_ (.A1(net5422),
    .A2(_06258_),
    .Y(_06260_),
    .B1(_08746_));
 sg13g2_o21ai_1 _22691_ (.B1(_06246_),
    .Y(_02147_),
    .A1(_06254_),
    .A2(_06260_));
 sg13g2_a21o_1 _22692_ (.A2(_08747_),
    .A1(net6318),
    .B1(_06255_),
    .X(_02148_));
 sg13g2_nand2b_2 _22693_ (.Y(_06261_),
    .B(net6609),
    .A_N(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[0] ));
 sg13g2_nand2_1 _22694_ (.Y(_06262_),
    .A(net6597),
    .B(net5146));
 sg13g2_nor2_2 _22695_ (.A(_06261_),
    .B(_06262_),
    .Y(_06263_));
 sg13g2_nor2_1 _22696_ (.A(net1732),
    .B(net4866),
    .Y(_06264_));
 sg13g2_a21oi_1 _22697_ (.A1(_04888_),
    .A2(net4866),
    .Y(_02149_),
    .B1(_06264_));
 sg13g2_mux2_1 _22698_ (.A0(net3134),
    .A1(_04896_),
    .S(net4866),
    .X(_02150_));
 sg13g2_mux2_1 _22699_ (.A0(net2703),
    .A1(_04901_),
    .S(net4866),
    .X(_02151_));
 sg13g2_mux2_1 _22700_ (.A0(net2937),
    .A1(_04906_),
    .S(net4866),
    .X(_02152_));
 sg13g2_mux2_1 _22701_ (.A0(net2298),
    .A1(_04911_),
    .S(_06263_),
    .X(_02153_));
 sg13g2_mux2_1 _22702_ (.A0(net2285),
    .A1(_04913_),
    .S(net4866),
    .X(_02154_));
 sg13g2_mux2_1 _22703_ (.A0(net2200),
    .A1(_04917_),
    .S(net4866),
    .X(_02155_));
 sg13g2_mux2_1 _22704_ (.A0(net2235),
    .A1(_04919_),
    .S(net4866),
    .X(_02156_));
 sg13g2_nor3_2 _22705_ (.A(net6590),
    .B(_06929_),
    .C(_03655_),
    .Y(_06265_));
 sg13g2_nor2_1 _22706_ (.A(net1837),
    .B(net4865),
    .Y(_06266_));
 sg13g2_a21oi_1 _22707_ (.A1(_04888_),
    .A2(net4865),
    .Y(_02157_),
    .B1(_06266_));
 sg13g2_mux2_1 _22708_ (.A0(net3323),
    .A1(_04896_),
    .S(net4865),
    .X(_02158_));
 sg13g2_mux2_1 _22709_ (.A0(net2313),
    .A1(_04901_),
    .S(net4865),
    .X(_02159_));
 sg13g2_mux2_1 _22710_ (.A0(net2229),
    .A1(_04906_),
    .S(net4865),
    .X(_02160_));
 sg13g2_mux2_1 _22711_ (.A0(net2452),
    .A1(_04911_),
    .S(_06265_),
    .X(_02161_));
 sg13g2_mux2_1 _22712_ (.A0(net2504),
    .A1(_04913_),
    .S(net4865),
    .X(_02162_));
 sg13g2_mux2_1 _22713_ (.A0(net2400),
    .A1(_04917_),
    .S(net4865),
    .X(_02163_));
 sg13g2_mux2_1 _22714_ (.A0(net3161),
    .A1(_04919_),
    .S(net4865),
    .X(_02164_));
 sg13g2_nor3_2 _22715_ (.A(net6589),
    .B(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[1] ),
    .C(_06262_),
    .Y(_06267_));
 sg13g2_nor2_1 _22716_ (.A(net1821),
    .B(net4864),
    .Y(_06268_));
 sg13g2_a21oi_1 _22717_ (.A1(_04888_),
    .A2(net4864),
    .Y(_02165_),
    .B1(net1822));
 sg13g2_mux2_1 _22718_ (.A0(net3544),
    .A1(_04896_),
    .S(net4864),
    .X(_02166_));
 sg13g2_mux2_1 _22719_ (.A0(net2423),
    .A1(_04901_),
    .S(net4864),
    .X(_02167_));
 sg13g2_mux2_1 _22720_ (.A0(net3178),
    .A1(_04906_),
    .S(net4864),
    .X(_02168_));
 sg13g2_mux2_1 _22721_ (.A0(net2951),
    .A1(_04911_),
    .S(_06267_),
    .X(_02169_));
 sg13g2_mux2_1 _22722_ (.A0(net2830),
    .A1(_04913_),
    .S(net4864),
    .X(_02170_));
 sg13g2_mux2_1 _22723_ (.A0(net2991),
    .A1(_04917_),
    .S(net4864),
    .X(_02171_));
 sg13g2_mux2_1 _22724_ (.A0(net2631),
    .A1(_04919_),
    .S(net4864),
    .X(_02172_));
 sg13g2_nor2_1 _22725_ (.A(net2020),
    .B(net4909),
    .Y(_06269_));
 sg13g2_a21oi_1 _22726_ (.A1(net4909),
    .A2(_04888_),
    .Y(_02173_),
    .B1(net2021));
 sg13g2_nand2_1 _22727_ (.Y(_06270_),
    .A(net4909),
    .B(_04896_));
 sg13g2_o21ai_1 _22728_ (.B1(_06270_),
    .Y(_02174_),
    .A1(_06851_),
    .A2(net4909));
 sg13g2_nand2_1 _22729_ (.Y(_06271_),
    .A(net4910),
    .B(_04901_));
 sg13g2_o21ai_1 _22730_ (.B1(_06271_),
    .Y(_02175_),
    .A1(_06853_),
    .A2(net4909));
 sg13g2_nand2_1 _22731_ (.Y(_06272_),
    .A(net4909),
    .B(_04906_));
 sg13g2_o21ai_1 _22732_ (.B1(_06272_),
    .Y(_02176_),
    .A1(_06856_),
    .A2(net4909));
 sg13g2_mux2_1 _22733_ (.A0(net2666),
    .A1(_04911_),
    .S(net4910),
    .X(_02177_));
 sg13g2_mux2_1 _22734_ (.A0(net3095),
    .A1(_04913_),
    .S(net4910),
    .X(_02178_));
 sg13g2_mux2_1 _22735_ (.A0(net2955),
    .A1(_04917_),
    .S(net4909),
    .X(_02179_));
 sg13g2_mux2_1 _22736_ (.A0(net2274),
    .A1(_04919_),
    .S(net4910),
    .X(_02180_));
 sg13g2_nor3_2 _22737_ (.A(net6592),
    .B(_03654_),
    .C(_06261_),
    .Y(_06273_));
 sg13g2_nor2_1 _22738_ (.A(net1880),
    .B(net4863),
    .Y(_06274_));
 sg13g2_a21oi_1 _22739_ (.A1(_04888_),
    .A2(net4863),
    .Y(_02181_),
    .B1(net1881));
 sg13g2_mux2_1 _22740_ (.A0(net3107),
    .A1(_04896_),
    .S(net4863),
    .X(_02182_));
 sg13g2_mux2_1 _22741_ (.A0(net3760),
    .A1(_04901_),
    .S(net4863),
    .X(_02183_));
 sg13g2_mux2_1 _22742_ (.A0(net2592),
    .A1(_04906_),
    .S(net4863),
    .X(_02184_));
 sg13g2_mux2_1 _22743_ (.A0(net2616),
    .A1(_04911_),
    .S(net4863),
    .X(_02185_));
 sg13g2_mux2_1 _22744_ (.A0(net2306),
    .A1(_04913_),
    .S(net4863),
    .X(_02186_));
 sg13g2_mux2_1 _22745_ (.A0(net2305),
    .A1(_04917_),
    .S(net4863),
    .X(_02187_));
 sg13g2_mux2_1 _22746_ (.A0(net2427),
    .A1(_04919_),
    .S(_06273_),
    .X(_02188_));
 sg13g2_nor3_2 _22747_ (.A(net6609),
    .B(net6592),
    .C(_03655_),
    .Y(_06275_));
 sg13g2_nor2_1 _22748_ (.A(net2025),
    .B(net4862),
    .Y(_06276_));
 sg13g2_a21oi_1 _22749_ (.A1(_04888_),
    .A2(net4862),
    .Y(_02189_),
    .B1(_06276_));
 sg13g2_nand2_1 _22750_ (.Y(_06277_),
    .A(_04896_),
    .B(net4862));
 sg13g2_o21ai_1 _22751_ (.B1(_06277_),
    .Y(_02190_),
    .A1(_06850_),
    .A2(net4862));
 sg13g2_mux2_1 _22752_ (.A0(net2923),
    .A1(_04901_),
    .S(net4862),
    .X(_02191_));
 sg13g2_nand2_1 _22753_ (.Y(_06278_),
    .A(_04906_),
    .B(net4862));
 sg13g2_o21ai_1 _22754_ (.B1(_06278_),
    .Y(_02192_),
    .A1(_06855_),
    .A2(_06275_));
 sg13g2_mux2_1 _22755_ (.A0(net2508),
    .A1(_04911_),
    .S(net4862),
    .X(_02193_));
 sg13g2_mux2_1 _22756_ (.A0(net2072),
    .A1(_04913_),
    .S(_06275_),
    .X(_02194_));
 sg13g2_mux2_1 _22757_ (.A0(net2167),
    .A1(_04917_),
    .S(net4862),
    .X(_02195_));
 sg13g2_mux2_1 _22758_ (.A0(net2983),
    .A1(_04919_),
    .S(_06275_),
    .X(_02196_));
 sg13g2_nor4_2 _22759_ (.A(net3032),
    .B(net6590),
    .C(net3356),
    .Y(_06279_),
    .D(_03654_));
 sg13g2_nor2_1 _22760_ (.A(net1868),
    .B(net4861),
    .Y(_06280_));
 sg13g2_a21oi_1 _22761_ (.A1(_04888_),
    .A2(net4861),
    .Y(_02197_),
    .B1(net1869));
 sg13g2_mux2_1 _22762_ (.A0(net1693),
    .A1(_04896_),
    .S(net4861),
    .X(_02198_));
 sg13g2_mux2_1 _22763_ (.A0(net3380),
    .A1(_04901_),
    .S(net4861),
    .X(_02199_));
 sg13g2_mux2_1 _22764_ (.A0(net3694),
    .A1(_04906_),
    .S(net3357),
    .X(_02200_));
 sg13g2_mux2_1 _22765_ (.A0(net2949),
    .A1(_04911_),
    .S(net4861),
    .X(_02201_));
 sg13g2_mux2_1 _22766_ (.A0(net2634),
    .A1(_04913_),
    .S(net4861),
    .X(_02202_));
 sg13g2_mux2_1 _22767_ (.A0(net2381),
    .A1(_04917_),
    .S(net4861),
    .X(_02203_));
 sg13g2_mux2_1 _22768_ (.A0(net2722),
    .A1(_04919_),
    .S(net4861),
    .X(_02204_));
 sg13g2_nand3_1 _22769_ (.B(net5668),
    .C(_03641_),
    .A(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[1] ),
    .Y(_06281_));
 sg13g2_mux2_1 _22770_ (.A0(net5612),
    .A1(net2152),
    .S(_06281_),
    .X(_02205_));
 sg13g2_mux2_1 _22771_ (.A0(net5611),
    .A1(net2287),
    .S(_06281_),
    .X(_02206_));
 sg13g2_mux2_1 _22772_ (.A0(net5610),
    .A1(net2520),
    .S(_06281_),
    .X(_02207_));
 sg13g2_mux2_1 _22773_ (.A0(net5609),
    .A1(net2430),
    .S(_06281_),
    .X(_02208_));
 sg13g2_mux2_1 _22774_ (.A0(net5608),
    .A1(net2360),
    .S(_06281_),
    .X(_02209_));
 sg13g2_mux2_1 _22775_ (.A0(net5607),
    .A1(net2187),
    .S(_06281_),
    .X(_02210_));
 sg13g2_mux2_1 _22776_ (.A0(net5606),
    .A1(net2259),
    .S(_06281_),
    .X(_02211_));
 sg13g2_mux2_1 _22777_ (.A0(net5605),
    .A1(net2165),
    .S(_06281_),
    .X(_02212_));
 sg13g2_mux4_1 _22778_ (.S0(net5678),
    .A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][0] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][0] ),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][0] ),
    .A3(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][0] ),
    .S1(net5674),
    .X(_06282_));
 sg13g2_nor2_1 _22779_ (.A(net5669),
    .B(_06282_),
    .Y(_06283_));
 sg13g2_nand2b_1 _22780_ (.Y(_06284_),
    .B(net5677),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][0] ));
 sg13g2_o21ai_1 _22781_ (.B1(_06284_),
    .Y(_06285_),
    .A1(net5677),
    .A2(net2696));
 sg13g2_mux2_1 _22782_ (.A0(net2667),
    .A1(net2152),
    .S(net5677),
    .X(_06286_));
 sg13g2_o21ai_1 _22783_ (.B1(net5669),
    .Y(_06287_),
    .A1(net5673),
    .A2(_06285_));
 sg13g2_a21oi_1 _22784_ (.A1(net5673),
    .A2(_06286_),
    .Y(_06288_),
    .B1(_06287_));
 sg13g2_nor3_1 _22785_ (.A(net5337),
    .B(_06283_),
    .C(_06288_),
    .Y(_06289_));
 sg13g2_a21o_1 _22786_ (.A2(net5336),
    .A1(net2724),
    .B1(_06289_),
    .X(_02213_));
 sg13g2_mux4_1 _22787_ (.S0(net5678),
    .A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][1] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][1] ),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][1] ),
    .A3(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][1] ),
    .S1(net5673),
    .X(_06290_));
 sg13g2_nor2_1 _22788_ (.A(net5669),
    .B(_06290_),
    .Y(_06291_));
 sg13g2_nand2b_1 _22789_ (.Y(_06292_),
    .B(net5677),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][1] ));
 sg13g2_o21ai_1 _22790_ (.B1(_06292_),
    .Y(_06293_),
    .A1(net5677),
    .A2(net2975));
 sg13g2_mux2_1 _22791_ (.A0(net2804),
    .A1(net2287),
    .S(net5678),
    .X(_06294_));
 sg13g2_o21ai_1 _22792_ (.B1(net5669),
    .Y(_06295_),
    .A1(net5673),
    .A2(_06293_));
 sg13g2_a21oi_1 _22793_ (.A1(net5673),
    .A2(_06294_),
    .Y(_06296_),
    .B1(_06295_));
 sg13g2_nor3_1 _22794_ (.A(net5337),
    .B(_06291_),
    .C(_06296_),
    .Y(_06297_));
 sg13g2_a21o_1 _22795_ (.A2(net5336),
    .A1(net3914),
    .B1(_06297_),
    .X(_02214_));
 sg13g2_mux4_1 _22796_ (.S0(net5679),
    .A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][2] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][2] ),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][2] ),
    .A3(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][2] ),
    .S1(net5672),
    .X(_06298_));
 sg13g2_nor2_1 _22797_ (.A(net5669),
    .B(_06298_),
    .Y(_06299_));
 sg13g2_nand2b_1 _22798_ (.Y(_06300_),
    .B(net5677),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][2] ));
 sg13g2_o21ai_1 _22799_ (.B1(_06300_),
    .Y(_06301_),
    .A1(net5677),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][2] ));
 sg13g2_mux2_1 _22800_ (.A0(net2774),
    .A1(net2520),
    .S(net5677),
    .X(_06302_));
 sg13g2_o21ai_1 _22801_ (.B1(net5669),
    .Y(_06303_),
    .A1(net5673),
    .A2(_06301_));
 sg13g2_a21oi_1 _22802_ (.A1(net5673),
    .A2(_06302_),
    .Y(_06304_),
    .B1(_06303_));
 sg13g2_nor3_1 _22803_ (.A(net5337),
    .B(_06299_),
    .C(_06304_),
    .Y(_06305_));
 sg13g2_a21o_1 _22804_ (.A2(net5336),
    .A1(net2852),
    .B1(_06305_),
    .X(_02215_));
 sg13g2_mux4_1 _22805_ (.S0(net5678),
    .A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][3] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][3] ),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][3] ),
    .A3(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][3] ),
    .S1(net5674),
    .X(_06306_));
 sg13g2_nor2_1 _22806_ (.A(net5669),
    .B(_06306_),
    .Y(_06307_));
 sg13g2_nand2b_1 _22807_ (.Y(_06308_),
    .B(net5676),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][3] ));
 sg13g2_o21ai_1 _22808_ (.B1(_06308_),
    .Y(_06309_),
    .A1(net5676),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][3] ));
 sg13g2_mux2_1 _22809_ (.A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][3] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][3] ),
    .S(net5679),
    .X(_06310_));
 sg13g2_o21ai_1 _22810_ (.B1(net5670),
    .Y(_06311_),
    .A1(net5672),
    .A2(_06309_));
 sg13g2_a21oi_1 _22811_ (.A1(net5672),
    .A2(_06310_),
    .Y(_06312_),
    .B1(_06311_));
 sg13g2_nor3_1 _22812_ (.A(net5337),
    .B(_06307_),
    .C(_06312_),
    .Y(_06313_));
 sg13g2_a21o_1 _22813_ (.A2(net5336),
    .A1(net3958),
    .B1(_06313_),
    .X(_02216_));
 sg13g2_mux4_1 _22814_ (.S0(net5678),
    .A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][4] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][4] ),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][4] ),
    .A3(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][4] ),
    .S1(net5674),
    .X(_06314_));
 sg13g2_nor2_1 _22815_ (.A(net5669),
    .B(_06314_),
    .Y(_06315_));
 sg13g2_nand2b_1 _22816_ (.Y(_06316_),
    .B(net5676),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][4] ));
 sg13g2_o21ai_1 _22817_ (.B1(_06316_),
    .Y(_06317_),
    .A1(net5676),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][4] ));
 sg13g2_mux2_1 _22818_ (.A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][4] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][4] ),
    .S(net5679),
    .X(_06318_));
 sg13g2_o21ai_1 _22819_ (.B1(net5670),
    .Y(_06319_),
    .A1(net5672),
    .A2(_06317_));
 sg13g2_a21oi_1 _22820_ (.A1(net5672),
    .A2(_06318_),
    .Y(_06320_),
    .B1(_06319_));
 sg13g2_nor3_1 _22821_ (.A(net5336),
    .B(_06315_),
    .C(_06320_),
    .Y(_06321_));
 sg13g2_a21o_1 _22822_ (.A2(net5336),
    .A1(net3623),
    .B1(_06321_),
    .X(_02217_));
 sg13g2_mux4_1 _22823_ (.S0(net5678),
    .A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][5] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][5] ),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][5] ),
    .A3(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][5] ),
    .S1(net5673),
    .X(_06322_));
 sg13g2_nor2_1 _22824_ (.A(\fpga_top.uart_top.uart_if.rx_fifo.radr[2] ),
    .B(_06322_),
    .Y(_06323_));
 sg13g2_nand2b_1 _22825_ (.Y(_06324_),
    .B(net5675),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][5] ));
 sg13g2_o21ai_1 _22826_ (.B1(_06324_),
    .Y(_06325_),
    .A1(net5676),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][5] ));
 sg13g2_mux2_1 _22827_ (.A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][5] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][5] ),
    .S(net5675),
    .X(_06326_));
 sg13g2_o21ai_1 _22828_ (.B1(net5670),
    .Y(_06327_),
    .A1(net5671),
    .A2(_06325_));
 sg13g2_a21oi_1 _22829_ (.A1(net5671),
    .A2(_06326_),
    .Y(_06328_),
    .B1(_06327_));
 sg13g2_nor3_1 _22830_ (.A(net5336),
    .B(_06323_),
    .C(_06328_),
    .Y(_06329_));
 sg13g2_a21o_1 _22831_ (.A2(net5336),
    .A1(net4002),
    .B1(_06329_),
    .X(_02218_));
 sg13g2_mux4_1 _22832_ (.S0(net5676),
    .A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][6] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][6] ),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][6] ),
    .A3(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][6] ),
    .S1(net5671),
    .X(_06330_));
 sg13g2_nor2_1 _22833_ (.A(net5670),
    .B(_06330_),
    .Y(_06331_));
 sg13g2_nand2b_1 _22834_ (.Y(_06332_),
    .B(net5675),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][6] ));
 sg13g2_o21ai_1 _22835_ (.B1(_06332_),
    .Y(_06333_),
    .A1(net5675),
    .A2(net2819));
 sg13g2_mux2_1 _22836_ (.A0(net3195),
    .A1(net2259),
    .S(net5675),
    .X(_06334_));
 sg13g2_o21ai_1 _22837_ (.B1(net5670),
    .Y(_06335_),
    .A1(net5671),
    .A2(_06333_));
 sg13g2_a21oi_1 _22838_ (.A1(net5671),
    .A2(_06334_),
    .Y(_06336_),
    .B1(_06335_));
 sg13g2_nor3_1 _22839_ (.A(net5338),
    .B(_06331_),
    .C(_06336_),
    .Y(_06337_));
 sg13g2_a21o_1 _22840_ (.A2(net5337),
    .A1(net6311),
    .B1(_06337_),
    .X(_02219_));
 sg13g2_mux4_1 _22841_ (.S0(net5676),
    .A0(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][7] ),
    .A1(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][7] ),
    .A2(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][7] ),
    .A3(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][7] ),
    .S1(net5671),
    .X(_06338_));
 sg13g2_nor2_1 _22842_ (.A(net5670),
    .B(_06338_),
    .Y(_06339_));
 sg13g2_nand2b_1 _22843_ (.Y(_06340_),
    .B(net5675),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][7] ));
 sg13g2_o21ai_1 _22844_ (.B1(_06340_),
    .Y(_06341_),
    .A1(net5675),
    .A2(net3162));
 sg13g2_mux2_1 _22845_ (.A0(net2536),
    .A1(net2165),
    .S(net5675),
    .X(_06342_));
 sg13g2_o21ai_1 _22846_ (.B1(net5670),
    .Y(_06343_),
    .A1(net5671),
    .A2(_06341_));
 sg13g2_a21oi_1 _22847_ (.A1(net5671),
    .A2(_06342_),
    .Y(_06344_),
    .B1(_06343_));
 sg13g2_nor3_1 _22848_ (.A(net5338),
    .B(_06339_),
    .C(_06344_),
    .Y(_06345_));
 sg13g2_a21o_1 _22849_ (.A2(net5338),
    .A1(net6310),
    .B1(_06345_),
    .X(_02220_));
 sg13g2_nor2b_1 _22850_ (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[0] ),
    .B_N(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[1] ),
    .Y(_06346_));
 sg13g2_nand3_1 _22851_ (.B(_03640_),
    .C(_06346_),
    .A(net5668),
    .Y(_06347_));
 sg13g2_mux2_1 _22852_ (.A0(net5612),
    .A1(net2667),
    .S(_06347_),
    .X(_02221_));
 sg13g2_mux2_1 _22853_ (.A0(net5611),
    .A1(net2804),
    .S(_06347_),
    .X(_02222_));
 sg13g2_mux2_1 _22854_ (.A0(net5610),
    .A1(net2774),
    .S(_06347_),
    .X(_02223_));
 sg13g2_mux2_1 _22855_ (.A0(net5609),
    .A1(net3343),
    .S(_06347_),
    .X(_02224_));
 sg13g2_mux2_1 _22856_ (.A0(net5608),
    .A1(net3447),
    .S(_06347_),
    .X(_02225_));
 sg13g2_mux2_1 _22857_ (.A0(net5607),
    .A1(net2905),
    .S(_06347_),
    .X(_02226_));
 sg13g2_mux2_1 _22858_ (.A0(net5606),
    .A1(net3195),
    .S(_06347_),
    .X(_02227_));
 sg13g2_mux2_1 _22859_ (.A0(net5605),
    .A1(net2536),
    .S(_06347_),
    .X(_02228_));
 sg13g2_nand3b_1 _22860_ (.B(net5668),
    .C(_03641_),
    .Y(_06348_),
    .A_N(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[1] ));
 sg13g2_mux2_1 _22861_ (.A0(net5612),
    .A1(net2120),
    .S(_06348_),
    .X(_02229_));
 sg13g2_mux2_1 _22862_ (.A0(net5611),
    .A1(net2280),
    .S(_06348_),
    .X(_02230_));
 sg13g2_mux2_1 _22863_ (.A0(net5610),
    .A1(net2203),
    .S(_06348_),
    .X(_02231_));
 sg13g2_mux2_1 _22864_ (.A0(net5609),
    .A1(net2249),
    .S(_06348_),
    .X(_02232_));
 sg13g2_mux2_1 _22865_ (.A0(net5608),
    .A1(net2148),
    .S(_06348_),
    .X(_02233_));
 sg13g2_mux2_1 _22866_ (.A0(net5607),
    .A1(net2107),
    .S(_06348_),
    .X(_02234_));
 sg13g2_mux2_1 _22867_ (.A0(net5606),
    .A1(net2133),
    .S(_06348_),
    .X(_02235_));
 sg13g2_mux2_1 _22868_ (.A0(net5605),
    .A1(net2573),
    .S(_06348_),
    .X(_02236_));
 sg13g2_nor4_1 _22869_ (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[0] ),
    .B(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[1] ),
    .C(_09541_),
    .D(_03639_),
    .Y(_06349_));
 sg13g2_nand2_2 _22870_ (.Y(_06350_),
    .A(net5668),
    .B(_06349_));
 sg13g2_mux2_1 _22871_ (.A0(net5612),
    .A1(net2696),
    .S(_06350_),
    .X(_02237_));
 sg13g2_mux2_1 _22872_ (.A0(net5611),
    .A1(net2975),
    .S(_06350_),
    .X(_02238_));
 sg13g2_mux2_1 _22873_ (.A0(net5610),
    .A1(net2740),
    .S(_06350_),
    .X(_02239_));
 sg13g2_mux2_1 _22874_ (.A0(net5609),
    .A1(net2961),
    .S(_06350_),
    .X(_02240_));
 sg13g2_mux2_1 _22875_ (.A0(net5608),
    .A1(net2550),
    .S(_06350_),
    .X(_02241_));
 sg13g2_mux2_1 _22876_ (.A0(net5607),
    .A1(net2590),
    .S(_06350_),
    .X(_02242_));
 sg13g2_mux2_1 _22877_ (.A0(net5606),
    .A1(net2819),
    .S(_06350_),
    .X(_02243_));
 sg13g2_mux2_1 _22878_ (.A0(net5605),
    .A1(net3162),
    .S(_06350_),
    .X(_02244_));
 sg13g2_mux2_1 _22879_ (.A0(net3556),
    .A1(net5612),
    .S(_03643_),
    .X(_02245_));
 sg13g2_mux2_1 _22880_ (.A0(net3585),
    .A1(net5611),
    .S(_03643_),
    .X(_02246_));
 sg13g2_mux2_1 _22881_ (.A0(net2626),
    .A1(net5610),
    .S(_03643_),
    .X(_02247_));
 sg13g2_mux2_1 _22882_ (.A0(net2945),
    .A1(net5609),
    .S(_03643_),
    .X(_02248_));
 sg13g2_mux2_1 _22883_ (.A0(net2755),
    .A1(net5608),
    .S(_03643_),
    .X(_02249_));
 sg13g2_mux2_1 _22884_ (.A0(net2294),
    .A1(net5607),
    .S(_03643_),
    .X(_02250_));
 sg13g2_mux2_1 _22885_ (.A0(net2530),
    .A1(net5606),
    .S(_03643_),
    .X(_02251_));
 sg13g2_mux2_1 _22886_ (.A0(net2546),
    .A1(net5605),
    .S(_03643_),
    .X(_02252_));
 sg13g2_nand3b_1 _22887_ (.B(_03640_),
    .C(_06346_),
    .Y(_06351_),
    .A_N(net5668));
 sg13g2_mux2_1 _22888_ (.A0(net5612),
    .A1(net3621),
    .S(_06351_),
    .X(_02253_));
 sg13g2_mux2_1 _22889_ (.A0(net5611),
    .A1(net3281),
    .S(_06351_),
    .X(_02254_));
 sg13g2_mux2_1 _22890_ (.A0(net5610),
    .A1(net3070),
    .S(_06351_),
    .X(_02255_));
 sg13g2_mux2_1 _22891_ (.A0(net5609),
    .A1(net2233),
    .S(_06351_),
    .X(_02256_));
 sg13g2_mux2_1 _22892_ (.A0(net5608),
    .A1(net2163),
    .S(_06351_),
    .X(_02257_));
 sg13g2_mux2_1 _22893_ (.A0(net5607),
    .A1(net3017),
    .S(_06351_),
    .X(_02258_));
 sg13g2_mux2_1 _22894_ (.A0(net5606),
    .A1(net3264),
    .S(_06351_),
    .X(_02259_));
 sg13g2_mux2_1 _22895_ (.A0(net5605),
    .A1(net2579),
    .S(_06351_),
    .X(_02260_));
 sg13g2_nor2_1 _22896_ (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[1] ),
    .B(net5668),
    .Y(_06352_));
 sg13g2_nand2_2 _22897_ (.Y(_06353_),
    .A(_03641_),
    .B(_06352_));
 sg13g2_mux2_1 _22898_ (.A0(net5612),
    .A1(net3498),
    .S(_06353_),
    .X(_02261_));
 sg13g2_mux2_1 _22899_ (.A0(\fpga_top.uart_top.uart_if.byte_data[1] ),
    .A1(net2450),
    .S(_06353_),
    .X(_02262_));
 sg13g2_mux2_1 _22900_ (.A0(\fpga_top.uart_top.uart_if.byte_data[2] ),
    .A1(net2456),
    .S(_06353_),
    .X(_02263_));
 sg13g2_mux2_1 _22901_ (.A0(\fpga_top.uart_top.uart_if.byte_data[3] ),
    .A1(net2800),
    .S(_06353_),
    .X(_02264_));
 sg13g2_mux2_1 _22902_ (.A0(\fpga_top.uart_top.uart_if.byte_data[4] ),
    .A1(net3310),
    .S(_06353_),
    .X(_02265_));
 sg13g2_mux2_1 _22903_ (.A0(net5607),
    .A1(net3507),
    .S(_06353_),
    .X(_02266_));
 sg13g2_mux2_1 _22904_ (.A0(net5606),
    .A1(net3555),
    .S(_06353_),
    .X(_02267_));
 sg13g2_mux2_1 _22905_ (.A0(net5605),
    .A1(net3172),
    .S(_06353_),
    .X(_02268_));
 sg13g2_nor2b_2 _22906_ (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[2] ),
    .B_N(_06349_),
    .Y(_06354_));
 sg13g2_mux2_1 _22907_ (.A0(net2566),
    .A1(\fpga_top.uart_top.uart_if.byte_data[0] ),
    .S(_06354_),
    .X(_02269_));
 sg13g2_mux2_1 _22908_ (.A0(net2918),
    .A1(\fpga_top.uart_top.uart_if.byte_data[1] ),
    .S(_06354_),
    .X(_02270_));
 sg13g2_mux2_1 _22909_ (.A0(net2338),
    .A1(\fpga_top.uart_top.uart_if.byte_data[2] ),
    .S(_06354_),
    .X(_02271_));
 sg13g2_mux2_1 _22910_ (.A0(net3308),
    .A1(\fpga_top.uart_top.uart_if.byte_data[3] ),
    .S(_06354_),
    .X(_02272_));
 sg13g2_mux2_1 _22911_ (.A0(net3040),
    .A1(\fpga_top.uart_top.uart_if.byte_data[4] ),
    .S(_06354_),
    .X(_02273_));
 sg13g2_mux2_1 _22912_ (.A0(net2174),
    .A1(\fpga_top.uart_top.uart_if.byte_data[5] ),
    .S(_06354_),
    .X(_02274_));
 sg13g2_mux2_1 _22913_ (.A0(net3670),
    .A1(net5606),
    .S(_06354_),
    .X(_02275_));
 sg13g2_mux2_1 _22914_ (.A0(net3631),
    .A1(net5605),
    .S(_06354_),
    .X(_02276_));
 sg13g2_nand3_1 _22915_ (.B(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[2] ),
    .C(_03029_),
    .A(net2062),
    .Y(_06355_));
 sg13g2_nand2_1 _22916_ (.Y(_06356_),
    .A(net1487),
    .B(net4412));
 sg13g2_o21ai_1 _22917_ (.B1(_06356_),
    .Y(_02277_),
    .A1(net4921),
    .A2(net4412));
 sg13g2_nand2_1 _22918_ (.Y(_06357_),
    .A(net1557),
    .B(net4413));
 sg13g2_o21ai_1 _22919_ (.B1(net1558),
    .Y(_02278_),
    .A1(net4916),
    .A2(net4413));
 sg13g2_nand2_1 _22920_ (.Y(_06358_),
    .A(net1472),
    .B(net4412));
 sg13g2_o21ai_1 _22921_ (.B1(_06358_),
    .Y(_02279_),
    .A1(net4849),
    .A2(net4412));
 sg13g2_mux2_1 _22922_ (.A0(net4841),
    .A1(net2291),
    .S(net4412),
    .X(_02280_));
 sg13g2_mux2_1 _22923_ (.A0(net4837),
    .A1(net3251),
    .S(net4413),
    .X(_02281_));
 sg13g2_nand2_1 _22924_ (.Y(_06359_),
    .A(net1419),
    .B(net4413));
 sg13g2_o21ai_1 _22925_ (.B1(net1420),
    .Y(_02282_),
    .A1(net4835),
    .A2(net4413));
 sg13g2_nand2_1 _22926_ (.Y(_06360_),
    .A(net1460),
    .B(net4412));
 sg13g2_o21ai_1 _22927_ (.B1(_06360_),
    .Y(_02283_),
    .A1(net4832),
    .A2(net4412));
 sg13g2_nand2_1 _22928_ (.Y(_06361_),
    .A(net1448),
    .B(net4412));
 sg13g2_o21ai_1 _22929_ (.B1(_06361_),
    .Y(_02284_),
    .A1(net4830),
    .A2(net4413));
 sg13g2_nor3_2 _22930_ (.A(net6598),
    .B(_06928_),
    .C(_03031_),
    .Y(_06362_));
 sg13g2_nor2_1 _22931_ (.A(net2056),
    .B(net4410),
    .Y(_06363_));
 sg13g2_a21oi_1 _22932_ (.A1(net4921),
    .A2(net4410),
    .Y(_02285_),
    .B1(net2057));
 sg13g2_nor2_1 _22933_ (.A(net1744),
    .B(net4411),
    .Y(_06364_));
 sg13g2_a21oi_1 _22934_ (.A1(net4916),
    .A2(net4411),
    .Y(_02286_),
    .B1(net1745));
 sg13g2_nor2_1 _22935_ (.A(net2351),
    .B(net4410),
    .Y(_06365_));
 sg13g2_a21oi_1 _22936_ (.A1(net4849),
    .A2(net4410),
    .Y(_02287_),
    .B1(net2352));
 sg13g2_mux2_1 _22937_ (.A0(net2393),
    .A1(net4841),
    .S(net4410),
    .X(_02288_));
 sg13g2_mux2_1 _22938_ (.A0(net2246),
    .A1(net4837),
    .S(net4411),
    .X(_02289_));
 sg13g2_nor2_1 _22939_ (.A(net1889),
    .B(net4411),
    .Y(_06366_));
 sg13g2_a21oi_1 _22940_ (.A1(net4835),
    .A2(net4411),
    .Y(_02290_),
    .B1(net1890));
 sg13g2_nor2_1 _22941_ (.A(net2029),
    .B(net4410),
    .Y(_06367_));
 sg13g2_a21oi_1 _22942_ (.A1(net4832),
    .A2(net4410),
    .Y(_02291_),
    .B1(net2030));
 sg13g2_nor2_1 _22943_ (.A(net2156),
    .B(net4411),
    .Y(_06368_));
 sg13g2_a21oi_1 _22944_ (.A1(net4830),
    .A2(net4410),
    .Y(_02292_),
    .B1(net2157));
 sg13g2_and3_1 _22945_ (.X(_06369_),
    .A(net6598),
    .B(net6601),
    .C(_03030_));
 sg13g2_nor2_1 _22946_ (.A(net1728),
    .B(net4425),
    .Y(_06370_));
 sg13g2_a21oi_1 _22947_ (.A1(net4921),
    .A2(net4425),
    .Y(_02293_),
    .B1(_06370_));
 sg13g2_nor2_1 _22948_ (.A(net1906),
    .B(net4426),
    .Y(_06371_));
 sg13g2_a21oi_1 _22949_ (.A1(net4916),
    .A2(net4426),
    .Y(_02294_),
    .B1(net1907));
 sg13g2_nor2_1 _22950_ (.A(net1804),
    .B(net4425),
    .Y(_06372_));
 sg13g2_a21oi_1 _22951_ (.A1(net4849),
    .A2(net4425),
    .Y(_02295_),
    .B1(_06372_));
 sg13g2_mux2_1 _22952_ (.A0(net3220),
    .A1(net4841),
    .S(net4425),
    .X(_02296_));
 sg13g2_mux2_1 _22953_ (.A0(net2864),
    .A1(net4837),
    .S(net4426),
    .X(_02297_));
 sg13g2_nor2_1 _22954_ (.A(net2051),
    .B(net4426),
    .Y(_06373_));
 sg13g2_a21oi_1 _22955_ (.A1(net4835),
    .A2(net4426),
    .Y(_02298_),
    .B1(_06373_));
 sg13g2_nor2_1 _22956_ (.A(net2145),
    .B(net4425),
    .Y(_06374_));
 sg13g2_a21oi_1 _22957_ (.A1(net4832),
    .A2(net4425),
    .Y(_02299_),
    .B1(_06374_));
 sg13g2_nor2_1 _22958_ (.A(net1870),
    .B(net4425),
    .Y(_06375_));
 sg13g2_a21oi_1 _22959_ (.A1(net4830),
    .A2(net4426),
    .Y(_02300_),
    .B1(_06375_));
 sg13g2_nand3b_1 _22960_ (.B(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[2] ),
    .C(_03030_),
    .Y(_06376_),
    .A_N(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[0] ));
 sg13g2_mux2_1 _22961_ (.A0(_10526_),
    .A1(net2748),
    .S(_06376_),
    .X(_02301_));
 sg13g2_mux2_1 _22962_ (.A0(net4845),
    .A1(net2434),
    .S(_06376_),
    .X(_02302_));
 sg13g2_mux2_1 _22963_ (.A0(_08915_),
    .A1(net2490),
    .S(_06376_),
    .X(_02303_));
 sg13g2_mux2_1 _22964_ (.A0(net4841),
    .A1(net3363),
    .S(_06376_),
    .X(_02304_));
 sg13g2_mux2_1 _22965_ (.A0(net4837),
    .A1(net2205),
    .S(_06376_),
    .X(_02305_));
 sg13g2_mux2_1 _22966_ (.A0(net4834),
    .A1(net2802),
    .S(_06376_),
    .X(_02306_));
 sg13g2_mux2_1 _22967_ (.A0(_02756_),
    .A1(net3077),
    .S(_06376_),
    .X(_02307_));
 sg13g2_mux2_1 _22968_ (.A0(_02760_),
    .A1(net3291),
    .S(_06376_),
    .X(_02308_));
 sg13g2_nand2_1 _22969_ (.Y(_06377_),
    .A(net1425),
    .B(net4421));
 sg13g2_o21ai_1 _22970_ (.B1(_06377_),
    .Y(_02309_),
    .A1(net4921),
    .A2(net4421));
 sg13g2_nand2_1 _22971_ (.Y(_06378_),
    .A(net1453),
    .B(net4422));
 sg13g2_o21ai_1 _22972_ (.B1(_06378_),
    .Y(_02310_),
    .A1(net4916),
    .A2(net4422));
 sg13g2_nand2_1 _22973_ (.Y(_06379_),
    .A(net1522),
    .B(net4422));
 sg13g2_o21ai_1 _22974_ (.B1(_06379_),
    .Y(_02311_),
    .A1(net4849),
    .A2(net4421));
 sg13g2_mux2_1 _22975_ (.A0(net4841),
    .A1(net2870),
    .S(net4422),
    .X(_02312_));
 sg13g2_mux2_1 _22976_ (.A0(net4837),
    .A1(net2941),
    .S(net4421),
    .X(_02313_));
 sg13g2_nand2_1 _22977_ (.Y(_06380_),
    .A(net1470),
    .B(net4422));
 sg13g2_o21ai_1 _22978_ (.B1(_06380_),
    .Y(_02314_),
    .A1(net4835),
    .A2(net4422));
 sg13g2_nand2_1 _22979_ (.Y(_06381_),
    .A(net1480),
    .B(net4421));
 sg13g2_o21ai_1 _22980_ (.B1(_06381_),
    .Y(_02315_),
    .A1(net4832),
    .A2(net4421));
 sg13g2_nand2_1 _22981_ (.Y(_06382_),
    .A(net1458),
    .B(net4421));
 sg13g2_o21ai_1 _22982_ (.B1(_06382_),
    .Y(_02316_),
    .A1(net4830),
    .A2(net4421));
 sg13g2_nor3_2 _22983_ (.A(net6617),
    .B(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[2] ),
    .C(_03031_),
    .Y(_06383_));
 sg13g2_nor2_1 _22984_ (.A(net1920),
    .B(net4408),
    .Y(_06384_));
 sg13g2_a21oi_1 _22985_ (.A1(net4921),
    .A2(net4408),
    .Y(_02317_),
    .B1(net1921));
 sg13g2_nor2_1 _22986_ (.A(net1747),
    .B(net4409),
    .Y(_06385_));
 sg13g2_a21oi_1 _22987_ (.A1(net4916),
    .A2(net4409),
    .Y(_02318_),
    .B1(net1748));
 sg13g2_nor2_1 _22988_ (.A(net1765),
    .B(net4409),
    .Y(_06386_));
 sg13g2_a21oi_1 _22989_ (.A1(net4849),
    .A2(net4408),
    .Y(_02319_),
    .B1(net1766));
 sg13g2_mux2_1 _22990_ (.A0(net2985),
    .A1(net4841),
    .S(net4409),
    .X(_02320_));
 sg13g2_mux2_1 _22991_ (.A0(net2296),
    .A1(net4837),
    .S(net4408),
    .X(_02321_));
 sg13g2_nor2_1 _22992_ (.A(net1798),
    .B(net4409),
    .Y(_06387_));
 sg13g2_a21oi_1 _22993_ (.A1(net4835),
    .A2(net4409),
    .Y(_02322_),
    .B1(net1799));
 sg13g2_nor2_1 _22994_ (.A(net1827),
    .B(net4408),
    .Y(_06388_));
 sg13g2_a21oi_1 _22995_ (.A1(net4832),
    .A2(net4408),
    .Y(_02323_),
    .B1(net1828));
 sg13g2_nor2_1 _22996_ (.A(net1652),
    .B(net4408),
    .Y(_06389_));
 sg13g2_a21oi_1 _22997_ (.A1(net4830),
    .A2(net4408),
    .Y(_02324_),
    .B1(net1653));
 sg13g2_and3_2 _22998_ (.X(_06390_),
    .A(net6598),
    .B(_06928_),
    .C(_03030_));
 sg13g2_nor2_1 _22999_ (.A(net2477),
    .B(net4423),
    .Y(_06391_));
 sg13g2_a21oi_1 _23000_ (.A1(net4921),
    .A2(net4423),
    .Y(_02325_),
    .B1(_06391_));
 sg13g2_nor2_1 _23001_ (.A(net1825),
    .B(net4424),
    .Y(_06392_));
 sg13g2_a21oi_1 _23002_ (.A1(net4916),
    .A2(net4424),
    .Y(_02326_),
    .B1(_06392_));
 sg13g2_nor2_1 _23003_ (.A(net1723),
    .B(net4424),
    .Y(_06393_));
 sg13g2_a21oi_1 _23004_ (.A1(net4849),
    .A2(net4423),
    .Y(_02327_),
    .B1(_06393_));
 sg13g2_mux2_1 _23005_ (.A0(net2762),
    .A1(net4841),
    .S(net4424),
    .X(_02328_));
 sg13g2_mux2_1 _23006_ (.A0(net3318),
    .A1(net4837),
    .S(net4423),
    .X(_02329_));
 sg13g2_nor2_1 _23007_ (.A(net1769),
    .B(net4424),
    .Y(_06394_));
 sg13g2_a21oi_1 _23008_ (.A1(net4835),
    .A2(net4424),
    .Y(_02330_),
    .B1(_06394_));
 sg13g2_nor2_1 _23009_ (.A(net1884),
    .B(net4423),
    .Y(_06395_));
 sg13g2_a21oi_1 _23010_ (.A1(net4832),
    .A2(net4423),
    .Y(_02331_),
    .B1(_06395_));
 sg13g2_nor2_1 _23011_ (.A(net1928),
    .B(net4423),
    .Y(_06396_));
 sg13g2_a21oi_1 _23012_ (.A1(net4830),
    .A2(net4423),
    .Y(_02332_),
    .B1(_06396_));
 sg13g2_nand3b_1 _23013_ (.B(_06928_),
    .C(_03030_),
    .Y(_06397_),
    .A_N(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[0] ));
 sg13g2_mux2_1 _23014_ (.A0(_10526_),
    .A1(net2224),
    .S(_06397_),
    .X(_02333_));
 sg13g2_mux2_1 _23015_ (.A0(net4845),
    .A1(net3522),
    .S(_06397_),
    .X(_02334_));
 sg13g2_mux2_1 _23016_ (.A0(_08915_),
    .A1(net3611),
    .S(_06397_),
    .X(_02335_));
 sg13g2_mux2_1 _23017_ (.A0(net4841),
    .A1(net3639),
    .S(_06397_),
    .X(_02336_));
 sg13g2_mux2_1 _23018_ (.A0(net4837),
    .A1(net2716),
    .S(_06397_),
    .X(_02337_));
 sg13g2_mux2_1 _23019_ (.A0(net4834),
    .A1(net3087),
    .S(_06397_),
    .X(_02338_));
 sg13g2_mux2_1 _23020_ (.A0(_02756_),
    .A1(net2877),
    .S(_06397_),
    .X(_02339_));
 sg13g2_mux2_1 _23021_ (.A0(_02760_),
    .A1(net2782),
    .S(_06397_),
    .X(_02340_));
 sg13g2_nor2b_1 _23022_ (.A(net5827),
    .B_N(\fpga_top.io_spi_lite.miso_byte_org[0] ),
    .Y(_06398_));
 sg13g2_a21oi_2 _23023_ (.B1(_06398_),
    .Y(_06399_),
    .A2(\fpga_top.io_spi_lite.miso_byte_org[7] ),
    .A1(net5827));
 sg13g2_nand2_1 _23024_ (.Y(_06400_),
    .A(net1564),
    .B(net5269));
 sg13g2_o21ai_1 _23025_ (.B1(_06400_),
    .Y(_02341_),
    .A1(net5269),
    .A2(_06399_));
 sg13g2_nor2b_1 _23026_ (.A(net5829),
    .B_N(\fpga_top.io_spi_lite.miso_byte_org[1] ),
    .Y(_06401_));
 sg13g2_a21oi_2 _23027_ (.B1(_06401_),
    .Y(_06402_),
    .A2(\fpga_top.io_spi_lite.miso_byte_org[6] ),
    .A1(net5829));
 sg13g2_nand2_1 _23028_ (.Y(_06403_),
    .A(net1526),
    .B(net5270));
 sg13g2_o21ai_1 _23029_ (.B1(_06403_),
    .Y(_02342_),
    .A1(net5270),
    .A2(_06402_));
 sg13g2_nor2b_1 _23030_ (.A(net5827),
    .B_N(\fpga_top.io_spi_lite.miso_byte_org[2] ),
    .Y(_06404_));
 sg13g2_a21oi_2 _23031_ (.B1(_06404_),
    .Y(_06405_),
    .A2(\fpga_top.io_spi_lite.miso_byte_org[5] ),
    .A1(net5827));
 sg13g2_nand2_1 _23032_ (.Y(_06406_),
    .A(net1398),
    .B(net5268));
 sg13g2_o21ai_1 _23033_ (.B1(_06406_),
    .Y(_02343_),
    .A1(net5268),
    .A2(_06405_));
 sg13g2_nor2b_1 _23034_ (.A(net5829),
    .B_N(\fpga_top.io_spi_lite.miso_byte_org[3] ),
    .Y(_06407_));
 sg13g2_a21oi_2 _23035_ (.B1(_06407_),
    .Y(_06408_),
    .A2(\fpga_top.io_spi_lite.miso_byte_org[4] ),
    .A1(net5829));
 sg13g2_nand2_1 _23036_ (.Y(_06409_),
    .A(net1483),
    .B(net5270));
 sg13g2_o21ai_1 _23037_ (.B1(_06409_),
    .Y(_02344_),
    .A1(net5270),
    .A2(_06408_));
 sg13g2_nor2b_1 _23038_ (.A(net5828),
    .B_N(\fpga_top.io_spi_lite.miso_byte_org[4] ),
    .Y(_06410_));
 sg13g2_a21oi_2 _23039_ (.B1(_06410_),
    .Y(_06411_),
    .A2(\fpga_top.io_spi_lite.miso_byte_org[3] ),
    .A1(net5828));
 sg13g2_nand2_1 _23040_ (.Y(_06412_),
    .A(net1413),
    .B(net5269));
 sg13g2_o21ai_1 _23041_ (.B1(_06412_),
    .Y(_02345_),
    .A1(net5269),
    .A2(_06411_));
 sg13g2_nor2b_1 _23042_ (.A(net5827),
    .B_N(\fpga_top.io_spi_lite.miso_byte_org[5] ),
    .Y(_06413_));
 sg13g2_a21oi_2 _23043_ (.B1(_06413_),
    .Y(_06414_),
    .A2(\fpga_top.io_spi_lite.miso_byte_org[2] ),
    .A1(net5827));
 sg13g2_nand2_1 _23044_ (.Y(_06415_),
    .A(net1434),
    .B(net5268));
 sg13g2_o21ai_1 _23045_ (.B1(_06415_),
    .Y(_02346_),
    .A1(net5268),
    .A2(_06414_));
 sg13g2_nor2b_1 _23046_ (.A(net5828),
    .B_N(\fpga_top.io_spi_lite.miso_byte_org[6] ),
    .Y(_06416_));
 sg13g2_a21oi_2 _23047_ (.B1(_06416_),
    .Y(_06417_),
    .A2(\fpga_top.io_spi_lite.miso_byte_org[1] ),
    .A1(net5828));
 sg13g2_nand2_1 _23048_ (.Y(_06418_),
    .A(net1422),
    .B(net5268));
 sg13g2_o21ai_1 _23049_ (.B1(_06418_),
    .Y(_02347_),
    .A1(net5268),
    .A2(_06417_));
 sg13g2_nor2b_1 _23050_ (.A(net5827),
    .B_N(\fpga_top.io_spi_lite.miso_byte_org[7] ),
    .Y(_06419_));
 sg13g2_a21oi_2 _23051_ (.B1(_06419_),
    .Y(_06420_),
    .A2(\fpga_top.io_spi_lite.miso_byte_org[0] ),
    .A1(net5827));
 sg13g2_nand2_1 _23052_ (.Y(_06421_),
    .A(net1493),
    .B(net5268));
 sg13g2_o21ai_1 _23053_ (.B1(_06421_),
    .Y(_02348_),
    .A1(net5268),
    .A2(_06420_));
 sg13g2_nor3_1 _23054_ (.A(_06786_),
    .B(_06787_),
    .C(_10578_),
    .Y(_06422_));
 sg13g2_nor2_1 _23055_ (.A(net1925),
    .B(net5251),
    .Y(_06423_));
 sg13g2_a21oi_1 _23056_ (.A1(_06399_),
    .A2(net5251),
    .Y(_02349_),
    .B1(_06423_));
 sg13g2_nor2_1 _23057_ (.A(net2059),
    .B(net5252),
    .Y(_06424_));
 sg13g2_a21oi_1 _23058_ (.A1(_06402_),
    .A2(net5252),
    .Y(_02350_),
    .B1(net2060));
 sg13g2_nor2_1 _23059_ (.A(net1754),
    .B(net5250),
    .Y(_06425_));
 sg13g2_a21oi_1 _23060_ (.A1(_06405_),
    .A2(net5250),
    .Y(_02351_),
    .B1(_06425_));
 sg13g2_nor2_1 _23061_ (.A(net2044),
    .B(net5252),
    .Y(_06426_));
 sg13g2_a21oi_1 _23062_ (.A1(_06408_),
    .A2(net5252),
    .Y(_02352_),
    .B1(net2045));
 sg13g2_nor2_1 _23063_ (.A(net1665),
    .B(net5251),
    .Y(_06427_));
 sg13g2_a21oi_1 _23064_ (.A1(_06411_),
    .A2(net5251),
    .Y(_02353_),
    .B1(_06427_));
 sg13g2_nor2_1 _23065_ (.A(net1627),
    .B(net5250),
    .Y(_06428_));
 sg13g2_a21oi_1 _23066_ (.A1(_06414_),
    .A2(net5250),
    .Y(_02354_),
    .B1(_06428_));
 sg13g2_nor2_1 _23067_ (.A(net1882),
    .B(net5250),
    .Y(_06429_));
 sg13g2_a21oi_1 _23068_ (.A1(_06417_),
    .A2(net5250),
    .Y(_02355_),
    .B1(_06429_));
 sg13g2_nor2_1 _23069_ (.A(net1912),
    .B(net5250),
    .Y(_06430_));
 sg13g2_a21oi_1 _23070_ (.A1(_06420_),
    .A2(net5250),
    .Y(_02356_),
    .B1(_06430_));
 sg13g2_nor3_1 _23071_ (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ),
    .B(_06787_),
    .C(_10576_),
    .Y(_06431_));
 sg13g2_nor2_1 _23072_ (.A(net2478),
    .B(net5248),
    .Y(_06432_));
 sg13g2_a21oi_1 _23073_ (.A1(_06399_),
    .A2(net5248),
    .Y(_02357_),
    .B1(_06432_));
 sg13g2_nor2_1 _23074_ (.A(net1965),
    .B(net5249),
    .Y(_06433_));
 sg13g2_a21oi_1 _23075_ (.A1(_06402_),
    .A2(net5249),
    .Y(_02358_),
    .B1(net1966));
 sg13g2_nor2_1 _23076_ (.A(net2093),
    .B(net5247),
    .Y(_06434_));
 sg13g2_a21oi_1 _23077_ (.A1(_06405_),
    .A2(net5247),
    .Y(_02359_),
    .B1(_06434_));
 sg13g2_nor2_1 _23078_ (.A(net1894),
    .B(net5249),
    .Y(_06435_));
 sg13g2_a21oi_1 _23079_ (.A1(_06408_),
    .A2(net5249),
    .Y(_02360_),
    .B1(net1895));
 sg13g2_nor2_1 _23080_ (.A(net1770),
    .B(net5248),
    .Y(_06436_));
 sg13g2_a21oi_1 _23081_ (.A1(_06411_),
    .A2(net5248),
    .Y(_02361_),
    .B1(_06436_));
 sg13g2_nor2_1 _23082_ (.A(net2052),
    .B(net5247),
    .Y(_06437_));
 sg13g2_a21oi_1 _23083_ (.A1(_06414_),
    .A2(net5247),
    .Y(_02362_),
    .B1(_06437_));
 sg13g2_nor2_1 _23084_ (.A(net1885),
    .B(net5247),
    .Y(_06438_));
 sg13g2_a21oi_1 _23085_ (.A1(_06417_),
    .A2(net5247),
    .Y(_02363_),
    .B1(_06438_));
 sg13g2_nor2_1 _23086_ (.A(net1805),
    .B(net5247),
    .Y(_06439_));
 sg13g2_a21oi_1 _23087_ (.A1(_06420_),
    .A2(net5247),
    .Y(_02364_),
    .B1(_06439_));
 sg13g2_nor3_1 _23088_ (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ),
    .B(_06787_),
    .C(_10578_),
    .Y(_06440_));
 sg13g2_nor2_1 _23089_ (.A(net1916),
    .B(net5245),
    .Y(_06441_));
 sg13g2_a21oi_1 _23090_ (.A1(_06399_),
    .A2(net5245),
    .Y(_02365_),
    .B1(_06441_));
 sg13g2_nor2_1 _23091_ (.A(net1875),
    .B(net5246),
    .Y(_06442_));
 sg13g2_a21oi_1 _23092_ (.A1(_06402_),
    .A2(net5246),
    .Y(_02366_),
    .B1(net1876));
 sg13g2_nor2_1 _23093_ (.A(net2150),
    .B(net5244),
    .Y(_06443_));
 sg13g2_a21oi_1 _23094_ (.A1(_06405_),
    .A2(net5244),
    .Y(_02367_),
    .B1(_06443_));
 sg13g2_nor2_1 _23095_ (.A(net1636),
    .B(net5246),
    .Y(_06444_));
 sg13g2_a21oi_1 _23096_ (.A1(_06408_),
    .A2(net5246),
    .Y(_02368_),
    .B1(net1637));
 sg13g2_nor2_1 _23097_ (.A(net2012),
    .B(net5245),
    .Y(_06445_));
 sg13g2_a21oi_1 _23098_ (.A1(_06411_),
    .A2(net5245),
    .Y(_02369_),
    .B1(_06445_));
 sg13g2_nor2_1 _23099_ (.A(net1649),
    .B(net5244),
    .Y(_06446_));
 sg13g2_a21oi_1 _23100_ (.A1(_06414_),
    .A2(net5244),
    .Y(_02370_),
    .B1(_06446_));
 sg13g2_nor2_1 _23101_ (.A(net1734),
    .B(net5244),
    .Y(_06447_));
 sg13g2_a21oi_1 _23102_ (.A1(_06417_),
    .A2(net5244),
    .Y(_02371_),
    .B1(_06447_));
 sg13g2_nor2_1 _23103_ (.A(net1671),
    .B(net5244),
    .Y(_06448_));
 sg13g2_a21oi_1 _23104_ (.A1(_06420_),
    .A2(net5244),
    .Y(_02372_),
    .B1(_06448_));
 sg13g2_nor2_1 _23105_ (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[2] ),
    .B(_10579_),
    .Y(_06449_));
 sg13g2_nor2_1 _23106_ (.A(net1729),
    .B(net5243),
    .Y(_06450_));
 sg13g2_a21oi_1 _23107_ (.A1(_06399_),
    .A2(net5243),
    .Y(_02373_),
    .B1(net1730));
 sg13g2_nor2_1 _23108_ (.A(net1607),
    .B(net5243),
    .Y(_06451_));
 sg13g2_a21oi_1 _23109_ (.A1(_06402_),
    .A2(net5243),
    .Y(_02374_),
    .B1(net1608));
 sg13g2_nor2_1 _23110_ (.A(net1952),
    .B(net5242),
    .Y(_06452_));
 sg13g2_a21oi_1 _23111_ (.A1(_06405_),
    .A2(net5242),
    .Y(_02375_),
    .B1(_06452_));
 sg13g2_nor2_1 _23112_ (.A(net1673),
    .B(net5243),
    .Y(_06453_));
 sg13g2_a21oi_1 _23113_ (.A1(_06408_),
    .A2(net5243),
    .Y(_02376_),
    .B1(net1674));
 sg13g2_nor2_1 _23114_ (.A(net2016),
    .B(net5243),
    .Y(_06454_));
 sg13g2_a21oi_1 _23115_ (.A1(_06411_),
    .A2(_06449_),
    .Y(_02377_),
    .B1(net2017));
 sg13g2_nor2_1 _23116_ (.A(net2036),
    .B(net5242),
    .Y(_06455_));
 sg13g2_a21oi_1 _23117_ (.A1(_06414_),
    .A2(net5242),
    .Y(_02378_),
    .B1(_06455_));
 sg13g2_nor2_1 _23118_ (.A(net1790),
    .B(net5242),
    .Y(_06456_));
 sg13g2_a21oi_1 _23119_ (.A1(_06417_),
    .A2(net5242),
    .Y(_02379_),
    .B1(_06456_));
 sg13g2_nor2_1 _23120_ (.A(net1761),
    .B(net5242),
    .Y(_06457_));
 sg13g2_a21oi_1 _23121_ (.A1(_06420_),
    .A2(net5242),
    .Y(_02380_),
    .B1(_06457_));
 sg13g2_nor3_1 _23122_ (.A(_06786_),
    .B(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[2] ),
    .C(_10578_),
    .Y(_06458_));
 sg13g2_nor2_1 _23123_ (.A(net1662),
    .B(net5241),
    .Y(_06459_));
 sg13g2_a21oi_1 _23124_ (.A1(_06399_),
    .A2(net5241),
    .Y(_02381_),
    .B1(net1663));
 sg13g2_nor2_1 _23125_ (.A(net1720),
    .B(net5241),
    .Y(_06460_));
 sg13g2_a21oi_1 _23126_ (.A1(_06402_),
    .A2(net5241),
    .Y(_02382_),
    .B1(net1721));
 sg13g2_nor2_1 _23127_ (.A(net1775),
    .B(net5240),
    .Y(_06461_));
 sg13g2_a21oi_1 _23128_ (.A1(_06405_),
    .A2(net5240),
    .Y(_02383_),
    .B1(_06461_));
 sg13g2_nor2_1 _23129_ (.A(net1708),
    .B(net5241),
    .Y(_06462_));
 sg13g2_a21oi_1 _23130_ (.A1(_06408_),
    .A2(net5241),
    .Y(_02384_),
    .B1(net1709));
 sg13g2_nor2_1 _23131_ (.A(net2524),
    .B(_06458_),
    .Y(_06463_));
 sg13g2_a21oi_1 _23132_ (.A1(_06411_),
    .A2(net5241),
    .Y(_02385_),
    .B1(net2525));
 sg13g2_nor2_1 _23133_ (.A(net1871),
    .B(net5240),
    .Y(_06464_));
 sg13g2_a21oi_1 _23134_ (.A1(_06414_),
    .A2(net5240),
    .Y(_02386_),
    .B1(_06464_));
 sg13g2_nor2_1 _23135_ (.A(net1701),
    .B(net5240),
    .Y(_06465_));
 sg13g2_a21oi_1 _23136_ (.A1(_06417_),
    .A2(net5240),
    .Y(_02387_),
    .B1(_06465_));
 sg13g2_nor2_1 _23137_ (.A(net1773),
    .B(net5240),
    .Y(_06466_));
 sg13g2_a21oi_1 _23138_ (.A1(_06420_),
    .A2(net5240),
    .Y(_02388_),
    .B1(_06466_));
 sg13g2_nor3_1 _23139_ (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ),
    .B(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[2] ),
    .C(_10576_),
    .Y(_06467_));
 sg13g2_nor2_1 _23140_ (.A(net1961),
    .B(net5239),
    .Y(_06468_));
 sg13g2_a21oi_1 _23141_ (.A1(_06399_),
    .A2(net5239),
    .Y(_02389_),
    .B1(net1962));
 sg13g2_nor2_1 _23142_ (.A(net1725),
    .B(net5239),
    .Y(_06469_));
 sg13g2_a21oi_1 _23143_ (.A1(_06402_),
    .A2(net5239),
    .Y(_02390_),
    .B1(net1726));
 sg13g2_nor2_1 _23144_ (.A(net2034),
    .B(net5238),
    .Y(_06470_));
 sg13g2_a21oi_1 _23145_ (.A1(_06405_),
    .A2(net5238),
    .Y(_02391_),
    .B1(_06470_));
 sg13g2_nor2_1 _23146_ (.A(net1848),
    .B(net5239),
    .Y(_06471_));
 sg13g2_a21oi_1 _23147_ (.A1(_06408_),
    .A2(net5239),
    .Y(_02392_),
    .B1(net1849));
 sg13g2_nor2_1 _23148_ (.A(net2192),
    .B(_06467_),
    .Y(_06472_));
 sg13g2_a21oi_1 _23149_ (.A1(_06411_),
    .A2(net5239),
    .Y(_02393_),
    .B1(net2193));
 sg13g2_nor2_1 _23150_ (.A(net1690),
    .B(net5238),
    .Y(_06473_));
 sg13g2_a21oi_1 _23151_ (.A1(_06414_),
    .A2(net5238),
    .Y(_02394_),
    .B1(_06473_));
 sg13g2_nor2_1 _23152_ (.A(net1815),
    .B(net5238),
    .Y(_06474_));
 sg13g2_a21oi_1 _23153_ (.A1(_06417_),
    .A2(net5238),
    .Y(_02395_),
    .B1(_06474_));
 sg13g2_nor2_1 _23154_ (.A(net1634),
    .B(net5238),
    .Y(_06475_));
 sg13g2_a21oi_1 _23155_ (.A1(_06420_),
    .A2(net5238),
    .Y(_02396_),
    .B1(_06475_));
 sg13g2_nor3_1 _23156_ (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ),
    .B(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[2] ),
    .C(_10578_),
    .Y(_06476_));
 sg13g2_nor2_1 _23157_ (.A(net1617),
    .B(net5237),
    .Y(_06477_));
 sg13g2_a21oi_1 _23158_ (.A1(_06399_),
    .A2(net5237),
    .Y(_02397_),
    .B1(net1618));
 sg13g2_nor2_1 _23159_ (.A(net1696),
    .B(net5237),
    .Y(_06478_));
 sg13g2_a21oi_1 _23160_ (.A1(_06402_),
    .A2(net5237),
    .Y(_02398_),
    .B1(net1697));
 sg13g2_nor2_1 _23161_ (.A(net1763),
    .B(net5236),
    .Y(_06479_));
 sg13g2_a21oi_1 _23162_ (.A1(_06405_),
    .A2(net5236),
    .Y(_02399_),
    .B1(_06479_));
 sg13g2_nor2_1 _23163_ (.A(net1758),
    .B(net5237),
    .Y(_06480_));
 sg13g2_a21oi_1 _23164_ (.A1(_06408_),
    .A2(net5237),
    .Y(_02400_),
    .B1(net1759));
 sg13g2_nor2_1 _23165_ (.A(net1840),
    .B(net5237),
    .Y(_06481_));
 sg13g2_a21oi_1 _23166_ (.A1(_06411_),
    .A2(_06476_),
    .Y(_02401_),
    .B1(net1841));
 sg13g2_nor2_1 _23167_ (.A(net1713),
    .B(net5236),
    .Y(_06482_));
 sg13g2_a21oi_1 _23168_ (.A1(_06414_),
    .A2(net5236),
    .Y(_02402_),
    .B1(_06482_));
 sg13g2_nor2_1 _23169_ (.A(net1750),
    .B(net5236),
    .Y(_06483_));
 sg13g2_a21oi_1 _23170_ (.A1(_06417_),
    .A2(net5236),
    .Y(_02403_),
    .B1(_06483_));
 sg13g2_nor2_1 _23171_ (.A(net1644),
    .B(net5236),
    .Y(_06484_));
 sg13g2_a21oi_1 _23172_ (.A1(_06420_),
    .A2(net5236),
    .Y(_02404_),
    .B1(_06484_));
 sg13g2_nand3_1 _23173_ (.B(_09658_),
    .C(_03179_),
    .A(_09655_),
    .Y(_06485_));
 sg13g2_mux2_1 _23174_ (.A0(net4362),
    .A1(net3111),
    .S(net4210),
    .X(_02405_));
 sg13g2_mux2_1 _23175_ (.A0(net4356),
    .A1(net3141),
    .S(net4212),
    .X(_02406_));
 sg13g2_mux2_1 _23176_ (.A0(net4349),
    .A1(net2159),
    .S(net4211),
    .X(_02407_));
 sg13g2_mux2_1 _23177_ (.A0(net4344),
    .A1(net2887),
    .S(net4210),
    .X(_02408_));
 sg13g2_mux2_1 _23178_ (.A0(net4340),
    .A1(net3294),
    .S(net4212),
    .X(_02409_));
 sg13g2_mux2_1 _23179_ (.A0(net4196),
    .A1(net2664),
    .S(net4212),
    .X(_02410_));
 sg13g2_mux2_1 _23180_ (.A0(net4334),
    .A1(net3673),
    .S(net4211),
    .X(_02411_));
 sg13g2_mux2_1 _23181_ (.A0(net4329),
    .A1(net3405),
    .S(net4213),
    .X(_02412_));
 sg13g2_mux2_1 _23182_ (.A0(net4324),
    .A1(net2719),
    .S(net4212),
    .X(_02413_));
 sg13g2_mux2_1 _23183_ (.A0(net4322),
    .A1(net2920),
    .S(net4211),
    .X(_02414_));
 sg13g2_mux2_1 _23184_ (.A0(net4190),
    .A1(net3396),
    .S(net4213),
    .X(_02415_));
 sg13g2_mux2_1 _23185_ (.A0(net4185),
    .A1(net3249),
    .S(net4210),
    .X(_02416_));
 sg13g2_mux2_1 _23186_ (.A0(net4312),
    .A1(net3202),
    .S(net4213),
    .X(_02417_));
 sg13g2_mux2_1 _23187_ (.A0(net4307),
    .A1(net3003),
    .S(net4210),
    .X(_02418_));
 sg13g2_mux2_1 _23188_ (.A0(net4301),
    .A1(net2273),
    .S(net4210),
    .X(_02419_));
 sg13g2_mux2_1 _23189_ (.A0(net4296),
    .A1(net2422),
    .S(net4213),
    .X(_02420_));
 sg13g2_mux2_1 _23190_ (.A0(net4290),
    .A1(net2272),
    .S(net4214),
    .X(_02421_));
 sg13g2_mux2_1 _23191_ (.A0(net4284),
    .A1(net3122),
    .S(net4210),
    .X(_02422_));
 sg13g2_mux2_1 _23192_ (.A0(net4279),
    .A1(net3412),
    .S(net4214),
    .X(_02423_));
 sg13g2_mux2_1 _23193_ (.A0(net4274),
    .A1(net2252),
    .S(net4212),
    .X(_02424_));
 sg13g2_mux2_1 _23194_ (.A0(net4269),
    .A1(net3609),
    .S(net4212),
    .X(_02425_));
 sg13g2_mux2_1 _23195_ (.A0(net4265),
    .A1(net2899),
    .S(net4210),
    .X(_02426_));
 sg13g2_mux2_1 _23196_ (.A0(net4260),
    .A1(net2467),
    .S(net4214),
    .X(_02427_));
 sg13g2_mux2_1 _23197_ (.A0(net4254),
    .A1(net2729),
    .S(net4213),
    .X(_02428_));
 sg13g2_mux2_1 _23198_ (.A0(net4404),
    .A1(net2513),
    .S(net4213),
    .X(_02429_));
 sg13g2_mux2_1 _23199_ (.A0(net4398),
    .A1(net3435),
    .S(net4212),
    .X(_02430_));
 sg13g2_mux2_1 _23200_ (.A0(net4394),
    .A1(net2686),
    .S(net4211),
    .X(_02431_));
 sg13g2_mux2_1 _23201_ (.A0(net4389),
    .A1(net3320),
    .S(net4210),
    .X(_02432_));
 sg13g2_mux2_1 _23202_ (.A0(net4387),
    .A1(net3290),
    .S(net4211),
    .X(_02433_));
 sg13g2_mux2_1 _23203_ (.A0(net4378),
    .A1(net2873),
    .S(net4213),
    .X(_02434_));
 sg13g2_mux2_1 _23204_ (.A0(net4373),
    .A1(net3300),
    .S(net4212),
    .X(_02435_));
 sg13g2_mux2_1 _23205_ (.A0(net4367),
    .A1(net2783),
    .S(net4213),
    .X(_02436_));
 sg13g2_nor2_2 _23206_ (.A(_08985_),
    .B(_02735_),
    .Y(_06486_));
 sg13g2_nor2_1 _23207_ (.A(net3792),
    .B(net4464),
    .Y(_06487_));
 sg13g2_a21oi_1 _23208_ (.A1(net4920),
    .A2(net4464),
    .Y(_02437_),
    .B1(_06487_));
 sg13g2_nor2_1 _23209_ (.A(net3921),
    .B(net4465),
    .Y(_06488_));
 sg13g2_a21oi_1 _23210_ (.A1(net4917),
    .A2(net4465),
    .Y(_02438_),
    .B1(_06488_));
 sg13g2_nor2_1 _23211_ (.A(net3908),
    .B(net4465),
    .Y(_06489_));
 sg13g2_a21oi_1 _23212_ (.A1(net4852),
    .A2(net4465),
    .Y(_02439_),
    .B1(_06489_));
 sg13g2_mux2_1 _23213_ (.A0(net3987),
    .A1(net4843),
    .S(net4465),
    .X(_02440_));
 sg13g2_mux2_1 _23214_ (.A0(net3931),
    .A1(net4839),
    .S(net4463),
    .X(_02441_));
 sg13g2_nor2_1 _23215_ (.A(net3847),
    .B(net4463),
    .Y(_06490_));
 sg13g2_a21oi_1 _23216_ (.A1(net4835),
    .A2(net4464),
    .Y(_02442_),
    .B1(_06490_));
 sg13g2_nor2_1 _23217_ (.A(net3907),
    .B(net4463),
    .Y(_06491_));
 sg13g2_a21oi_1 _23218_ (.A1(net4832),
    .A2(net4464),
    .Y(_02443_),
    .B1(_06491_));
 sg13g2_nor2_1 _23219_ (.A(net1621),
    .B(net4463),
    .Y(_06492_));
 sg13g2_a21oi_1 _23220_ (.A1(net4830),
    .A2(net4464),
    .Y(_02444_),
    .B1(_06492_));
 sg13g2_nor2_1 _23221_ (.A(net3026),
    .B(net4463),
    .Y(_06493_));
 sg13g2_a21oi_1 _23222_ (.A1(_02763_),
    .A2(net4463),
    .Y(_02445_),
    .B1(_06493_));
 sg13g2_nor2_1 _23223_ (.A(net2047),
    .B(net4463),
    .Y(_06494_));
 sg13g2_a21oi_1 _23224_ (.A1(_02767_),
    .A2(net4463),
    .Y(_02446_),
    .B1(_06494_));
 sg13g2_xor2_1 _23225_ (.B(net5076),
    .A(net1369),
    .X(_02447_));
 sg13g2_or2_1 _23226_ (.X(_06495_),
    .B(_05319_),
    .A(_09659_));
 sg13g2_mux2_1 _23227_ (.A0(net4364),
    .A1(net3189),
    .S(net4080),
    .X(_02448_));
 sg13g2_mux2_1 _23228_ (.A0(net4359),
    .A1(net3430),
    .S(net4082),
    .X(_02449_));
 sg13g2_mux2_1 _23229_ (.A0(net4353),
    .A1(net2218),
    .S(net4081),
    .X(_02450_));
 sg13g2_mux2_1 _23230_ (.A0(net4345),
    .A1(net2406),
    .S(net4080),
    .X(_02451_));
 sg13g2_mux2_1 _23231_ (.A0(net4341),
    .A1(net3229),
    .S(net4082),
    .X(_02452_));
 sg13g2_mux2_1 _23232_ (.A0(net4198),
    .A1(net3149),
    .S(net4082),
    .X(_02453_));
 sg13g2_mux2_1 _23233_ (.A0(net4338),
    .A1(net3287),
    .S(net4080),
    .X(_02454_));
 sg13g2_mux2_1 _23234_ (.A0(net4333),
    .A1(net2844),
    .S(net4083),
    .X(_02455_));
 sg13g2_mux2_1 _23235_ (.A0(net4326),
    .A1(net3603),
    .S(net4084),
    .X(_02456_));
 sg13g2_mux2_1 _23236_ (.A0(net4319),
    .A1(net2217),
    .S(net4081),
    .X(_02457_));
 sg13g2_mux2_1 _23237_ (.A0(net4192),
    .A1(net3000),
    .S(net4083),
    .X(_02458_));
 sg13g2_mux2_1 _23238_ (.A0(net4187),
    .A1(net2581),
    .S(net4081),
    .X(_02459_));
 sg13g2_mux2_1 _23239_ (.A0(net4315),
    .A1(net3089),
    .S(net4083),
    .X(_02460_));
 sg13g2_mux2_1 _23240_ (.A0(net4311),
    .A1(net3440),
    .S(net4081),
    .X(_02461_));
 sg13g2_mux2_1 _23241_ (.A0(net4301),
    .A1(net3257),
    .S(net4080),
    .X(_02462_));
 sg13g2_mux2_1 _23242_ (.A0(net4299),
    .A1(net3233),
    .S(net4084),
    .X(_02463_));
 sg13g2_mux2_1 _23243_ (.A0(net4295),
    .A1(net3060),
    .S(net4083),
    .X(_02464_));
 sg13g2_mux2_1 _23244_ (.A0(net4287),
    .A1(net2670),
    .S(net4080),
    .X(_02465_));
 sg13g2_mux2_1 _23245_ (.A0(net4282),
    .A1(net2403),
    .S(net4083),
    .X(_02466_));
 sg13g2_mux2_1 _23246_ (.A0(net4277),
    .A1(net3478),
    .S(net4080),
    .X(_02467_));
 sg13g2_mux2_1 _23247_ (.A0(net4271),
    .A1(net2610),
    .S(net4082),
    .X(_02468_));
 sg13g2_mux2_1 _23248_ (.A0(net4265),
    .A1(net2482),
    .S(net4080),
    .X(_02469_));
 sg13g2_mux2_1 _23249_ (.A0(net4262),
    .A1(net2387),
    .S(net4082),
    .X(_02470_));
 sg13g2_mux2_1 _23250_ (.A0(net4258),
    .A1(net2168),
    .S(net4083),
    .X(_02471_));
 sg13g2_mux2_1 _23251_ (.A0(net4406),
    .A1(net2779),
    .S(net4083),
    .X(_02472_));
 sg13g2_mux2_1 _23252_ (.A0(net4401),
    .A1(net2401),
    .S(net4082),
    .X(_02473_));
 sg13g2_mux2_1 _23253_ (.A0(net4396),
    .A1(net2996),
    .S(net4081),
    .X(_02474_));
 sg13g2_mux2_1 _23254_ (.A0(net4390),
    .A1(net2921),
    .S(net4080),
    .X(_02475_));
 sg13g2_mux2_1 _23255_ (.A0(net4382),
    .A1(net2196),
    .S(net4081),
    .X(_02476_));
 sg13g2_mux2_1 _23256_ (.A0(net4380),
    .A1(net2583),
    .S(net4083),
    .X(_02477_));
 sg13g2_mux2_1 _23257_ (.A0(net4375),
    .A1(net2220),
    .S(net4082),
    .X(_02478_));
 sg13g2_mux2_1 _23258_ (.A0(net4369),
    .A1(net2458),
    .S(net4082),
    .X(_02479_));
 sg13g2_or2_1 _23259_ (.X(_06496_),
    .B(_05319_),
    .A(_02993_));
 sg13g2_mux2_1 _23260_ (.A0(net4364),
    .A1(net2365),
    .S(net4075),
    .X(_02480_));
 sg13g2_mux2_1 _23261_ (.A0(net4359),
    .A1(net2198),
    .S(net4077),
    .X(_02481_));
 sg13g2_mux2_1 _23262_ (.A0(net4353),
    .A1(net2871),
    .S(net4076),
    .X(_02482_));
 sg13g2_mux2_1 _23263_ (.A0(net4345),
    .A1(net3321),
    .S(net4075),
    .X(_02483_));
 sg13g2_mux2_1 _23264_ (.A0(net4341),
    .A1(net2840),
    .S(net4077),
    .X(_02484_));
 sg13g2_mux2_1 _23265_ (.A0(net4198),
    .A1(net2658),
    .S(net4077),
    .X(_02485_));
 sg13g2_mux2_1 _23266_ (.A0(net4338),
    .A1(net3022),
    .S(net4075),
    .X(_02486_));
 sg13g2_mux2_1 _23267_ (.A0(net4333),
    .A1(net3083),
    .S(net4078),
    .X(_02487_));
 sg13g2_mux2_1 _23268_ (.A0(net4326),
    .A1(net3501),
    .S(net4079),
    .X(_02488_));
 sg13g2_mux2_1 _23269_ (.A0(net4319),
    .A1(net2578),
    .S(net4076),
    .X(_02489_));
 sg13g2_mux2_1 _23270_ (.A0(net4192),
    .A1(net2509),
    .S(net4078),
    .X(_02490_));
 sg13g2_mux2_1 _23271_ (.A0(net4187),
    .A1(net2943),
    .S(net4076),
    .X(_02491_));
 sg13g2_mux2_1 _23272_ (.A0(net4315),
    .A1(net2538),
    .S(net4078),
    .X(_02492_));
 sg13g2_mux2_1 _23273_ (.A0(net4311),
    .A1(net2917),
    .S(net4076),
    .X(_02493_));
 sg13g2_mux2_1 _23274_ (.A0(net4301),
    .A1(net3152),
    .S(net4075),
    .X(_02494_));
 sg13g2_mux2_1 _23275_ (.A0(net4298),
    .A1(net2181),
    .S(net4079),
    .X(_02495_));
 sg13g2_mux2_1 _23276_ (.A0(net4295),
    .A1(net3044),
    .S(net4078),
    .X(_02496_));
 sg13g2_mux2_1 _23277_ (.A0(net4288),
    .A1(net3369),
    .S(net4075),
    .X(_02497_));
 sg13g2_mux2_1 _23278_ (.A0(net4282),
    .A1(net3053),
    .S(net4078),
    .X(_02498_));
 sg13g2_mux2_1 _23279_ (.A0(net4277),
    .A1(net2440),
    .S(net4075),
    .X(_02499_));
 sg13g2_mux2_1 _23280_ (.A0(net4271),
    .A1(net2673),
    .S(net4077),
    .X(_02500_));
 sg13g2_mux2_1 _23281_ (.A0(net4265),
    .A1(net2304),
    .S(net4075),
    .X(_02501_));
 sg13g2_mux2_1 _23282_ (.A0(net4262),
    .A1(net2794),
    .S(net4077),
    .X(_02502_));
 sg13g2_mux2_1 _23283_ (.A0(net4258),
    .A1(net2582),
    .S(net4078),
    .X(_02503_));
 sg13g2_mux2_1 _23284_ (.A0(net4406),
    .A1(net2549),
    .S(net4078),
    .X(_02504_));
 sg13g2_mux2_1 _23285_ (.A0(net4401),
    .A1(net2466),
    .S(net4077),
    .X(_02505_));
 sg13g2_mux2_1 _23286_ (.A0(net4396),
    .A1(net2315),
    .S(net4076),
    .X(_02506_));
 sg13g2_mux2_1 _23287_ (.A0(net4390),
    .A1(net2925),
    .S(net4075),
    .X(_02507_));
 sg13g2_mux2_1 _23288_ (.A0(net4382),
    .A1(net3350),
    .S(net4076),
    .X(_02508_));
 sg13g2_mux2_1 _23289_ (.A0(net4380),
    .A1(net2928),
    .S(net4078),
    .X(_02509_));
 sg13g2_mux2_1 _23290_ (.A0(net4375),
    .A1(net2988),
    .S(net4077),
    .X(_02510_));
 sg13g2_mux2_1 _23291_ (.A0(net4369),
    .A1(net3165),
    .S(net4077),
    .X(_02511_));
 sg13g2_mux2_1 _23292_ (.A0(net4363),
    .A1(net2195),
    .S(net4205),
    .X(_02512_));
 sg13g2_mux2_1 _23293_ (.A0(net4355),
    .A1(net3496),
    .S(net4207),
    .X(_02513_));
 sg13g2_mux2_1 _23294_ (.A0(net4351),
    .A1(net2202),
    .S(net4206),
    .X(_02514_));
 sg13g2_mux2_1 _23295_ (.A0(net4344),
    .A1(net2665),
    .S(net4205),
    .X(_02515_));
 sg13g2_mux2_1 _23296_ (.A0(net4340),
    .A1(net2967),
    .S(net4207),
    .X(_02516_));
 sg13g2_mux2_1 _23297_ (.A0(net4195),
    .A1(net2333),
    .S(net4207),
    .X(_02517_));
 sg13g2_mux2_1 _23298_ (.A0(net4335),
    .A1(net2270),
    .S(net4206),
    .X(_02518_));
 sg13g2_mux2_1 _23299_ (.A0(net4330),
    .A1(net2319),
    .S(net4209),
    .X(_02519_));
 sg13g2_mux2_1 _23300_ (.A0(net4325),
    .A1(net3594),
    .S(net4207),
    .X(_02520_));
 sg13g2_mux2_1 _23301_ (.A0(net4320),
    .A1(net3151),
    .S(net4206),
    .X(_02521_));
 sg13g2_mux2_1 _23302_ (.A0(net4191),
    .A1(net2255),
    .S(net4208),
    .X(_02522_));
 sg13g2_mux2_1 _23303_ (.A0(net4187),
    .A1(net2335),
    .S(net4205),
    .X(_02523_));
 sg13g2_mux2_1 _23304_ (.A0(net4312),
    .A1(net2325),
    .S(net4208),
    .X(_02524_));
 sg13g2_mux2_1 _23305_ (.A0(net4309),
    .A1(net3072),
    .S(net4205),
    .X(_02525_));
 sg13g2_mux2_1 _23306_ (.A0(net4303),
    .A1(net2344),
    .S(net4205),
    .X(_02526_));
 sg13g2_mux2_1 _23307_ (.A0(net4297),
    .A1(net2878),
    .S(net4208),
    .X(_02527_));
 sg13g2_mux2_1 _23308_ (.A0(net4292),
    .A1(net2331),
    .S(net4208),
    .X(_02528_));
 sg13g2_mux2_1 _23309_ (.A0(net4285),
    .A1(net3221),
    .S(net4205),
    .X(_02529_));
 sg13g2_mux2_1 _23310_ (.A0(net4280),
    .A1(net2620),
    .S(net4209),
    .X(_02530_));
 sg13g2_mux2_1 _23311_ (.A0(net4274),
    .A1(net2995),
    .S(net4207),
    .X(_02531_));
 sg13g2_mux2_1 _23312_ (.A0(net4270),
    .A1(net3219),
    .S(net4207),
    .X(_02532_));
 sg13g2_mux2_1 _23313_ (.A0(net4266),
    .A1(net3453),
    .S(net4205),
    .X(_02533_));
 sg13g2_mux2_1 _23314_ (.A0(net4259),
    .A1(net3121),
    .S(net4209),
    .X(_02534_));
 sg13g2_mux2_1 _23315_ (.A0(net4255),
    .A1(net2947),
    .S(net4208),
    .X(_02535_));
 sg13g2_buf_1 _23316_ (.A(net1374),
    .X(_00147_));
 sg13g2_buf_1 _23317_ (.A(net1685),
    .X(_00144_));
 sg13g2_buf_1 _23318_ (.A(net1389),
    .X(_00143_));
 sg13g2_buf_1 _23319_ (.A(net1395),
    .X(_00142_));
 sg13g2_buf_1 _23320_ (.A(net1394),
    .X(_00140_));
 sg13g2_buf_1 _23321_ (.A(net1383),
    .X(_00139_));
 sg13g2_buf_1 _23322_ (.A(net1372),
    .X(_00138_));
 sg13g2_buf_1 _23323_ (.A(net2105),
    .X(_00137_));
 sg13g2_buf_1 _23324_ (.A(net1620),
    .X(_00136_));
 sg13g2_buf_1 _23325_ (.A(net1499),
    .X(_00135_));
 sg13g2_buf_1 _23326_ (.A(net1516),
    .X(_00131_));
 sg13g2_buf_1 _23327_ (.A(net1539),
    .X(_00130_));
 sg13g2_buf_1 _23328_ (.A(net1384),
    .X(_00129_));
 sg13g2_buf_1 _23329_ (.A(net1545),
    .X(_00128_));
 sg13g2_nor3_1 _23330_ (.A(net1396),
    .B(_09638_),
    .C(_09640_),
    .Y(_01301_));
 sg13g2_dfrbpq_1 _23331_ (.RESET_B(net49),
    .D(_00148_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][24] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _23332_ (.RESET_B(net697),
    .D(_00149_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][25] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _23333_ (.RESET_B(net696),
    .D(_00150_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][26] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _23334_ (.RESET_B(net695),
    .D(_00151_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][27] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _23335_ (.RESET_B(net694),
    .D(_00152_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][28] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _23336_ (.RESET_B(net693),
    .D(_00153_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][29] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _23337_ (.RESET_B(net692),
    .D(_00154_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][30] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _23338_ (.RESET_B(net691),
    .D(_00155_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][31] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _23339_ (.RESET_B(net690),
    .D(_00156_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][0] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _23340_ (.RESET_B(net689),
    .D(_00157_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][1] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _23341_ (.RESET_B(net688),
    .D(_00158_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][2] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _23342_ (.RESET_B(net687),
    .D(_00159_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][3] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _23343_ (.RESET_B(net686),
    .D(_00160_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][4] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _23344_ (.RESET_B(net685),
    .D(_00161_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][5] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _23345_ (.RESET_B(net684),
    .D(_00162_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][6] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _23346_ (.RESET_B(net683),
    .D(_00163_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][7] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _23347_ (.RESET_B(net682),
    .D(_00164_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][8] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _23348_ (.RESET_B(net681),
    .D(_00165_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][9] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _23349_ (.RESET_B(net680),
    .D(_00166_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _23350_ (.RESET_B(net679),
    .D(_00167_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][11] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _23351_ (.RESET_B(net678),
    .D(_00168_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][12] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _23352_ (.RESET_B(net677),
    .D(_00169_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][13] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _23353_ (.RESET_B(net676),
    .D(_00170_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][14] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _23354_ (.RESET_B(net675),
    .D(_00171_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][15] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _23355_ (.RESET_B(net674),
    .D(_00172_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][16] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _23356_ (.RESET_B(net673),
    .D(_00173_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][17] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _23357_ (.RESET_B(net672),
    .D(_00174_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][18] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _23358_ (.RESET_B(net671),
    .D(_00175_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _23359_ (.RESET_B(net670),
    .D(_00176_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _23360_ (.RESET_B(net669),
    .D(_00177_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][21] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _23361_ (.RESET_B(net668),
    .D(_00178_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][22] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _23362_ (.RESET_B(net667),
    .D(_00179_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][23] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _23363_ (.RESET_B(net666),
    .D(_00180_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][24] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _23364_ (.RESET_B(net665),
    .D(_00181_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][25] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _23365_ (.RESET_B(net664),
    .D(_00182_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][26] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _23366_ (.RESET_B(net663),
    .D(_00183_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][27] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _23367_ (.RESET_B(net662),
    .D(_00184_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][28] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _23368_ (.RESET_B(net661),
    .D(_00185_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][29] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _23369_ (.RESET_B(net660),
    .D(_00186_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][30] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _23370_ (.RESET_B(net659),
    .D(_00187_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][31] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _23371_ (.RESET_B(net5930),
    .D(_00188_),
    .Q(\fpga_top.io_led.led_value[0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _23372_ (.RESET_B(net5930),
    .D(_00189_),
    .Q(\fpga_top.io_led.led_value[1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _23373_ (.RESET_B(net5929),
    .D(_00190_),
    .Q(\fpga_top.io_led.led_value[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _23374_ (.RESET_B(net5844),
    .D(net6193),
    .Q(\fpga_top.io_spi_lite.spi_state[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _23375_ (.RESET_B(net5844),
    .D(net3828),
    .Q(\fpga_top.io_spi_lite.spi_state[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _23376_ (.RESET_B(net5924),
    .D(\fpga_top.io_spi_lite.re_spi_mode ),
    .Q(\fpga_top.io_spi_lite.re_spi_value_dly[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _23377_ (.RESET_B(net5888),
    .D(\fpga_top.io_spi_lite.re_spi_sdiv ),
    .Q(\fpga_top.io_spi_lite.re_spi_value_dly[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _23378_ (.RESET_B(net5889),
    .D(\fpga_top.io_spi_lite.re_spi_mosi ),
    .Q(\fpga_top.io_spi_lite.re_spi_value_dly[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _23379_ (.RESET_B(net5898),
    .D(\fpga_top.io_spi_lite.re_spi_miso ),
    .Q(\fpga_top.io_spi_lite.miso_fifo.rnext ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _23380_ (.RESET_B(net5846),
    .D(\fpga_top.io_spi_lite.miso_read_next_byte ),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wen ),
    .CLK(clknet_leaf_321_clk));
 sg13g2_dfrbpq_1 _23381_ (.RESET_B(net5889),
    .D(\fpga_top.io_spi_lite.org_spi_sck ),
    .Q(\fpga_top.io_spi_lite.sel_sck[1] ),
    .CLK(clknet_leaf_320_clk));
 sg13g2_dfrbpq_1 _23382_ (.RESET_B(net5896),
    .D(net1349),
    .Q(\fpga_top.io_spi_lite.sel_sck[2] ),
    .CLK(clknet_leaf_320_clk));
 sg13g2_dfrbpq_1 _23383_ (.RESET_B(net5896),
    .D(net1354),
    .Q(\fpga_top.io_spi_lite.sel_sck[3] ),
    .CLK(clknet_leaf_320_clk));
 sg13g2_dfrbpq_1 _23384_ (.RESET_B(net5900),
    .D(net1351),
    .Q(\fpga_top.io_spi_lite.sel_sck[4] ),
    .CLK(clknet_leaf_322_clk));
 sg13g2_dfrbpq_1 _23385_ (.RESET_B(net5900),
    .D(net1352),
    .Q(\fpga_top.io_spi_lite.sel_sck[5] ),
    .CLK(clknet_leaf_322_clk));
 sg13g2_dfrbpq_1 _23386_ (.RESET_B(net5900),
    .D(net1355),
    .Q(\fpga_top.io_spi_lite.sel_sck[6] ),
    .CLK(clknet_leaf_322_clk));
 sg13g2_dfrbpq_1 _23387_ (.RESET_B(net5900),
    .D(net1336),
    .Q(\fpga_top.io_spi_lite.sel_sck[7] ),
    .CLK(clknet_leaf_319_clk));
 sg13g2_dfrbpq_2 _23388_ (.RESET_B(net5840),
    .D(_00193_),
    .Q(\fpga_top.io_spi_lite.miso_byte_org[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _23389_ (.RESET_B(net5843),
    .D(_00194_),
    .Q(\fpga_top.io_spi_lite.miso_byte_org[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _23390_ (.RESET_B(net5843),
    .D(_00195_),
    .Q(\fpga_top.io_spi_lite.miso_byte_org[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _23391_ (.RESET_B(net5843),
    .D(_00196_),
    .Q(\fpga_top.io_spi_lite.miso_byte_org[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _23392_ (.RESET_B(net5843),
    .D(_00197_),
    .Q(\fpga_top.io_spi_lite.miso_byte_org[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _23393_ (.RESET_B(net5843),
    .D(_00198_),
    .Q(\fpga_top.io_spi_lite.miso_byte_org[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _23394_ (.RESET_B(net5843),
    .D(_00199_),
    .Q(\fpga_top.io_spi_lite.miso_byte_org[6] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _23395_ (.RESET_B(net5843),
    .D(_00200_),
    .Q(\fpga_top.io_spi_lite.miso_byte_org[7] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _23396_ (.RESET_B(net5860),
    .D(net1371),
    .Q(\fpga_top.io_spi_lite.miso_lat[2] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _23397_ (.RESET_B(net5861),
    .D(net1357),
    .Q(\fpga_top.io_spi_lite.miso_lat[3] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _23398_ (.RESET_B(net5860),
    .D(net1360),
    .Q(\fpga_top.io_spi_lite.miso_lat[4] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _23399_ (.RESET_B(net5861),
    .D(net1358),
    .Q(\fpga_top.io_spi_lite.miso_lat[5] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _23400_ (.RESET_B(net5861),
    .D(net1345),
    .Q(\fpga_top.io_spi_lite.miso_lat[6] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _23401_ (.RESET_B(net5861),
    .D(net1356),
    .Q(\fpga_top.io_spi_lite.miso_lat[7] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _23402_ (.RESET_B(net5892),
    .D(_00028_),
    .Q(\fpga_top.io_spi_lite.sck_div[0] ),
    .CLK(clknet_leaf_324_clk));
 sg13g2_dfrbpq_2 _23403_ (.RESET_B(net5892),
    .D(_00029_),
    .Q(\fpga_top.io_spi_lite.sck_div[1] ),
    .CLK(clknet_leaf_324_clk));
 sg13g2_dfrbpq_1 _23404_ (.RESET_B(net5892),
    .D(net1901),
    .Q(\fpga_top.io_spi_lite.sck_div[2] ),
    .CLK(clknet_leaf_325_clk));
 sg13g2_dfrbpq_1 _23405_ (.RESET_B(net5893),
    .D(_00031_),
    .Q(\fpga_top.io_spi_lite.sck_div[3] ),
    .CLK(clknet_leaf_325_clk));
 sg13g2_dfrbpq_2 _23406_ (.RESET_B(net5892),
    .D(net3873),
    .Q(\fpga_top.io_spi_lite.sck_div[4] ),
    .CLK(clknet_leaf_324_clk));
 sg13g2_dfrbpq_2 _23407_ (.RESET_B(net5892),
    .D(_00033_),
    .Q(\fpga_top.io_spi_lite.sck_div[5] ),
    .CLK(clknet_leaf_324_clk));
 sg13g2_dfrbpq_2 _23408_ (.RESET_B(net5892),
    .D(_00034_),
    .Q(\fpga_top.io_spi_lite.sck_div[6] ),
    .CLK(clknet_leaf_324_clk));
 sg13g2_dfrbpq_1 _23409_ (.RESET_B(net5892),
    .D(net3727),
    .Q(\fpga_top.io_spi_lite.sck_div[7] ),
    .CLK(clknet_leaf_324_clk));
 sg13g2_dfrbpq_2 _23410_ (.RESET_B(net5892),
    .D(_00036_),
    .Q(\fpga_top.io_spi_lite.sck_div[8] ),
    .CLK(clknet_leaf_323_clk));
 sg13g2_dfrbpq_2 _23411_ (.RESET_B(net5891),
    .D(_00037_),
    .Q(\fpga_top.io_spi_lite.sck_div[9] ),
    .CLK(clknet_leaf_323_clk));
 sg13g2_dfrbpq_1 _23412_ (.RESET_B(net5926),
    .D(\fpga_top.io_spi_lite.cs_all_status ),
    .Q(\fpga_top.io_spi_lite.sel_cs[1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23413_ (.RESET_B(net5927),
    .D(net1353),
    .Q(\fpga_top.io_spi_lite.sel_cs[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23414_ (.RESET_B(net5933),
    .D(net1347),
    .Q(\fpga_top.io_spi_lite.sel_cs[3] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23415_ (.RESET_B(net5933),
    .D(net1344),
    .Q(\fpga_top.io_spi_lite.sel_cs[4] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23416_ (.RESET_B(net5933),
    .D(net1340),
    .Q(\fpga_top.io_spi_lite.sel_cs[5] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23417_ (.RESET_B(net5933),
    .D(net1359),
    .Q(\fpga_top.io_spi_lite.sel_cs[6] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23418_ (.RESET_B(net5934),
    .D(net1341),
    .Q(\fpga_top.io_spi_lite.sel_cs[7] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23419_ (.RESET_B(net5930),
    .D(\fpga_top.io_spi_lite.spi_mosi_pre ),
    .Q(\fpga_top.io_spi_lite.spi_mosi ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _23420_ (.RESET_B(net5927),
    .D(\fpga_top.io_spi_lite.org_mosi ),
    .Q(\fpga_top.io_spi_lite.sel_mosi[1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23421_ (.RESET_B(net5933),
    .D(net1348),
    .Q(\fpga_top.io_spi_lite.sel_mosi[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23422_ (.RESET_B(net5934),
    .D(net1324),
    .Q(\fpga_top.io_spi_lite.sel_mosi[3] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _23423_ (.RESET_B(net5938),
    .D(net1363),
    .Q(\fpga_top.io_spi_lite.sel_mosi[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23424_ (.RESET_B(net5938),
    .D(net1342),
    .Q(\fpga_top.io_spi_lite.sel_mosi[5] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23425_ (.RESET_B(net5938),
    .D(net1350),
    .Q(\fpga_top.io_spi_lite.sel_mosi[6] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _23426_ (.RESET_B(net5937),
    .D(net1343),
    .Q(\fpga_top.io_spi_lite.sel_mosi[7] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _23427_ (.RESET_B(net5842),
    .D(_00201_),
    .Q(\fpga_top.io_spi_lite.mosi_pp_cntr[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _23428_ (.RESET_B(net5842),
    .D(net1757),
    .Q(\fpga_top.io_spi_lite.mosi_pp_cntr[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _23429_ (.RESET_B(net5842),
    .D(net1581),
    .Q(\fpga_top.io_spi_lite.mosi_pp_cntr[2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _23430_ (.RESET_B(net5842),
    .D(net1682),
    .Q(\fpga_top.io_spi_lite.mosi_pp_cntr[3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _23431_ (.RESET_B(net5846),
    .D(net1656),
    .Q(\fpga_top.io_spi_lite.miso_bit_cntr[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23432_ (.RESET_B(net5846),
    .D(net1429),
    .Q(\fpga_top.io_spi_lite.miso_bit_cntr[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23433_ (.RESET_B(net5846),
    .D(net1409),
    .Q(\fpga_top.io_spi_lite.miso_bit_cntr[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23434_ (.RESET_B(net5887),
    .D(net1369),
    .Q(\fpga_top.io_spi_lite.org_sck_dly ),
    .CLK(clknet_leaf_320_clk));
 sg13g2_dfrbpq_2 _23435_ (.RESET_B(net5842),
    .D(net1704),
    .Q(\fpga_top.io_spi_lite.bit_sel_org[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _23436_ (.RESET_B(net5857),
    .D(net1977),
    .Q(\fpga_top.io_spi_lite.bit_sel_org[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _23437_ (.RESET_B(net5841),
    .D(_00210_),
    .Q(\fpga_top.io_spi_lite.bit_sel_org[2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _23438_ (.RESET_B(net5839),
    .D(net1893),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.radr[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _23439_ (.RESET_B(net5839),
    .D(\fpga_top.io_spi_lite.mosi_fifo.radr_early[1] ),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.radr[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _23440_ (.RESET_B(net5839),
    .D(net1573),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.radr[2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _23441_ (.RESET_B(net5887),
    .D(net6416),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[0] ),
    .CLK(clknet_leaf_325_clk));
 sg13g2_dfrbpq_2 _23442_ (.RESET_B(net5846),
    .D(net6492),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ),
    .CLK(clknet_leaf_325_clk));
 sg13g2_dfrbpq_2 _23443_ (.RESET_B(net5846),
    .D(_00213_),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[2] ),
    .CLK(clknet_leaf_326_clk));
 sg13g2_dfrbpq_1 _23444_ (.RESET_B(net658),
    .D(_00214_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][0] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _23445_ (.RESET_B(net657),
    .D(_00215_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][1] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _23446_ (.RESET_B(net656),
    .D(_00216_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][2] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _23447_ (.RESET_B(net655),
    .D(_00217_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][3] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _23448_ (.RESET_B(net654),
    .D(_00218_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][4] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _23449_ (.RESET_B(net653),
    .D(_00219_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][5] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _23450_ (.RESET_B(net652),
    .D(_00220_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][6] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _23451_ (.RESET_B(net651),
    .D(_00221_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][7] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _23452_ (.RESET_B(net650),
    .D(_00222_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][8] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _23453_ (.RESET_B(net649),
    .D(_00223_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][9] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _23454_ (.RESET_B(net648),
    .D(_00224_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _23455_ (.RESET_B(net647),
    .D(_00225_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][11] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _23456_ (.RESET_B(net646),
    .D(_00226_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][12] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _23457_ (.RESET_B(net645),
    .D(_00227_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][13] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _23458_ (.RESET_B(net644),
    .D(_00228_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][14] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _23459_ (.RESET_B(net643),
    .D(_00229_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][15] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _23460_ (.RESET_B(net642),
    .D(_00230_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][16] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _23461_ (.RESET_B(net641),
    .D(_00231_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][17] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _23462_ (.RESET_B(net640),
    .D(_00232_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][18] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _23463_ (.RESET_B(net639),
    .D(_00233_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][19] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _23464_ (.RESET_B(net638),
    .D(_00234_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][20] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _23465_ (.RESET_B(net637),
    .D(_00235_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][21] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _23466_ (.RESET_B(net636),
    .D(_00236_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][22] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _23467_ (.RESET_B(net635),
    .D(_00237_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][23] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _23468_ (.RESET_B(net634),
    .D(_00238_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][24] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _23469_ (.RESET_B(net633),
    .D(_00239_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _23470_ (.RESET_B(net632),
    .D(_00240_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][26] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _23471_ (.RESET_B(net631),
    .D(_00241_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][27] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _23472_ (.RESET_B(net630),
    .D(_00242_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][28] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _23473_ (.RESET_B(net629),
    .D(_00243_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][29] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _23474_ (.RESET_B(net628),
    .D(_00244_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][30] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _23475_ (.RESET_B(net57),
    .D(_00245_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][31] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _23476_ (.RESET_B(net5887),
    .D(_00038_),
    .Q(\fpga_top.io_spi_lite.miso_fifo.radr[0] ),
    .CLK(clknet_leaf_321_clk));
 sg13g2_dfrbpq_2 _23477_ (.RESET_B(net5887),
    .D(_00039_),
    .Q(\fpga_top.io_spi_lite.miso_fifo.radr[1] ),
    .CLK(clknet_leaf_325_clk));
 sg13g2_dfrbpq_1 _23478_ (.RESET_B(net5887),
    .D(_00040_),
    .Q(\fpga_top.io_spi_lite.miso_fifo.radr[2] ),
    .CLK(clknet_leaf_325_clk));
 sg13g2_dfrbpq_2 _23479_ (.RESET_B(net5930),
    .D(_00246_),
    .Q(\fpga_top.io_spi_lite.spi_mode[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23480_ (.RESET_B(net5890),
    .D(_00247_),
    .Q(\fpga_top.io_spi_lite.spi_mode[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _23481_ (.RESET_B(net5890),
    .D(_00248_),
    .Q(\fpga_top.io_spi_lite.spi_mode[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _23482_ (.RESET_B(net5890),
    .D(_00249_),
    .Q(_00085_),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _23483_ (.RESET_B(net5943),
    .D(_00250_),
    .Q(\fpga_top.io_spi_lite.spi_mode[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _23484_ (.RESET_B(net5931),
    .D(_00251_),
    .Q(\fpga_top.io_spi_lite.spi_mode[5] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23485_ (.RESET_B(net5931),
    .D(_00252_),
    .Q(\fpga_top.io_spi_lite.spi_mode[6] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23486_ (.RESET_B(net5897),
    .D(_00253_),
    .Q(\fpga_top.io_spi_lite.spi_mode[7] ),
    .CLK(clknet_leaf_319_clk));
 sg13g2_dfrbpq_2 _23487_ (.RESET_B(net5900),
    .D(_00254_),
    .Q(\fpga_top.io_spi_lite.spi_mode[8] ),
    .CLK(clknet_leaf_320_clk));
 sg13g2_dfrbpq_2 _23488_ (.RESET_B(net5900),
    .D(_00255_),
    .Q(\fpga_top.io_spi_lite.spi_mode[9] ),
    .CLK(clknet_leaf_319_clk));
 sg13g2_dfrbpq_2 _23489_ (.RESET_B(net5931),
    .D(_00256_),
    .Q(\fpga_top.io_spi_lite.spi_mode[10] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23490_ (.RESET_B(net5943),
    .D(_00257_),
    .Q(\fpga_top.io_spi_lite.spi_mode[11] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _23491_ (.RESET_B(net5930),
    .D(_00258_),
    .Q(\fpga_top.io_spi_lite.spi_mode[12] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _23492_ (.RESET_B(net5898),
    .D(net1373),
    .Q(\fpga_top.interrupter.int0_3lat ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _23493_ (.RESET_B(net5904),
    .D(\fpga_top.interrupter.re_int_enable ),
    .Q(\fpga_top.interrupter.re_int_dly[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _23494_ (.RESET_B(net5898),
    .D(\fpga_top.interrupter.re_int_status ),
    .Q(\fpga_top.interrupter.re_int_dly[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _23495_ (.RESET_B(net5989),
    .D(\fpga_top.cpu_top.execution.csr_array.g_interrupt ),
    .Q(\fpga_top.interrupter.g_interrupt_dly ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _23496_ (.RESET_B(net6065),
    .D(_00259_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[0] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _23497_ (.RESET_B(net6067),
    .D(_00260_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[1] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _23498_ (.RESET_B(net6077),
    .D(_00261_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[2] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _23499_ (.RESET_B(net6066),
    .D(_00262_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[3] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _23500_ (.RESET_B(net6066),
    .D(_00263_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[4] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _23501_ (.RESET_B(net6066),
    .D(_00264_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[5] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _23502_ (.RESET_B(net6067),
    .D(_00265_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[6] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _23503_ (.RESET_B(net6076),
    .D(_00266_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[7] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _23504_ (.RESET_B(net6077),
    .D(_00267_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[8] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _23505_ (.RESET_B(net6076),
    .D(_00268_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[9] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _23506_ (.RESET_B(net6075),
    .D(_00269_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[10] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _23507_ (.RESET_B(net6077),
    .D(_00270_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[11] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _23508_ (.RESET_B(net6075),
    .D(_00271_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[12] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _23509_ (.RESET_B(net6075),
    .D(_00272_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[13] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _23510_ (.RESET_B(net6062),
    .D(_00273_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[14] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _23511_ (.RESET_B(net6073),
    .D(_00274_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[15] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _23512_ (.RESET_B(net6074),
    .D(_00275_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[16] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _23513_ (.RESET_B(net6062),
    .D(_00276_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[17] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _23514_ (.RESET_B(net6076),
    .D(_00277_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[18] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _23515_ (.RESET_B(net6073),
    .D(_00278_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[19] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _23516_ (.RESET_B(net6073),
    .D(_00279_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[20] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _23517_ (.RESET_B(net6070),
    .D(_00280_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[21] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _23518_ (.RESET_B(net6074),
    .D(_00281_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[22] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _23519_ (.RESET_B(net6076),
    .D(_00282_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[23] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _23520_ (.RESET_B(net6076),
    .D(_00283_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[24] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _23521_ (.RESET_B(net6070),
    .D(_00284_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[25] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _23522_ (.RESET_B(net6076),
    .D(_00285_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[26] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _23523_ (.RESET_B(net6070),
    .D(_00286_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[27] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _23524_ (.RESET_B(net6074),
    .D(_00287_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[28] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _23525_ (.RESET_B(net6074),
    .D(_00288_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[29] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _23526_ (.RESET_B(net6073),
    .D(_00289_),
    .Q(\fpga_top.cpu_top.execution.csr_array.rs1_sel[30] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _23527_ (.RESET_B(net6075),
    .D(_00290_),
    .Q(\fpga_top.cpu_top.execution.alu_sra[31] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _23528_ (.RESET_B(net5936),
    .D(net1320),
    .Q(\fpga_top.interrupter.int0_2lat ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _23529_ (.RESET_B(net5899),
    .D(net3970),
    .Q(\fpga_top.interrupter.int_status_int0 ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _23530_ (.RESET_B(net5935),
    .D(net2),
    .Q(\fpga_top.interrupter.int0_1lat ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _23531_ (.RESET_B(net5899),
    .D(net2836),
    .Q(\fpga_top.interrupter.int_status_rx ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _23532_ (.RESET_B(net5898),
    .D(_00293_),
    .Q(\fpga_top.io_frc.frc_cmp_val[32] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _23533_ (.RESET_B(net5898),
    .D(_00294_),
    .Q(\fpga_top.io_frc.frc_cmp_val[33] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _23534_ (.RESET_B(net5922),
    .D(_00295_),
    .Q(\fpga_top.io_frc.frc_cmp_val[34] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _23535_ (.RESET_B(net5924),
    .D(_00296_),
    .Q(\fpga_top.io_frc.frc_cmp_val[35] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _23536_ (.RESET_B(net5924),
    .D(_00297_),
    .Q(\fpga_top.io_frc.frc_cmp_val[36] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _23537_ (.RESET_B(net5922),
    .D(_00298_),
    .Q(\fpga_top.io_frc.frc_cmp_val[37] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _23538_ (.RESET_B(net5898),
    .D(_00299_),
    .Q(\fpga_top.io_frc.frc_cmp_val[38] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _23539_ (.RESET_B(net5898),
    .D(_00300_),
    .Q(\fpga_top.io_frc.frc_cmp_val[39] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _23540_ (.RESET_B(net5895),
    .D(_00301_),
    .Q(\fpga_top.io_frc.frc_cmp_val[40] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23541_ (.RESET_B(net5894),
    .D(_00302_),
    .Q(\fpga_top.io_frc.frc_cmp_val[41] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _23542_ (.RESET_B(net5895),
    .D(_00303_),
    .Q(\fpga_top.io_frc.frc_cmp_val[42] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _23543_ (.RESET_B(net5901),
    .D(_00304_),
    .Q(\fpga_top.io_frc.frc_cmp_val[43] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23544_ (.RESET_B(net5917),
    .D(_00305_),
    .Q(\fpga_top.io_frc.frc_cmp_val[44] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _23545_ (.RESET_B(net5917),
    .D(_00306_),
    .Q(\fpga_top.io_frc.frc_cmp_val[45] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _23546_ (.RESET_B(net5917),
    .D(_00307_),
    .Q(\fpga_top.io_frc.frc_cmp_val[46] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23547_ (.RESET_B(net5942),
    .D(_00308_),
    .Q(\fpga_top.io_frc.frc_cmp_val[47] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _23548_ (.RESET_B(net5905),
    .D(_00309_),
    .Q(\fpga_top.io_frc.frc_cmp_val[48] ),
    .CLK(clknet_leaf_324_clk));
 sg13g2_dfrbpq_1 _23549_ (.RESET_B(net5905),
    .D(_00310_),
    .Q(\fpga_top.io_frc.frc_cmp_val[49] ),
    .CLK(clknet_leaf_323_clk));
 sg13g2_dfrbpq_2 _23550_ (.RESET_B(net5906),
    .D(_00311_),
    .Q(\fpga_top.io_frc.frc_cmp_val[50] ),
    .CLK(clknet_leaf_323_clk));
 sg13g2_dfrbpq_2 _23551_ (.RESET_B(net5906),
    .D(_00312_),
    .Q(\fpga_top.io_frc.frc_cmp_val[51] ),
    .CLK(clknet_leaf_323_clk));
 sg13g2_dfrbpq_1 _23552_ (.RESET_B(net5907),
    .D(_00313_),
    .Q(\fpga_top.io_frc.frc_cmp_val[52] ),
    .CLK(clknet_leaf_323_clk));
 sg13g2_dfrbpq_2 _23553_ (.RESET_B(net5907),
    .D(_00314_),
    .Q(\fpga_top.io_frc.frc_cmp_val[53] ),
    .CLK(clknet_leaf_323_clk));
 sg13g2_dfrbpq_2 _23554_ (.RESET_B(net5918),
    .D(_00315_),
    .Q(\fpga_top.io_frc.frc_cmp_val[54] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _23555_ (.RESET_B(net5915),
    .D(_00316_),
    .Q(\fpga_top.io_frc.frc_cmp_val[55] ),
    .CLK(clknet_leaf_318_clk));
 sg13g2_dfrbpq_2 _23556_ (.RESET_B(net5943),
    .D(_00317_),
    .Q(\fpga_top.io_frc.frc_cmp_val[56] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23557_ (.RESET_B(net5944),
    .D(_00318_),
    .Q(\fpga_top.io_frc.frc_cmp_val[57] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23558_ (.RESET_B(net5944),
    .D(_00319_),
    .Q(\fpga_top.io_frc.frc_cmp_val[58] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _23559_ (.RESET_B(net5944),
    .D(_00320_),
    .Q(\fpga_top.io_frc.frc_cmp_val[59] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23560_ (.RESET_B(net5944),
    .D(_00321_),
    .Q(\fpga_top.io_frc.frc_cmp_val[60] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _23561_ (.RESET_B(net5943),
    .D(_00322_),
    .Q(\fpga_top.io_frc.frc_cmp_val[61] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _23562_ (.RESET_B(net5942),
    .D(_00323_),
    .Q(\fpga_top.io_frc.frc_cmp_val[62] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _23563_ (.RESET_B(net5942),
    .D(_00324_),
    .Q(\fpga_top.io_frc.frc_cmp_val[63] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _23564_ (.RESET_B(net5922),
    .D(\fpga_top.io_frc.re_frc_vallo ),
    .Q(\fpga_top.io_frc.re_frc_dly[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _23565_ (.RESET_B(net5922),
    .D(\fpga_top.io_frc.re_frc_valhi ),
    .Q(\fpga_top.io_frc.re_frc_dly[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _23566_ (.RESET_B(net5922),
    .D(\fpga_top.io_frc.re_frc_cmplo ),
    .Q(\fpga_top.io_frc.re_frc_dly[2] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _23567_ (.RESET_B(net5922),
    .D(\fpga_top.io_frc.re_frc_cmphi ),
    .Q(\fpga_top.io_frc.re_frc_dly[3] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _23568_ (.RESET_B(net5925),
    .D(\fpga_top.io_frc.re_frc_cntrl ),
    .Q(\fpga_top.io_frc.re_frc_dly[4] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _23569_ (.RESET_B(net5904),
    .D(_00325_),
    .Q(\fpga_top.interrupter.int_enable_rx ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _23570_ (.RESET_B(net5899),
    .D(_00326_),
    .Q(\fpga_top.interrupter.int_enable_int0 ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _23571_ (.RESET_B(net5903),
    .D(\fpga_top.io_frc.frc_cntr_val_rst_pre ),
    .Q(\fpga_top.io_frc.frc_cntr_val_rst_lat ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23572_ (.RESET_B(net5903),
    .D(_00327_),
    .Q(\fpga_top.io_frc.frc_cntrl_val ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23573_ (.RESET_B(net5918),
    .D(net1382),
    .Q(\fpga_top.cpu_top.execution.csr_array.frc_cntr_val_leq ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _23574_ (.RESET_B(net622),
    .D(_00329_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][0] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _23575_ (.RESET_B(net621),
    .D(_00330_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][1] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _23576_ (.RESET_B(net620),
    .D(_00331_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][2] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _23577_ (.RESET_B(net619),
    .D(_00332_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][3] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _23578_ (.RESET_B(net618),
    .D(_00333_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][4] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _23579_ (.RESET_B(net617),
    .D(_00334_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _23580_ (.RESET_B(net616),
    .D(_00335_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][6] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _23581_ (.RESET_B(net615),
    .D(_00336_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][7] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _23582_ (.RESET_B(net614),
    .D(_00337_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][8] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _23583_ (.RESET_B(net613),
    .D(_00338_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][9] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _23584_ (.RESET_B(net612),
    .D(_00339_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _23585_ (.RESET_B(net611),
    .D(_00340_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][11] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _23586_ (.RESET_B(net610),
    .D(_00341_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][12] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _23587_ (.RESET_B(net609),
    .D(_00342_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][13] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _23588_ (.RESET_B(net608),
    .D(_00343_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][14] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _23589_ (.RESET_B(net607),
    .D(_00344_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][15] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _23590_ (.RESET_B(net606),
    .D(_00345_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][16] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _23591_ (.RESET_B(net605),
    .D(_00346_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][17] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _23592_ (.RESET_B(net604),
    .D(_00347_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][18] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _23593_ (.RESET_B(net603),
    .D(_00348_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _23594_ (.RESET_B(net602),
    .D(_00349_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _23595_ (.RESET_B(net601),
    .D(_00350_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][21] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _23596_ (.RESET_B(net600),
    .D(_00351_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][22] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _23597_ (.RESET_B(net599),
    .D(_00352_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][23] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _23598_ (.RESET_B(net598),
    .D(_00353_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][24] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _23599_ (.RESET_B(net597),
    .D(_00354_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _23600_ (.RESET_B(net596),
    .D(_00355_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][26] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _23601_ (.RESET_B(net595),
    .D(_00356_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][27] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _23602_ (.RESET_B(net594),
    .D(_00357_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][28] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _23603_ (.RESET_B(net593),
    .D(_00358_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][29] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _23604_ (.RESET_B(net592),
    .D(_00359_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][30] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _23605_ (.RESET_B(net591),
    .D(_00360_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][31] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _23606_ (.RESET_B(net5877),
    .D(_00361_),
    .Q(\fpga_top.io_uart_out.uart_term[0] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _23607_ (.RESET_B(net5877),
    .D(_00362_),
    .Q(\fpga_top.io_uart_out.uart_term[1] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _23608_ (.RESET_B(net5877),
    .D(_00363_),
    .Q(\fpga_top.io_uart_out.uart_term[2] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _23609_ (.RESET_B(net5877),
    .D(_00364_),
    .Q(\fpga_top.io_uart_out.uart_term[3] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _23610_ (.RESET_B(net5878),
    .D(_00365_),
    .Q(\fpga_top.io_uart_out.uart_term[4] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _23611_ (.RESET_B(net5877),
    .D(_00366_),
    .Q(\fpga_top.io_uart_out.uart_term[5] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _23612_ (.RESET_B(net5877),
    .D(_00367_),
    .Q(\fpga_top.io_uart_out.uart_term[6] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _23613_ (.RESET_B(net5877),
    .D(_00368_),
    .Q(\fpga_top.io_uart_out.uart_term[7] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _23614_ (.RESET_B(net5881),
    .D(_00369_),
    .Q(\fpga_top.io_uart_out.uart_term[8] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _23615_ (.RESET_B(net5923),
    .D(_00370_),
    .Q(\fpga_top.io_uart_out.uart_term[9] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _23616_ (.RESET_B(net5881),
    .D(_00371_),
    .Q(\fpga_top.io_uart_out.uart_term[10] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23617_ (.RESET_B(net5924),
    .D(_00372_),
    .Q(\fpga_top.io_uart_out.uart_term[11] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _23618_ (.RESET_B(net5930),
    .D(_00373_),
    .Q(\fpga_top.io_uart_out.uart_term[12] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23619_ (.RESET_B(net5931),
    .D(_00374_),
    .Q(\fpga_top.io_uart_out.uart_term[13] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23620_ (.RESET_B(net5929),
    .D(_00375_),
    .Q(\fpga_top.io_uart_out.uart_term[14] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _23621_ (.RESET_B(net5930),
    .D(_00376_),
    .Q(\fpga_top.io_uart_out.uart_term[15] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23622_ (.RESET_B(net5923),
    .D(\fpga_top.io_uart_out.re_uart_char ),
    .Q(\fpga_top.io_uart_out.re_uart_rdflg_dly[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _23623_ (.RESET_B(net5924),
    .D(\fpga_top.io_uart_out.re_uart_full ),
    .Q(\fpga_top.io_uart_out.re_uart_rdflg_dly[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _23624_ (.RESET_B(net5922),
    .D(\fpga_top.io_uart_out.re_uart_term ),
    .Q(\fpga_top.io_uart_out.re_uart_rdflg_dly[2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _23625_ (.RESET_B(net5924),
    .D(\fpga_top.io_uart_out.re_uart_rxch ),
    .Q(\fpga_top.io_uart_out.re_uart_rdflg_dly[3] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _23626_ (.RESET_B(net5924),
    .D(\fpga_top.io_uart_out.re_uart_rxec ),
    .Q(\fpga_top.io_uart_out.re_uart_rdflg_dly[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _23627_ (.RESET_B(net5839),
    .D(_00377_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _23628_ (.RESET_B(net5858),
    .D(net2063),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _23629_ (.RESET_B(net5858),
    .D(_00379_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _23630_ (.RESET_B(net5933),
    .D(_00380_),
    .Q(\fpga_top.io_uart_out.rx_disable_echoback_value ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _23631_ (.RESET_B(net5881),
    .D(_00041_),
    .Q(\fpga_top.io_uart_out.uart_io_we ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _23632_ (.RESET_B(net5927),
    .D(_00381_),
    .Q(\fpga_top.io_uart_out.rx_write_error ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _23633_ (.RESET_B(net5930),
    .D(net1388),
    .Q(\fpga_top.io_uart_out.rx_first_read ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _23634_ (.RESET_B(net5933),
    .D(net1687),
    .Q(\fpga_top.io_uart_out.rx_data_latch[0] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _23635_ (.RESET_B(net5884),
    .D(net3884),
    .Q(\fpga_top.io_uart_out.rx_data_latch[1] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _23636_ (.RESET_B(net5884),
    .D(_00385_),
    .Q(\fpga_top.io_uart_out.rx_data_latch[2] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _23637_ (.RESET_B(net5934),
    .D(net3816),
    .Q(\fpga_top.io_uart_out.rx_data_latch[3] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23638_ (.RESET_B(net5933),
    .D(_00387_),
    .Q(\fpga_top.io_uart_out.rx_data_latch[4] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23639_ (.RESET_B(net5934),
    .D(net3736),
    .Q(\fpga_top.io_uart_out.rx_data_latch[5] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _23640_ (.RESET_B(net5934),
    .D(net3596),
    .Q(\fpga_top.io_uart_out.rx_data_latch[6] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _23641_ (.RESET_B(net5926),
    .D(net1712),
    .Q(\fpga_top.io_uart_out.rx_data_latch[7] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _23642_ (.RESET_B(net5902),
    .D(net4013),
    .Q(\fpga_top.io_led.dbg_smpl_trgsig ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _23643_ (.RESET_B(net5924),
    .D(\fpga_top.io_led.re_led_value ),
    .Q(\fpga_top.io_led.re_led_value_dly ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _23644_ (.RESET_B(net5875),
    .D(net1346),
    .Q(\fpga_top.io_led.gpi_init_lat2[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23645_ (.RESET_B(net5875),
    .D(net1332),
    .Q(\fpga_top.io_led.gpi_init_lat2[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _23646_ (.RESET_B(net5862),
    .D(net1318),
    .Q(\fpga_top.io_led.gpi_init_lat2[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _23647_ (.RESET_B(net5935),
    .D(net1337),
    .Q(\fpga_top.io_led.gpi_init_lat2[3] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _23648_ (.RESET_B(net5881),
    .D(net1327),
    .Q(\fpga_top.io_led.gpi_init_lat2[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _23649_ (.RESET_B(net5872),
    .D(net1322),
    .Q(\fpga_top.io_led.gpi_init_lat2[5] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _23650_ (.RESET_B(net5869),
    .D(_00392_),
    .Q(uio_out[4]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _23651_ (.RESET_B(net5868),
    .D(_00393_),
    .Q(uio_out[5]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _23652_ (.RESET_B(net5869),
    .D(_00394_),
    .Q(uio_out[6]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _23653_ (.RESET_B(net5869),
    .D(_00395_),
    .Q(uio_out[7]),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _23654_ (.RESET_B(net5865),
    .D(net1334),
    .Q(\fpga_top.io_led.gpio_in_lat2[0] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _23655_ (.RESET_B(net5868),
    .D(net1330),
    .Q(\fpga_top.io_led.gpio_in_lat2[1] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _23656_ (.RESET_B(net5864),
    .D(net1338),
    .Q(\fpga_top.io_led.gpio_in_lat2[2] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _23657_ (.RESET_B(net5864),
    .D(net1333),
    .Q(\fpga_top.io_led.gpio_in_lat2[3] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _23658_ (.RESET_B(net5899),
    .D(_00396_),
    .Q(\fpga_top.io_frc.frc_cntr_val[0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _23659_ (.RESET_B(net5899),
    .D(_00397_),
    .Q(\fpga_top.io_frc.frc_cntr_val[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _23660_ (.RESET_B(net5899),
    .D(_00398_),
    .Q(\fpga_top.io_frc.frc_cntr_val[2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _23661_ (.RESET_B(net5889),
    .D(net6180),
    .Q(\fpga_top.io_frc.frc_cntr_val[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _23662_ (.RESET_B(net5888),
    .D(net6322),
    .Q(\fpga_top.io_frc.frc_cntr_val[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _23663_ (.RESET_B(net5896),
    .D(_00401_),
    .Q(\fpga_top.io_frc.frc_cntr_val[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _23664_ (.RESET_B(net5896),
    .D(_00402_),
    .Q(\fpga_top.io_frc.frc_cntr_val[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _23665_ (.RESET_B(net5896),
    .D(net6198),
    .Q(\fpga_top.io_frc.frc_cntr_val[7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _23666_ (.RESET_B(net5895),
    .D(_00404_),
    .Q(\fpga_top.io_frc.frc_cntr_val[8] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _23667_ (.RESET_B(net5895),
    .D(net4029),
    .Q(\fpga_top.io_frc.frc_cntr_val[9] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _23668_ (.RESET_B(net5908),
    .D(net4017),
    .Q(\fpga_top.io_frc.frc_cntr_val[10] ),
    .CLK(clknet_leaf_319_clk));
 sg13g2_dfrbpq_2 _23669_ (.RESET_B(net5915),
    .D(_00407_),
    .Q(\fpga_top.io_frc.frc_cntr_val[11] ),
    .CLK(clknet_leaf_318_clk));
 sg13g2_dfrbpq_1 _23670_ (.RESET_B(net5916),
    .D(_00408_),
    .Q(\fpga_top.io_frc.frc_cntr_val[12] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _23671_ (.RESET_B(net5916),
    .D(net3746),
    .Q(\fpga_top.io_frc.frc_cntr_val[13] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _23672_ (.RESET_B(net5916),
    .D(_00410_),
    .Q(\fpga_top.io_frc.frc_cntr_val[14] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _23673_ (.RESET_B(net5917),
    .D(net3903),
    .Q(\fpga_top.io_frc.frc_cntr_val[15] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _23674_ (.RESET_B(net5908),
    .D(_00412_),
    .Q(\fpga_top.io_frc.frc_cntr_val[16] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_2 _23675_ (.RESET_B(net5908),
    .D(_00413_),
    .Q(\fpga_top.io_frc.frc_cntr_val[17] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_2 _23676_ (.RESET_B(net5907),
    .D(_00414_),
    .Q(\fpga_top.io_frc.frc_cntr_val[18] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _23677_ (.RESET_B(net5908),
    .D(net3804),
    .Q(\fpga_top.io_frc.frc_cntr_val[19] ),
    .CLK(clknet_leaf_318_clk));
 sg13g2_dfrbpq_2 _23678_ (.RESET_B(net5908),
    .D(net3757),
    .Q(\fpga_top.io_frc.frc_cntr_val[20] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_2 _23679_ (.RESET_B(net5908),
    .D(_00417_),
    .Q(\fpga_top.io_frc.frc_cntr_val[21] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_2 _23680_ (.RESET_B(net5915),
    .D(_00418_),
    .Q(\fpga_top.io_frc.frc_cntr_val[22] ),
    .CLK(clknet_leaf_318_clk));
 sg13g2_dfrbpq_1 _23681_ (.RESET_B(net5903),
    .D(_00419_),
    .Q(\fpga_top.io_frc.frc_cntr_val[23] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _23682_ (.RESET_B(net5928),
    .D(net4006),
    .Q(\fpga_top.io_frc.frc_cntr_val[24] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _23683_ (.RESET_B(net5929),
    .D(net6182),
    .Q(\fpga_top.io_frc.frc_cntr_val[25] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _23684_ (.RESET_B(net5928),
    .D(net4041),
    .Q(\fpga_top.io_frc.frc_cntr_val[26] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23685_ (.RESET_B(net5928),
    .D(net3863),
    .Q(\fpga_top.io_frc.frc_cntr_val[27] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _23686_ (.RESET_B(net5928),
    .D(_00424_),
    .Q(\fpga_top.io_frc.frc_cntr_val[28] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _23687_ (.RESET_B(net5928),
    .D(net6137),
    .Q(\fpga_top.io_frc.frc_cntr_val[29] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _23688_ (.RESET_B(net5928),
    .D(_00426_),
    .Q(\fpga_top.io_frc.frc_cntr_val[30] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _23689_ (.RESET_B(net5929),
    .D(net6087),
    .Q(\fpga_top.io_frc.frc_cntr_val[31] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _23690_ (.RESET_B(net5875),
    .D(net3),
    .Q(\fpga_top.io_led.gpi_init_lat1[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23691_ (.RESET_B(net5874),
    .D(net4),
    .Q(\fpga_top.io_led.gpi_init_lat1[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _23692_ (.RESET_B(net5862),
    .D(net5),
    .Q(\fpga_top.io_led.gpi_init_lat1[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23693_ (.RESET_B(net5935),
    .D(net6),
    .Q(\fpga_top.io_led.gpi_init_lat1[3] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _23694_ (.RESET_B(net5874),
    .D(net7),
    .Q(\fpga_top.io_led.gpi_init_lat1[4] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _23695_ (.RESET_B(net5872),
    .D(net8),
    .Q(\fpga_top.io_led.gpi_init_lat1[5] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _23696_ (.RESET_B(net5865),
    .D(net13),
    .Q(\fpga_top.io_led.gpio_in_lat1[0] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _23697_ (.RESET_B(net5864),
    .D(net14),
    .Q(\fpga_top.io_led.gpio_in_lat1[1] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _23698_ (.RESET_B(net5864),
    .D(net15),
    .Q(\fpga_top.io_led.gpio_in_lat1[2] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _23699_ (.RESET_B(net5864),
    .D(net16),
    .Q(\fpga_top.io_led.gpio_in_lat1[3] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _23700_ (.RESET_B(net5866),
    .D(_00428_),
    .Q(uio_oe[4]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _23701_ (.RESET_B(net5869),
    .D(_00429_),
    .Q(uio_oe[5]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _23702_ (.RESET_B(net5866),
    .D(_00430_),
    .Q(uio_oe[6]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _23703_ (.RESET_B(net5866),
    .D(_00431_),
    .Q(uio_oe[7]),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _23704_ (.RESET_B(net5922),
    .D(\fpga_top.io_led.re_gpi_value ),
    .Q(\fpga_top.io_led.re_gpio_value_dly[0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _23705_ (.RESET_B(net5877),
    .D(\fpga_top.io_led.re_gpio_out_value ),
    .Q(\fpga_top.io_led.re_gpio_value_dly[1] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _23706_ (.RESET_B(net5880),
    .D(\fpga_top.io_led.re_gpio_in_value ),
    .Q(\fpga_top.io_led.re_gpio_value_dly[2] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _23707_ (.RESET_B(net5880),
    .D(\fpga_top.io_led.re_gpio_en_value ),
    .Q(\fpga_top.io_led.re_gpio_value_dly[3] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _23708_ (.RESET_B(net5882),
    .D(net1328),
    .Q(\fpga_top.qspi_if.sio_in_mt1[0] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _23709_ (.RESET_B(net5868),
    .D(net1316),
    .Q(\fpga_top.qspi_if.sio_in_mt1[1] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _23710_ (.RESET_B(net5885),
    .D(net1319),
    .Q(\fpga_top.qspi_if.sio_in_mt1[2] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _23711_ (.RESET_B(net5868),
    .D(net1339),
    .Q(\fpga_top.qspi_if.sio_in_mt1[3] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _23712_ (.RESET_B(net590),
    .D(_00432_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][0] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _23713_ (.RESET_B(net589),
    .D(_00433_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][1] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _23714_ (.RESET_B(net588),
    .D(_00434_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][2] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _23715_ (.RESET_B(net587),
    .D(_00435_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][3] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _23716_ (.RESET_B(net586),
    .D(_00436_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][4] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _23717_ (.RESET_B(net585),
    .D(_00437_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][5] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _23718_ (.RESET_B(net584),
    .D(_00438_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][6] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _23719_ (.RESET_B(net583),
    .D(_00439_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][7] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _23720_ (.RESET_B(net582),
    .D(_00440_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][8] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _23721_ (.RESET_B(net581),
    .D(_00441_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][9] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _23722_ (.RESET_B(net580),
    .D(_00442_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][10] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _23723_ (.RESET_B(net579),
    .D(_00443_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][11] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _23724_ (.RESET_B(net578),
    .D(_00444_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][12] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _23725_ (.RESET_B(net577),
    .D(_00445_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][13] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _23726_ (.RESET_B(net576),
    .D(_00446_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][14] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _23727_ (.RESET_B(net575),
    .D(_00447_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][15] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _23728_ (.RESET_B(net574),
    .D(_00448_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][16] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _23729_ (.RESET_B(net573),
    .D(_00449_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][17] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _23730_ (.RESET_B(net572),
    .D(_00450_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][18] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _23731_ (.RESET_B(net571),
    .D(_00451_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _23732_ (.RESET_B(net570),
    .D(_00452_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][20] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _23733_ (.RESET_B(net569),
    .D(_00453_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][21] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _23734_ (.RESET_B(net568),
    .D(_00454_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][22] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _23735_ (.RESET_B(net567),
    .D(_00455_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][23] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _23736_ (.RESET_B(net566),
    .D(_00456_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][24] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _23737_ (.RESET_B(net565),
    .D(_00457_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _23738_ (.RESET_B(net564),
    .D(_00458_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][26] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _23739_ (.RESET_B(net563),
    .D(_00459_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][27] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _23740_ (.RESET_B(net562),
    .D(_00460_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][28] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _23741_ (.RESET_B(net561),
    .D(_00461_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][29] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _23742_ (.RESET_B(net560),
    .D(_00462_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][30] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _23743_ (.RESET_B(net559),
    .D(_00463_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][31] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _23744_ (.RESET_B(net558),
    .D(_00464_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][0] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _23745_ (.RESET_B(net557),
    .D(_00465_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][1] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _23746_ (.RESET_B(net556),
    .D(_00466_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][2] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _23747_ (.RESET_B(net555),
    .D(_00467_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][3] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _23748_ (.RESET_B(net554),
    .D(_00468_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][4] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _23749_ (.RESET_B(net553),
    .D(_00469_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][5] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _23750_ (.RESET_B(net552),
    .D(_00470_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][6] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _23751_ (.RESET_B(net551),
    .D(_00471_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][7] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _23752_ (.RESET_B(net550),
    .D(_00472_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][8] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _23753_ (.RESET_B(net549),
    .D(_00473_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][9] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _23754_ (.RESET_B(net548),
    .D(_00474_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][10] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _23755_ (.RESET_B(net547),
    .D(_00475_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][11] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _23756_ (.RESET_B(net546),
    .D(_00476_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][12] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _23757_ (.RESET_B(net545),
    .D(_00477_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][13] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _23758_ (.RESET_B(net544),
    .D(_00478_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][14] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _23759_ (.RESET_B(net543),
    .D(_00479_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][15] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _23760_ (.RESET_B(net542),
    .D(_00480_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][16] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _23761_ (.RESET_B(net541),
    .D(_00481_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][17] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _23762_ (.RESET_B(net540),
    .D(_00482_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][18] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _23763_ (.RESET_B(net539),
    .D(_00483_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _23764_ (.RESET_B(net538),
    .D(_00484_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][20] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _23765_ (.RESET_B(net537),
    .D(_00485_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][21] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _23766_ (.RESET_B(net536),
    .D(_00486_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][22] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _23767_ (.RESET_B(net535),
    .D(_00487_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][23] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _23768_ (.RESET_B(net534),
    .D(_00488_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][24] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _23769_ (.RESET_B(net533),
    .D(_00489_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][25] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _23770_ (.RESET_B(net532),
    .D(_00490_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][26] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _23771_ (.RESET_B(net531),
    .D(_00491_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][27] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _23772_ (.RESET_B(net530),
    .D(_00492_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][28] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _23773_ (.RESET_B(net529),
    .D(_00493_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][29] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _23774_ (.RESET_B(net528),
    .D(_00494_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][30] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _23775_ (.RESET_B(net527),
    .D(_00495_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][31] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _23776_ (.RESET_B(net526),
    .D(_00496_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][0] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _23777_ (.RESET_B(net525),
    .D(_00497_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][1] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _23778_ (.RESET_B(net524),
    .D(_00498_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][2] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _23779_ (.RESET_B(net523),
    .D(_00499_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][3] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _23780_ (.RESET_B(net522),
    .D(_00500_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][4] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _23781_ (.RESET_B(net521),
    .D(_00501_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][5] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _23782_ (.RESET_B(net520),
    .D(_00502_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][6] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _23783_ (.RESET_B(net519),
    .D(_00503_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][7] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _23784_ (.RESET_B(net518),
    .D(_00504_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][8] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _23785_ (.RESET_B(net517),
    .D(_00505_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][9] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _23786_ (.RESET_B(net516),
    .D(_00506_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][10] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _23787_ (.RESET_B(net515),
    .D(_00507_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][11] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _23788_ (.RESET_B(net514),
    .D(_00508_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][12] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _23789_ (.RESET_B(net513),
    .D(_00509_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][13] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _23790_ (.RESET_B(net512),
    .D(_00510_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][14] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _23791_ (.RESET_B(net511),
    .D(_00511_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][15] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _23792_ (.RESET_B(net510),
    .D(_00512_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][16] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _23793_ (.RESET_B(net509),
    .D(_00513_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][17] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _23794_ (.RESET_B(net508),
    .D(_00514_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][18] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _23795_ (.RESET_B(net507),
    .D(_00515_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _23796_ (.RESET_B(net506),
    .D(_00516_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _23797_ (.RESET_B(net505),
    .D(_00517_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][21] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _23798_ (.RESET_B(net504),
    .D(_00518_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][22] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _23799_ (.RESET_B(net503),
    .D(_00519_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][23] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _23800_ (.RESET_B(net502),
    .D(_00520_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][24] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _23801_ (.RESET_B(net501),
    .D(_00521_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _23802_ (.RESET_B(net500),
    .D(_00522_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][26] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _23803_ (.RESET_B(net499),
    .D(_00523_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][27] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _23804_ (.RESET_B(net498),
    .D(_00524_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][28] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _23805_ (.RESET_B(net497),
    .D(_00525_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][29] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _23806_ (.RESET_B(net496),
    .D(_00526_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][30] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _23807_ (.RESET_B(net124),
    .D(_00527_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][31] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _23808_ (.RESET_B(net5870),
    .D(net9),
    .Q(\fpga_top.qspi_if.sio_in_mt0[0] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _23809_ (.RESET_B(net5870),
    .D(net10),
    .Q(\fpga_top.qspi_if.sio_in_mt0[1] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _23810_ (.RESET_B(net5868),
    .D(net11),
    .Q(\fpga_top.qspi_if.sio_in_mt0[2] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _23811_ (.RESET_B(net5868),
    .D(net12),
    .Q(\fpga_top.qspi_if.sio_in_mt0[3] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _23812_ (.RESET_B(net5847),
    .D(_00042_),
    .Q(\fpga_top.qspi_if.sck_cntr[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _23813_ (.RESET_B(net5847),
    .D(_00043_),
    .Q(\fpga_top.qspi_if.sck_cntr[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _23814_ (.RESET_B(net5847),
    .D(_00044_),
    .Q(\fpga_top.qspi_if.sck_cntr[2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _23815_ (.RESET_B(net5841),
    .D(_00045_),
    .Q(\fpga_top.qspi_if.sck_cntr[3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _23816_ (.RESET_B(net5841),
    .D(_00046_),
    .Q(\fpga_top.qspi_if.sck_cntr[4] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _23817_ (.RESET_B(net5840),
    .D(_00047_),
    .Q(\fpga_top.qspi_if.sck_cntr[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _23818_ (.RESET_B(net5841),
    .D(net2005),
    .Q(\fpga_top.qspi_if.sck_cntr[6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _23819_ (.RESET_B(net5840),
    .D(_00049_),
    .Q(\fpga_top.qspi_if.sck_cntr[7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _23820_ (.RESET_B(net5840),
    .D(_00050_),
    .Q(\fpga_top.qspi_if.sck_cntr[8] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _23821_ (.RESET_B(net5840),
    .D(_00051_),
    .Q(\fpga_top.qspi_if.sck_cntr[9] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _23822_ (.RESET_B(net5884),
    .D(\fpga_top.qspi_if.sio_out_enbl_pre ),
    .Q(\fpga_top.qspi_if.sio_out_enbl_dly ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _23823_ (.RESET_B(net5927),
    .D(_00528_),
    .Q(\fpga_top.qspi_if.cmd_ofs[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _23824_ (.RESET_B(net5927),
    .D(_00529_),
    .Q(\fpga_top.qspi_if.cmd_ofs[1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _23825_ (.RESET_B(net5938),
    .D(_00530_),
    .Q(\fpga_top.qspi_if.cmd_ofs[2] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _23826_ (.RESET_B(net495),
    .D(_00531_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][0] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _23827_ (.RESET_B(net494),
    .D(_00532_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][1] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _23828_ (.RESET_B(net493),
    .D(_00533_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][2] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _23829_ (.RESET_B(net492),
    .D(_00534_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][3] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _23830_ (.RESET_B(net491),
    .D(_00535_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][4] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _23831_ (.RESET_B(net490),
    .D(_00536_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][5] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _23832_ (.RESET_B(net489),
    .D(_00537_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][6] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _23833_ (.RESET_B(net488),
    .D(_00538_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][7] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _23834_ (.RESET_B(net487),
    .D(_00539_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][8] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _23835_ (.RESET_B(net486),
    .D(_00540_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][9] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _23836_ (.RESET_B(net485),
    .D(_00541_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _23837_ (.RESET_B(net484),
    .D(_00542_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][11] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _23838_ (.RESET_B(net483),
    .D(_00543_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][12] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _23839_ (.RESET_B(net482),
    .D(_00544_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][13] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _23840_ (.RESET_B(net481),
    .D(_00545_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][14] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _23841_ (.RESET_B(net480),
    .D(_00546_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][15] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _23842_ (.RESET_B(net479),
    .D(_00547_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][16] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _23843_ (.RESET_B(net478),
    .D(_00548_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][17] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _23844_ (.RESET_B(net477),
    .D(_00549_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][18] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _23845_ (.RESET_B(net476),
    .D(_00550_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][19] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _23846_ (.RESET_B(net475),
    .D(_00551_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _23847_ (.RESET_B(net474),
    .D(_00552_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _23848_ (.RESET_B(net473),
    .D(_00553_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][22] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _23849_ (.RESET_B(net472),
    .D(_00554_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][23] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _23850_ (.RESET_B(net471),
    .D(_00555_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][24] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _23851_ (.RESET_B(net470),
    .D(_00556_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][25] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _23852_ (.RESET_B(net469),
    .D(_00557_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][26] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _23853_ (.RESET_B(net468),
    .D(_00558_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][27] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _23854_ (.RESET_B(net467),
    .D(_00559_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][28] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _23855_ (.RESET_B(net466),
    .D(_00560_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][29] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _23856_ (.RESET_B(net465),
    .D(_00561_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][30] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _23857_ (.RESET_B(net464),
    .D(_00562_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][31] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _23858_ (.RESET_B(net463),
    .D(_00563_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][0] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _23859_ (.RESET_B(net462),
    .D(_00564_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][1] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _23860_ (.RESET_B(net461),
    .D(_00565_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][2] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _23861_ (.RESET_B(net460),
    .D(_00566_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][3] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _23862_ (.RESET_B(net459),
    .D(_00567_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][4] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _23863_ (.RESET_B(net458),
    .D(_00568_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][5] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _23864_ (.RESET_B(net457),
    .D(_00569_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][6] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _23865_ (.RESET_B(net456),
    .D(_00570_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][7] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _23866_ (.RESET_B(net455),
    .D(_00571_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][8] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _23867_ (.RESET_B(net454),
    .D(_00572_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][9] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _23868_ (.RESET_B(net453),
    .D(_00573_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _23869_ (.RESET_B(net452),
    .D(_00574_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][11] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _23870_ (.RESET_B(net451),
    .D(_00575_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][12] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _23871_ (.RESET_B(net450),
    .D(_00576_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][13] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_1 _23872_ (.RESET_B(net449),
    .D(_00577_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][14] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _23873_ (.RESET_B(net448),
    .D(_00578_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][15] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _23874_ (.RESET_B(net447),
    .D(_00579_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][16] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _23875_ (.RESET_B(net446),
    .D(_00580_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][17] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _23876_ (.RESET_B(net445),
    .D(_00581_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][18] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _23877_ (.RESET_B(net444),
    .D(_00582_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _23878_ (.RESET_B(net443),
    .D(_00583_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][20] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _23879_ (.RESET_B(net442),
    .D(_00584_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][21] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _23880_ (.RESET_B(net441),
    .D(_00585_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][22] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _23881_ (.RESET_B(net440),
    .D(_00586_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][23] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _23882_ (.RESET_B(net439),
    .D(_00587_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][24] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _23883_ (.RESET_B(net438),
    .D(_00588_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][25] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _23884_ (.RESET_B(net437),
    .D(_00589_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][26] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _23885_ (.RESET_B(net436),
    .D(_00590_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][27] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _23886_ (.RESET_B(net435),
    .D(_00591_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][28] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _23887_ (.RESET_B(net434),
    .D(_00592_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][29] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _23888_ (.RESET_B(net433),
    .D(_00593_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][30] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _23889_ (.RESET_B(net192),
    .D(_00594_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][31] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _23890_ (.RESET_B(net5885),
    .D(net1315),
    .Q(\fpga_top.qspi_if.sio_in_sync[0] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _23891_ (.RESET_B(net5940),
    .D(net1323),
    .Q(\fpga_top.qspi_if.sio_in_sync[1] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _23892_ (.RESET_B(net5950),
    .D(net1361),
    .Q(\fpga_top.qspi_if.sio_in_sync[2] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _23893_ (.RESET_B(net5885),
    .D(net1366),
    .Q(\fpga_top.qspi_if.sio_in_sync[3] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _23894_ (.RESET_B(net432),
    .D(_00595_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][0] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _23895_ (.RESET_B(net431),
    .D(_00596_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][1] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _23896_ (.RESET_B(net430),
    .D(_00597_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][2] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _23897_ (.RESET_B(net429),
    .D(_00598_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][3] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _23898_ (.RESET_B(net428),
    .D(_00599_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][4] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _23899_ (.RESET_B(net427),
    .D(_00600_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][5] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _23900_ (.RESET_B(net426),
    .D(_00601_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][6] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _23901_ (.RESET_B(net425),
    .D(_00602_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][7] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _23902_ (.RESET_B(net424),
    .D(_00603_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][8] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _23903_ (.RESET_B(net423),
    .D(_00604_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][9] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _23904_ (.RESET_B(net422),
    .D(_00605_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _23905_ (.RESET_B(net421),
    .D(_00606_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][11] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _23906_ (.RESET_B(net420),
    .D(_00607_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][12] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _23907_ (.RESET_B(net419),
    .D(_00608_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][13] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _23908_ (.RESET_B(net418),
    .D(_00609_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][14] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _23909_ (.RESET_B(net417),
    .D(_00610_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][15] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _23910_ (.RESET_B(net416),
    .D(_00611_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][16] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _23911_ (.RESET_B(net415),
    .D(_00612_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][17] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _23912_ (.RESET_B(net414),
    .D(_00613_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][18] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _23913_ (.RESET_B(net413),
    .D(_00614_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][19] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _23914_ (.RESET_B(net412),
    .D(_00615_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _23915_ (.RESET_B(net411),
    .D(_00616_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _23916_ (.RESET_B(net410),
    .D(_00617_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][22] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _23917_ (.RESET_B(net409),
    .D(_00618_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][23] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _23918_ (.RESET_B(net408),
    .D(_00619_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][24] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _23919_ (.RESET_B(net407),
    .D(_00620_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][25] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _23920_ (.RESET_B(net406),
    .D(_00621_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][26] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _23921_ (.RESET_B(net405),
    .D(_00622_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][27] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _23922_ (.RESET_B(net404),
    .D(_00623_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][28] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _23923_ (.RESET_B(net403),
    .D(_00624_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][29] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _23924_ (.RESET_B(net402),
    .D(_00625_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][30] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _23925_ (.RESET_B(net401),
    .D(_00626_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][31] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _23926_ (.RESET_B(net400),
    .D(_00627_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][0] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_1 _23927_ (.RESET_B(net399),
    .D(_00628_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][1] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _23928_ (.RESET_B(net398),
    .D(_00629_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][2] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _23929_ (.RESET_B(net397),
    .D(_00630_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][3] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _23930_ (.RESET_B(net396),
    .D(_00631_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][4] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _23931_ (.RESET_B(net395),
    .D(_00632_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][5] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _23932_ (.RESET_B(net394),
    .D(_00633_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][6] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _23933_ (.RESET_B(net393),
    .D(_00634_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][7] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _23934_ (.RESET_B(net392),
    .D(_00635_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][8] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _23935_ (.RESET_B(net391),
    .D(_00636_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][9] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _23936_ (.RESET_B(net390),
    .D(_00637_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][10] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _23937_ (.RESET_B(net389),
    .D(_00638_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][11] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _23938_ (.RESET_B(net388),
    .D(_00639_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][12] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _23939_ (.RESET_B(net387),
    .D(_00640_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][13] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _23940_ (.RESET_B(net386),
    .D(_00641_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][14] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _23941_ (.RESET_B(net385),
    .D(_00642_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][15] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _23942_ (.RESET_B(net383),
    .D(_00643_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][16] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _23943_ (.RESET_B(net382),
    .D(_00644_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][17] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _23944_ (.RESET_B(net381),
    .D(_00645_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][18] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _23945_ (.RESET_B(net380),
    .D(_00646_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][19] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _23946_ (.RESET_B(net379),
    .D(_00647_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][20] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _23947_ (.RESET_B(net378),
    .D(_00648_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][21] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _23948_ (.RESET_B(net377),
    .D(_00649_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][22] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _23949_ (.RESET_B(net376),
    .D(_00650_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][23] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _23950_ (.RESET_B(net375),
    .D(_00651_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][24] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _23951_ (.RESET_B(net374),
    .D(_00652_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][25] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _23952_ (.RESET_B(net373),
    .D(_00653_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][26] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _23953_ (.RESET_B(net372),
    .D(_00654_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][27] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _23954_ (.RESET_B(net371),
    .D(_00655_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][28] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _23955_ (.RESET_B(net370),
    .D(_00656_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][29] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _23956_ (.RESET_B(net369),
    .D(_00657_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][30] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _23957_ (.RESET_B(net368),
    .D(_00658_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][31] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _23958_ (.RESET_B(net367),
    .D(_00659_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][0] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _23959_ (.RESET_B(net366),
    .D(_00660_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][1] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _23960_ (.RESET_B(net365),
    .D(_00661_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][2] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _23961_ (.RESET_B(net364),
    .D(_00662_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][3] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _23962_ (.RESET_B(net363),
    .D(_00663_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][4] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _23963_ (.RESET_B(net362),
    .D(_00664_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][5] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _23964_ (.RESET_B(net361),
    .D(_00665_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][6] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _23965_ (.RESET_B(net360),
    .D(_00666_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][7] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _23966_ (.RESET_B(net359),
    .D(_00667_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][8] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _23967_ (.RESET_B(net358),
    .D(_00668_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][9] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _23968_ (.RESET_B(net357),
    .D(_00669_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][10] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _23969_ (.RESET_B(net356),
    .D(_00670_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][11] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _23970_ (.RESET_B(net355),
    .D(_00671_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][12] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _23971_ (.RESET_B(net354),
    .D(_00672_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][13] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _23972_ (.RESET_B(net353),
    .D(_00673_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][14] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _23973_ (.RESET_B(net352),
    .D(_00674_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][15] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _23974_ (.RESET_B(net351),
    .D(_00675_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][16] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _23975_ (.RESET_B(net350),
    .D(_00676_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][17] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _23976_ (.RESET_B(net349),
    .D(_00677_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][18] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _23977_ (.RESET_B(net348),
    .D(_00678_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][19] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _23978_ (.RESET_B(net347),
    .D(_00679_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _23979_ (.RESET_B(net346),
    .D(_00680_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _23980_ (.RESET_B(net345),
    .D(_00681_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][22] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _23981_ (.RESET_B(net344),
    .D(_00682_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][23] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _23982_ (.RESET_B(net343),
    .D(_00683_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][24] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _23983_ (.RESET_B(net342),
    .D(_00684_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][25] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _23984_ (.RESET_B(net341),
    .D(_00685_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][26] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _23985_ (.RESET_B(net340),
    .D(_00686_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][27] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _23986_ (.RESET_B(net339),
    .D(_00687_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][28] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _23987_ (.RESET_B(net338),
    .D(_00688_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][29] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _23988_ (.RESET_B(net337),
    .D(_00689_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][30] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _23989_ (.RESET_B(net336),
    .D(_00690_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][31] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _23990_ (.RESET_B(net335),
    .D(_00691_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][0] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _23991_ (.RESET_B(net334),
    .D(_00692_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][1] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _23992_ (.RESET_B(net333),
    .D(_00693_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][2] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _23993_ (.RESET_B(net332),
    .D(_00694_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][3] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _23994_ (.RESET_B(net331),
    .D(_00695_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][4] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _23995_ (.RESET_B(net330),
    .D(_00696_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][5] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _23996_ (.RESET_B(net329),
    .D(_00697_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][6] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _23997_ (.RESET_B(net328),
    .D(_00698_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][7] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _23998_ (.RESET_B(net327),
    .D(_00699_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][8] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _23999_ (.RESET_B(net326),
    .D(_00700_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][9] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _24000_ (.RESET_B(net325),
    .D(_00701_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _24001_ (.RESET_B(net324),
    .D(_00702_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][11] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _24002_ (.RESET_B(net323),
    .D(_00703_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][12] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _24003_ (.RESET_B(net322),
    .D(_00704_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][13] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _24004_ (.RESET_B(net321),
    .D(_00705_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][14] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _24005_ (.RESET_B(net320),
    .D(_00706_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][15] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _24006_ (.RESET_B(net319),
    .D(_00707_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][16] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _24007_ (.RESET_B(net318),
    .D(_00708_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][17] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _24008_ (.RESET_B(net317),
    .D(_00709_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][18] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _24009_ (.RESET_B(net316),
    .D(_00710_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][19] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _24010_ (.RESET_B(net315),
    .D(_00711_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _24011_ (.RESET_B(net314),
    .D(_00712_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _24012_ (.RESET_B(net313),
    .D(_00713_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][22] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _24013_ (.RESET_B(net312),
    .D(_00714_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][23] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _24014_ (.RESET_B(net311),
    .D(_00715_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][24] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _24015_ (.RESET_B(net310),
    .D(_00716_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][25] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _24016_ (.RESET_B(net309),
    .D(_00717_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][26] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _24017_ (.RESET_B(net308),
    .D(_00718_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][27] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _24018_ (.RESET_B(net307),
    .D(_00719_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][28] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _24019_ (.RESET_B(net306),
    .D(_00720_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][29] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _24020_ (.RESET_B(net305),
    .D(_00721_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][30] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _24021_ (.RESET_B(net304),
    .D(_00722_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][31] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _24022_ (.RESET_B(net303),
    .D(_00723_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][0] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _24023_ (.RESET_B(net302),
    .D(_00724_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][1] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _24024_ (.RESET_B(net301),
    .D(_00725_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][2] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _24025_ (.RESET_B(net300),
    .D(_00726_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][3] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _24026_ (.RESET_B(net299),
    .D(_00727_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][4] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _24027_ (.RESET_B(net298),
    .D(_00728_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][5] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _24028_ (.RESET_B(net297),
    .D(_00729_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][6] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _24029_ (.RESET_B(net296),
    .D(_00730_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][7] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _24030_ (.RESET_B(net295),
    .D(_00731_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][8] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _24031_ (.RESET_B(net294),
    .D(_00732_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][9] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _24032_ (.RESET_B(net293),
    .D(_00733_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][10] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _24033_ (.RESET_B(net292),
    .D(_00734_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][11] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _24034_ (.RESET_B(net291),
    .D(_00735_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][12] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _24035_ (.RESET_B(net290),
    .D(_00736_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][13] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _24036_ (.RESET_B(net289),
    .D(_00737_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][14] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _24037_ (.RESET_B(net288),
    .D(_00738_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][15] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _24038_ (.RESET_B(net287),
    .D(_00739_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][16] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _24039_ (.RESET_B(net286),
    .D(_00740_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][17] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _24040_ (.RESET_B(net285),
    .D(_00741_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][18] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _24041_ (.RESET_B(net284),
    .D(_00742_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][19] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _24042_ (.RESET_B(net283),
    .D(_00743_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][20] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _24043_ (.RESET_B(net282),
    .D(_00744_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _24044_ (.RESET_B(net281),
    .D(_00745_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][22] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _24045_ (.RESET_B(net280),
    .D(_00746_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][23] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _24046_ (.RESET_B(net279),
    .D(_00747_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][24] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _24047_ (.RESET_B(net278),
    .D(_00748_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][25] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _24048_ (.RESET_B(net277),
    .D(_00749_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][26] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _24049_ (.RESET_B(net276),
    .D(_00750_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][27] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _24050_ (.RESET_B(net275),
    .D(_00751_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][28] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _24051_ (.RESET_B(net274),
    .D(_00752_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][29] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _24052_ (.RESET_B(net273),
    .D(_00753_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][30] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _24053_ (.RESET_B(net272),
    .D(_00754_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][31] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _24054_ (.RESET_B(net271),
    .D(_00755_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][0] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _24055_ (.RESET_B(net270),
    .D(_00756_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][1] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _24056_ (.RESET_B(net269),
    .D(_00757_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][2] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _24057_ (.RESET_B(net268),
    .D(_00758_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][3] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _24058_ (.RESET_B(net267),
    .D(_00759_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][4] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _24059_ (.RESET_B(net266),
    .D(_00760_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][5] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _24060_ (.RESET_B(net265),
    .D(_00761_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][6] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _24061_ (.RESET_B(net264),
    .D(_00762_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][7] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _24062_ (.RESET_B(net263),
    .D(_00763_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][8] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _24063_ (.RESET_B(net262),
    .D(_00764_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][9] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _24064_ (.RESET_B(net261),
    .D(_00765_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _24065_ (.RESET_B(net260),
    .D(_00766_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][11] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _24066_ (.RESET_B(net259),
    .D(_00767_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][12] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _24067_ (.RESET_B(net258),
    .D(_00768_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][13] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _24068_ (.RESET_B(net257),
    .D(_00769_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][14] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _24069_ (.RESET_B(net256),
    .D(_00770_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][15] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _24070_ (.RESET_B(net255),
    .D(_00771_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][16] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _24071_ (.RESET_B(net254),
    .D(_00772_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][17] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _24072_ (.RESET_B(net253),
    .D(_00773_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][18] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _24073_ (.RESET_B(net252),
    .D(_00774_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][19] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _24074_ (.RESET_B(net251),
    .D(_00775_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][20] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _24075_ (.RESET_B(net250),
    .D(_00776_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _24076_ (.RESET_B(net249),
    .D(_00777_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][22] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _24077_ (.RESET_B(net248),
    .D(_00778_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][23] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _24078_ (.RESET_B(net247),
    .D(_00779_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][24] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _24079_ (.RESET_B(net246),
    .D(_00780_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][25] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _24080_ (.RESET_B(net245),
    .D(_00781_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][26] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _24081_ (.RESET_B(net244),
    .D(_00782_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][27] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _24082_ (.RESET_B(net243),
    .D(_00783_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][28] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _24083_ (.RESET_B(net242),
    .D(_00784_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][29] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _24084_ (.RESET_B(net241),
    .D(_00785_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][30] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _24085_ (.RESET_B(net384),
    .D(_00786_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][31] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _24086_ (.RESET_B(net5955),
    .D(\fpga_top.qspi_if.sio_out_pre[0] ),
    .Q(\fpga_top.qspi_if.sio_out_dly[0] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24087_ (.RESET_B(net5954),
    .D(net6339),
    .Q(\fpga_top.qspi_if.sio_out_dly[1] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _24088_ (.RESET_B(net5936),
    .D(\fpga_top.qspi_if.sio_out_pre[2] ),
    .Q(\fpga_top.qspi_if.sio_out_dly[2] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24089_ (.RESET_B(net5940),
    .D(\fpga_top.qspi_if.sio_out_pre[3] ),
    .Q(\fpga_top.qspi_if.sio_out_dly[3] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24090_ (.RESET_B(net240),
    .D(_00787_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][0] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _24091_ (.RESET_B(net239),
    .D(_00788_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][1] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _24092_ (.RESET_B(net238),
    .D(_00789_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][2] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _24093_ (.RESET_B(net237),
    .D(_00790_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][3] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _24094_ (.RESET_B(net236),
    .D(_00791_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][4] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _24095_ (.RESET_B(net235),
    .D(_00792_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][5] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _24096_ (.RESET_B(net234),
    .D(_00793_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][6] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _24097_ (.RESET_B(net233),
    .D(_00794_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][7] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _24098_ (.RESET_B(net232),
    .D(_00795_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][8] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _24099_ (.RESET_B(net231),
    .D(_00796_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][9] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _24100_ (.RESET_B(net230),
    .D(_00797_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _24101_ (.RESET_B(net229),
    .D(_00798_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][11] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _24102_ (.RESET_B(net228),
    .D(_00799_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][12] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _24103_ (.RESET_B(net227),
    .D(_00800_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][13] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _24104_ (.RESET_B(net226),
    .D(_00801_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][14] ),
    .CLK(clknet_leaf_263_clk));
 sg13g2_dfrbpq_1 _24105_ (.RESET_B(net225),
    .D(_00802_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][15] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _24106_ (.RESET_B(net224),
    .D(_00803_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][16] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _24107_ (.RESET_B(net223),
    .D(_00804_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][17] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _24108_ (.RESET_B(net222),
    .D(_00805_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][18] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _24109_ (.RESET_B(net221),
    .D(_00806_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][19] ),
    .CLK(clknet_leaf_249_clk));
 sg13g2_dfrbpq_1 _24110_ (.RESET_B(net220),
    .D(_00807_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][20] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _24111_ (.RESET_B(net219),
    .D(_00808_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][21] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _24112_ (.RESET_B(net218),
    .D(_00809_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][22] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _24113_ (.RESET_B(net217),
    .D(_00810_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][23] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _24114_ (.RESET_B(net216),
    .D(_00811_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][24] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _24115_ (.RESET_B(net215),
    .D(_00812_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][25] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _24116_ (.RESET_B(net214),
    .D(_00813_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][26] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _24117_ (.RESET_B(net213),
    .D(_00814_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][27] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _24118_ (.RESET_B(net212),
    .D(_00815_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][28] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _24119_ (.RESET_B(net211),
    .D(_00816_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][29] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _24120_ (.RESET_B(net210),
    .D(_00817_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][30] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_1 _24121_ (.RESET_B(net209),
    .D(_00818_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][31] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _24122_ (.RESET_B(net208),
    .D(_00819_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][0] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _24123_ (.RESET_B(net207),
    .D(_00820_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][1] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_1 _24124_ (.RESET_B(net206),
    .D(_00821_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][2] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _24125_ (.RESET_B(net205),
    .D(_00822_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][3] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _24126_ (.RESET_B(net204),
    .D(_00823_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][4] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _24127_ (.RESET_B(net203),
    .D(_00824_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][5] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _24128_ (.RESET_B(net202),
    .D(_00825_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][6] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _24129_ (.RESET_B(net201),
    .D(_00826_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][7] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _24130_ (.RESET_B(net200),
    .D(_00827_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][8] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _24131_ (.RESET_B(net199),
    .D(_00828_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][9] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _24132_ (.RESET_B(net198),
    .D(_00829_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][10] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _24133_ (.RESET_B(net197),
    .D(_00830_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][11] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _24134_ (.RESET_B(net196),
    .D(_00831_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][12] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _24135_ (.RESET_B(net195),
    .D(_00832_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][13] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _24136_ (.RESET_B(net194),
    .D(_00833_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][14] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _24137_ (.RESET_B(net193),
    .D(_00834_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][15] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _24138_ (.RESET_B(net191),
    .D(_00835_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][16] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _24139_ (.RESET_B(net190),
    .D(_00836_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][17] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _24140_ (.RESET_B(net189),
    .D(_00837_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][18] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _24141_ (.RESET_B(net188),
    .D(_00838_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][19] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _24142_ (.RESET_B(net187),
    .D(_00839_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][20] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _24143_ (.RESET_B(net186),
    .D(_00840_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][21] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _24144_ (.RESET_B(net185),
    .D(_00841_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][22] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _24145_ (.RESET_B(net184),
    .D(_00842_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][23] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _24146_ (.RESET_B(net183),
    .D(_00843_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][24] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _24147_ (.RESET_B(net182),
    .D(_00844_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _24148_ (.RESET_B(net181),
    .D(_00845_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][26] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _24149_ (.RESET_B(net180),
    .D(_00846_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][27] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _24150_ (.RESET_B(net179),
    .D(_00847_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][28] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _24151_ (.RESET_B(net178),
    .D(_00848_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][29] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _24152_ (.RESET_B(net177),
    .D(_00849_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][30] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _24153_ (.RESET_B(net176),
    .D(_00850_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][31] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _24154_ (.RESET_B(net175),
    .D(_00851_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][0] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _24155_ (.RESET_B(net174),
    .D(_00852_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][1] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _24156_ (.RESET_B(net173),
    .D(_00853_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][2] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _24157_ (.RESET_B(net172),
    .D(_00854_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][3] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _24158_ (.RESET_B(net171),
    .D(_00855_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][4] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _24159_ (.RESET_B(net170),
    .D(_00856_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _24160_ (.RESET_B(net169),
    .D(_00857_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][6] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _24161_ (.RESET_B(net168),
    .D(_00858_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][7] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _24162_ (.RESET_B(net167),
    .D(_00859_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][8] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _24163_ (.RESET_B(net166),
    .D(_00860_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][9] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _24164_ (.RESET_B(net165),
    .D(_00861_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][10] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _24165_ (.RESET_B(net164),
    .D(_00862_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][11] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _24166_ (.RESET_B(net163),
    .D(_00863_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][12] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _24167_ (.RESET_B(net162),
    .D(_00864_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][13] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _24168_ (.RESET_B(net161),
    .D(_00865_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][14] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _24169_ (.RESET_B(net160),
    .D(_00866_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][15] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _24170_ (.RESET_B(net159),
    .D(_00867_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][16] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _24171_ (.RESET_B(net158),
    .D(_00868_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][17] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _24172_ (.RESET_B(net157),
    .D(_00869_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][18] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _24173_ (.RESET_B(net156),
    .D(_00870_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][19] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _24174_ (.RESET_B(net155),
    .D(_00871_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][20] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _24175_ (.RESET_B(net154),
    .D(_00872_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][21] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _24176_ (.RESET_B(net153),
    .D(_00873_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][22] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _24177_ (.RESET_B(net152),
    .D(_00874_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][23] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _24178_ (.RESET_B(net151),
    .D(_00875_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][24] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _24179_ (.RESET_B(net150),
    .D(_00876_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][25] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _24180_ (.RESET_B(net149),
    .D(_00877_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][26] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _24181_ (.RESET_B(net148),
    .D(_00878_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][27] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _24182_ (.RESET_B(net147),
    .D(_00879_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _24183_ (.RESET_B(net146),
    .D(_00880_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][29] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _24184_ (.RESET_B(net145),
    .D(_00881_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][30] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _24185_ (.RESET_B(net144),
    .D(_00882_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _24186_ (.RESET_B(net143),
    .D(_00883_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][0] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _24187_ (.RESET_B(net142),
    .D(_00884_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][1] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _24188_ (.RESET_B(net141),
    .D(_00885_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][2] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _24189_ (.RESET_B(net140),
    .D(_00886_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][3] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _24190_ (.RESET_B(net139),
    .D(_00887_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][4] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _24191_ (.RESET_B(net138),
    .D(_00888_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _24192_ (.RESET_B(net137),
    .D(_00889_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][6] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _24193_ (.RESET_B(net136),
    .D(_00890_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][7] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _24194_ (.RESET_B(net135),
    .D(_00891_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][8] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _24195_ (.RESET_B(net134),
    .D(_00892_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][9] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _24196_ (.RESET_B(net133),
    .D(_00893_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][10] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _24197_ (.RESET_B(net132),
    .D(_00894_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][11] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _24198_ (.RESET_B(net131),
    .D(_00895_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][12] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _24199_ (.RESET_B(net130),
    .D(_00896_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][13] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _24200_ (.RESET_B(net129),
    .D(_00897_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][14] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _24201_ (.RESET_B(net128),
    .D(_00898_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][15] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _24202_ (.RESET_B(net127),
    .D(_00899_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][16] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _24203_ (.RESET_B(net126),
    .D(_00900_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][17] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _24204_ (.RESET_B(net125),
    .D(_00901_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][18] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _24205_ (.RESET_B(net123),
    .D(_00902_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][19] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _24206_ (.RESET_B(net122),
    .D(_00903_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][20] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _24207_ (.RESET_B(net121),
    .D(_00904_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][21] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _24208_ (.RESET_B(net120),
    .D(_00905_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][22] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _24209_ (.RESET_B(net119),
    .D(_00906_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][23] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _24210_ (.RESET_B(net118),
    .D(_00907_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][24] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _24211_ (.RESET_B(net117),
    .D(_00908_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _24212_ (.RESET_B(net116),
    .D(_00909_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][26] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _24213_ (.RESET_B(net115),
    .D(_00910_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][27] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _24214_ (.RESET_B(net114),
    .D(_00911_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _24215_ (.RESET_B(net113),
    .D(_00912_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][29] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _24216_ (.RESET_B(net112),
    .D(_00913_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][30] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _24217_ (.RESET_B(net111),
    .D(_00914_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _24218_ (.RESET_B(net5854),
    .D(_00128_),
    .Q(_00086_),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _24219_ (.RESET_B(net5934),
    .D(_00915_),
    .Q(\fpga_top.io_uart_out.uart_io_char[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _24220_ (.RESET_B(net5884),
    .D(_00916_),
    .Q(\fpga_top.io_uart_out.uart_io_char[1] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _24221_ (.RESET_B(net5884),
    .D(_00917_),
    .Q(\fpga_top.io_uart_out.uart_io_char[2] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _24222_ (.RESET_B(net5934),
    .D(_00918_),
    .Q(\fpga_top.io_uart_out.uart_io_char[3] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _24223_ (.RESET_B(net5923),
    .D(_00919_),
    .Q(\fpga_top.io_uart_out.uart_io_char[4] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _24224_ (.RESET_B(net5926),
    .D(_00920_),
    .Q(\fpga_top.io_uart_out.uart_io_char[5] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _24225_ (.RESET_B(net5926),
    .D(_00921_),
    .Q(\fpga_top.io_uart_out.uart_io_char[6] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _24226_ (.RESET_B(net5923),
    .D(_00922_),
    .Q(\fpga_top.io_uart_out.uart_io_char[7] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _24227_ (.RESET_B(net5937),
    .D(net1375),
    .Q(\fpga_top.qspi_if.dbg_2div_cew_lat ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24228_ (.RESET_B(net5948),
    .D(_00923_),
    .Q(\fpga_top.qspi_if.wdata[0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _24229_ (.RESET_B(net5948),
    .D(_00924_),
    .Q(\fpga_top.qspi_if.wdata[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24230_ (.RESET_B(net5953),
    .D(net2797),
    .Q(\fpga_top.qspi_if.wdata[2] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24231_ (.RESET_B(net5953),
    .D(_00926_),
    .Q(\fpga_top.qspi_if.wdata[3] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _24232_ (.RESET_B(net6000),
    .D(_00927_),
    .Q(\fpga_top.qspi_if.wdata[4] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _24233_ (.RESET_B(net5947),
    .D(_00928_),
    .Q(\fpga_top.qspi_if.wdata[5] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _24234_ (.RESET_B(net5953),
    .D(net1783),
    .Q(\fpga_top.qspi_if.wdata[6] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24235_ (.RESET_B(net5953),
    .D(net1905),
    .Q(\fpga_top.qspi_if.wdata[7] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _24236_ (.RESET_B(net5947),
    .D(net1839),
    .Q(\fpga_top.qspi_if.wdata[8] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _24237_ (.RESET_B(net5953),
    .D(net1668),
    .Q(\fpga_top.qspi_if.wdata[9] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _24238_ (.RESET_B(net5953),
    .D(_00933_),
    .Q(\fpga_top.qspi_if.wdata[10] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _24239_ (.RESET_B(net6005),
    .D(net2116),
    .Q(\fpga_top.qspi_if.wdata[11] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _24240_ (.RESET_B(net6000),
    .D(net6245),
    .Q(\fpga_top.qspi_if.wdata[12] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _24241_ (.RESET_B(net5953),
    .D(net6237),
    .Q(\fpga_top.qspi_if.wdata[13] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _24242_ (.RESET_B(net6005),
    .D(net6185),
    .Q(\fpga_top.qspi_if.wdata[14] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _24243_ (.RESET_B(net5999),
    .D(_00938_),
    .Q(\fpga_top.qspi_if.wdata[15] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _24244_ (.RESET_B(net5948),
    .D(_00939_),
    .Q(\fpga_top.qspi_if.wdata[16] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24245_ (.RESET_B(net5948),
    .D(net6223),
    .Q(\fpga_top.qspi_if.wdata[17] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24246_ (.RESET_B(net6006),
    .D(net6128),
    .Q(\fpga_top.qspi_if.wdata[18] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _24247_ (.RESET_B(net6000),
    .D(net4032),
    .Q(\fpga_top.qspi_if.wdata[19] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _24248_ (.RESET_B(net5948),
    .D(_00943_),
    .Q(\fpga_top.qspi_if.wdata[20] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24249_ (.RESET_B(net6000),
    .D(net3963),
    .Q(\fpga_top.qspi_if.wdata[21] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _24250_ (.RESET_B(net6000),
    .D(net3992),
    .Q(\fpga_top.qspi_if.wdata[22] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _24251_ (.RESET_B(net5999),
    .D(net4060),
    .Q(\fpga_top.qspi_if.wdata[23] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _24252_ (.RESET_B(net5999),
    .D(net6105),
    .Q(\fpga_top.qspi_if.wdata[24] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _24253_ (.RESET_B(net6006),
    .D(net6146),
    .Q(\fpga_top.qspi_if.wdata[25] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _24254_ (.RESET_B(net6005),
    .D(net4064),
    .Q(\fpga_top.qspi_if.wdata[26] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _24255_ (.RESET_B(net5947),
    .D(net3984),
    .Q(\fpga_top.qspi_if.wdata[27] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _24256_ (.RESET_B(net5948),
    .D(net4071),
    .Q(\fpga_top.qspi_if.wdata[28] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24257_ (.RESET_B(net5947),
    .D(net6178),
    .Q(\fpga_top.qspi_if.wdata[29] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _24258_ (.RESET_B(net5947),
    .D(net6114),
    .Q(\fpga_top.qspi_if.wdata[30] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _24259_ (.RESET_B(net5999),
    .D(net3877),
    .Q(\fpga_top.qspi_if.wdata[31] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _24260_ (.RESET_B(net6006),
    .D(net6578),
    .Q(\fpga_top.qspi_if.word_w ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _24261_ (.RESET_B(net5854),
    .D(_00129_),
    .Q(_00087_),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _24262_ (.RESET_B(net6005),
    .D(net6328),
    .Q(\fpga_top.qspi_if.word_hw ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _24263_ (.RESET_B(net5951),
    .D(net3738),
    .Q(\fpga_top.qspi_if.word_data[0] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _24264_ (.RESET_B(net6007),
    .D(net3766),
    .Q(\fpga_top.qspi_if.word_data[1] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _24265_ (.RESET_B(net5955),
    .D(net1630),
    .Q(\fpga_top.qspi_if.word_data[2] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _24266_ (.RESET_B(net5955),
    .D(net3744),
    .Q(\fpga_top.qspi_if.word_data[3] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _24267_ (.RESET_B(net6012),
    .D(net3289),
    .Q(\fpga_top.qspi_if.word_data[4] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _24268_ (.RESET_B(net6023),
    .D(net2096),
    .Q(\fpga_top.qspi_if.word_data[5] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24269_ (.RESET_B(net6023),
    .D(net3880),
    .Q(\fpga_top.qspi_if.word_data[6] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _24270_ (.RESET_B(net6025),
    .D(net3791),
    .Q(\fpga_top.qspi_if.word_data[7] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _24271_ (.RESET_B(net6012),
    .D(_00965_),
    .Q(\fpga_top.qspi_if.word_data[8] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _24272_ (.RESET_B(net6025),
    .D(_00966_),
    .Q(\fpga_top.qspi_if.word_data[9] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _24273_ (.RESET_B(net6024),
    .D(net1864),
    .Q(\fpga_top.qspi_if.word_data[10] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _24274_ (.RESET_B(net6012),
    .D(net2000),
    .Q(\fpga_top.qspi_if.word_data[11] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _24275_ (.RESET_B(net6012),
    .D(net3729),
    .Q(\fpga_top.qspi_if.word_data[12] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _24276_ (.RESET_B(net6025),
    .D(net1719),
    .Q(\fpga_top.qspi_if.word_data[13] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24277_ (.RESET_B(net6025),
    .D(_00971_),
    .Q(\fpga_top.qspi_if.word_data[14] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _24278_ (.RESET_B(net6012),
    .D(net1911),
    .Q(\fpga_top.qspi_if.word_data[15] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _24279_ (.RESET_B(net6012),
    .D(net2007),
    .Q(\fpga_top.qspi_if.word_data[16] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _24280_ (.RESET_B(net6023),
    .D(net1611),
    .Q(\fpga_top.qspi_if.word_data[17] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _24281_ (.RESET_B(net6023),
    .D(net1785),
    .Q(\fpga_top.qspi_if.word_data[18] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _24282_ (.RESET_B(net6025),
    .D(net1847),
    .Q(\fpga_top.qspi_if.word_data[19] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _24283_ (.RESET_B(net6025),
    .D(net1658),
    .Q(\fpga_top.qspi_if.word_data[20] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _24284_ (.RESET_B(net6023),
    .D(_00978_),
    .Q(\fpga_top.qspi_if.word_data[21] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _24285_ (.RESET_B(net6023),
    .D(net1670),
    .Q(\fpga_top.qspi_if.word_data[22] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _24286_ (.RESET_B(net6025),
    .D(_00980_),
    .Q(\fpga_top.qspi_if.word_data[23] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _24287_ (.RESET_B(net6012),
    .D(_00981_),
    .Q(\fpga_top.qspi_if.word_data[24] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _24288_ (.RESET_B(net6024),
    .D(_00982_),
    .Q(\fpga_top.qspi_if.word_data[25] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _24289_ (.RESET_B(net6023),
    .D(_00983_),
    .Q(\fpga_top.qspi_if.word_data[26] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _24290_ (.RESET_B(net6025),
    .D(net1684),
    .Q(\fpga_top.qspi_if.word_data[27] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _24291_ (.RESET_B(net6012),
    .D(net1498),
    .Q(\fpga_top.qspi_if.word_data[28] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _24292_ (.RESET_B(net6024),
    .D(net1616),
    .Q(\fpga_top.qspi_if.word_data[29] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _24293_ (.RESET_B(net6023),
    .D(net1443),
    .Q(\fpga_top.qspi_if.word_data[30] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _24294_ (.RESET_B(net6013),
    .D(net1403),
    .Q(\fpga_top.qspi_if.word_data[31] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _24295_ (.RESET_B(net5950),
    .D(\fpga_top.qspi_if.inner_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/qspi_if.v:768$329.$result[0] ),
    .Q(\fpga_top.qspi_if.inner_state[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _24296_ (.RESET_B(net5950),
    .D(net1808),
    .Q(\fpga_top.qspi_if.inner_state[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _24297_ (.RESET_B(net6006),
    .D(_00989_),
    .Q(\fpga_top.qspi_if.adr_rw[0] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _24298_ (.RESET_B(net6006),
    .D(_00990_),
    .Q(\fpga_top.qspi_if.adr_rw[1] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _24299_ (.RESET_B(net5999),
    .D(net6296),
    .Q(\fpga_top.qspi_if.adr_rw[2] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _24300_ (.RESET_B(net5998),
    .D(net6249),
    .Q(\fpga_top.qspi_if.adr_rw[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24301_ (.RESET_B(net5998),
    .D(net6278),
    .Q(\fpga_top.qspi_if.adr_rw[4] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _24302_ (.RESET_B(net5997),
    .D(net6454),
    .Q(\fpga_top.qspi_if.adr_rw[5] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _24303_ (.RESET_B(net5997),
    .D(_00995_),
    .Q(\fpga_top.qspi_if.adr_rw[6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _24304_ (.RESET_B(net5997),
    .D(net6268),
    .Q(\fpga_top.qspi_if.adr_rw[7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _24305_ (.RESET_B(net5998),
    .D(_00997_),
    .Q(\fpga_top.qspi_if.adr_rw[8] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _24306_ (.RESET_B(net5997),
    .D(net6254),
    .Q(\fpga_top.qspi_if.adr_rw[9] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _24307_ (.RESET_B(net5920),
    .D(_00999_),
    .Q(\fpga_top.qspi_if.adr_rw[10] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _24308_ (.RESET_B(net5973),
    .D(_01000_),
    .Q(\fpga_top.qspi_if.adr_rw[11] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _24309_ (.RESET_B(net5973),
    .D(net3174),
    .Q(\fpga_top.qspi_if.adr_rw[12] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _24310_ (.RESET_B(net5973),
    .D(net6131),
    .Q(\fpga_top.qspi_if.adr_rw[13] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _24311_ (.RESET_B(net5974),
    .D(net6272),
    .Q(\fpga_top.qspi_if.adr_rw[14] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _24312_ (.RESET_B(net5974),
    .D(_01004_),
    .Q(\fpga_top.qspi_if.adr_rw[15] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _24313_ (.RESET_B(net5974),
    .D(_01005_),
    .Q(\fpga_top.qspi_if.adr_rw[16] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _24314_ (.RESET_B(net5974),
    .D(_01006_),
    .Q(\fpga_top.qspi_if.adr_rw[17] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_1 _24315_ (.RESET_B(net5998),
    .D(_01007_),
    .Q(\fpga_top.qspi_if.adr_rw[18] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _24316_ (.RESET_B(net5974),
    .D(_01008_),
    .Q(\fpga_top.qspi_if.adr_rw[19] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _24317_ (.RESET_B(net5974),
    .D(net6398),
    .Q(\fpga_top.qspi_if.adr_rw[20] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _24318_ (.RESET_B(net5975),
    .D(net6502),
    .Q(\fpga_top.qspi_if.adr_rw[21] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _24319_ (.RESET_B(net5973),
    .D(_01011_),
    .Q(\fpga_top.qspi_if.adr_rw[22] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _24320_ (.RESET_B(net5971),
    .D(_01012_),
    .Q(\fpga_top.qspi_if.adr_rw[23] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _24321_ (.RESET_B(net5973),
    .D(_01013_),
    .Q(\fpga_top.qspi_if.word_adr[24] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _24322_ (.RESET_B(net5973),
    .D(_01014_),
    .Q(\fpga_top.qspi_if.word_adr[25] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _24323_ (.RESET_B(net5854),
    .D(_00130_),
    .Q(_00088_),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _24324_ (.RESET_B(net5938),
    .D(_01015_),
    .Q(\fpga_top.qspi_if.read_cntr[0] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24325_ (.RESET_B(net5939),
    .D(net3912),
    .Q(\fpga_top.qspi_if.read_cntr[1] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24326_ (.RESET_B(net5938),
    .D(_01017_),
    .Q(\fpga_top.qspi_if.read_cntr[2] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24327_ (.RESET_B(net5940),
    .D(net1490),
    .Q(\fpga_top.qspi_if.read_cntr[3] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _24328_ (.RESET_B(net5881),
    .D(\fpga_top.qspi_if.re_qspi_latency0 ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _24329_ (.RESET_B(net5881),
    .D(\fpga_top.qspi_if.re_qspi_latency1 ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _24330_ (.RESET_B(net5855),
    .D(\fpga_top.qspi_if.re_qspi_latency2 ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _24331_ (.RESET_B(net5898),
    .D(\fpga_top.qspi_if.re_qspi_sckdiv ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _24332_ (.RESET_B(net5855),
    .D(\fpga_top.qspi_if.re_qspi_rdcmd0 ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _24333_ (.RESET_B(net5855),
    .D(\fpga_top.qspi_if.re_qspi_rdcmd1 ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24334_ (.RESET_B(net5855),
    .D(\fpga_top.qspi_if.re_qspi_wrcmd0 ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _24335_ (.RESET_B(net5855),
    .D(\fpga_top.qspi_if.re_qspi_wrcmd1 ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[7] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _24336_ (.RESET_B(net5855),
    .D(\fpga_top.qspi_if.re_qspi_rdwrch ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _24337_ (.RESET_B(net5855),
    .D(\fpga_top.qspi_if.re_qspi_rdedge ),
    .Q(\fpga_top.qspi_if.re_qspi_latency_dly[9] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _24338_ (.RESET_B(net5872),
    .D(_01019_),
    .Q(\fpga_top.qspi_if.rwait_cntr[0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _24339_ (.RESET_B(net5839),
    .D(_01020_),
    .Q(\fpga_top.qspi_if.rwait_cntr[1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _24340_ (.RESET_B(net5872),
    .D(_01021_),
    .Q(\fpga_top.qspi_if.rwait_cntr[2] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _24341_ (.RESET_B(net5848),
    .D(net2399),
    .Q(\fpga_top.qspi_if.rwait_cntr[3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _24342_ (.RESET_B(net5854),
    .D(_00131_),
    .Q(_00089_),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _24343_ (.RESET_B(net5855),
    .D(_01023_),
    .Q(\fpga_top.qspi_if.rdedge[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _24344_ (.RESET_B(net5854),
    .D(_01024_),
    .Q(_00090_),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _24345_ (.RESET_B(net5854),
    .D(_01025_),
    .Q(\fpga_top.qspi_if.rdedge[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _24346_ (.RESET_B(net5866),
    .D(net6263),
    .Q(_00091_),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _24347_ (.RESET_B(net5868),
    .D(_00133_),
    .Q(_00092_),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _24348_ (.RESET_B(net5870),
    .D(_00134_),
    .Q(_00093_),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _24349_ (.RESET_B(net5849),
    .D(_01026_),
    .Q(\fpga_top.qspi_if.wredge[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24350_ (.RESET_B(net5854),
    .D(_01027_),
    .Q(_00094_),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24351_ (.RESET_B(net5881),
    .D(_01028_),
    .Q(\fpga_top.qspi_if.wredge[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _24352_ (.RESET_B(net5847),
    .D(_01029_),
    .Q(\fpga_top.qspi_if.rdwrch[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _24353_ (.RESET_B(net5849),
    .D(_01030_),
    .Q(\fpga_top.qspi_if.rdwrch[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24354_ (.RESET_B(net5850),
    .D(_01031_),
    .Q(\fpga_top.qspi_if.rdwrch[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24355_ (.RESET_B(net5848),
    .D(_01032_),
    .Q(\fpga_top.qspi_if.rdwrch[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _24356_ (.RESET_B(net5851),
    .D(_01033_),
    .Q(\fpga_top.qspi_if.rdwrch[4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24357_ (.RESET_B(net5851),
    .D(_01034_),
    .Q(\fpga_top.qspi_if.rdwrch[5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _24358_ (.RESET_B(net5854),
    .D(_00135_),
    .Q(_00095_),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _24359_ (.RESET_B(net5853),
    .D(_01035_),
    .Q(\fpga_top.qspi_if.wrcmd1[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24360_ (.RESET_B(net5844),
    .D(_01036_),
    .Q(\fpga_top.qspi_if.wrcmd1[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _24361_ (.RESET_B(net5852),
    .D(_01037_),
    .Q(\fpga_top.qspi_if.wrcmd1[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _24362_ (.RESET_B(net5853),
    .D(_01038_),
    .Q(_00096_),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _24363_ (.RESET_B(net5844),
    .D(_01039_),
    .Q(_00097_),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _24364_ (.RESET_B(net5851),
    .D(_01040_),
    .Q(_00098_),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _24365_ (.RESET_B(net5845),
    .D(_01041_),
    .Q(\fpga_top.qspi_if.wrcmd1[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _24366_ (.RESET_B(net5845),
    .D(_01042_),
    .Q(\fpga_top.qspi_if.wrcmd1[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _24367_ (.RESET_B(net5952),
    .D(_01043_),
    .Q(\fpga_top.qspi_if.wdata_ofs[0] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24368_ (.RESET_B(net5952),
    .D(_01044_),
    .Q(\fpga_top.qspi_if.wdata_ofs[1] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24369_ (.RESET_B(net5952),
    .D(_01045_),
    .Q(\fpga_top.qspi_if.wdata_ofs[2] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24370_ (.RESET_B(net5844),
    .D(_01046_),
    .Q(\fpga_top.qspi_if.wrcmd0[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _24371_ (.RESET_B(net5844),
    .D(_01047_),
    .Q(\fpga_top.qspi_if.wrcmd0[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _24372_ (.RESET_B(net5852),
    .D(_01048_),
    .Q(\fpga_top.qspi_if.wrcmd0[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _24373_ (.RESET_B(net5853),
    .D(_01049_),
    .Q(_00099_),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _24374_ (.RESET_B(net5846),
    .D(_01050_),
    .Q(_00100_),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _24375_ (.RESET_B(net5851),
    .D(_01051_),
    .Q(_00101_),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _24376_ (.RESET_B(net5845),
    .D(_01052_),
    .Q(\fpga_top.qspi_if.wrcmd0[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _24377_ (.RESET_B(net5845),
    .D(_01053_),
    .Q(\fpga_top.qspi_if.wrcmd0[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _24378_ (.RESET_B(net5852),
    .D(_01054_),
    .Q(_00102_),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _24379_ (.RESET_B(net5852),
    .D(_01055_),
    .Q(_00103_),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _24380_ (.RESET_B(net5845),
    .D(_01056_),
    .Q(\fpga_top.qspi_if.rdcmd1[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _24381_ (.RESET_B(net5844),
    .D(_01057_),
    .Q(_00104_),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _24382_ (.RESET_B(net5845),
    .D(_01058_),
    .Q(\fpga_top.qspi_if.rdcmd1[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _24383_ (.RESET_B(net5851),
    .D(_01059_),
    .Q(_00105_),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _24384_ (.RESET_B(net5851),
    .D(_01060_),
    .Q(_00106_),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _24385_ (.RESET_B(net5851),
    .D(_01061_),
    .Q(\fpga_top.qspi_if.rdcmd1[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _24386_ (.RESET_B(net5849),
    .D(_00136_),
    .Q(_00107_),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _24387_ (.RESET_B(net5852),
    .D(_01062_),
    .Q(_00108_),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _24388_ (.RESET_B(net5852),
    .D(_01063_),
    .Q(_00109_),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _24389_ (.RESET_B(net5850),
    .D(_01064_),
    .Q(\fpga_top.qspi_if.rdcmd0[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _24390_ (.RESET_B(net5844),
    .D(_01065_),
    .Q(_00110_),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _24391_ (.RESET_B(net5845),
    .D(_01066_),
    .Q(\fpga_top.qspi_if.rdcmd0[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _24392_ (.RESET_B(net5851),
    .D(_01067_),
    .Q(_00111_),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _24393_ (.RESET_B(net5850),
    .D(_01068_),
    .Q(_00112_),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _24394_ (.RESET_B(net5847),
    .D(_01069_),
    .Q(_00113_),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _24395_ (.RESET_B(net5915),
    .D(_01070_),
    .Q(\fpga_top.qspi_if.dbg_2div_wirte_half_end ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _24396_ (.RESET_B(net5901),
    .D(_01071_),
    .Q(\fpga_top.qspi_if.dbg_2div_read_half_end ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _24397_ (.RESET_B(net5901),
    .D(_01072_),
    .Q(\fpga_top.qspi_if.dbg_reg_2div_cec_write ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _24398_ (.RESET_B(net5900),
    .D(_01073_),
    .Q(\fpga_top.qspi_if.dbg_reg_2div_cec_read ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _24399_ (.RESET_B(net5896),
    .D(_01074_),
    .Q(\fpga_top.qspi_if.dbg_2div_trt ),
    .CLK(clknet_leaf_319_clk));
 sg13g2_dfrbpq_1 _24400_ (.RESET_B(net5902),
    .D(_01075_),
    .Q(\fpga_top.dbg_bpoint_en[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _24401_ (.RESET_B(net5917),
    .D(_01076_),
    .Q(\fpga_top.dbg_bpoint_en[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _24402_ (.RESET_B(net5902),
    .D(_01077_),
    .Q(\fpga_top.dbg_bpoint_en[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _24403_ (.RESET_B(net5847),
    .D(_01078_),
    .Q(_00114_),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _24404_ (.RESET_B(net5847),
    .D(_01079_),
    .Q(\fpga_top.qspi_if.sck_div[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _24405_ (.RESET_B(net5842),
    .D(_01080_),
    .Q(\fpga_top.qspi_if.sck_div[2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _24406_ (.RESET_B(net5847),
    .D(_01081_),
    .Q(\fpga_top.qspi_if.sck_div[3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _24407_ (.RESET_B(net5841),
    .D(_01082_),
    .Q(\fpga_top.qspi_if.sck_div[4] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _24408_ (.RESET_B(net5840),
    .D(_01083_),
    .Q(\fpga_top.qspi_if.sck_div[5] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _24409_ (.RESET_B(net5840),
    .D(_01084_),
    .Q(\fpga_top.qspi_if.sck_div[6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _24410_ (.RESET_B(net5840),
    .D(_01085_),
    .Q(\fpga_top.qspi_if.sck_div[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _24411_ (.RESET_B(net5890),
    .D(_01086_),
    .Q(\fpga_top.qspi_if.sck_div[8] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _24412_ (.RESET_B(net5888),
    .D(_01087_),
    .Q(\fpga_top.qspi_if.sck_div[9] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _24413_ (.RESET_B(net5849),
    .D(_00137_),
    .Q(_00115_),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _24414_ (.RESET_B(net5873),
    .D(_01088_),
    .Q(\fpga_top.qspi_if.read_latency_2[0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _24415_ (.RESET_B(net5849),
    .D(_01089_),
    .Q(\fpga_top.qspi_if.read_latency_2[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _24416_ (.RESET_B(net5848),
    .D(_01090_),
    .Q(\fpga_top.qspi_if.read_latency_2[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _24417_ (.RESET_B(net5848),
    .D(_01091_),
    .Q(\fpga_top.qspi_if.read_latency_2[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _24418_ (.RESET_B(net5873),
    .D(_01092_),
    .Q(\fpga_top.qspi_if.read_latency_1[0] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _24419_ (.RESET_B(net5873),
    .D(_01093_),
    .Q(\fpga_top.qspi_if.read_latency_1[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _24420_ (.RESET_B(net5848),
    .D(_01094_),
    .Q(\fpga_top.qspi_if.read_latency_1[2] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _24421_ (.RESET_B(net5848),
    .D(_01095_),
    .Q(\fpga_top.qspi_if.read_latency_1[3] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _24422_ (.RESET_B(net5872),
    .D(_01096_),
    .Q(\fpga_top.qspi_if.read_latency_0[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _24423_ (.RESET_B(net5873),
    .D(_01097_),
    .Q(\fpga_top.qspi_if.read_latency_0[1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _24424_ (.RESET_B(net5848),
    .D(_01098_),
    .Q(\fpga_top.qspi_if.read_latency_0[2] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _24425_ (.RESET_B(net5848),
    .D(_01099_),
    .Q(\fpga_top.qspi_if.read_latency_0[3] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _24426_ (.RESET_B(net5947),
    .D(net6465),
    .Q(\fpga_top.qspi_if.adr_ofs[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _24427_ (.RESET_B(net5947),
    .D(net6159),
    .Q(\fpga_top.qspi_if.adr_ofs[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _24428_ (.RESET_B(net5947),
    .D(_01102_),
    .Q(\fpga_top.qspi_if.adr_ofs[2] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _24429_ (.RESET_B(net5905),
    .D(_01103_),
    .Q(\fpga_top.qspi_if.rst_cntr[0] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _24430_ (.RESET_B(net5905),
    .D(net3526),
    .Q(\fpga_top.qspi_if.rst_cntr[1] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _24431_ (.RESET_B(net5905),
    .D(net3789),
    .Q(\fpga_top.qspi_if.rst_cntr[2] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _24432_ (.RESET_B(net5905),
    .D(_01106_),
    .Q(\fpga_top.qspi_if.rst_cntr[3] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _24433_ (.RESET_B(net5866),
    .D(net1321),
    .Q(\fpga_top.qspi_if.sio_en ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _24434_ (.RESET_B(net5938),
    .D(\fpga_top.qspi_if.dbg_2div_cec_pre ),
    .Q(\fpga_top.qspi_if.dbg_2div_cec_lat ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _24435_ (.RESET_B(net5864),
    .D(net1317),
    .Q(uio_out[0]),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24436_ (.RESET_B(net5865),
    .D(net1325),
    .Q(uio_out[1]),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24437_ (.RESET_B(net5864),
    .D(net1335),
    .Q(uio_out[2]),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _24438_ (.RESET_B(net5864),
    .D(net1331),
    .Q(uio_out[3]),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _24439_ (.RESET_B(net623),
    .D(net1370),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.radr[0] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _24440_ (.RESET_B(net624),
    .D(net1367),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.radr[1] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _24441_ (.RESET_B(net625),
    .D(net1364),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.radr[2] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _24442_ (.RESET_B(net5879),
    .D(_00052_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _24443_ (.RESET_B(net5879),
    .D(_00059_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _24444_ (.RESET_B(net5884),
    .D(_00060_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[2] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _24445_ (.RESET_B(net5879),
    .D(net3974),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[3] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _24446_ (.RESET_B(net5878),
    .D(_00062_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[4] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _24447_ (.RESET_B(net5878),
    .D(_00063_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[5] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _24448_ (.RESET_B(net5879),
    .D(_00064_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[6] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _24449_ (.RESET_B(net5878),
    .D(_00065_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[7] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _24450_ (.RESET_B(net5926),
    .D(net3997),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[8] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _24451_ (.RESET_B(net5926),
    .D(_00067_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[9] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _24452_ (.RESET_B(net5926),
    .D(net6209),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[10] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _24453_ (.RESET_B(net5926),
    .D(net6176),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[11] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _24454_ (.RESET_B(net5878),
    .D(_00055_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[12] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _24455_ (.RESET_B(net5878),
    .D(_00056_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[13] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _24456_ (.RESET_B(net5878),
    .D(net6148),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[14] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _24457_ (.RESET_B(net5878),
    .D(_00058_),
    .Q(\fpga_top.uart_top.uart_if.sample_cntr[15] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _24458_ (.RESET_B(net5936),
    .D(_00138_),
    .Q(_00116_),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _24459_ (.RESET_B(net5939),
    .D(net6190),
    .Q(\fpga_top.uart_top.uart_if.rx_state[0] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _24460_ (.RESET_B(net5939),
    .D(\fpga_top.uart_top.uart_if.next_rx_state[1] ),
    .Q(\fpga_top.uart_top.uart_if.rx_state[1] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _24461_ (.RESET_B(net5939),
    .D(\fpga_top.uart_top.uart_if.next_rx_state[2] ),
    .Q(\fpga_top.uart_top.uart_if.rx_state[2] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _24462_ (.RESET_B(net5939),
    .D(net1603),
    .Q(\fpga_top.uart_top.uart_if.rx_state[3] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _24463_ (.RESET_B(net5940),
    .D(_00139_),
    .Q(_00117_),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _24464_ (.RESET_B(net5868),
    .D(_01107_),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[0] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _24465_ (.RESET_B(net5882),
    .D(_01108_),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[1] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24466_ (.RESET_B(net5882),
    .D(_01109_),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[2] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _24467_ (.RESET_B(net5869),
    .D(_01110_),
    .Q(\fpga_top.uart_top.rx_fifo_rcntr[0] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _24468_ (.RESET_B(net5869),
    .D(_01111_),
    .Q(\fpga_top.uart_top.rx_fifo_rcntr[1] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _24469_ (.RESET_B(net5869),
    .D(_01112_),
    .Q(\fpga_top.uart_top.rx_fifo_rcntr[2] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _24470_ (.RESET_B(net5865),
    .D(_01113_),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[0] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _24471_ (.RESET_B(net5865),
    .D(_01114_),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[1] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _24472_ (.RESET_B(net5865),
    .D(_01115_),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[2] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _24473_ (.RESET_B(net5865),
    .D(net1898),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[3] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _24474_ (.RESET_B(net5951),
    .D(_00140_),
    .Q(_00118_),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _24475_ (.RESET_B(net5867),
    .D(_01117_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[0] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _24476_ (.RESET_B(net5867),
    .D(_01118_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[1] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _24477_ (.RESET_B(net5867),
    .D(_01119_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[2] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _24478_ (.RESET_B(net5859),
    .D(_01120_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram_radr[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _24479_ (.RESET_B(net5859),
    .D(_01121_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram_radr[1] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _24480_ (.RESET_B(net5859),
    .D(_01122_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram_radr[2] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _24481_ (.RESET_B(net5936),
    .D(_00141_),
    .Q(_00119_),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _24482_ (.RESET_B(net5839),
    .D(net1537),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24483_ (.RESET_B(net5839),
    .D(_01124_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _24484_ (.RESET_B(net5839),
    .D(net3387),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[2] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _24485_ (.RESET_B(net5859),
    .D(_01126_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[3] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _24486_ (.RESET_B(net5951),
    .D(_00142_),
    .Q(_00120_),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _24487_ (.RESET_B(net5859),
    .D(_01127_),
    .Q(\fpga_top.uart_top.uart_if.tx_out_cntr[0] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _24488_ (.RESET_B(net5867),
    .D(_01128_),
    .Q(\fpga_top.uart_top.uart_if.tx_out_cntr[1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _24489_ (.RESET_B(net5867),
    .D(net3732),
    .Q(\fpga_top.uart_top.uart_if.tx_out_cntr[2] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _24490_ (.RESET_B(net5867),
    .D(net3445),
    .Q(\fpga_top.uart_top.uart_if.tx_out_cntr[3] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _24491_ (.RESET_B(net5859),
    .D(net1386),
    .Q(_00121_),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _24492_ (.RESET_B(net5859),
    .D(net1632),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _24493_ (.RESET_B(net5860),
    .D(_01133_),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[2] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _24494_ (.RESET_B(net5860),
    .D(net1492),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[3] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _24495_ (.RESET_B(net5860),
    .D(net1957),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[4] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _24496_ (.RESET_B(net5860),
    .D(net1515),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[5] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _24497_ (.RESET_B(net5860),
    .D(net1577),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[6] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _24498_ (.RESET_B(net5860),
    .D(net1412),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[7] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _24499_ (.RESET_B(net5859),
    .D(net1605),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[8] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _24500_ (.RESET_B(net5862),
    .D(_01140_),
    .Q(\fpga_top.uart_top.uart_if.tx_out_data[9] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _24501_ (.RESET_B(net5875),
    .D(net1903),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[0] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _24502_ (.RESET_B(net5875),
    .D(net1974),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[1] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _24503_ (.RESET_B(net5875),
    .D(net2124),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[2] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _24504_ (.RESET_B(net5875),
    .D(net2114),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[3] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _24505_ (.RESET_B(net5875),
    .D(_00078_),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[4] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _24506_ (.RESET_B(net5876),
    .D(net2374),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[5] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _24507_ (.RESET_B(net5876),
    .D(net3143),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[6] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _24508_ (.RESET_B(net5876),
    .D(net3607),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[7] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _24509_ (.RESET_B(net5873),
    .D(net3966),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[8] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _24510_ (.RESET_B(net5872),
    .D(net3306),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[9] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _24511_ (.RESET_B(net5872),
    .D(net3989),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[10] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _24512_ (.RESET_B(net5872),
    .D(net6168),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[11] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _24513_ (.RESET_B(net5873),
    .D(net4023),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[12] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24514_ (.RESET_B(net5873),
    .D(net4044),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[13] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24515_ (.RESET_B(net5873),
    .D(net6112),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[14] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24516_ (.RESET_B(net5881),
    .D(net1936),
    .Q(\fpga_top.uart_top.uart_if.tx_cycle_cntr[15] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _24517_ (.RESET_B(net5950),
    .D(_00143_),
    .Q(_00122_),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _24518_ (.RESET_B(net5863),
    .D(\fpga_top.uart_top.uart_if.next_tx_state[0] ),
    .Q(\fpga_top.uart_top.uart_if.tx_state[0] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _24519_ (.RESET_B(net5863),
    .D(\fpga_top.uart_top.uart_if.next_tx_state[1] ),
    .Q(\fpga_top.uart_top.uart_if.tx_state[1] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _24520_ (.RESET_B(net5849),
    .D(_01141_),
    .Q(_00123_),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _24521_ (.RESET_B(net6033),
    .D(_01142_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[0] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_1 _24522_ (.RESET_B(net5980),
    .D(_01143_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[1] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _24523_ (.RESET_B(net6032),
    .D(_01144_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[2] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_1 _24524_ (.RESET_B(net5982),
    .D(_01145_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[3] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _24525_ (.RESET_B(net5979),
    .D(_01146_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[6] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _24526_ (.RESET_B(net5981),
    .D(net1624),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[7] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_1 _24527_ (.RESET_B(net5984),
    .D(_01148_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[8] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _24528_ (.RESET_B(net6036),
    .D(_01149_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[9] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _24529_ (.RESET_B(net6050),
    .D(_01150_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[10] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _24530_ (.RESET_B(net5981),
    .D(net1787),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[11] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_1 _24531_ (.RESET_B(net5984),
    .D(net1797),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[12] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_1 _24532_ (.RESET_B(net6036),
    .D(_01153_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[13] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _24533_ (.RESET_B(net6036),
    .D(_01154_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[14] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _24534_ (.RESET_B(net6037),
    .D(_01155_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[15] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _24535_ (.RESET_B(net6039),
    .D(_01156_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[16] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _24536_ (.RESET_B(net6050),
    .D(_01157_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[17] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _24537_ (.RESET_B(net6048),
    .D(_01158_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[18] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_1 _24538_ (.RESET_B(net6051),
    .D(_01159_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[19] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _24539_ (.RESET_B(net6046),
    .D(_01160_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[20] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _24540_ (.RESET_B(net6054),
    .D(_01161_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[21] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _24541_ (.RESET_B(net6045),
    .D(_01162_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[22] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _24542_ (.RESET_B(net6055),
    .D(net1984),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[23] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _24543_ (.RESET_B(net6047),
    .D(_01164_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[24] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _24544_ (.RESET_B(net6047),
    .D(_01165_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[25] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_1 _24545_ (.RESET_B(net6051),
    .D(_01166_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[26] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _24546_ (.RESET_B(net6053),
    .D(_01167_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[27] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_1 _24547_ (.RESET_B(net6050),
    .D(_01168_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[28] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _24548_ (.RESET_B(net6052),
    .D(_01169_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[29] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _24549_ (.RESET_B(net6045),
    .D(_01170_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[30] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _24550_ (.RESET_B(net6032),
    .D(_01171_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[31] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _24551_ (.RESET_B(net5951),
    .D(_00144_),
    .Q(_00124_),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _24552_ (.RESET_B(net47),
    .D(_01172_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][0] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _24553_ (.RESET_B(net46),
    .D(_01173_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][1] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _24554_ (.RESET_B(net45),
    .D(_01174_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][2] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _24555_ (.RESET_B(net44),
    .D(_01175_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][3] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _24556_ (.RESET_B(net43),
    .D(_01176_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][4] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _24557_ (.RESET_B(net42),
    .D(_01177_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _24558_ (.RESET_B(net41),
    .D(_01178_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][6] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_1 _24559_ (.RESET_B(net40),
    .D(_01179_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][7] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _24560_ (.RESET_B(net39),
    .D(_01180_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][8] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _24561_ (.RESET_B(net38),
    .D(_01181_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][9] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _24562_ (.RESET_B(net37),
    .D(_01182_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _24563_ (.RESET_B(net36),
    .D(_01183_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][11] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _24564_ (.RESET_B(net35),
    .D(_01184_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][12] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _24565_ (.RESET_B(net34),
    .D(_01185_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][13] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _24566_ (.RESET_B(net33),
    .D(_01186_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][14] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _24567_ (.RESET_B(net32),
    .D(_01187_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][15] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _24568_ (.RESET_B(net31),
    .D(_01188_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][16] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _24569_ (.RESET_B(net30),
    .D(_01189_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][17] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _24570_ (.RESET_B(net29),
    .D(_01190_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][18] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _24571_ (.RESET_B(net28),
    .D(_01191_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _24572_ (.RESET_B(net27),
    .D(_01192_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _24573_ (.RESET_B(net26),
    .D(_01193_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][21] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _24574_ (.RESET_B(net25),
    .D(_01194_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][22] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _24575_ (.RESET_B(net24),
    .D(_01195_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][23] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _24576_ (.RESET_B(net23),
    .D(_01196_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][24] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _24577_ (.RESET_B(net22),
    .D(_01197_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _24578_ (.RESET_B(net21),
    .D(_01198_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][26] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _24579_ (.RESET_B(net20),
    .D(_01199_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][27] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _24580_ (.RESET_B(net19),
    .D(_01200_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][28] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _24581_ (.RESET_B(net18),
    .D(_01201_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][29] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _24582_ (.RESET_B(net17),
    .D(_01202_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][30] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _24583_ (.RESET_B(net699),
    .D(_01203_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][31] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _24584_ (.RESET_B(net5869),
    .D(\fpga_top.uart_top.rx_fifo_dvalid ),
    .Q(\fpga_top.io_uart_out.rout_en ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _24585_ (.RESET_B(net5946),
    .D(net6576),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _24586_ (.RESET_B(net5946),
    .D(net6403),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _24587_ (.RESET_B(net5946),
    .D(net6435),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[2] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _24588_ (.RESET_B(net5949),
    .D(_01207_),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[3] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _24589_ (.RESET_B(net5949),
    .D(net6371),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[4] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _24590_ (.RESET_B(net5920),
    .D(_01209_),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[5] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _24591_ (.RESET_B(net5920),
    .D(_01210_),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[6] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _24592_ (.RESET_B(net5919),
    .D(_01211_),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _24593_ (.RESET_B(net5919),
    .D(_01212_),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _24594_ (.RESET_B(net5919),
    .D(_01213_),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[9] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _24595_ (.RESET_B(net5919),
    .D(net4037),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[10] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _24596_ (.RESET_B(net5919),
    .D(_01215_),
    .Q(\fpga_top.cpu_top.csr_wadr_mon[11] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _24597_ (.RESET_B(net5919),
    .D(net6275),
    .Q(\fpga_top.dma_io_wadr_u[14] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _24598_ (.RESET_B(net5919),
    .D(net6367),
    .Q(\fpga_top.dma_io_wadr_u[15] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _24599_ (.RESET_B(net5971),
    .D(net6152),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[16] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _24600_ (.RESET_B(net5972),
    .D(net6170),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[17] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _24601_ (.RESET_B(net5971),
    .D(net6096),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[18] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _24602_ (.RESET_B(net5971),
    .D(net6142),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[19] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _24603_ (.RESET_B(net5971),
    .D(_01222_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[20] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _24604_ (.RESET_B(net5971),
    .D(net6116),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[21] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _24605_ (.RESET_B(net5971),
    .D(net6110),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[22] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _24606_ (.RESET_B(net5971),
    .D(net6083),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[23] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _24607_ (.RESET_B(net5963),
    .D(net6164),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[24] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_2 _24608_ (.RESET_B(net5963),
    .D(_01227_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[25] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _24609_ (.RESET_B(net5963),
    .D(net4050),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[26] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _24610_ (.RESET_B(net5963),
    .D(net4008),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[27] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _24611_ (.RESET_B(net5913),
    .D(_01230_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[28] ),
    .CLK(clknet_leaf_318_clk));
 sg13g2_dfrbpq_1 _24612_ (.RESET_B(net5963),
    .D(net6079),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[29] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_1 _24613_ (.RESET_B(net5972),
    .D(net3982),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[30] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _24614_ (.RESET_B(net5972),
    .D(_01233_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[31] ),
    .CLK(clknet_leaf_295_clk));
 sg13g2_dfrbpq_2 _24615_ (.RESET_B(net5953),
    .D(_01234_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint_ld ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24616_ (.RESET_B(net5911),
    .D(_01235_),
    .Q(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _24617_ (.RESET_B(net5912),
    .D(net6487),
    .Q(\fpga_top.cpu_top.csr_wdata_mon[1] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _24618_ (.RESET_B(net5912),
    .D(_01237_),
    .Q(\fpga_top.cpu_start_adr[2] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_2 _24619_ (.RESET_B(net5912),
    .D(_01238_),
    .Q(\fpga_top.cpu_start_adr[3] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _24620_ (.RESET_B(net5911),
    .D(net3799),
    .Q(\fpga_top.cpu_start_adr[4] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _24621_ (.RESET_B(net5911),
    .D(_01240_),
    .Q(\fpga_top.cpu_start_adr[5] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _24622_ (.RESET_B(net5968),
    .D(net1856),
    .Q(\fpga_top.cpu_start_adr[6] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _24623_ (.RESET_B(net5968),
    .D(_01242_),
    .Q(\fpga_top.cpu_start_adr[7] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_2 _24624_ (.RESET_B(net5910),
    .D(_01243_),
    .Q(\fpga_top.cpu_start_adr[8] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_2 _24625_ (.RESET_B(net5910),
    .D(_01244_),
    .Q(\fpga_top.cpu_start_adr[9] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _24626_ (.RESET_B(net5963),
    .D(_01245_),
    .Q(\fpga_top.cpu_start_adr[10] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_2 _24627_ (.RESET_B(net5964),
    .D(_01246_),
    .Q(\fpga_top.cpu_start_adr[11] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_2 _24628_ (.RESET_B(net5909),
    .D(_01247_),
    .Q(\fpga_top.cpu_start_adr[12] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _24629_ (.RESET_B(net5909),
    .D(_01248_),
    .Q(\fpga_top.cpu_start_adr[13] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_2 _24630_ (.RESET_B(net5961),
    .D(net2015),
    .Q(\fpga_top.cpu_start_adr[14] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_2 _24631_ (.RESET_B(net5961),
    .D(_01250_),
    .Q(\fpga_top.cpu_start_adr[15] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_2 _24632_ (.RESET_B(net5909),
    .D(_01251_),
    .Q(\fpga_top.cpu_start_adr[16] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _24633_ (.RESET_B(net5909),
    .D(_01252_),
    .Q(\fpga_top.cpu_start_adr[17] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24634_ (.RESET_B(net5969),
    .D(net1780),
    .Q(\fpga_top.cpu_start_adr[18] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_2 _24635_ (.RESET_B(net5961),
    .D(net1648),
    .Q(\fpga_top.cpu_start_adr[19] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_2 _24636_ (.RESET_B(net5910),
    .D(_01255_),
    .Q(\fpga_top.cpu_start_adr[20] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24637_ (.RESET_B(net5967),
    .D(_01256_),
    .Q(\fpga_top.cpu_start_adr[21] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_2 _24638_ (.RESET_B(net5966),
    .D(net1813),
    .Q(\fpga_top.cpu_start_adr[22] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_2 _24639_ (.RESET_B(net5966),
    .D(_01258_),
    .Q(\fpga_top.cpu_start_adr[23] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_2 _24640_ (.RESET_B(net5960),
    .D(net1836),
    .Q(\fpga_top.cpu_start_adr[24] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24641_ (.RESET_B(net5983),
    .D(net2118),
    .Q(\fpga_top.cpu_start_adr[25] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _24642_ (.RESET_B(net5969),
    .D(net1579),
    .Q(\fpga_top.cpu_start_adr[26] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_2 _24643_ (.RESET_B(net5983),
    .D(_01262_),
    .Q(\fpga_top.cpu_start_adr[27] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _24644_ (.RESET_B(net5960),
    .D(_01263_),
    .Q(\fpga_top.cpu_start_adr[28] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_2 _24645_ (.RESET_B(net5966),
    .D(_01264_),
    .Q(\fpga_top.cpu_start_adr[29] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_2 _24646_ (.RESET_B(net5966),
    .D(_01265_),
    .Q(\fpga_top.cpu_start_adr[30] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_2 _24647_ (.RESET_B(net5965),
    .D(_01266_),
    .Q(\fpga_top.cpu_start_adr[31] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_1 _24648_ (.RESET_B(net5955),
    .D(\fpga_top.uart_top.uart_rec_char.word_valid_pre ),
    .Q(\fpga_top.uart_top.uart_rec_char.word_valid ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _24649_ (.RESET_B(net5955),
    .D(\fpga_top.uart_top.uart_rec_char.next_cmd_status[0] ),
    .Q(\fpga_top.uart_top.uart_rec_char.cmd_status[0] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _24650_ (.RESET_B(net5954),
    .D(\fpga_top.uart_top.uart_rec_char.next_cmd_status[1] ),
    .Q(\fpga_top.uart_top.uart_rec_char.cmd_status[1] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _24651_ (.RESET_B(net5954),
    .D(\fpga_top.uart_top.uart_rec_char.next_cmd_status[2] ),
    .Q(\fpga_top.uart_top.uart_rec_char.cmd_status[2] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _24652_ (.RESET_B(net5954),
    .D(\fpga_top.uart_top.uart_rec_char.next_cmd_status[3] ),
    .Q(\fpga_top.uart_top.uart_rec_char.cmd_status[3] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _24653_ (.RESET_B(net5954),
    .D(\fpga_top.uart_top.uart_rec_char.next_cmd_status[4] ),
    .Q(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _24654_ (.RESET_B(net6003),
    .D(net2070),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint_en ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _24655_ (.RESET_B(net5975),
    .D(_01268_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[2] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _24656_ (.RESET_B(net6001),
    .D(net1960),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _24657_ (.RESET_B(net6001),
    .D(net3960),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _24658_ (.RESET_B(net5991),
    .D(net4046),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[5] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _24659_ (.RESET_B(net5991),
    .D(net2100),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _24660_ (.RESET_B(net5975),
    .D(net1971),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[7] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _24661_ (.RESET_B(net5975),
    .D(net2769),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[8] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _24662_ (.RESET_B(net5975),
    .D(_01275_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[9] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_1 _24663_ (.RESET_B(net5991),
    .D(_01276_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[10] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _24664_ (.RESET_B(net5976),
    .D(_01277_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[11] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_2 _24665_ (.RESET_B(net5975),
    .D(_01278_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[12] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24666_ (.RESET_B(net5975),
    .D(_01279_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[13] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _24667_ (.RESET_B(net5989),
    .D(net2144),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[14] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _24668_ (.RESET_B(net5976),
    .D(_01281_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[15] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_1 _24669_ (.RESET_B(net5976),
    .D(net3352),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[16] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_2 _24670_ (.RESET_B(net5976),
    .D(_01283_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[17] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _24671_ (.RESET_B(net5976),
    .D(net2721),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[18] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_2 _24672_ (.RESET_B(net5989),
    .D(net2088),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[19] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24673_ (.RESET_B(net5991),
    .D(_01286_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[20] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _24674_ (.RESET_B(net5977),
    .D(_01287_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[21] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24675_ (.RESET_B(net5976),
    .D(net2876),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[22] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_1 _24676_ (.RESET_B(net5989),
    .D(net2994),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[23] ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _24677_ (.RESET_B(net5991),
    .D(net2009),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[24] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _24678_ (.RESET_B(net5977),
    .D(net2892),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[25] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_2 _24679_ (.RESET_B(net6001),
    .D(_01292_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[26] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _24680_ (.RESET_B(net5991),
    .D(_01293_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[27] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _24681_ (.RESET_B(net5975),
    .D(_01294_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[28] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _24682_ (.RESET_B(net5976),
    .D(_01295_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[29] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_1 _24683_ (.RESET_B(net5992),
    .D(_01296_),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[30] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_2 _24684_ (.RESET_B(net6001),
    .D(net1982),
    .Q(\fpga_top.uart_top.uart_rec_char.bpoint[31] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _24685_ (.RESET_B(net5950),
    .D(net5667),
    .Q(\fpga_top.uart_top.uart_rec_char.data_en ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _24686_ (.RESET_B(net6007),
    .D(net1329),
    .Q(\fpga_top.uart_top.uart_rec_char.g_crlf_dly2 ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _24687_ (.RESET_B(net6007),
    .D(net6469),
    .Q(\fpga_top.uart_top.uart_rec_char.g_crlf_dly ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _24688_ (.RESET_B(net6008),
    .D(_01298_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_cntr[0] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _24689_ (.RESET_B(net6008),
    .D(net2791),
    .Q(\fpga_top.uart_top.uart_rec_char.data_cntr[1] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _24690_ (.RESET_B(net6008),
    .D(net2142),
    .Q(\fpga_top.uart_top.uart_rec_char.data_cntr[2] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _24691_ (.RESET_B(net6008),
    .D(net1397),
    .Q(\fpga_top.uart_top.uart_rec_char.data_cntr[3] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _24692_ (.RESET_B(net6008),
    .D(net1326),
    .Q(\fpga_top.cpu_start ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _24693_ (.RESET_B(net5905),
    .D(_01302_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[0] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _24694_ (.RESET_B(net5911),
    .D(net1866),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[1] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _24695_ (.RESET_B(net5912),
    .D(_01304_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[2] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _24696_ (.RESET_B(net5909),
    .D(_01305_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[3] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_1 _24697_ (.RESET_B(net5911),
    .D(_01306_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[4] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _24698_ (.RESET_B(net5910),
    .D(_01307_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[5] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _24699_ (.RESET_B(net5962),
    .D(_01308_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[6] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _24700_ (.RESET_B(net5960),
    .D(_01309_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[7] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_1 _24701_ (.RESET_B(net5911),
    .D(_01310_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[8] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _24702_ (.RESET_B(net5910),
    .D(_01311_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[9] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_2 _24703_ (.RESET_B(net5960),
    .D(_01312_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[10] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _24704_ (.RESET_B(net5960),
    .D(_01313_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[11] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_2 _24705_ (.RESET_B(net5911),
    .D(_01314_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[12] ),
    .CLK(clknet_leaf_312_clk));
 sg13g2_dfrbpq_1 _24706_ (.RESET_B(net5910),
    .D(_01315_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[13] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _24707_ (.RESET_B(net5967),
    .D(_01316_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[14] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_1 _24708_ (.RESET_B(net5967),
    .D(_01317_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[15] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_1 _24709_ (.RESET_B(net5910),
    .D(_01318_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[16] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_2 _24710_ (.RESET_B(net5960),
    .D(_01319_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[17] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _24711_ (.RESET_B(net5965),
    .D(_01320_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[18] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_1 _24712_ (.RESET_B(net5967),
    .D(_01321_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[19] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_1 _24713_ (.RESET_B(net5962),
    .D(_01322_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[20] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _24714_ (.RESET_B(net5965),
    .D(_01323_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[21] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_1 _24715_ (.RESET_B(net5965),
    .D(_01324_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[22] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_1 _24716_ (.RESET_B(net5965),
    .D(_01325_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[23] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_1 _24717_ (.RESET_B(net5960),
    .D(_01326_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[24] ),
    .CLK(clknet_leaf_311_clk));
 sg13g2_dfrbpq_1 _24718_ (.RESET_B(net5965),
    .D(_01327_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[25] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_1 _24719_ (.RESET_B(net5965),
    .D(_01328_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[26] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_1 _24720_ (.RESET_B(net5965),
    .D(_01329_),
    .Q(\fpga_top.uart_top.uart_rec_char.data_word[27] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_1 _24721_ (.RESET_B(net5937),
    .D(net1401),
    .Q(_00125_),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _24722_ (.RESET_B(net5952),
    .D(net1535),
    .Q(\fpga_top.qspi_if.qspi_state[1] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _24723_ (.RESET_B(net5937),
    .D(_00017_),
    .Q(\fpga_top.qspi_if.qspi_state[2] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24724_ (.RESET_B(net5937),
    .D(net3900),
    .Q(\fpga_top.qspi_if.qspi_state[3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _24725_ (.RESET_B(net5952),
    .D(net3327),
    .Q(\fpga_top.qspi_if.qspi_state[4] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24726_ (.RESET_B(net5952),
    .D(_00020_),
    .Q(\fpga_top.qspi_if.dbg_2div_cew_pre ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _24727_ (.RESET_B(net5937),
    .D(net3977),
    .Q(\fpga_top.qspi_if.qspi_state[6] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _24728_ (.RESET_B(net5952),
    .D(_00022_),
    .Q(\fpga_top.qspi_if.qspi_state[7] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24729_ (.RESET_B(net5937),
    .D(net3763),
    .Q(\fpga_top.qspi_if.qspi_state[8] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _24730_ (.RESET_B(net5952),
    .D(_00014_),
    .Q(\fpga_top.qspi_if.qspi_state[10] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _24731_ (.RESET_B(net5937),
    .D(_00015_),
    .Q(\fpga_top.qspi_if.qspi_state[11] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _24732_ (.RESET_B(net5950),
    .D(net2726),
    .Q(\fpga_top.uart_top.uart_rec_char.pdata[0] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _24733_ (.RESET_B(net5939),
    .D(net3915),
    .Q(\fpga_top.uart_top.uart_rec_char.pdata[1] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _24734_ (.RESET_B(net5950),
    .D(net2854),
    .Q(\fpga_top.uart_top.uart_rec_char.pdata[2] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _24735_ (.RESET_B(net5936),
    .D(net3919),
    .Q(\fpga_top.uart_top.uart_rec_char.pdata[3] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _24736_ (.RESET_B(net5950),
    .D(net3625),
    .Q(\fpga_top.uart_top.uart_rec_char.pdata[4] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _24737_ (.RESET_B(net5939),
    .D(net3986),
    .Q(\fpga_top.uart_top.uart_rec_char.pdata[5] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _24738_ (.RESET_B(net5940),
    .D(net4021),
    .Q(\fpga_top.uart_top.uart_rec_char.pdata[6] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _24739_ (.RESET_B(net5939),
    .D(net4034),
    .Q(\fpga_top.uart_top.uart_rec_char.pdata[7] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _24740_ (.RESET_B(net6007),
    .D(net6460),
    .Q(\fpga_top.uart_top.uart_logics.status_dump[0] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _24741_ (.RESET_B(net6007),
    .D(net6526),
    .Q(\fpga_top.uart_top.uart_logics.status_dump[1] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _24742_ (.RESET_B(net6007),
    .D(\fpga_top.uart_top.uart_logics.next_status_dump[2] ),
    .Q(\fpga_top.uart_top.uart_logics.status_dump[2] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _24743_ (.RESET_B(net6002),
    .D(_01338_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _24744_ (.RESET_B(net6001),
    .D(net3028),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _24745_ (.RESET_B(net5999),
    .D(net3823),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[4] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _24746_ (.RESET_B(net5999),
    .D(net3139),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[5] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _24747_ (.RESET_B(net6001),
    .D(net2279),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _24748_ (.RESET_B(net5997),
    .D(net3538),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _24749_ (.RESET_B(net5920),
    .D(net1955),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[8] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _24750_ (.RESET_B(net5973),
    .D(net2760),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[9] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _24751_ (.RESET_B(net5972),
    .D(_01346_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[10] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _24752_ (.RESET_B(net5972),
    .D(_01347_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _24753_ (.RESET_B(net5919),
    .D(_01348_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[12] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _24754_ (.RESET_B(net5963),
    .D(_01349_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[13] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_1 _24755_ (.RESET_B(net5963),
    .D(net2560),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[14] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _24756_ (.RESET_B(net5964),
    .D(_01351_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[15] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_1 _24757_ (.RESET_B(net5969),
    .D(net1803),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[16] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _24758_ (.RESET_B(net5968),
    .D(_01353_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[17] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _24759_ (.RESET_B(net5968),
    .D(net2420),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[18] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_1 _24760_ (.RESET_B(net5968),
    .D(net1949),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[19] ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _24761_ (.RESET_B(net5967),
    .D(_01356_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[20] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24762_ (.RESET_B(net5967),
    .D(net3689),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[21] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24763_ (.RESET_B(net5967),
    .D(net1874),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[22] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24764_ (.RESET_B(net5960),
    .D(_01359_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[23] ),
    .CLK(clknet_leaf_309_clk));
 sg13g2_dfrbpq_1 _24765_ (.RESET_B(net5961),
    .D(net3434),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[24] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_1 _24766_ (.RESET_B(net5961),
    .D(net2269),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[25] ),
    .CLK(clknet_leaf_310_clk));
 sg13g2_dfrbpq_1 _24767_ (.RESET_B(net5909),
    .D(net2328),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[26] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_1 _24768_ (.RESET_B(net5911),
    .D(net3834),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[27] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_1 _24769_ (.RESET_B(net5912),
    .D(_01364_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[28] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_1 _24770_ (.RESET_B(net5912),
    .D(_01365_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[29] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_1 _24771_ (.RESET_B(net5946),
    .D(net1689),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[30] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _24772_ (.RESET_B(net5946),
    .D(_01367_),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_end[31] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _24773_ (.RESET_B(net6001),
    .D(net5285),
    .Q(\fpga_top.uart_top.uart_logics.dma_io_data_en ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _24774_ (.RESET_B(net6010),
    .D(_01368_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[0] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _24775_ (.RESET_B(net6010),
    .D(_01369_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[1] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _24776_ (.RESET_B(net6010),
    .D(_01370_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[2] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _24777_ (.RESET_B(net6014),
    .D(_01371_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[3] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24778_ (.RESET_B(net6010),
    .D(_01372_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[4] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _24779_ (.RESET_B(net6003),
    .D(_01373_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[5] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24780_ (.RESET_B(net6015),
    .D(_01374_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[6] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _24781_ (.RESET_B(net6002),
    .D(_01375_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[7] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24782_ (.RESET_B(net6010),
    .D(_01376_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[8] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _24783_ (.RESET_B(net6022),
    .D(_01377_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[9] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _24784_ (.RESET_B(net6014),
    .D(_01378_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[10] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24785_ (.RESET_B(net6014),
    .D(_01379_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[11] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _24786_ (.RESET_B(net6019),
    .D(_01380_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[12] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _24787_ (.RESET_B(net6019),
    .D(_01381_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[13] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _24788_ (.RESET_B(net6015),
    .D(_01382_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[14] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _24789_ (.RESET_B(net6015),
    .D(_01383_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[15] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24790_ (.RESET_B(net6002),
    .D(net1987),
    .Q(\fpga_top.uart_top.uart_logics.data_0[16] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _24791_ (.RESET_B(net6010),
    .D(_01385_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[17] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _24792_ (.RESET_B(net6002),
    .D(_01386_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[18] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _24793_ (.RESET_B(net6015),
    .D(_01387_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[19] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24794_ (.RESET_B(net6010),
    .D(net2563),
    .Q(\fpga_top.uart_top.uart_logics.data_0[20] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _24795_ (.RESET_B(net6019),
    .D(_01389_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[21] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _24796_ (.RESET_B(net6001),
    .D(net1969),
    .Q(\fpga_top.uart_top.uart_logics.data_0[22] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _24797_ (.RESET_B(net6003),
    .D(_01391_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[23] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24798_ (.RESET_B(net6010),
    .D(net2065),
    .Q(\fpga_top.uart_top.uart_logics.data_0[24] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _24799_ (.RESET_B(net6011),
    .D(net2553),
    .Q(\fpga_top.uart_top.uart_logics.data_0[25] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _24800_ (.RESET_B(net6002),
    .D(net2186),
    .Q(\fpga_top.uart_top.uart_logics.data_0[26] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _24801_ (.RESET_B(net6014),
    .D(_01395_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[27] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _24802_ (.RESET_B(net6019),
    .D(net2136),
    .Q(\fpga_top.uart_top.uart_logics.data_0[28] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _24803_ (.RESET_B(net6019),
    .D(_01397_),
    .Q(\fpga_top.uart_top.uart_logics.data_0[29] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _24804_ (.RESET_B(net6014),
    .D(net2083),
    .Q(\fpga_top.uart_top.uart_logics.data_0[30] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _24805_ (.RESET_B(net6002),
    .D(net3481),
    .Q(\fpga_top.uart_top.uart_logics.data_0[31] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _24806_ (.RESET_B(net5954),
    .D(net6380),
    .Q(\fpga_top.uart_top.trush_running ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _24807_ (.RESET_B(net6005),
    .D(_01401_),
    .Q(\fpga_top.bus_gather.u_read_adr[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _24808_ (.RESET_B(net6005),
    .D(net3852),
    .Q(\fpga_top.bus_gather.u_read_adr[3] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _24809_ (.RESET_B(net5999),
    .D(net6450),
    .Q(\fpga_top.bus_gather.u_read_adr[4] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _24810_ (.RESET_B(net5997),
    .D(_01404_),
    .Q(\fpga_top.bus_gather.u_read_adr[5] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _24811_ (.RESET_B(net5997),
    .D(net6316),
    .Q(\fpga_top.bus_gather.u_read_adr[6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _24812_ (.RESET_B(net5997),
    .D(net6150),
    .Q(\fpga_top.bus_gather.u_read_adr[7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _24813_ (.RESET_B(net5973),
    .D(_01407_),
    .Q(\fpga_top.bus_gather.u_read_adr[8] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _24814_ (.RESET_B(net5920),
    .D(net6121),
    .Q(\fpga_top.bus_gather.u_read_adr[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _24815_ (.RESET_B(net5920),
    .D(net6342),
    .Q(\fpga_top.bus_gather.u_read_adr[10] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _24816_ (.RESET_B(net5920),
    .D(_01410_),
    .Q(\fpga_top.bus_gather.u_read_adr[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _24817_ (.RESET_B(net5972),
    .D(_01411_),
    .Q(\fpga_top.bus_gather.u_read_adr[12] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _24818_ (.RESET_B(net5972),
    .D(net6287),
    .Q(\fpga_top.bus_gather.u_read_adr[13] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _24819_ (.RESET_B(net5964),
    .D(net6258),
    .Q(\fpga_top.bus_gather.u_read_adr[14] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_2 _24820_ (.RESET_B(net5964),
    .D(net6226),
    .Q(\fpga_top.bus_gather.u_read_adr[15] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_2 _24821_ (.RESET_B(net5964),
    .D(net6232),
    .Q(\fpga_top.bus_gather.u_read_adr[16] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_2 _24822_ (.RESET_B(net5976),
    .D(net6256),
    .Q(\fpga_top.bus_gather.u_read_adr[17] ),
    .CLK(clknet_leaf_294_clk));
 sg13g2_dfrbpq_2 _24823_ (.RESET_B(net5968),
    .D(net6290),
    .Q(\fpga_top.bus_gather.u_read_adr[18] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_2 _24824_ (.RESET_B(net5968),
    .D(net6265),
    .Q(\fpga_top.bus_gather.u_read_adr[19] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_2 _24825_ (.RESET_B(net5964),
    .D(net6292),
    .Q(\fpga_top.bus_gather.u_read_adr[20] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_2 _24826_ (.RESET_B(net5968),
    .D(net6528),
    .Q(\fpga_top.bus_gather.u_read_adr[21] ),
    .CLK(clknet_leaf_296_clk));
 sg13g2_dfrbpq_2 _24827_ (.RESET_B(net5964),
    .D(net6234),
    .Q(\fpga_top.bus_gather.u_read_adr[22] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_2 _24828_ (.RESET_B(net5964),
    .D(_01422_),
    .Q(\fpga_top.bus_gather.u_read_adr[23] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_2 _24829_ (.RESET_B(net5961),
    .D(net6320),
    .Q(\fpga_top.bus_gather.u_read_adr[24] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _24830_ (.RESET_B(net5961),
    .D(net6240),
    .Q(\fpga_top.bus_gather.u_read_adr[25] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _24831_ (.RESET_B(net5962),
    .D(net3955),
    .Q(\fpga_top.bus_gather.u_read_adr[26] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _24832_ (.RESET_B(net5909),
    .D(_01426_),
    .Q(\fpga_top.bus_gather.u_read_adr[27] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_2 _24833_ (.RESET_B(net5909),
    .D(_01427_),
    .Q(\fpga_top.bus_gather.u_read_adr[28] ),
    .CLK(clknet_leaf_315_clk));
 sg13g2_dfrbpq_1 _24834_ (.RESET_B(net5912),
    .D(_01428_),
    .Q(\fpga_top.bus_gather.u_read_adr[29] ),
    .CLK(clknet_leaf_316_clk));
 sg13g2_dfrbpq_2 _24835_ (.RESET_B(net5912),
    .D(_01429_),
    .Q(\fpga_top.bus_gather.u_read_adr[30] ),
    .CLK(clknet_leaf_297_clk));
 sg13g2_dfrbpq_2 _24836_ (.RESET_B(net5946),
    .D(_01430_),
    .Q(\fpga_top.bus_gather.u_read_adr[31] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _24837_ (.RESET_B(net5946),
    .D(net1642),
    .Q(\fpga_top.uart_top.uart_logics.cmd_read_adr[32] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _24838_ (.RESET_B(net5884),
    .D(_01432_),
    .Q(\fpga_top.uart_top.uart_if.byte_data[0] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _24839_ (.RESET_B(net5885),
    .D(net6405),
    .Q(\fpga_top.uart_top.uart_if.byte_data[1] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24840_ (.RESET_B(net5882),
    .D(_01434_),
    .Q(\fpga_top.uart_top.uart_if.byte_data[2] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24841_ (.RESET_B(net5882),
    .D(net6409),
    .Q(\fpga_top.uart_top.uart_if.byte_data[3] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24842_ (.RESET_B(net5882),
    .D(net3660),
    .Q(\fpga_top.uart_top.uart_if.byte_data[4] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _24843_ (.RESET_B(net5883),
    .D(_01437_),
    .Q(\fpga_top.uart_top.uart_if.byte_data[5] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _24844_ (.RESET_B(net5882),
    .D(_01438_),
    .Q(\fpga_top.uart_top.uart_if.byte_data[6] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _24845_ (.RESET_B(net5882),
    .D(_01439_),
    .Q(\fpga_top.uart_top.uart_if.byte_data[7] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _24846_ (.RESET_B(net5954),
    .D(net1379),
    .Q(\fpga_top.uart_top.uart_logics.trash_cond_dly ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _24847_ (.RESET_B(net6007),
    .D(net1852),
    .Q(\fpga_top.uart_top.uart_logics.rdata_snd_wait_dly ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _24848_ (.RESET_B(net5956),
    .D(net3316),
    .Q(\fpga_top.uart_top.uart_logics.write_stat ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _24849_ (.RESET_B(net1309),
    .D(_01441_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _24850_ (.RESET_B(net1308),
    .D(_01442_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][1] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _24851_ (.RESET_B(net1307),
    .D(_01443_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][2] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _24852_ (.RESET_B(net1306),
    .D(_01444_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _24853_ (.RESET_B(net1305),
    .D(_01445_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][4] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _24854_ (.RESET_B(net1304),
    .D(_01446_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _24855_ (.RESET_B(net1303),
    .D(_01447_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _24856_ (.RESET_B(net1302),
    .D(_01448_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][7] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _24857_ (.RESET_B(net6007),
    .D(net1314),
    .Q(_00126_),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _24858_ (.RESET_B(net5954),
    .D(_00147_),
    .Q(_00127_),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _24859_ (.RESET_B(net6028),
    .D(\fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[0] ),
    .Q(\fpga_top.cpu_top.cpu_state_machine.cpu_state[0] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _24860_ (.RESET_B(net6028),
    .D(\fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[1] ),
    .Q(\fpga_top.cpu_top.cpu_state_machine.cpu_state[1] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _24861_ (.RESET_B(net6028),
    .D(\fpga_top.cpu_top.cpu_state_machine.cpu_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/sequencer.v:70$1116.$result[2] ),
    .Q(\fpga_top.cpu_top.cpu_state_machine.cpu_state[2] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _24862_ (.RESET_B(net5993),
    .D(net1811),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[2] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24863_ (.RESET_B(net5993),
    .D(net1700),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[3] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24864_ (.RESET_B(net5994),
    .D(net3368),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[4] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24865_ (.RESET_B(net5993),
    .D(net1521),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[5] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_1 _24866_ (.RESET_B(net5993),
    .D(net1476),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[6] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_1 _24867_ (.RESET_B(net6042),
    .D(net1542),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[7] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_1 _24868_ (.RESET_B(net5993),
    .D(_01455_),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[8] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_1 _24869_ (.RESET_B(net6041),
    .D(net1478),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[9] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24870_ (.RESET_B(net6043),
    .D(net1418),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[10] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24871_ (.RESET_B(net6034),
    .D(net1510),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[11] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24872_ (.RESET_B(net6041),
    .D(net1532),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[12] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24873_ (.RESET_B(net6041),
    .D(net1496),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[13] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24874_ (.RESET_B(net6041),
    .D(net1551),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[14] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24875_ (.RESET_B(net6041),
    .D(net1447),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[15] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_1 _24876_ (.RESET_B(net6057),
    .D(net3754),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[16] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_1 _24877_ (.RESET_B(net6059),
    .D(net1441),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[17] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _24878_ (.RESET_B(net6043),
    .D(net1525),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[18] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_1 _24879_ (.RESET_B(net6062),
    .D(net1583),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[19] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _24880_ (.RESET_B(net6043),
    .D(net1513),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[20] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _24881_ (.RESET_B(net6060),
    .D(net1507),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[21] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _24882_ (.RESET_B(net6060),
    .D(net3780),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[22] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _24883_ (.RESET_B(net6060),
    .D(net1556),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[23] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _24884_ (.RESET_B(net6059),
    .D(net1547),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[24] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _24885_ (.RESET_B(net6043),
    .D(net1945),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[25] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_1 _24886_ (.RESET_B(net6062),
    .D(net1601),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[26] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _24887_ (.RESET_B(net6062),
    .D(net1592),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[27] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _24888_ (.RESET_B(net6060),
    .D(net3648),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[28] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_1 _24889_ (.RESET_B(net6057),
    .D(net2028),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[29] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _24890_ (.RESET_B(net6062),
    .D(net1677),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[30] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _24891_ (.RESET_B(net6044),
    .D(net1439),
    .Q(\fpga_top.cpu_top.execution.csr_array.pc_excep2[31] ),
    .CLK(clknet_leaf_285_clk));
 sg13g2_dfrbpq_2 _24892_ (.RESET_B(net5987),
    .D(_01479_),
    .Q(\fpga_top.cpu_top.pc_stage.pc_int_ecall_syn_state ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _24893_ (.RESET_B(net5994),
    .D(_01480_),
    .Q(\fpga_top.bus_gather.i_read_adr[2] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _24894_ (.RESET_B(net5989),
    .D(_01481_),
    .Q(\fpga_top.bus_gather.i_read_adr[3] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_1 _24895_ (.RESET_B(net5995),
    .D(net6499),
    .Q(\fpga_top.bus_gather.i_read_adr[4] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _24896_ (.RESET_B(net5995),
    .D(_01483_),
    .Q(\fpga_top.bus_gather.i_read_adr[5] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_1 _24897_ (.RESET_B(net5989),
    .D(net6541),
    .Q(\fpga_top.bus_gather.i_read_adr[6] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _24898_ (.RESET_B(net5991),
    .D(_01485_),
    .Q(\fpga_top.bus_gather.i_read_adr[7] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _24899_ (.RESET_B(net5994),
    .D(net2542),
    .Q(\fpga_top.bus_gather.i_read_adr[8] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _24900_ (.RESET_B(net6042),
    .D(_01487_),
    .Q(\fpga_top.bus_gather.i_read_adr[9] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _24901_ (.RESET_B(net6041),
    .D(_01488_),
    .Q(\fpga_top.bus_gather.i_read_adr[10] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24902_ (.RESET_B(net5994),
    .D(_01489_),
    .Q(\fpga_top.bus_gather.i_read_adr[11] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _24903_ (.RESET_B(net6042),
    .D(_01490_),
    .Q(\fpga_top.bus_gather.i_read_adr[12] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _24904_ (.RESET_B(net6042),
    .D(_01491_),
    .Q(\fpga_top.bus_gather.i_read_adr[13] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24905_ (.RESET_B(net6042),
    .D(net6505),
    .Q(\fpga_top.bus_gather.i_read_adr[14] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24906_ (.RESET_B(net6041),
    .D(_01493_),
    .Q(\fpga_top.bus_gather.i_read_adr[15] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_1 _24907_ (.RESET_B(net6044),
    .D(net6553),
    .Q(\fpga_top.bus_gather.i_read_adr[16] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _24908_ (.RESET_B(net6041),
    .D(_01495_),
    .Q(\fpga_top.bus_gather.i_read_adr[17] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24909_ (.RESET_B(net6043),
    .D(_01496_),
    .Q(\fpga_top.bus_gather.i_read_adr[18] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24910_ (.RESET_B(net5995),
    .D(net6580),
    .Q(\fpga_top.bus_gather.i_read_adr[19] ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_2 _24911_ (.RESET_B(net6057),
    .D(_01498_),
    .Q(\fpga_top.bus_gather.i_read_adr[20] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _24912_ (.RESET_B(net6058),
    .D(_01499_),
    .Q(\fpga_top.bus_gather.i_read_adr[21] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_1 _24913_ (.RESET_B(net6058),
    .D(_01500_),
    .Q(\fpga_top.bus_gather.i_read_adr[22] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _24914_ (.RESET_B(net6057),
    .D(net6476),
    .Q(\fpga_top.bus_gather.i_read_adr[23] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _24915_ (.RESET_B(net6043),
    .D(net6550),
    .Q(\fpga_top.bus_gather.i_read_adr[24] ),
    .CLK(clknet_leaf_286_clk));
 sg13g2_dfrbpq_2 _24916_ (.RESET_B(net6044),
    .D(_01503_),
    .Q(\fpga_top.bus_gather.i_read_adr[25] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _24917_ (.RESET_B(net6057),
    .D(_01504_),
    .Q(\fpga_top.bus_gather.i_read_adr[26] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _24918_ (.RESET_B(net6058),
    .D(_01505_),
    .Q(\fpga_top.bus_gather.i_read_adr[27] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _24919_ (.RESET_B(net6058),
    .D(_01506_),
    .Q(\fpga_top.bus_gather.i_read_adr[28] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _24920_ (.RESET_B(net6057),
    .D(_01507_),
    .Q(\fpga_top.bus_gather.i_read_adr[29] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _24921_ (.RESET_B(net5994),
    .D(_01508_),
    .Q(\fpga_top.bus_gather.i_read_adr[30] ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_2 _24922_ (.RESET_B(net5991),
    .D(_01509_),
    .Q(\fpga_top.bus_gather.i_read_adr[31] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _24923_ (.RESET_B(net5990),
    .D(net1377),
    .Q(\fpga_top.cpu_top.pc_stage.g_interrupt_latch ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_2 _24924_ (.RESET_B(net5992),
    .D(_01511_),
    .Q(\fpga_top.cpu_top.pc_stage.cpu_adr_ld ),
    .CLK(clknet_leaf_288_clk));
 sg13g2_dfrbpq_1 _24925_ (.RESET_B(net5990),
    .D(_01512_),
    .Q(\fpga_top.cpu_top.pc_stage.frc_cntr_val_leq_latch ),
    .CLK(clknet_leaf_293_clk));
 sg13g2_dfrbpq_1 _24926_ (.RESET_B(net5989),
    .D(net6354),
    .Q(\fpga_top.cpu_top.pc_stage.frc_cntr_val_leq_lat ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _24927_ (.RESET_B(net6024),
    .D(_01513_),
    .Q(\fpga_top.cpu_top.inst_mem_read.imr_stat ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _24928_ (.RESET_B(net5995),
    .D(net1845),
    .Q(\fpga_top.cpu_top.pc_stage.cmd_ebreak_pc_pre ),
    .CLK(clknet_leaf_287_clk));
 sg13g2_dfrbpq_1 _24929_ (.RESET_B(net1296),
    .D(_01515_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][0] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _24930_ (.RESET_B(net1295),
    .D(_01516_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][1] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _24931_ (.RESET_B(net1294),
    .D(_01517_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][2] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _24932_ (.RESET_B(net1293),
    .D(_01518_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][3] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _24933_ (.RESET_B(net1292),
    .D(_01519_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][4] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _24934_ (.RESET_B(net1291),
    .D(_01520_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][5] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _24935_ (.RESET_B(net1290),
    .D(_01521_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][6] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _24936_ (.RESET_B(net1289),
    .D(_01522_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][7] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _24937_ (.RESET_B(net1288),
    .D(_01523_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][8] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _24938_ (.RESET_B(net1287),
    .D(_01524_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][9] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _24939_ (.RESET_B(net1286),
    .D(_01525_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _24940_ (.RESET_B(net1285),
    .D(_01526_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][11] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _24941_ (.RESET_B(net1284),
    .D(_01527_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][12] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _24942_ (.RESET_B(net1283),
    .D(_01528_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][13] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _24943_ (.RESET_B(net1282),
    .D(_01529_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][14] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _24944_ (.RESET_B(net1281),
    .D(_01530_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][15] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _24945_ (.RESET_B(net1280),
    .D(_01531_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][16] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _24946_ (.RESET_B(net1279),
    .D(_01532_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][17] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _24947_ (.RESET_B(net1278),
    .D(_01533_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][18] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _24948_ (.RESET_B(net1277),
    .D(_01534_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][19] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _24949_ (.RESET_B(net1276),
    .D(_01535_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][20] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _24950_ (.RESET_B(net1275),
    .D(_01536_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][21] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _24951_ (.RESET_B(net1274),
    .D(_01537_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][22] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _24952_ (.RESET_B(net1273),
    .D(_01538_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][23] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _24953_ (.RESET_B(net1272),
    .D(_01539_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][24] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _24954_ (.RESET_B(net1271),
    .D(_01540_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][25] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _24955_ (.RESET_B(net1270),
    .D(_01541_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][26] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _24956_ (.RESET_B(net1269),
    .D(_01542_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][27] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _24957_ (.RESET_B(net1268),
    .D(_01543_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][28] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _24958_ (.RESET_B(net1267),
    .D(_01544_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][29] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _24959_ (.RESET_B(net1266),
    .D(_01545_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][30] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _24960_ (.RESET_B(net1265),
    .D(_01546_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _24961_ (.RESET_B(net1264),
    .D(_01547_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][0] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _24962_ (.RESET_B(net1263),
    .D(_01548_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][1] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _24963_ (.RESET_B(net1262),
    .D(_01549_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][2] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _24964_ (.RESET_B(net1261),
    .D(_01550_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][3] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _24965_ (.RESET_B(net1260),
    .D(_01551_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][4] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _24966_ (.RESET_B(net1259),
    .D(_01552_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][5] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _24967_ (.RESET_B(net1258),
    .D(_01553_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][6] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _24968_ (.RESET_B(net1257),
    .D(_01554_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][7] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _24969_ (.RESET_B(net1256),
    .D(_01555_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][8] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _24970_ (.RESET_B(net1255),
    .D(_01556_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][9] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _24971_ (.RESET_B(net1254),
    .D(_01557_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _24972_ (.RESET_B(net1253),
    .D(_01558_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][11] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _24973_ (.RESET_B(net1252),
    .D(_01559_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][12] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _24974_ (.RESET_B(net1251),
    .D(_01560_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][13] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _24975_ (.RESET_B(net1250),
    .D(_01561_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][14] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _24976_ (.RESET_B(net1249),
    .D(_01562_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][15] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _24977_ (.RESET_B(net1248),
    .D(_01563_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][16] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _24978_ (.RESET_B(net1247),
    .D(_01564_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][17] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _24979_ (.RESET_B(net1246),
    .D(_01565_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][18] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _24980_ (.RESET_B(net1245),
    .D(_01566_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][19] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _24981_ (.RESET_B(net1244),
    .D(_01567_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][20] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _24982_ (.RESET_B(net1243),
    .D(_01568_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][21] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _24983_ (.RESET_B(net1242),
    .D(_01569_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][22] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _24984_ (.RESET_B(net1241),
    .D(_01570_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][23] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _24985_ (.RESET_B(net1240),
    .D(_01571_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][24] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _24986_ (.RESET_B(net1239),
    .D(_01572_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][25] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _24987_ (.RESET_B(net1238),
    .D(_01573_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][26] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _24988_ (.RESET_B(net1237),
    .D(_01574_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][27] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _24989_ (.RESET_B(net1236),
    .D(_01575_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][28] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _24990_ (.RESET_B(net1235),
    .D(_01576_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][29] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _24991_ (.RESET_B(net1234),
    .D(_01577_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][30] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _24992_ (.RESET_B(net1003),
    .D(_01578_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _24993_ (.RESET_B(net6024),
    .D(net1380),
    .Q(\fpga_top.cpu_top.inst_mem_read.imr_stat_dly ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _24994_ (.RESET_B(net6027),
    .D(net3584),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[0] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _24995_ (.RESET_B(net6016),
    .D(_01580_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[1] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _24996_ (.RESET_B(net6027),
    .D(_01581_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[2] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _24997_ (.RESET_B(net6017),
    .D(net1456),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[3] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _24998_ (.RESET_B(net6017),
    .D(net3156),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[4] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _24999_ (.RESET_B(net6017),
    .D(net1529),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[5] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _25000_ (.RESET_B(net6017),
    .D(_01585_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[6] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _25001_ (.RESET_B(net6017),
    .D(_01586_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[7] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _25002_ (.RESET_B(net6017),
    .D(_01587_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[8] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _25003_ (.RESET_B(net6069),
    .D(_01588_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[9] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _25004_ (.RESET_B(net6065),
    .D(_01589_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[10] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _25005_ (.RESET_B(net6017),
    .D(net1640),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[11] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _25006_ (.RESET_B(net6065),
    .D(net1795),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[12] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _25007_ (.RESET_B(net6066),
    .D(_01592_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[13] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _25008_ (.RESET_B(net6065),
    .D(_01593_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[14] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _25009_ (.RESET_B(net6066),
    .D(_01594_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[15] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _25010_ (.RESET_B(net6066),
    .D(_01595_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[16] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _25011_ (.RESET_B(net6066),
    .D(_01596_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[17] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _25012_ (.RESET_B(net6068),
    .D(_01597_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[18] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _25013_ (.RESET_B(net6070),
    .D(_01598_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[19] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _25014_ (.RESET_B(net6071),
    .D(net1833),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[20] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _25015_ (.RESET_B(net6070),
    .D(_01600_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[21] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _25016_ (.RESET_B(net6071),
    .D(net1743),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[22] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _25017_ (.RESET_B(net6071),
    .D(_01602_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[23] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _25018_ (.RESET_B(net6068),
    .D(_01603_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[24] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _25019_ (.RESET_B(net6071),
    .D(_01604_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[25] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _25020_ (.RESET_B(net6071),
    .D(_01605_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[26] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _25021_ (.RESET_B(net6072),
    .D(_01606_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[27] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_1 _25022_ (.RESET_B(net6070),
    .D(_01607_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[28] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _25023_ (.RESET_B(net6071),
    .D(_01608_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[29] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _25024_ (.RESET_B(net6071),
    .D(net2033),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[30] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _25025_ (.RESET_B(net6067),
    .D(_01610_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[31] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _25026_ (.RESET_B(net6020),
    .D(_01611_),
    .Q(\fpga_top.cpu_top.decoder.illegal_ops_inst[0] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _25027_ (.RESET_B(net6020),
    .D(_01612_),
    .Q(\fpga_top.cpu_top.decoder.illegal_ops_inst[1] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _25028_ (.RESET_B(net6014),
    .D(_01613_),
    .Q(\fpga_top.cpu_top.decoder.illegal_ops_inst[2] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _25029_ (.RESET_B(net6016),
    .D(_01614_),
    .Q(\fpga_top.cpu_top.decoder.illegal_ops_inst[3] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25030_ (.RESET_B(net6016),
    .D(_01615_),
    .Q(\fpga_top.cpu_top.decoder.illegal_ops_inst[4] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25031_ (.RESET_B(net6020),
    .D(_01616_),
    .Q(\fpga_top.cpu_top.decoder.illegal_ops_inst[5] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _25032_ (.RESET_B(net6016),
    .D(_01617_),
    .Q(\fpga_top.cpu_top.decoder.illegal_ops_inst[6] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25033_ (.RESET_B(net6014),
    .D(_01618_),
    .Q(\fpga_top.cpu_top.br_ofs[11] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25034_ (.RESET_B(net6020),
    .D(_01619_),
    .Q(\fpga_top.cpu_top.br_ofs[1] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _25035_ (.RESET_B(net6026),
    .D(_01620_),
    .Q(\fpga_top.cpu_top.br_ofs[2] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _25036_ (.RESET_B(net6020),
    .D(_01621_),
    .Q(\fpga_top.cpu_top.br_ofs[3] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _25037_ (.RESET_B(net6020),
    .D(_01622_),
    .Q(\fpga_top.cpu_top.br_ofs[4] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _25038_ (.RESET_B(net6026),
    .D(_01623_),
    .Q(\fpga_top.cpu_top.alu_code[0] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _25039_ (.RESET_B(net6026),
    .D(_01624_),
    .Q(\fpga_top.cpu_top.alu_code[1] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _25040_ (.RESET_B(net6026),
    .D(_01625_),
    .Q(\fpga_top.cpu_top.alu_code[2] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25041_ (.RESET_B(net6017),
    .D(_01626_),
    .Q(\fpga_top.cpu_top.csr_uimm[0] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _25042_ (.RESET_B(net6016),
    .D(_01627_),
    .Q(\fpga_top.cpu_top.csr_uimm[1] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25043_ (.RESET_B(net6016),
    .D(_01628_),
    .Q(\fpga_top.cpu_top.csr_uimm[2] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25044_ (.RESET_B(net6018),
    .D(_01629_),
    .Q(\fpga_top.cpu_top.csr_uimm[3] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25045_ (.RESET_B(net6016),
    .D(_01630_),
    .Q(\fpga_top.cpu_top.csr_uimm[4] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _25046_ (.RESET_B(net6011),
    .D(_01631_),
    .Q(\fpga_top.cpu_top.alui_shamt[0] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25047_ (.RESET_B(net6019),
    .D(_01632_),
    .Q(\fpga_top.cpu_top.alui_shamt[1] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25048_ (.RESET_B(net6002),
    .D(_01633_),
    .Q(\fpga_top.cpu_top.alui_shamt[2] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25049_ (.RESET_B(net6011),
    .D(_01634_),
    .Q(\fpga_top.cpu_top.alui_shamt[3] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _25050_ (.RESET_B(net6011),
    .D(net6518),
    .Q(\fpga_top.cpu_top.alui_shamt[4] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25051_ (.RESET_B(net6015),
    .D(net6446),
    .Q(\fpga_top.cpu_top.br_ofs[5] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _25052_ (.RESET_B(net6011),
    .D(net6556),
    .Q(\fpga_top.cpu_top.br_ofs[6] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _25053_ (.RESET_B(net6027),
    .D(net6426),
    .Q(\fpga_top.cpu_top.br_ofs[7] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _25054_ (.RESET_B(net6026),
    .D(_01639_),
    .Q(\fpga_top.cpu_top.br_ofs[8] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _25055_ (.RESET_B(net6021),
    .D(_01640_),
    .Q(\fpga_top.cpu_top.br_ofs[9] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _25056_ (.RESET_B(net6014),
    .D(_01641_),
    .Q(\fpga_top.cpu_top.br_ofs[10] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _25057_ (.RESET_B(net6015),
    .D(_01642_),
    .Q(\fpga_top.cpu_top.br_ofs[12] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _25058_ (.RESET_B(net6066),
    .D(_01643_),
    .Q(\fpga_top.bus_gather.d_write_data[0] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _25059_ (.RESET_B(net6018),
    .D(_01644_),
    .Q(\fpga_top.bus_gather.d_write_data[1] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25060_ (.RESET_B(net6027),
    .D(_01645_),
    .Q(\fpga_top.bus_gather.d_write_data[2] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25061_ (.RESET_B(net6018),
    .D(_01646_),
    .Q(\fpga_top.bus_gather.d_write_data[3] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25062_ (.RESET_B(net6016),
    .D(_01647_),
    .Q(\fpga_top.bus_gather.d_write_data[4] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _25063_ (.RESET_B(net6069),
    .D(_01648_),
    .Q(\fpga_top.bus_gather.d_write_data[5] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _25064_ (.RESET_B(net6065),
    .D(_01649_),
    .Q(\fpga_top.bus_gather.d_write_data[6] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _25065_ (.RESET_B(net6027),
    .D(_01650_),
    .Q(\fpga_top.bus_gather.d_write_data[7] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25066_ (.RESET_B(net6069),
    .D(_01651_),
    .Q(\fpga_top.bus_gather.d_write_data[8] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _25067_ (.RESET_B(net6026),
    .D(_01652_),
    .Q(\fpga_top.bus_gather.d_write_data[9] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25068_ (.RESET_B(net6027),
    .D(_01653_),
    .Q(\fpga_top.bus_gather.d_write_data[10] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25069_ (.RESET_B(net6065),
    .D(_01654_),
    .Q(\fpga_top.bus_gather.d_write_data[11] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _25070_ (.RESET_B(net6067),
    .D(_01655_),
    .Q(\fpga_top.bus_gather.d_write_data[12] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _25071_ (.RESET_B(net6065),
    .D(_01656_),
    .Q(\fpga_top.bus_gather.d_write_data[13] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _25072_ (.RESET_B(net6073),
    .D(_01657_),
    .Q(\fpga_top.bus_gather.d_write_data[14] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _25073_ (.RESET_B(net6067),
    .D(_01658_),
    .Q(\fpga_top.bus_gather.d_write_data[15] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _25074_ (.RESET_B(net6067),
    .D(_01659_),
    .Q(\fpga_top.bus_gather.d_write_data[16] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _25075_ (.RESET_B(net6073),
    .D(_01660_),
    .Q(\fpga_top.bus_gather.d_write_data[17] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _25076_ (.RESET_B(net6067),
    .D(_01661_),
    .Q(\fpga_top.bus_gather.d_write_data[18] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _25077_ (.RESET_B(net6070),
    .D(_01662_),
    .Q(\fpga_top.bus_gather.d_write_data[19] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _25078_ (.RESET_B(net6073),
    .D(_01663_),
    .Q(\fpga_top.bus_gather.d_write_data[20] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _25079_ (.RESET_B(net6070),
    .D(_01664_),
    .Q(\fpga_top.bus_gather.d_write_data[21] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _25080_ (.RESET_B(net6072),
    .D(_01665_),
    .Q(\fpga_top.bus_gather.d_write_data[22] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _25081_ (.RESET_B(net6074),
    .D(_01666_),
    .Q(\fpga_top.bus_gather.d_write_data[23] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _25082_ (.RESET_B(net6072),
    .D(_01667_),
    .Q(\fpga_top.bus_gather.d_write_data[24] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _25083_ (.RESET_B(net6074),
    .D(_01668_),
    .Q(\fpga_top.bus_gather.d_write_data[25] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _25084_ (.RESET_B(net6026),
    .D(_01669_),
    .Q(\fpga_top.bus_gather.d_write_data[26] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25085_ (.RESET_B(net6074),
    .D(_01670_),
    .Q(\fpga_top.bus_gather.d_write_data[27] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _25086_ (.RESET_B(net6074),
    .D(_01671_),
    .Q(\fpga_top.bus_gather.d_write_data[28] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _25087_ (.RESET_B(net6067),
    .D(_01672_),
    .Q(\fpga_top.bus_gather.d_write_data[29] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _25088_ (.RESET_B(net6073),
    .D(_01673_),
    .Q(\fpga_top.bus_gather.d_write_data[30] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _25089_ (.RESET_B(net6065),
    .D(_01674_),
    .Q(\fpga_top.bus_gather.d_write_data[31] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _25090_ (.RESET_B(net5993),
    .D(net1940),
    .Q(\fpga_top.cpu_top.pc_stage.cmd_ecall_pc_pre ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_2 _25091_ (.RESET_B(net6028),
    .D(net6221),
    .Q(\fpga_top.cpu_top.register_file.rfr_state[0] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _25092_ (.RESET_B(net6028),
    .D(\fpga_top.cpu_top.register_file.next_rfr_state[1] ),
    .Q(\fpga_top.cpu_top.register_file.rfr_state[1] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _25093_ (.RESET_B(net6028),
    .D(net3896),
    .Q(\fpga_top.cpu_top.register_file.rfr_state[2] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _25094_ (.RESET_B(net1231),
    .D(_01676_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][0] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _25095_ (.RESET_B(net1230),
    .D(_01677_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][1] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25096_ (.RESET_B(net1229),
    .D(_01678_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][2] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25097_ (.RESET_B(net1228),
    .D(_01679_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][3] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _25098_ (.RESET_B(net1227),
    .D(_01680_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][4] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25099_ (.RESET_B(net1226),
    .D(_01681_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _25100_ (.RESET_B(net1225),
    .D(_01682_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][6] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _25101_ (.RESET_B(net1224),
    .D(_01683_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][7] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25102_ (.RESET_B(net1223),
    .D(_01684_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][8] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25103_ (.RESET_B(net1222),
    .D(_01685_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][9] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _25104_ (.RESET_B(net1221),
    .D(_01686_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][10] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _25105_ (.RESET_B(net1220),
    .D(_01687_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][11] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _25106_ (.RESET_B(net1219),
    .D(_01688_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][12] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25107_ (.RESET_B(net1218),
    .D(_01689_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][13] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _25108_ (.RESET_B(net1217),
    .D(_01690_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][14] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _25109_ (.RESET_B(net1216),
    .D(_01691_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][15] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25110_ (.RESET_B(net1215),
    .D(_01692_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][16] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25111_ (.RESET_B(net1214),
    .D(_01693_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][17] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25112_ (.RESET_B(net1213),
    .D(_01694_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][18] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _25113_ (.RESET_B(net1212),
    .D(_01695_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][19] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _25114_ (.RESET_B(net1211),
    .D(_01696_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _25115_ (.RESET_B(net1210),
    .D(_01697_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][21] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _25116_ (.RESET_B(net1209),
    .D(_01698_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][22] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _25117_ (.RESET_B(net1208),
    .D(_01699_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][23] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25118_ (.RESET_B(net1207),
    .D(_01700_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][24] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25119_ (.RESET_B(net1206),
    .D(_01701_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][25] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25120_ (.RESET_B(net1205),
    .D(_01702_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][26] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25121_ (.RESET_B(net1204),
    .D(_01703_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][27] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _25122_ (.RESET_B(net1203),
    .D(_01704_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][28] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _25123_ (.RESET_B(net1202),
    .D(_01705_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][29] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25124_ (.RESET_B(net1201),
    .D(_01706_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][30] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _25125_ (.RESET_B(net1200),
    .D(_01707_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][31] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25126_ (.RESET_B(net1199),
    .D(_01708_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][0] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _25127_ (.RESET_B(net1198),
    .D(_01709_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][1] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25128_ (.RESET_B(net1197),
    .D(_01710_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][2] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25129_ (.RESET_B(net1196),
    .D(_01711_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][3] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _25130_ (.RESET_B(net1195),
    .D(_01712_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][4] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25131_ (.RESET_B(net1194),
    .D(_01713_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][5] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25132_ (.RESET_B(net1193),
    .D(_01714_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][6] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _25133_ (.RESET_B(net1192),
    .D(_01715_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][7] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _25134_ (.RESET_B(net1191),
    .D(_01716_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][8] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25135_ (.RESET_B(net1190),
    .D(_01717_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][9] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _25136_ (.RESET_B(net1189),
    .D(_01718_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25137_ (.RESET_B(net1188),
    .D(_01719_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][11] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25138_ (.RESET_B(net1187),
    .D(_01720_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][12] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25139_ (.RESET_B(net1186),
    .D(_01721_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][13] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _25140_ (.RESET_B(net1185),
    .D(_01722_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][14] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _25141_ (.RESET_B(net1184),
    .D(_01723_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][15] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25142_ (.RESET_B(net1183),
    .D(_01724_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][16] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25143_ (.RESET_B(net1182),
    .D(_01725_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][17] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _25144_ (.RESET_B(net1181),
    .D(_01726_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][18] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _25145_ (.RESET_B(net1180),
    .D(_01727_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][19] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _25146_ (.RESET_B(net1179),
    .D(_01728_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _25147_ (.RESET_B(net1178),
    .D(_01729_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][21] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _25148_ (.RESET_B(net1177),
    .D(_01730_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][22] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _25149_ (.RESET_B(net1176),
    .D(_01731_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][23] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25150_ (.RESET_B(net1175),
    .D(_01732_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][24] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25151_ (.RESET_B(net1174),
    .D(_01733_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][25] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _25152_ (.RESET_B(net1173),
    .D(_01734_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][26] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25153_ (.RESET_B(net1172),
    .D(_01735_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][27] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _25154_ (.RESET_B(net1171),
    .D(_01736_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][28] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _25155_ (.RESET_B(net1170),
    .D(_01737_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][29] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25156_ (.RESET_B(net1169),
    .D(_01738_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][30] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _25157_ (.RESET_B(net1168),
    .D(_01739_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][31] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25158_ (.RESET_B(net1167),
    .D(_01740_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][0] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _25159_ (.RESET_B(net1166),
    .D(_01741_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][1] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25160_ (.RESET_B(net1165),
    .D(_01742_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][2] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _25161_ (.RESET_B(net1164),
    .D(_01743_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][3] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _25162_ (.RESET_B(net1163),
    .D(_01744_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][4] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _25163_ (.RESET_B(net1162),
    .D(_01745_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][5] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _25164_ (.RESET_B(net1161),
    .D(_01746_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][6] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25165_ (.RESET_B(net1160),
    .D(_01747_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][7] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _25166_ (.RESET_B(net1159),
    .D(_01748_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][8] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _25167_ (.RESET_B(net1158),
    .D(_01749_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][9] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25168_ (.RESET_B(net1157),
    .D(_01750_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25169_ (.RESET_B(net1156),
    .D(_01751_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][11] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_1 _25170_ (.RESET_B(net1155),
    .D(_01752_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][12] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _25171_ (.RESET_B(net1154),
    .D(_01753_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][13] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _25172_ (.RESET_B(net1153),
    .D(_01754_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][14] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _25173_ (.RESET_B(net1152),
    .D(_01755_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][15] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25174_ (.RESET_B(net1151),
    .D(_01756_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][16] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25175_ (.RESET_B(net1150),
    .D(_01757_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][17] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_1 _25176_ (.RESET_B(net1149),
    .D(_01758_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][18] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25177_ (.RESET_B(net1148),
    .D(_01759_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][19] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _25178_ (.RESET_B(net1147),
    .D(_01760_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][20] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25179_ (.RESET_B(net1146),
    .D(_01761_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _25180_ (.RESET_B(net1145),
    .D(_01762_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][22] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _25181_ (.RESET_B(net1144),
    .D(_01763_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][23] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _25182_ (.RESET_B(net1143),
    .D(_01764_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][24] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _25183_ (.RESET_B(net1142),
    .D(_01765_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][25] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25184_ (.RESET_B(net1141),
    .D(_01766_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][26] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _25185_ (.RESET_B(net1140),
    .D(_01767_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][27] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _25186_ (.RESET_B(net1139),
    .D(_01768_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][28] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _25187_ (.RESET_B(net1138),
    .D(_01769_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][29] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25188_ (.RESET_B(net1137),
    .D(_01770_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][30] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _25189_ (.RESET_B(net1136),
    .D(_01771_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][31] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _25190_ (.RESET_B(net1135),
    .D(_01772_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][0] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25191_ (.RESET_B(net1134),
    .D(_01773_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][1] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25192_ (.RESET_B(net1133),
    .D(_01774_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][2] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25193_ (.RESET_B(net1132),
    .D(_01775_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][3] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _25194_ (.RESET_B(net1131),
    .D(_01776_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][4] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _25195_ (.RESET_B(net1130),
    .D(_01777_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _25196_ (.RESET_B(net1129),
    .D(_01778_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][6] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25197_ (.RESET_B(net1128),
    .D(_01779_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][7] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25198_ (.RESET_B(net1127),
    .D(_01780_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][8] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_1 _25199_ (.RESET_B(net1126),
    .D(_01781_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][9] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _25200_ (.RESET_B(net1125),
    .D(_01782_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][10] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25201_ (.RESET_B(net1124),
    .D(_01783_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][11] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _25202_ (.RESET_B(net1123),
    .D(_01784_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][12] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25203_ (.RESET_B(net1122),
    .D(_01785_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][13] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25204_ (.RESET_B(net1121),
    .D(_01786_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][14] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _25205_ (.RESET_B(net1120),
    .D(_01787_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][15] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_1 _25206_ (.RESET_B(net1119),
    .D(_01788_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][16] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25207_ (.RESET_B(net1118),
    .D(_01789_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][17] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _25208_ (.RESET_B(net1117),
    .D(_01790_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][18] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25209_ (.RESET_B(net1116),
    .D(_01791_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][19] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _25210_ (.RESET_B(net1115),
    .D(_01792_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][20] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25211_ (.RESET_B(net1114),
    .D(_01793_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][21] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _25212_ (.RESET_B(net1113),
    .D(_01794_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][22] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _25213_ (.RESET_B(net1112),
    .D(_01795_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][23] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _25214_ (.RESET_B(net1111),
    .D(_01796_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][24] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _25215_ (.RESET_B(net1110),
    .D(_01797_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][25] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25216_ (.RESET_B(net1109),
    .D(_01798_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][26] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _25217_ (.RESET_B(net1108),
    .D(_01799_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][27] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_1 _25218_ (.RESET_B(net1107),
    .D(_01800_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25219_ (.RESET_B(net1106),
    .D(_01801_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][29] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25220_ (.RESET_B(net1105),
    .D(_01802_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][30] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25221_ (.RESET_B(net1004),
    .D(_01803_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][31] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25222_ (.RESET_B(net1005),
    .D(\fpga_top.cpu_top.register_file.inst_rs[8] ),
    .Q(_00000_),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_1 _25223_ (.RESET_B(net1006),
    .D(\fpga_top.cpu_top.register_file.inst_rs[7] ),
    .Q(_00001_),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _25224_ (.RESET_B(net1007),
    .D(\fpga_top.cpu_top.register_file.inst_rs[6] ),
    .Q(_00002_),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _25225_ (.RESET_B(net1232),
    .D(\fpga_top.cpu_top.register_file.inst_rs[5] ),
    .Q(_00003_),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _25226_ (.RESET_B(net1104),
    .D(\fpga_top.cpu_top.register_file.inst_rs[4] ),
    .Q(_00004_),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_1 _25227_ (.RESET_B(net1103),
    .D(_01804_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][0] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25228_ (.RESET_B(net1102),
    .D(_01805_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][1] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25229_ (.RESET_B(net1101),
    .D(_01806_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][2] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25230_ (.RESET_B(net1100),
    .D(_01807_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][3] ),
    .CLK(clknet_leaf_255_clk));
 sg13g2_dfrbpq_1 _25231_ (.RESET_B(net1099),
    .D(_01808_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][4] ),
    .CLK(clknet_leaf_241_clk));
 sg13g2_dfrbpq_1 _25232_ (.RESET_B(net1098),
    .D(_01809_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][5] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25233_ (.RESET_B(net1097),
    .D(_01810_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][6] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25234_ (.RESET_B(net1096),
    .D(_01811_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][7] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25235_ (.RESET_B(net1095),
    .D(_01812_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][8] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_1 _25236_ (.RESET_B(net1094),
    .D(_01813_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][9] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_1 _25237_ (.RESET_B(net1093),
    .D(_01814_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][10] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _25238_ (.RESET_B(net1092),
    .D(_01815_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][11] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_1 _25239_ (.RESET_B(net1091),
    .D(_01816_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][12] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _25240_ (.RESET_B(net1090),
    .D(_01817_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][13] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _25241_ (.RESET_B(net1089),
    .D(_01818_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][14] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _25242_ (.RESET_B(net1088),
    .D(_01819_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][15] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25243_ (.RESET_B(net1087),
    .D(_01820_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][16] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _25244_ (.RESET_B(net1086),
    .D(_01821_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][17] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _25245_ (.RESET_B(net1085),
    .D(_01822_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][18] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25246_ (.RESET_B(net1084),
    .D(_01823_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][19] ),
    .CLK(clknet_leaf_253_clk));
 sg13g2_dfrbpq_1 _25247_ (.RESET_B(net1083),
    .D(_01824_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][20] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25248_ (.RESET_B(net1082),
    .D(_01825_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][21] ),
    .CLK(clknet_leaf_254_clk));
 sg13g2_dfrbpq_1 _25249_ (.RESET_B(net1081),
    .D(_01826_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][22] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _25250_ (.RESET_B(net1080),
    .D(_01827_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][23] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _25251_ (.RESET_B(net1079),
    .D(_01828_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][24] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25252_ (.RESET_B(net1078),
    .D(_01829_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _25253_ (.RESET_B(net1077),
    .D(_01830_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][26] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25254_ (.RESET_B(net1076),
    .D(_01831_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][27] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _25255_ (.RESET_B(net1075),
    .D(_01832_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25256_ (.RESET_B(net1074),
    .D(_01833_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][29] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _25257_ (.RESET_B(net1073),
    .D(_01834_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][30] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _25258_ (.RESET_B(net1072),
    .D(_01835_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25259_ (.RESET_B(net1071),
    .D(_01836_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][0] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25260_ (.RESET_B(net1070),
    .D(_01837_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][1] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25261_ (.RESET_B(net1069),
    .D(_01838_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][2] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _25262_ (.RESET_B(net1068),
    .D(_01839_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][3] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _25263_ (.RESET_B(net1067),
    .D(_01840_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][4] ),
    .CLK(clknet_leaf_239_clk));
 sg13g2_dfrbpq_1 _25264_ (.RESET_B(net1066),
    .D(_01841_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _25265_ (.RESET_B(net1065),
    .D(_01842_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][6] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_1 _25266_ (.RESET_B(net1064),
    .D(_01843_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][7] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _25267_ (.RESET_B(net1063),
    .D(_01844_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][8] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_1 _25268_ (.RESET_B(net1062),
    .D(_01845_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][9] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_1 _25269_ (.RESET_B(net1061),
    .D(_01846_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][10] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25270_ (.RESET_B(net1060),
    .D(_01847_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][11] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _25271_ (.RESET_B(net1059),
    .D(_01848_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][12] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25272_ (.RESET_B(net1058),
    .D(_01849_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][13] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _25273_ (.RESET_B(net1057),
    .D(_01850_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][14] ),
    .CLK(clknet_leaf_280_clk));
 sg13g2_dfrbpq_1 _25274_ (.RESET_B(net1056),
    .D(_01851_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][15] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25275_ (.RESET_B(net1055),
    .D(_01852_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][16] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _25276_ (.RESET_B(net1054),
    .D(_01853_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][17] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _25277_ (.RESET_B(net1053),
    .D(_01854_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][18] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25278_ (.RESET_B(net1052),
    .D(_01855_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][19] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _25279_ (.RESET_B(net1051),
    .D(_01856_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][20] ),
    .CLK(clknet_leaf_240_clk));
 sg13g2_dfrbpq_1 _25280_ (.RESET_B(net1050),
    .D(_01857_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][21] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_1 _25281_ (.RESET_B(net1049),
    .D(_01858_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][22] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_1 _25282_ (.RESET_B(net1048),
    .D(_01859_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][23] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _25283_ (.RESET_B(net1047),
    .D(_01860_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][24] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25284_ (.RESET_B(net1046),
    .D(_01861_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][25] ),
    .CLK(clknet_leaf_238_clk));
 sg13g2_dfrbpq_1 _25285_ (.RESET_B(net1045),
    .D(_01862_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][26] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _25286_ (.RESET_B(net1044),
    .D(_01863_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][27] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _25287_ (.RESET_B(net1043),
    .D(_01864_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][28] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_1 _25288_ (.RESET_B(net1042),
    .D(_01865_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][29] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _25289_ (.RESET_B(net1041),
    .D(_01866_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][30] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25290_ (.RESET_B(net1040),
    .D(_01867_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][31] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25291_ (.RESET_B(net1039),
    .D(_01868_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][0] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _25292_ (.RESET_B(net1038),
    .D(_01869_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][1] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _25293_ (.RESET_B(net1037),
    .D(_01870_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][2] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _25294_ (.RESET_B(net1036),
    .D(_01871_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][3] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _25295_ (.RESET_B(net1035),
    .D(_01872_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][4] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _25296_ (.RESET_B(net1034),
    .D(_01873_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][5] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25297_ (.RESET_B(net1033),
    .D(_01874_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][6] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _25298_ (.RESET_B(net1032),
    .D(_01875_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][7] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _25299_ (.RESET_B(net1031),
    .D(_01876_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][8] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _25300_ (.RESET_B(net1030),
    .D(_01877_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][9] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25301_ (.RESET_B(net1029),
    .D(_01878_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][10] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _25302_ (.RESET_B(net1028),
    .D(_01879_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][11] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _25303_ (.RESET_B(net1027),
    .D(_01880_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][12] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _25304_ (.RESET_B(net1026),
    .D(_01881_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][13] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _25305_ (.RESET_B(net1025),
    .D(_01882_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][14] ),
    .CLK(clknet_leaf_258_clk));
 sg13g2_dfrbpq_1 _25306_ (.RESET_B(net1024),
    .D(_01883_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][15] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _25307_ (.RESET_B(net1023),
    .D(_01884_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][16] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_1 _25308_ (.RESET_B(net1022),
    .D(_01885_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][17] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _25309_ (.RESET_B(net1021),
    .D(_01886_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][18] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _25310_ (.RESET_B(net1020),
    .D(_01887_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][19] ),
    .CLK(clknet_leaf_247_clk));
 sg13g2_dfrbpq_1 _25311_ (.RESET_B(net1019),
    .D(_01888_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][20] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _25312_ (.RESET_B(net1018),
    .D(_01889_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][21] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _25313_ (.RESET_B(net1017),
    .D(_01890_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][22] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _25314_ (.RESET_B(net1016),
    .D(_01891_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][23] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _25315_ (.RESET_B(net1015),
    .D(_01892_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][24] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25316_ (.RESET_B(net1014),
    .D(_01893_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][25] ),
    .CLK(clknet_leaf_237_clk));
 sg13g2_dfrbpq_1 _25317_ (.RESET_B(net1013),
    .D(_01894_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][26] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _25318_ (.RESET_B(net1012),
    .D(_01895_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][27] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_1 _25319_ (.RESET_B(net1011),
    .D(_01896_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][28] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _25320_ (.RESET_B(net1010),
    .D(_01897_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][29] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _25321_ (.RESET_B(net1009),
    .D(_01898_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][30] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_1 _25322_ (.RESET_B(net1008),
    .D(_01899_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][31] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _25323_ (.RESET_B(net5990),
    .D(_01900_),
    .Q(\fpga_top.cpu_top.csr_rmie ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_1 _25324_ (.RESET_B(net6019),
    .D(net1469),
    .Q(\fpga_top.cpu_top.data_rw_mem.unsigned_bit_dly ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _25325_ (.RESET_B(net5981),
    .D(_01902_),
    .Q(\fpga_top.cpu_top.csr_msie ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_2 _25326_ (.RESET_B(net5981),
    .D(_01903_),
    .Q(\fpga_top.cpu_top.csr_mtie ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_2 _25327_ (.RESET_B(net5981),
    .D(_01904_),
    .Q(\fpga_top.cpu_top.csr_meie ),
    .CLK(clknet_leaf_298_clk));
 sg13g2_dfrbpq_1 _25328_ (.RESET_B(net5990),
    .D(net2067),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mpie ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_1 _25329_ (.RESET_B(net5985),
    .D(net2081),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[0] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _25330_ (.RESET_B(net5982),
    .D(net1570),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[1] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _25331_ (.RESET_B(net6033),
    .D(_01908_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[2] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _25332_ (.RESET_B(net5981),
    .D(_01909_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[3] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _25333_ (.RESET_B(net5985),
    .D(_01910_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[4] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _25334_ (.RESET_B(net5985),
    .D(_01911_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[5] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_1 _25335_ (.RESET_B(net5978),
    .D(net1567),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[6] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _25336_ (.RESET_B(net5989),
    .D(_01913_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[7] ),
    .CLK(clknet_leaf_292_clk));
 sg13g2_dfrbpq_1 _25337_ (.RESET_B(net5978),
    .D(_01914_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[8] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_1 _25338_ (.RESET_B(net6035),
    .D(_01915_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[9] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _25339_ (.RESET_B(net6049),
    .D(_01916_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[10] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _25340_ (.RESET_B(net5981),
    .D(_01917_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[11] ),
    .CLK(clknet_leaf_299_clk));
 sg13g2_dfrbpq_1 _25341_ (.RESET_B(net5984),
    .D(_01918_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[12] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _25342_ (.RESET_B(net6038),
    .D(_01919_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[13] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_1 _25343_ (.RESET_B(net6032),
    .D(_01920_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[14] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_1 _25344_ (.RESET_B(net6038),
    .D(_01921_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[15] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_1 _25345_ (.RESET_B(net6039),
    .D(_01922_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[16] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_1 _25346_ (.RESET_B(net6057),
    .D(_01923_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[17] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_1 _25347_ (.RESET_B(net6048),
    .D(_01924_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[18] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _25348_ (.RESET_B(net6054),
    .D(_01925_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[19] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_1 _25349_ (.RESET_B(net6049),
    .D(_01926_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[20] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _25350_ (.RESET_B(net6054),
    .D(_01927_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[21] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _25351_ (.RESET_B(net6049),
    .D(_01928_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[22] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _25352_ (.RESET_B(net6054),
    .D(_01929_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[23] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _25353_ (.RESET_B(net6048),
    .D(_01930_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[24] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_1 _25354_ (.RESET_B(net6039),
    .D(_01931_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[25] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_1 _25355_ (.RESET_B(net6053),
    .D(_01932_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[26] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _25356_ (.RESET_B(net6053),
    .D(_01933_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[27] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _25357_ (.RESET_B(net6045),
    .D(_01934_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[28] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _25358_ (.RESET_B(net6054),
    .D(_01935_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[29] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _25359_ (.RESET_B(net6049),
    .D(_01936_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[30] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_1 _25360_ (.RESET_B(net6033),
    .D(net1789),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtval[31] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_1 _25361_ (.RESET_B(net5985),
    .D(net3494),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mcause[0] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _25362_ (.RESET_B(net5986),
    .D(net1706),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mcause[1] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_1 _25363_ (.RESET_B(net5988),
    .D(net3782),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mcause[2] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _25364_ (.RESET_B(net5987),
    .D(net3490),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mcause[3] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _25365_ (.RESET_B(net5986),
    .D(_01942_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mcause[4] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _25366_ (.RESET_B(net5988),
    .D(_01943_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mcause[5] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _25367_ (.RESET_B(net6034),
    .D(net3599),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mcause[6] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_1 _25368_ (.RESET_B(net5987),
    .D(_01945_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[2] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _25369_ (.RESET_B(net5987),
    .D(net1753),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[3] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _25370_ (.RESET_B(net5994),
    .D(net1879),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[4] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_2 _25371_ (.RESET_B(net5994),
    .D(_01948_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[5] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_2 _25372_ (.RESET_B(net5993),
    .D(_01949_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[6] ),
    .CLK(clknet_leaf_290_clk));
 sg13g2_dfrbpq_2 _25373_ (.RESET_B(net5993),
    .D(_01950_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[7] ),
    .CLK(clknet_leaf_289_clk));
 sg13g2_dfrbpq_1 _25374_ (.RESET_B(net5987),
    .D(net2128),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[8] ),
    .CLK(clknet_leaf_291_clk));
 sg13g2_dfrbpq_2 _25375_ (.RESET_B(net6035),
    .D(_01952_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[9] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25376_ (.RESET_B(net6038),
    .D(_01953_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[10] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _25377_ (.RESET_B(net6034),
    .D(net1820),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[11] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_1 _25378_ (.RESET_B(net6034),
    .D(_01955_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[12] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_2 _25379_ (.RESET_B(net6034),
    .D(_01956_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[13] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25380_ (.RESET_B(net6034),
    .D(net1980),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[14] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25381_ (.RESET_B(net6043),
    .D(net1818),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[15] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_2 _25382_ (.RESET_B(net6048),
    .D(net3349),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[16] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _25383_ (.RESET_B(net6061),
    .D(_01960_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[17] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_2 _25384_ (.RESET_B(net6039),
    .D(_01961_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[18] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _25385_ (.RESET_B(net6061),
    .D(_01962_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[19] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_1 _25386_ (.RESET_B(net6057),
    .D(net2211),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[20] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_2 _25387_ (.RESET_B(net6061),
    .D(_01964_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[21] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_2 _25388_ (.RESET_B(net6059),
    .D(net3338),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[22] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _25389_ (.RESET_B(net6059),
    .D(_01966_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[23] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _25390_ (.RESET_B(net6048),
    .D(_01967_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[24] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _25391_ (.RESET_B(net6038),
    .D(net1997),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[25] ),
    .CLK(clknet_leaf_275_clk));
 sg13g2_dfrbpq_2 _25392_ (.RESET_B(net6059),
    .D(_01969_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[26] ),
    .CLK(clknet_leaf_283_clk));
 sg13g2_dfrbpq_2 _25393_ (.RESET_B(net6060),
    .D(_01970_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[27] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _25394_ (.RESET_B(net6059),
    .D(net2049),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[28] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _25395_ (.RESET_B(net6059),
    .D(net1793),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[29] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _25396_ (.RESET_B(net6059),
    .D(_01973_),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[30] ),
    .CLK(clknet_leaf_282_clk));
 sg13g2_dfrbpq_2 _25397_ (.RESET_B(net6043),
    .D(net2011),
    .Q(\fpga_top.cpu_top.csr_mepc_ex[31] ),
    .CLK(clknet_leaf_284_clk));
 sg13g2_dfrbpq_1 _25398_ (.RESET_B(net5982),
    .D(_01975_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mpp[0] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_2 _25399_ (.RESET_B(net5981),
    .D(_01976_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mpp[1] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_1 _25400_ (.RESET_B(net6033),
    .D(_01977_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[0] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_1 _25401_ (.RESET_B(net5980),
    .D(_01978_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[1] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_1 _25402_ (.RESET_B(net6032),
    .D(_01979_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[2] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_1 _25403_ (.RESET_B(net5978),
    .D(_01980_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[3] ),
    .CLK(clknet_leaf_307_clk));
 sg13g2_dfrbpq_1 _25404_ (.RESET_B(net6033),
    .D(_01981_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[4] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _25405_ (.RESET_B(net5985),
    .D(_01982_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[5] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _25406_ (.RESET_B(net5979),
    .D(_01983_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[6] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _25407_ (.RESET_B(net5978),
    .D(_01984_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[7] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _25408_ (.RESET_B(net5984),
    .D(_01985_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[8] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _25409_ (.RESET_B(net6036),
    .D(net1553),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[9] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_1 _25410_ (.RESET_B(net6050),
    .D(_01987_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[10] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _25411_ (.RESET_B(net5978),
    .D(_01988_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[11] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _25412_ (.RESET_B(net5984),
    .D(_01989_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[12] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _25413_ (.RESET_B(net6036),
    .D(_01990_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[13] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _25414_ (.RESET_B(net6038),
    .D(_01991_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[14] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _25415_ (.RESET_B(net6036),
    .D(_01992_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[15] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _25416_ (.RESET_B(net6037),
    .D(net1613),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[16] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _25417_ (.RESET_B(net6052),
    .D(net2112),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[17] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _25418_ (.RESET_B(net6047),
    .D(_01995_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[18] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _25419_ (.RESET_B(net6051),
    .D(_01996_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[19] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _25420_ (.RESET_B(net6046),
    .D(_01997_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[20] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _25421_ (.RESET_B(net6055),
    .D(_01998_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[21] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _25422_ (.RESET_B(net6045),
    .D(_01999_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[22] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _25423_ (.RESET_B(net6051),
    .D(net2039),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[23] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _25424_ (.RESET_B(net6040),
    .D(_02001_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[24] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _25425_ (.RESET_B(net6037),
    .D(_02002_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[25] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _25426_ (.RESET_B(net6051),
    .D(_02003_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[26] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _25427_ (.RESET_B(net6053),
    .D(_02004_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[27] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_1 _25428_ (.RESET_B(net6050),
    .D(_02005_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[28] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _25429_ (.RESET_B(net6052),
    .D(_02006_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[29] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _25430_ (.RESET_B(net6045),
    .D(_02007_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[30] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _25431_ (.RESET_B(net6032),
    .D(_02008_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[31] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_1 _25432_ (.RESET_B(net5986),
    .D(_02009_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_spie ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_1 _25433_ (.RESET_B(net6033),
    .D(_02010_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[0] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _25434_ (.RESET_B(net5980),
    .D(_02011_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[1] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _25435_ (.RESET_B(net6032),
    .D(_02012_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[2] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_1 _25436_ (.RESET_B(net5978),
    .D(_02013_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[3] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _25437_ (.RESET_B(net6033),
    .D(_02014_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[4] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _25438_ (.RESET_B(net5985),
    .D(_02015_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[5] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _25439_ (.RESET_B(net5979),
    .D(_02016_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[6] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _25440_ (.RESET_B(net5978),
    .D(_02017_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[7] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_1 _25441_ (.RESET_B(net5984),
    .D(_02018_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[8] ),
    .CLK(clknet_leaf_306_clk));
 sg13g2_dfrbpq_1 _25442_ (.RESET_B(net6036),
    .D(net1586),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[9] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_1 _25443_ (.RESET_B(net6050),
    .D(_02020_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[10] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _25444_ (.RESET_B(net5978),
    .D(_02021_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[11] ),
    .CLK(clknet_leaf_308_clk));
 sg13g2_dfrbpq_1 _25445_ (.RESET_B(net6033),
    .D(_02022_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[12] ),
    .CLK(clknet_leaf_305_clk));
 sg13g2_dfrbpq_1 _25446_ (.RESET_B(net6037),
    .D(_02023_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[13] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _25447_ (.RESET_B(net6032),
    .D(_02024_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[14] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _25448_ (.RESET_B(net6037),
    .D(_02025_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[15] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _25449_ (.RESET_B(net6037),
    .D(net1518),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[16] ),
    .CLK(clknet_leaf_271_clk));
 sg13g2_dfrbpq_1 _25450_ (.RESET_B(net6050),
    .D(net1590),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[17] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _25451_ (.RESET_B(net6047),
    .D(_02028_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[18] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _25452_ (.RESET_B(net6051),
    .D(_02029_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[19] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _25453_ (.RESET_B(net6046),
    .D(_02030_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[20] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _25454_ (.RESET_B(net6055),
    .D(_02031_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[21] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_1 _25455_ (.RESET_B(net6045),
    .D(_02032_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[22] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _25456_ (.RESET_B(net6052),
    .D(net1943),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[23] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_1 _25457_ (.RESET_B(net6037),
    .D(_02034_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[24] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _25458_ (.RESET_B(net6047),
    .D(_02035_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[25] ),
    .CLK(clknet_leaf_268_clk));
 sg13g2_dfrbpq_1 _25459_ (.RESET_B(net6051),
    .D(_02036_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[26] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _25460_ (.RESET_B(net6053),
    .D(net1502),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[27] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_1 _25461_ (.RESET_B(net6050),
    .D(_02038_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[28] ),
    .CLK(clknet_leaf_267_clk));
 sg13g2_dfrbpq_1 _25462_ (.RESET_B(net6051),
    .D(_02039_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[29] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _25463_ (.RESET_B(net6045),
    .D(_02040_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[30] ),
    .CLK(clknet_leaf_266_clk));
 sg13g2_dfrbpq_1 _25464_ (.RESET_B(net6032),
    .D(_02041_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[31] ),
    .CLK(clknet_leaf_270_clk));
 sg13g2_dfrbpq_2 _25465_ (.RESET_B(net5985),
    .D(_02042_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[0] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _25466_ (.RESET_B(net5984),
    .D(_02043_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[1] ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_2 _25467_ (.RESET_B(net6034),
    .D(_02044_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[2] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_2 _25468_ (.RESET_B(net5987),
    .D(net6081),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[3] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_2 _25469_ (.RESET_B(net5985),
    .D(_02046_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[4] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _25470_ (.RESET_B(net5987),
    .D(_02047_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[5] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_2 _25471_ (.RESET_B(net5982),
    .D(_02048_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[6] ),
    .CLK(clknet_leaf_301_clk));
 sg13g2_dfrbpq_2 _25472_ (.RESET_B(net5982),
    .D(_02049_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[7] ),
    .CLK(clknet_leaf_302_clk));
 sg13g2_dfrbpq_1 _25473_ (.RESET_B(net5987),
    .D(_02050_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[8] ),
    .CLK(clknet_leaf_300_clk));
 sg13g2_dfrbpq_2 _25474_ (.RESET_B(net6035),
    .D(net4015),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[9] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25475_ (.RESET_B(net6046),
    .D(_02052_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[10] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _25476_ (.RESET_B(net5988),
    .D(_02053_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[11] ),
    .CLK(clknet_leaf_304_clk));
 sg13g2_dfrbpq_2 _25477_ (.RESET_B(net6034),
    .D(_02054_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[12] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_2 _25478_ (.RESET_B(net6038),
    .D(net3951),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[13] ),
    .CLK(clknet_leaf_274_clk));
 sg13g2_dfrbpq_2 _25479_ (.RESET_B(net6038),
    .D(net6200),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[14] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_2 _25480_ (.RESET_B(net6038),
    .D(_02057_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[15] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_2 _25481_ (.RESET_B(net6039),
    .D(net4019),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[16] ),
    .CLK(clknet_leaf_273_clk));
 sg13g2_dfrbpq_2 _25482_ (.RESET_B(net6049),
    .D(net3942),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[17] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _25483_ (.RESET_B(net6039),
    .D(_02060_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[18] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _25484_ (.RESET_B(net6052),
    .D(_02061_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[19] ),
    .CLK(clknet_leaf_265_clk));
 sg13g2_dfrbpq_2 _25485_ (.RESET_B(net6048),
    .D(net3887),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[20] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _25486_ (.RESET_B(net6054),
    .D(_02063_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_2 _25487_ (.RESET_B(net6049),
    .D(net6107),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[22] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _25488_ (.RESET_B(net6054),
    .D(net6202),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[23] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _25489_ (.RESET_B(net6048),
    .D(net3844),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[24] ),
    .CLK(clknet_leaf_276_clk));
 sg13g2_dfrbpq_2 _25490_ (.RESET_B(net6048),
    .D(_02067_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[25] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _25491_ (.RESET_B(net6053),
    .D(_02068_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[26] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _25492_ (.RESET_B(net6053),
    .D(net2002),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[27] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _25493_ (.RESET_B(net6049),
    .D(_02070_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[28] ),
    .CLK(clknet_leaf_277_clk));
 sg13g2_dfrbpq_2 _25494_ (.RESET_B(net6053),
    .D(_02071_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[29] ),
    .CLK(clknet_leaf_278_clk));
 sg13g2_dfrbpq_2 _25495_ (.RESET_B(net6045),
    .D(net3740),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[30] ),
    .CLK(clknet_leaf_272_clk));
 sg13g2_dfrbpq_2 _25496_ (.RESET_B(net6036),
    .D(_02073_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[31] ),
    .CLK(clknet_leaf_269_clk));
 sg13g2_dfrbpq_1 _25497_ (.RESET_B(net5979),
    .D(_02074_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_sie ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_1 _25498_ (.RESET_B(net5984),
    .D(_02075_),
    .Q(\fpga_top.cpu_top.execution.csr_array.csr_spp ),
    .CLK(clknet_leaf_303_clk));
 sg13g2_dfrbpq_2 _25499_ (.RESET_B(net6020),
    .D(_00025_),
    .Q(\fpga_top.cmd_st_ma ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _25500_ (.RESET_B(net6020),
    .D(net6309),
    .Q(\fpga_top.cmd_ld_ma ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _25501_ (.RESET_B(net6026),
    .D(net3866),
    .Q(\fpga_top.cpu_top.data_rw_mem.wbk_rd_reg_ma ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _25502_ (.RESET_B(net6019),
    .D(net2303),
    .Q(\fpga_top.cpu_top.data_rw_mem.req_hw_dly ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _25503_ (.RESET_B(net6011),
    .D(_02077_),
    .Q(\fpga_top.cpu_top.data_rw_mem.req_w_dly ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _25504_ (.RESET_B(net6002),
    .D(\fpga_top.cpu_top.data_rw_mem.dma_io_radr_en ),
    .Q(\fpga_top.cpu_top.data_rw_mem.dma_io_ren_wb ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _25505_ (.RESET_B(net5955),
    .D(_02078_),
    .Q(\fpga_top.cpu_run_state ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _25506_ (.RESET_B(net6021),
    .D(\fpga_top.cpu_top.data_rw_mem.next_data_state[0] ),
    .Q(\fpga_top.cpu_top.data_rw_mem.data_state[0] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _25507_ (.RESET_B(net6021),
    .D(\fpga_top.cpu_top.data_rw_mem.next_data_state[1] ),
    .Q(\fpga_top.cpu_top.data_rw_mem.data_state[1] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _25508_ (.RESET_B(net6021),
    .D(net3935),
    .Q(\fpga_top.cpu_top.data_rw_mem.data_state[2] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _25509_ (.RESET_B(net5941),
    .D(net3080),
    .Q(\fpga_top.qspi_if.qspi_state[9] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _25510_ (.RESET_B(net5899),
    .D(_02080_),
    .Q(\fpga_top.io_frc.frc_cmp_val[0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _25511_ (.RESET_B(net5888),
    .D(_02081_),
    .Q(\fpga_top.io_frc.frc_cmp_val[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _25512_ (.RESET_B(net5888),
    .D(_02082_),
    .Q(\fpga_top.io_frc.frc_cmp_val[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _25513_ (.RESET_B(net5889),
    .D(_02083_),
    .Q(\fpga_top.io_frc.frc_cmp_val[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _25514_ (.RESET_B(net5888),
    .D(_02084_),
    .Q(\fpga_top.io_frc.frc_cmp_val[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _25515_ (.RESET_B(net5888),
    .D(_02085_),
    .Q(\fpga_top.io_frc.frc_cmp_val[5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _25516_ (.RESET_B(net5888),
    .D(_02086_),
    .Q(\fpga_top.io_frc.frc_cmp_val[6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _25517_ (.RESET_B(net5895),
    .D(_02087_),
    .Q(\fpga_top.io_frc.frc_cmp_val[7] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _25518_ (.RESET_B(net5894),
    .D(_02088_),
    .Q(\fpga_top.io_frc.frc_cmp_val[8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _25519_ (.RESET_B(net5894),
    .D(_02089_),
    .Q(\fpga_top.io_frc.frc_cmp_val[9] ),
    .CLK(clknet_leaf_319_clk));
 sg13g2_dfrbpq_1 _25520_ (.RESET_B(net5906),
    .D(_02090_),
    .Q(\fpga_top.io_frc.frc_cmp_val[10] ),
    .CLK(clknet_leaf_319_clk));
 sg13g2_dfrbpq_1 _25521_ (.RESET_B(net5915),
    .D(_02091_),
    .Q(\fpga_top.io_frc.frc_cmp_val[11] ),
    .CLK(clknet_leaf_318_clk));
 sg13g2_dfrbpq_2 _25522_ (.RESET_B(net5920),
    .D(_02092_),
    .Q(\fpga_top.io_frc.frc_cmp_val[12] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _25523_ (.RESET_B(net5916),
    .D(_02093_),
    .Q(\fpga_top.io_frc.frc_cmp_val[13] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _25524_ (.RESET_B(net5916),
    .D(_02094_),
    .Q(\fpga_top.io_frc.frc_cmp_val[14] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _25525_ (.RESET_B(net5942),
    .D(_02095_),
    .Q(\fpga_top.io_frc.frc_cmp_val[15] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _25526_ (.RESET_B(net5905),
    .D(_02096_),
    .Q(\fpga_top.io_frc.frc_cmp_val[16] ),
    .CLK(clknet_leaf_324_clk));
 sg13g2_dfrbpq_2 _25527_ (.RESET_B(net5906),
    .D(_02097_),
    .Q(\fpga_top.io_frc.frc_cmp_val[17] ),
    .CLK(clknet_leaf_323_clk));
 sg13g2_dfrbpq_2 _25528_ (.RESET_B(net5908),
    .D(_02098_),
    .Q(\fpga_top.io_frc.frc_cmp_val[18] ),
    .CLK(clknet_leaf_322_clk));
 sg13g2_dfrbpq_2 _25529_ (.RESET_B(net5906),
    .D(_02099_),
    .Q(\fpga_top.io_frc.frc_cmp_val[19] ),
    .CLK(clknet_leaf_322_clk));
 sg13g2_dfrbpq_2 _25530_ (.RESET_B(net5907),
    .D(_02100_),
    .Q(\fpga_top.io_frc.frc_cmp_val[20] ),
    .CLK(clknet_leaf_322_clk));
 sg13g2_dfrbpq_2 _25531_ (.RESET_B(net5914),
    .D(_02101_),
    .Q(\fpga_top.io_frc.frc_cmp_val[21] ),
    .CLK(clknet_leaf_317_clk));
 sg13g2_dfrbpq_2 _25532_ (.RESET_B(net5915),
    .D(_02102_),
    .Q(\fpga_top.io_frc.frc_cmp_val[22] ),
    .CLK(clknet_leaf_318_clk));
 sg13g2_dfrbpq_2 _25533_ (.RESET_B(net5915),
    .D(_02103_),
    .Q(\fpga_top.io_frc.frc_cmp_val[23] ),
    .CLK(clknet_leaf_319_clk));
 sg13g2_dfrbpq_1 _25534_ (.RESET_B(net5929),
    .D(_02104_),
    .Q(\fpga_top.io_frc.frc_cmp_val[24] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _25535_ (.RESET_B(net5943),
    .D(_02105_),
    .Q(\fpga_top.io_frc.frc_cmp_val[25] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _25536_ (.RESET_B(net5929),
    .D(_02106_),
    .Q(\fpga_top.io_frc.frc_cmp_val[26] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _25537_ (.RESET_B(net5944),
    .D(_02107_),
    .Q(\fpga_top.io_frc.frc_cmp_val[27] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _25538_ (.RESET_B(net5931),
    .D(_02108_),
    .Q(\fpga_top.io_frc.frc_cmp_val[28] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _25539_ (.RESET_B(net5943),
    .D(_02109_),
    .Q(\fpga_top.io_frc.frc_cmp_val[29] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _25540_ (.RESET_B(net5946),
    .D(_02110_),
    .Q(\fpga_top.io_frc.frc_cmp_val[30] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _25541_ (.RESET_B(net5928),
    .D(_02111_),
    .Q(\fpga_top.io_frc.frc_cmp_val[31] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _25542_ (.RESET_B(net5902),
    .D(_02112_),
    .Q(\fpga_top.io_frc.frc_cntr_val[32] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _25543_ (.RESET_B(net5902),
    .D(net2183),
    .Q(\fpga_top.io_frc.frc_cntr_val[33] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _25544_ (.RESET_B(net5902),
    .D(net3126),
    .Q(\fpga_top.io_frc.frc_cntr_val[34] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _25545_ (.RESET_B(net5902),
    .D(net3972),
    .Q(\fpga_top.io_frc.frc_cntr_val[35] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _25546_ (.RESET_B(net5902),
    .D(net2213),
    .Q(\fpga_top.io_frc.frc_cntr_val[36] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _25547_ (.RESET_B(net5901),
    .D(_02117_),
    .Q(\fpga_top.io_frc.frc_cntr_val[37] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _25548_ (.RESET_B(net5901),
    .D(net3450),
    .Q(\fpga_top.io_frc.frc_cntr_val[38] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _25549_ (.RESET_B(net5901),
    .D(_02119_),
    .Q(\fpga_top.io_frc.frc_cntr_val[39] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _25550_ (.RESET_B(net5895),
    .D(_02120_),
    .Q(\fpga_top.io_frc.frc_cntr_val[40] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _25551_ (.RESET_B(net5895),
    .D(net2075),
    .Q(\fpga_top.io_frc.frc_cntr_val[41] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _25552_ (.RESET_B(net5895),
    .D(net3710),
    .Q(\fpga_top.io_frc.frc_cntr_val[42] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _25553_ (.RESET_B(net5900),
    .D(net3114),
    .Q(\fpga_top.io_frc.frc_cntr_val[43] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _25554_ (.RESET_B(net5916),
    .D(net3619),
    .Q(\fpga_top.io_frc.frc_cntr_val[44] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _25555_ (.RESET_B(net5916),
    .D(_02125_),
    .Q(\fpga_top.io_frc.frc_cntr_val[45] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _25556_ (.RESET_B(net5916),
    .D(net2079),
    .Q(\fpga_top.io_frc.frc_cntr_val[46] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _25557_ (.RESET_B(net5945),
    .D(_02127_),
    .Q(\fpga_top.io_frc.frc_cntr_val[47] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _25558_ (.RESET_B(net5907),
    .D(_02128_),
    .Q(\fpga_top.io_frc.frc_cntr_val[48] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _25559_ (.RESET_B(net5907),
    .D(net3775),
    .Q(\fpga_top.io_frc.frc_cntr_val[49] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _25560_ (.RESET_B(net5906),
    .D(_02130_),
    .Q(\fpga_top.io_frc.frc_cntr_val[50] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _25561_ (.RESET_B(net5906),
    .D(_02131_),
    .Q(\fpga_top.io_frc.frc_cntr_val[51] ),
    .CLK(clknet_leaf_313_clk));
 sg13g2_dfrbpq_2 _25562_ (.RESET_B(net5907),
    .D(_02132_),
    .Q(\fpga_top.io_frc.frc_cntr_val[52] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_1 _25563_ (.RESET_B(net5907),
    .D(_02133_),
    .Q(\fpga_top.io_frc.frc_cntr_val[53] ),
    .CLK(clknet_leaf_314_clk));
 sg13g2_dfrbpq_2 _25564_ (.RESET_B(net5915),
    .D(_02134_),
    .Q(\fpga_top.io_frc.frc_cntr_val[54] ),
    .CLK(clknet_leaf_318_clk));
 sg13g2_dfrbpq_2 _25565_ (.RESET_B(net5917),
    .D(_02135_),
    .Q(\fpga_top.io_frc.frc_cntr_val[55] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _25566_ (.RESET_B(net5942),
    .D(_02136_),
    .Q(\fpga_top.io_frc.frc_cntr_val[56] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _25567_ (.RESET_B(net5942),
    .D(_02137_),
    .Q(\fpga_top.io_frc.frc_cntr_val[57] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _25568_ (.RESET_B(net5943),
    .D(_02138_),
    .Q(\fpga_top.io_frc.frc_cntr_val[58] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _25569_ (.RESET_B(net5945),
    .D(_02139_),
    .Q(\fpga_top.io_frc.frc_cntr_val[59] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _25570_ (.RESET_B(net5943),
    .D(net3924),
    .Q(\fpga_top.io_frc.frc_cntr_val[60] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _25571_ (.RESET_B(net5942),
    .D(_02141_),
    .Q(\fpga_top.io_frc.frc_cntr_val[61] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _25572_ (.RESET_B(net5928),
    .D(net3408),
    .Q(\fpga_top.io_frc.frc_cntr_val[62] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _25573_ (.RESET_B(net5942),
    .D(net2131),
    .Q(\fpga_top.io_frc.frc_cntr_val[63] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _25574_ (.RESET_B(net6005),
    .D(_02144_),
    .Q(\fpga_top.uart_top.uart_send_char.send_cntr[0] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _25575_ (.RESET_B(net6008),
    .D(net6509),
    .Q(\fpga_top.uart_top.uart_send_char.send_cntr[1] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _25576_ (.RESET_B(net6008),
    .D(net6298),
    .Q(\fpga_top.uart_top.uart_send_char.send_cntr[2] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _25577_ (.RESET_B(net6008),
    .D(net3999),
    .Q(\fpga_top.uart_top.uart_send_char.send_cntr[3] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _25578_ (.RESET_B(net6005),
    .D(_02148_),
    .Q(\fpga_top.uart_top.uart_send_char.send_cntr[4] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _25579_ (.RESET_B(net1233),
    .D(net1368),
    .Q(_00011_),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _25580_ (.RESET_B(net1297),
    .D(net1365),
    .Q(_00012_),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _25581_ (.RESET_B(net1002),
    .D(net1362),
    .Q(_00013_),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _25582_ (.RESET_B(net1001),
    .D(_02149_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _25583_ (.RESET_B(net1000),
    .D(_02150_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][1] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _25584_ (.RESET_B(net999),
    .D(_02151_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][2] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _25585_ (.RESET_B(net998),
    .D(_02152_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _25586_ (.RESET_B(net997),
    .D(net2299),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][4] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _25587_ (.RESET_B(net996),
    .D(_02154_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][5] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _25588_ (.RESET_B(net995),
    .D(_02155_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _25589_ (.RESET_B(net994),
    .D(_02156_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][7] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _25590_ (.RESET_B(net993),
    .D(_02157_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _25591_ (.RESET_B(net992),
    .D(_02158_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _25592_ (.RESET_B(net991),
    .D(_02159_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][2] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _25593_ (.RESET_B(net990),
    .D(_02160_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _25594_ (.RESET_B(net989),
    .D(net2453),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _25595_ (.RESET_B(net988),
    .D(_02162_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _25596_ (.RESET_B(net987),
    .D(_02163_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _25597_ (.RESET_B(net986),
    .D(_02164_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _25598_ (.RESET_B(net985),
    .D(net1823),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _25599_ (.RESET_B(net984),
    .D(net3545),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][1] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _25600_ (.RESET_B(net983),
    .D(_02167_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][2] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _25601_ (.RESET_B(net982),
    .D(net3179),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _25602_ (.RESET_B(net981),
    .D(net2952),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][4] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _25603_ (.RESET_B(net980),
    .D(_02170_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _25604_ (.RESET_B(net979),
    .D(_02171_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _25605_ (.RESET_B(net978),
    .D(_02172_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _25606_ (.RESET_B(net977),
    .D(net2022),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _25607_ (.RESET_B(net976),
    .D(net1831),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][1] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _25608_ (.RESET_B(net975),
    .D(_02175_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][2] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _25609_ (.RESET_B(net974),
    .D(net1854),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _25610_ (.RESET_B(net973),
    .D(_02177_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][4] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _25611_ (.RESET_B(net972),
    .D(_02178_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][5] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _25612_ (.RESET_B(net971),
    .D(_02179_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][6] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _25613_ (.RESET_B(net970),
    .D(_02180_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][7] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _25614_ (.RESET_B(net969),
    .D(_02181_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _25615_ (.RESET_B(net968),
    .D(_02182_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][1] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _25616_ (.RESET_B(net967),
    .D(net3761),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][2] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _25617_ (.RESET_B(net966),
    .D(_02184_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _25618_ (.RESET_B(net965),
    .D(_02185_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][4] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _25619_ (.RESET_B(net964),
    .D(_02186_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][5] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _25620_ (.RESET_B(net963),
    .D(_02187_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _25621_ (.RESET_B(net962),
    .D(net2428),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][7] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _25622_ (.RESET_B(net961),
    .D(_02189_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _25623_ (.RESET_B(net960),
    .D(_02190_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][1] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _25624_ (.RESET_B(net959),
    .D(_02191_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][2] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _25625_ (.RESET_B(net958),
    .D(net1739),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _25626_ (.RESET_B(net957),
    .D(_02193_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][4] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _25627_ (.RESET_B(net956),
    .D(net2073),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][5] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _25628_ (.RESET_B(net955),
    .D(_02195_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][6] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _25629_ (.RESET_B(net954),
    .D(net2984),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][7] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _25630_ (.RESET_B(net953),
    .D(_02197_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _25631_ (.RESET_B(net952),
    .D(_02198_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][1] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _25632_ (.RESET_B(net951),
    .D(_02199_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][2] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _25633_ (.RESET_B(net950),
    .D(_02200_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][3] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _25634_ (.RESET_B(net949),
    .D(_02201_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _25635_ (.RESET_B(net948),
    .D(_02202_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][5] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _25636_ (.RESET_B(net947),
    .D(_02203_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][6] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _25637_ (.RESET_B(net946),
    .D(_02204_),
    .Q(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][7] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _25638_ (.RESET_B(net945),
    .D(net2153),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][0] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _25639_ (.RESET_B(net944),
    .D(net2288),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][1] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _25640_ (.RESET_B(net943),
    .D(net2521),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][2] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _25641_ (.RESET_B(net942),
    .D(net2431),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][3] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _25642_ (.RESET_B(net941),
    .D(net2361),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][4] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _25643_ (.RESET_B(net940),
    .D(net2188),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _25644_ (.RESET_B(net939),
    .D(net2260),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][6] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _25645_ (.RESET_B(net938),
    .D(net2166),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][7] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _25646_ (.RESET_B(net5935),
    .D(_02213_),
    .Q(\fpga_top.io_uart_out.rout[0] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _25647_ (.RESET_B(net5935),
    .D(_02214_),
    .Q(\fpga_top.io_uart_out.rout[1] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _25648_ (.RESET_B(net5884),
    .D(_02215_),
    .Q(\fpga_top.io_uart_out.rout[2] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _25649_ (.RESET_B(net5935),
    .D(_02216_),
    .Q(\fpga_top.io_uart_out.rout[3] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _25650_ (.RESET_B(net5935),
    .D(_02217_),
    .Q(\fpga_top.io_uart_out.rout[4] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _25651_ (.RESET_B(net5935),
    .D(net4003),
    .Q(\fpga_top.io_uart_out.rout[5] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _25652_ (.RESET_B(net5883),
    .D(_02219_),
    .Q(\fpga_top.io_uart_out.rout[6] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _25653_ (.RESET_B(net5883),
    .D(_02220_),
    .Q(\fpga_top.io_uart_out.rout[7] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _25654_ (.RESET_B(net937),
    .D(net2668),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][0] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _25655_ (.RESET_B(net936),
    .D(net2805),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][1] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _25656_ (.RESET_B(net935),
    .D(net2775),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][2] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _25657_ (.RESET_B(net934),
    .D(net3344),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][3] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _25658_ (.RESET_B(net933),
    .D(net3448),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][4] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _25659_ (.RESET_B(net932),
    .D(net2906),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _25660_ (.RESET_B(net931),
    .D(net3196),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][6] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _25661_ (.RESET_B(net930),
    .D(net2537),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][7] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _25662_ (.RESET_B(net929),
    .D(net2121),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][0] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _25663_ (.RESET_B(net928),
    .D(net2281),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][1] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _25664_ (.RESET_B(net927),
    .D(net2204),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][2] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _25665_ (.RESET_B(net926),
    .D(net2250),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][3] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _25666_ (.RESET_B(net925),
    .D(net2149),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][4] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _25667_ (.RESET_B(net924),
    .D(net2108),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][5] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _25668_ (.RESET_B(net923),
    .D(net2134),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][6] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _25669_ (.RESET_B(net922),
    .D(net2574),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][7] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _25670_ (.RESET_B(net921),
    .D(net2697),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][0] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _25671_ (.RESET_B(net920),
    .D(net2976),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][1] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _25672_ (.RESET_B(net919),
    .D(net2741),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][2] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _25673_ (.RESET_B(net918),
    .D(net2962),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][3] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _25674_ (.RESET_B(net917),
    .D(net2551),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][4] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _25675_ (.RESET_B(net916),
    .D(net2591),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][5] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _25676_ (.RESET_B(net915),
    .D(net2820),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][6] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _25677_ (.RESET_B(net914),
    .D(net3163),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][7] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _25678_ (.RESET_B(net913),
    .D(net3557),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][0] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _25679_ (.RESET_B(net912),
    .D(net3586),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][1] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _25680_ (.RESET_B(net911),
    .D(net2627),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][2] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _25681_ (.RESET_B(net910),
    .D(net2946),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][3] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _25682_ (.RESET_B(net909),
    .D(net2756),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][4] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _25683_ (.RESET_B(net908),
    .D(net2295),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][5] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _25684_ (.RESET_B(net907),
    .D(net2531),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _25685_ (.RESET_B(net906),
    .D(net2547),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][7] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _25686_ (.RESET_B(net905),
    .D(net3622),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][0] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _25687_ (.RESET_B(net904),
    .D(net3282),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][1] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _25688_ (.RESET_B(net903),
    .D(net3071),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][2] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _25689_ (.RESET_B(net902),
    .D(net2234),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][3] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _25690_ (.RESET_B(net901),
    .D(net2164),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][4] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _25691_ (.RESET_B(net900),
    .D(net3018),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _25692_ (.RESET_B(net899),
    .D(net3265),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _25693_ (.RESET_B(net898),
    .D(net2580),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][7] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _25694_ (.RESET_B(net897),
    .D(net3499),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][0] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _25695_ (.RESET_B(net896),
    .D(net2451),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][1] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _25696_ (.RESET_B(net895),
    .D(net2457),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][2] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _25697_ (.RESET_B(net894),
    .D(net2801),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][3] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _25698_ (.RESET_B(net893),
    .D(net3311),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][4] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _25699_ (.RESET_B(net892),
    .D(net3508),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][5] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _25700_ (.RESET_B(net891),
    .D(_02267_),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _25701_ (.RESET_B(net890),
    .D(_02268_),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][7] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _25702_ (.RESET_B(net889),
    .D(net2567),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][0] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _25703_ (.RESET_B(net888),
    .D(net2919),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][1] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _25704_ (.RESET_B(net887),
    .D(net2339),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][2] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _25705_ (.RESET_B(net886),
    .D(net3309),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][3] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _25706_ (.RESET_B(net885),
    .D(net3041),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][4] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _25707_ (.RESET_B(net884),
    .D(net2175),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][5] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _25708_ (.RESET_B(net883),
    .D(net3671),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _25709_ (.RESET_B(net882),
    .D(net3632),
    .Q(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][7] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _25710_ (.RESET_B(net881),
    .D(net1488),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _25711_ (.RESET_B(net880),
    .D(net1559),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _25712_ (.RESET_B(net879),
    .D(_02279_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25713_ (.RESET_B(net878),
    .D(_02280_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25714_ (.RESET_B(net877),
    .D(net3252),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _25715_ (.RESET_B(net876),
    .D(net1421),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _25716_ (.RESET_B(net875),
    .D(net1461),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _25717_ (.RESET_B(net1298),
    .D(net1449),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][7] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _25718_ (.RESET_B(net1299),
    .D(net1893),
    .Q(_00008_),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _25719_ (.RESET_B(net1310),
    .D(\fpga_top.io_spi_lite.mosi_fifo.radr_early[1] ),
    .Q(_00009_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _25720_ (.RESET_B(net874),
    .D(net1573),
    .Q(_00010_),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _25721_ (.RESET_B(net873),
    .D(net2058),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _25722_ (.RESET_B(net872),
    .D(net1746),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _25723_ (.RESET_B(net871),
    .D(net2353),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25724_ (.RESET_B(net870),
    .D(_02288_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25725_ (.RESET_B(net869),
    .D(net2247),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _25726_ (.RESET_B(net868),
    .D(net1891),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _25727_ (.RESET_B(net867),
    .D(net2031),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _25728_ (.RESET_B(net866),
    .D(net2158),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][7] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _25729_ (.RESET_B(net865),
    .D(_02293_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _25730_ (.RESET_B(net864),
    .D(net1908),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][1] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _25731_ (.RESET_B(net863),
    .D(_02295_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25732_ (.RESET_B(net862),
    .D(_02296_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25733_ (.RESET_B(net861),
    .D(_02297_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _25734_ (.RESET_B(net860),
    .D(_02298_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _25735_ (.RESET_B(net859),
    .D(_02299_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _25736_ (.RESET_B(net858),
    .D(_02300_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][7] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _25737_ (.RESET_B(net857),
    .D(_02301_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _25738_ (.RESET_B(net856),
    .D(_02302_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _25739_ (.RESET_B(net855),
    .D(_02303_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25740_ (.RESET_B(net854),
    .D(_02304_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _25741_ (.RESET_B(net853),
    .D(_02305_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _25742_ (.RESET_B(net852),
    .D(_02306_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _25743_ (.RESET_B(net851),
    .D(_02307_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _25744_ (.RESET_B(net850),
    .D(_02308_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _25745_ (.RESET_B(net849),
    .D(net1426),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25746_ (.RESET_B(net848),
    .D(net1454),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _25747_ (.RESET_B(net847),
    .D(net1523),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25748_ (.RESET_B(net846),
    .D(_02312_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25749_ (.RESET_B(net845),
    .D(_02313_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _25750_ (.RESET_B(net844),
    .D(net1471),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _25751_ (.RESET_B(net843),
    .D(net1481),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][6] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _25752_ (.RESET_B(net842),
    .D(net1459),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _25753_ (.RESET_B(net841),
    .D(net1922),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25754_ (.RESET_B(net840),
    .D(net1749),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25755_ (.RESET_B(net839),
    .D(net1767),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25756_ (.RESET_B(net838),
    .D(_02320_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25757_ (.RESET_B(net837),
    .D(net2297),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _25758_ (.RESET_B(net836),
    .D(net1800),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25759_ (.RESET_B(net835),
    .D(net1829),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _25760_ (.RESET_B(net834),
    .D(net1654),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _25761_ (.RESET_B(net833),
    .D(_02325_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25762_ (.RESET_B(net832),
    .D(_02326_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _25763_ (.RESET_B(net831),
    .D(_02327_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25764_ (.RESET_B(net830),
    .D(_02328_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25765_ (.RESET_B(net829),
    .D(_02329_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _25766_ (.RESET_B(net828),
    .D(_02330_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _25767_ (.RESET_B(net827),
    .D(_02331_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _25768_ (.RESET_B(net826),
    .D(_02332_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _25769_ (.RESET_B(net825),
    .D(_02333_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25770_ (.RESET_B(net824),
    .D(_02334_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _25771_ (.RESET_B(net823),
    .D(_02335_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _25772_ (.RESET_B(net822),
    .D(_02336_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25773_ (.RESET_B(net821),
    .D(_02337_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _25774_ (.RESET_B(net820),
    .D(_02338_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _25775_ (.RESET_B(net819),
    .D(_02339_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _25776_ (.RESET_B(net818),
    .D(_02340_),
    .Q(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _25777_ (.RESET_B(net817),
    .D(net1565),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][0] ),
    .CLK(clknet_leaf_329_clk));
 sg13g2_dfrbpq_1 _25778_ (.RESET_B(net816),
    .D(net1527),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][1] ),
    .CLK(clknet_leaf_326_clk));
 sg13g2_dfrbpq_1 _25779_ (.RESET_B(net815),
    .D(net1399),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][2] ),
    .CLK(clknet_leaf_330_clk));
 sg13g2_dfrbpq_1 _25780_ (.RESET_B(net814),
    .D(net1484),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][3] ),
    .CLK(clknet_leaf_329_clk));
 sg13g2_dfrbpq_1 _25781_ (.RESET_B(net813),
    .D(net1414),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][4] ),
    .CLK(clknet_leaf_328_clk));
 sg13g2_dfrbpq_1 _25782_ (.RESET_B(net812),
    .D(net1435),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _25783_ (.RESET_B(net811),
    .D(net1423),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][6] ),
    .CLK(clknet_leaf_330_clk));
 sg13g2_dfrbpq_1 _25784_ (.RESET_B(net1311),
    .D(net1494),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _25785_ (.RESET_B(net1312),
    .D(net1862),
    .Q(_00005_),
    .CLK(clknet_leaf_326_clk));
 sg13g2_dfrbpq_2 _25786_ (.RESET_B(net1300),
    .D(\fpga_top.io_spi_lite.miso_fifo.radr_early[1] ),
    .Q(_00006_),
    .CLK(clknet_leaf_325_clk));
 sg13g2_dfrbpq_2 _25787_ (.RESET_B(net810),
    .D(net1992),
    .Q(_00007_),
    .CLK(clknet_leaf_325_clk));
 sg13g2_dfrbpq_1 _25788_ (.RESET_B(net809),
    .D(net1926),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][0] ),
    .CLK(clknet_leaf_329_clk));
 sg13g2_dfrbpq_1 _25789_ (.RESET_B(net808),
    .D(net2061),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][1] ),
    .CLK(clknet_leaf_326_clk));
 sg13g2_dfrbpq_1 _25790_ (.RESET_B(net807),
    .D(net1755),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][2] ),
    .CLK(clknet_leaf_330_clk));
 sg13g2_dfrbpq_1 _25791_ (.RESET_B(net806),
    .D(net2046),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][3] ),
    .CLK(clknet_leaf_328_clk));
 sg13g2_dfrbpq_1 _25792_ (.RESET_B(net805),
    .D(net1666),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][4] ),
    .CLK(clknet_leaf_328_clk));
 sg13g2_dfrbpq_1 _25793_ (.RESET_B(net804),
    .D(net1628),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _25794_ (.RESET_B(net803),
    .D(net1883),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][6] ),
    .CLK(clknet_leaf_330_clk));
 sg13g2_dfrbpq_1 _25795_ (.RESET_B(net802),
    .D(net1913),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _25796_ (.RESET_B(net801),
    .D(net2479),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][0] ),
    .CLK(clknet_leaf_329_clk));
 sg13g2_dfrbpq_1 _25797_ (.RESET_B(net800),
    .D(net1967),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][1] ),
    .CLK(clknet_leaf_326_clk));
 sg13g2_dfrbpq_1 _25798_ (.RESET_B(net799),
    .D(net2094),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][2] ),
    .CLK(clknet_leaf_331_clk));
 sg13g2_dfrbpq_1 _25799_ (.RESET_B(net798),
    .D(net1896),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][3] ),
    .CLK(clknet_leaf_329_clk));
 sg13g2_dfrbpq_1 _25800_ (.RESET_B(net797),
    .D(net1771),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][4] ),
    .CLK(clknet_leaf_329_clk));
 sg13g2_dfrbpq_1 _25801_ (.RESET_B(net796),
    .D(net2053),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][5] ),
    .CLK(clknet_leaf_331_clk));
 sg13g2_dfrbpq_1 _25802_ (.RESET_B(net795),
    .D(net1886),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][6] ),
    .CLK(clknet_leaf_330_clk));
 sg13g2_dfrbpq_1 _25803_ (.RESET_B(net794),
    .D(net1806),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _25804_ (.RESET_B(net793),
    .D(net1917),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][0] ),
    .CLK(clknet_leaf_329_clk));
 sg13g2_dfrbpq_1 _25805_ (.RESET_B(net792),
    .D(net1877),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][1] ),
    .CLK(clknet_leaf_326_clk));
 sg13g2_dfrbpq_1 _25806_ (.RESET_B(net791),
    .D(net2151),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][2] ),
    .CLK(clknet_leaf_330_clk));
 sg13g2_dfrbpq_1 _25807_ (.RESET_B(net790),
    .D(net1638),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][3] ),
    .CLK(clknet_leaf_328_clk));
 sg13g2_dfrbpq_1 _25808_ (.RESET_B(net789),
    .D(net2013),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][4] ),
    .CLK(clknet_leaf_328_clk));
 sg13g2_dfrbpq_1 _25809_ (.RESET_B(net788),
    .D(net1650),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _25810_ (.RESET_B(net787),
    .D(net1735),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][6] ),
    .CLK(clknet_leaf_330_clk));
 sg13g2_dfrbpq_1 _25811_ (.RESET_B(net786),
    .D(net1672),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _25812_ (.RESET_B(net785),
    .D(net1731),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][0] ),
    .CLK(clknet_leaf_329_clk));
 sg13g2_dfrbpq_1 _25813_ (.RESET_B(net784),
    .D(net1609),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][1] ),
    .CLK(clknet_leaf_328_clk));
 sg13g2_dfrbpq_1 _25814_ (.RESET_B(net783),
    .D(net1953),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][2] ),
    .CLK(clknet_leaf_331_clk));
 sg13g2_dfrbpq_1 _25815_ (.RESET_B(net782),
    .D(net1675),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][3] ),
    .CLK(clknet_leaf_328_clk));
 sg13g2_dfrbpq_1 _25816_ (.RESET_B(net781),
    .D(net2018),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][4] ),
    .CLK(clknet_leaf_326_clk));
 sg13g2_dfrbpq_1 _25817_ (.RESET_B(net780),
    .D(net2037),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _25818_ (.RESET_B(net779),
    .D(net1791),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][6] ),
    .CLK(clknet_leaf_331_clk));
 sg13g2_dfrbpq_1 _25819_ (.RESET_B(net778),
    .D(net1762),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _25820_ (.RESET_B(net777),
    .D(net1664),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][0] ),
    .CLK(clknet_leaf_328_clk));
 sg13g2_dfrbpq_1 _25821_ (.RESET_B(net776),
    .D(net1722),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][1] ),
    .CLK(clknet_leaf_327_clk));
 sg13g2_dfrbpq_1 _25822_ (.RESET_B(net775),
    .D(net1776),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _25823_ (.RESET_B(net774),
    .D(net1710),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][3] ),
    .CLK(clknet_leaf_327_clk));
 sg13g2_dfrbpq_1 _25824_ (.RESET_B(net773),
    .D(net2526),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][4] ),
    .CLK(clknet_leaf_327_clk));
 sg13g2_dfrbpq_1 _25825_ (.RESET_B(net772),
    .D(net1872),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _25826_ (.RESET_B(net771),
    .D(net1702),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][6] ),
    .CLK(clknet_leaf_331_clk));
 sg13g2_dfrbpq_1 _25827_ (.RESET_B(net770),
    .D(net1774),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _25828_ (.RESET_B(net769),
    .D(net1963),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _25829_ (.RESET_B(net768),
    .D(net1727),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][1] ),
    .CLK(clknet_leaf_327_clk));
 sg13g2_dfrbpq_1 _25830_ (.RESET_B(net767),
    .D(net2035),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][2] ),
    .CLK(clknet_leaf_331_clk));
 sg13g2_dfrbpq_1 _25831_ (.RESET_B(net766),
    .D(net1850),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][3] ),
    .CLK(clknet_leaf_327_clk));
 sg13g2_dfrbpq_1 _25832_ (.RESET_B(net765),
    .D(net2194),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][4] ),
    .CLK(clknet_leaf_326_clk));
 sg13g2_dfrbpq_1 _25833_ (.RESET_B(net764),
    .D(net1691),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _25834_ (.RESET_B(net763),
    .D(net1816),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][6] ),
    .CLK(clknet_leaf_330_clk));
 sg13g2_dfrbpq_1 _25835_ (.RESET_B(net762),
    .D(net1635),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _25836_ (.RESET_B(net761),
    .D(net1619),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _25837_ (.RESET_B(net760),
    .D(net1698),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][1] ),
    .CLK(clknet_leaf_327_clk));
 sg13g2_dfrbpq_1 _25838_ (.RESET_B(net759),
    .D(net1764),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _25839_ (.RESET_B(net758),
    .D(net1760),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][3] ),
    .CLK(clknet_leaf_327_clk));
 sg13g2_dfrbpq_1 _25840_ (.RESET_B(net757),
    .D(net1842),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][4] ),
    .CLK(clknet_leaf_327_clk));
 sg13g2_dfrbpq_1 _25841_ (.RESET_B(net756),
    .D(net1714),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _25842_ (.RESET_B(net755),
    .D(net1751),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][6] ),
    .CLK(clknet_leaf_331_clk));
 sg13g2_dfrbpq_1 _25843_ (.RESET_B(net754),
    .D(net1645),
    .Q(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _25844_ (.RESET_B(net753),
    .D(_02405_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][0] ),
    .CLK(clknet_leaf_279_clk));
 sg13g2_dfrbpq_1 _25845_ (.RESET_B(net752),
    .D(_02406_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][1] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _25846_ (.RESET_B(net751),
    .D(_02407_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][2] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _25847_ (.RESET_B(net750),
    .D(_02408_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][3] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _25848_ (.RESET_B(net749),
    .D(_02409_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][4] ),
    .CLK(clknet_leaf_245_clk));
 sg13g2_dfrbpq_1 _25849_ (.RESET_B(net748),
    .D(_02410_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][5] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25850_ (.RESET_B(net747),
    .D(_02411_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][6] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _25851_ (.RESET_B(net746),
    .D(_02412_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][7] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _25852_ (.RESET_B(net745),
    .D(_02413_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][8] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_1 _25853_ (.RESET_B(net744),
    .D(_02414_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][9] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _25854_ (.RESET_B(net743),
    .D(_02415_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][10] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _25855_ (.RESET_B(net742),
    .D(_02416_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][11] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _25856_ (.RESET_B(net741),
    .D(_02417_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][12] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _25857_ (.RESET_B(net740),
    .D(_02418_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][13] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_1 _25858_ (.RESET_B(net739),
    .D(_02419_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][14] ),
    .CLK(clknet_leaf_260_clk));
 sg13g2_dfrbpq_1 _25859_ (.RESET_B(net738),
    .D(_02420_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][15] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _25860_ (.RESET_B(net737),
    .D(_02421_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][16] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25861_ (.RESET_B(net736),
    .D(_02422_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][17] ),
    .CLK(clknet_leaf_264_clk));
 sg13g2_dfrbpq_1 _25862_ (.RESET_B(net735),
    .D(_02423_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][18] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _25863_ (.RESET_B(net734),
    .D(_02424_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][19] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _25864_ (.RESET_B(net733),
    .D(_02425_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][20] ),
    .CLK(clknet_leaf_248_clk));
 sg13g2_dfrbpq_1 _25865_ (.RESET_B(net732),
    .D(_02426_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][21] ),
    .CLK(clknet_leaf_256_clk));
 sg13g2_dfrbpq_1 _25866_ (.RESET_B(net731),
    .D(_02427_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][22] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _25867_ (.RESET_B(net730),
    .D(_02428_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][23] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _25868_ (.RESET_B(net729),
    .D(_02429_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][24] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _25869_ (.RESET_B(net728),
    .D(_02430_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][25] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_1 _25870_ (.RESET_B(net727),
    .D(_02431_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][26] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _25871_ (.RESET_B(net726),
    .D(_02432_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][27] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _25872_ (.RESET_B(net725),
    .D(_02433_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][28] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_1 _25873_ (.RESET_B(net724),
    .D(_02434_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][29] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _25874_ (.RESET_B(net723),
    .D(_02435_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][30] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _25875_ (.RESET_B(net722),
    .D(_02436_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][31] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _25876_ (.RESET_B(net5896),
    .D(_02437_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[0] ),
    .CLK(clknet_leaf_320_clk));
 sg13g2_dfrbpq_2 _25877_ (.RESET_B(net5887),
    .D(_02438_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[1] ),
    .CLK(clknet_leaf_321_clk));
 sg13g2_dfrbpq_2 _25878_ (.RESET_B(net5891),
    .D(_02439_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[2] ),
    .CLK(clknet_leaf_320_clk));
 sg13g2_dfrbpq_2 _25879_ (.RESET_B(net5887),
    .D(_02440_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[3] ),
    .CLK(clknet_leaf_321_clk));
 sg13g2_dfrbpq_2 _25880_ (.RESET_B(net5893),
    .D(_02441_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[4] ),
    .CLK(clknet_leaf_322_clk));
 sg13g2_dfrbpq_2 _25881_ (.RESET_B(net5893),
    .D(_02442_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[5] ),
    .CLK(clknet_leaf_321_clk));
 sg13g2_dfrbpq_2 _25882_ (.RESET_B(net5893),
    .D(_02443_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[6] ),
    .CLK(clknet_leaf_321_clk));
 sg13g2_dfrbpq_2 _25883_ (.RESET_B(net5893),
    .D(_02444_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[7] ),
    .CLK(clknet_leaf_321_clk));
 sg13g2_dfrbpq_1 _25884_ (.RESET_B(net5893),
    .D(_02445_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[8] ),
    .CLK(clknet_leaf_322_clk));
 sg13g2_dfrbpq_1 _25885_ (.RESET_B(net5893),
    .D(_02446_),
    .Q(\fpga_top.io_spi_lite.spi_sck_div[9] ),
    .CLK(clknet_leaf_321_clk));
 sg13g2_dfrbpq_2 _25886_ (.RESET_B(net5887),
    .D(_02447_),
    .Q(\fpga_top.io_spi_lite.org_sck ),
    .CLK(clknet_leaf_320_clk));
 sg13g2_dfrbpq_1 _25887_ (.RESET_B(net721),
    .D(_02448_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][0] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25888_ (.RESET_B(net720),
    .D(_02449_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][1] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25889_ (.RESET_B(net719),
    .D(_02450_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][2] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25890_ (.RESET_B(net718),
    .D(_02451_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][3] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _25891_ (.RESET_B(net717),
    .D(_02452_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][4] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25892_ (.RESET_B(net716),
    .D(_02453_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][5] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25893_ (.RESET_B(net715),
    .D(_02454_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][6] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _25894_ (.RESET_B(net714),
    .D(_02455_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][7] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25895_ (.RESET_B(net713),
    .D(_02456_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][8] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25896_ (.RESET_B(net712),
    .D(_02457_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][9] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25897_ (.RESET_B(net711),
    .D(_02458_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][10] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _25898_ (.RESET_B(net710),
    .D(_02459_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][11] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25899_ (.RESET_B(net709),
    .D(_02460_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][12] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25900_ (.RESET_B(net708),
    .D(_02461_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][13] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25901_ (.RESET_B(net707),
    .D(_02462_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][14] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _25902_ (.RESET_B(net706),
    .D(_02463_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][15] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25903_ (.RESET_B(net705),
    .D(_02464_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][16] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25904_ (.RESET_B(net704),
    .D(_02465_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][17] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25905_ (.RESET_B(net703),
    .D(_02466_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][18] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _25906_ (.RESET_B(net702),
    .D(_02467_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][19] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _25907_ (.RESET_B(net701),
    .D(_02468_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _25908_ (.RESET_B(net700),
    .D(_02469_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][21] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _25909_ (.RESET_B(net698),
    .D(_02470_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][22] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_1 _25910_ (.RESET_B(net627),
    .D(_02471_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][23] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25911_ (.RESET_B(net626),
    .D(_02472_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][24] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _25912_ (.RESET_B(net110),
    .D(_02473_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][25] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25913_ (.RESET_B(net109),
    .D(_02474_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][26] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25914_ (.RESET_B(net108),
    .D(_02475_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][27] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25915_ (.RESET_B(net107),
    .D(_02476_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][28] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_1 _25916_ (.RESET_B(net106),
    .D(_02477_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][29] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25917_ (.RESET_B(net105),
    .D(_02478_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][30] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _25918_ (.RESET_B(net104),
    .D(_02479_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][31] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25919_ (.RESET_B(net103),
    .D(_02480_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][0] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_1 _25920_ (.RESET_B(net102),
    .D(_02481_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][1] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_1 _25921_ (.RESET_B(net101),
    .D(_02482_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][2] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _25922_ (.RESET_B(net100),
    .D(_02483_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][3] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _25923_ (.RESET_B(net99),
    .D(_02484_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][4] ),
    .CLK(clknet_leaf_243_clk));
 sg13g2_dfrbpq_1 _25924_ (.RESET_B(net98),
    .D(_02485_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][5] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _25925_ (.RESET_B(net97),
    .D(_02486_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][6] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_1 _25926_ (.RESET_B(net96),
    .D(_02487_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][7] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _25927_ (.RESET_B(net95),
    .D(_02488_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][8] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_1 _25928_ (.RESET_B(net94),
    .D(_02489_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][9] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _25929_ (.RESET_B(net93),
    .D(_02490_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][10] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _25930_ (.RESET_B(net92),
    .D(_02491_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][11] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _25931_ (.RESET_B(net91),
    .D(_02492_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][12] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _25932_ (.RESET_B(net90),
    .D(_02493_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][13] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _25933_ (.RESET_B(net89),
    .D(_02494_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][14] ),
    .CLK(clknet_leaf_262_clk));
 sg13g2_dfrbpq_1 _25934_ (.RESET_B(net88),
    .D(_02495_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][15] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _25935_ (.RESET_B(net87),
    .D(_02496_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][16] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _25936_ (.RESET_B(net86),
    .D(_02497_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][17] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_1 _25937_ (.RESET_B(net85),
    .D(_02498_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][18] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25938_ (.RESET_B(net84),
    .D(_02499_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][19] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _25939_ (.RESET_B(net83),
    .D(_02500_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][20] ),
    .CLK(clknet_leaf_244_clk));
 sg13g2_dfrbpq_1 _25940_ (.RESET_B(net82),
    .D(_02501_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][21] ),
    .CLK(clknet_leaf_257_clk));
 sg13g2_dfrbpq_1 _25941_ (.RESET_B(net81),
    .D(_02502_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][22] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_1 _25942_ (.RESET_B(net80),
    .D(_02503_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][23] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _25943_ (.RESET_B(net79),
    .D(_02504_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][24] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _25944_ (.RESET_B(net78),
    .D(_02505_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][25] ),
    .CLK(clknet_leaf_242_clk));
 sg13g2_dfrbpq_1 _25945_ (.RESET_B(net77),
    .D(_02506_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][26] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _25946_ (.RESET_B(net76),
    .D(_02507_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][27] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_1 _25947_ (.RESET_B(net75),
    .D(_02508_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][28] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_1 _25948_ (.RESET_B(net74),
    .D(_02509_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][29] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _25949_ (.RESET_B(net73),
    .D(_02510_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][30] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_1 _25950_ (.RESET_B(net72),
    .D(_02511_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][31] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_1 _25951_ (.RESET_B(net71),
    .D(_02512_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][0] ),
    .CLK(clknet_leaf_281_clk));
 sg13g2_dfrbpq_1 _25952_ (.RESET_B(net70),
    .D(_02513_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][1] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _25953_ (.RESET_B(net69),
    .D(_02514_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][2] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _25954_ (.RESET_B(net68),
    .D(_02515_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][3] ),
    .CLK(clknet_leaf_250_clk));
 sg13g2_dfrbpq_1 _25955_ (.RESET_B(net67),
    .D(_02516_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][4] ),
    .CLK(clknet_leaf_246_clk));
 sg13g2_dfrbpq_1 _25956_ (.RESET_B(net66),
    .D(_02517_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][5] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_1 _25957_ (.RESET_B(net65),
    .D(_02518_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][6] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _25958_ (.RESET_B(net64),
    .D(_02519_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][7] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _25959_ (.RESET_B(net63),
    .D(_02520_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][8] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _25960_ (.RESET_B(net62),
    .D(_02521_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][9] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_1 _25961_ (.RESET_B(net61),
    .D(_02522_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][10] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _25962_ (.RESET_B(net60),
    .D(_02523_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][11] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _25963_ (.RESET_B(net59),
    .D(_02524_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][12] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _25964_ (.RESET_B(net58),
    .D(_02525_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][13] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _25965_ (.RESET_B(net56),
    .D(_02526_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][14] ),
    .CLK(clknet_leaf_259_clk));
 sg13g2_dfrbpq_1 _25966_ (.RESET_B(net55),
    .D(_02527_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][15] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_1 _25967_ (.RESET_B(net54),
    .D(_02528_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][16] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _25968_ (.RESET_B(net53),
    .D(_02529_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][17] ),
    .CLK(clknet_leaf_261_clk));
 sg13g2_dfrbpq_1 _25969_ (.RESET_B(net52),
    .D(_02530_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][18] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _25970_ (.RESET_B(net51),
    .D(_02531_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][19] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _25971_ (.RESET_B(net50),
    .D(_02532_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][20] ),
    .CLK(clknet_leaf_252_clk));
 sg13g2_dfrbpq_1 _25972_ (.RESET_B(net48),
    .D(_02533_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][21] ),
    .CLK(clknet_leaf_251_clk));
 sg13g2_dfrbpq_1 _25973_ (.RESET_B(net1313),
    .D(_02534_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][22] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _25974_ (.RESET_B(net1301),
    .D(_02535_),
    .Q(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][23] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_tiehi _24581__18 (.L_HI(net18));
 sg13g2_tiehi _24580__19 (.L_HI(net19));
 sg13g2_tiehi _24579__20 (.L_HI(net20));
 sg13g2_tiehi _24578__21 (.L_HI(net21));
 sg13g2_tiehi _24577__22 (.L_HI(net22));
 sg13g2_tiehi _24576__23 (.L_HI(net23));
 sg13g2_tiehi _24575__24 (.L_HI(net24));
 sg13g2_tiehi _24574__25 (.L_HI(net25));
 sg13g2_tiehi _24573__26 (.L_HI(net26));
 sg13g2_tiehi _24572__27 (.L_HI(net27));
 sg13g2_tiehi _24571__28 (.L_HI(net28));
 sg13g2_tiehi _24570__29 (.L_HI(net29));
 sg13g2_tiehi _24569__30 (.L_HI(net30));
 sg13g2_tiehi _24568__31 (.L_HI(net31));
 sg13g2_tiehi _24567__32 (.L_HI(net32));
 sg13g2_tiehi _24566__33 (.L_HI(net33));
 sg13g2_tiehi _24565__34 (.L_HI(net34));
 sg13g2_tiehi _24564__35 (.L_HI(net35));
 sg13g2_tiehi _24563__36 (.L_HI(net36));
 sg13g2_tiehi _24562__37 (.L_HI(net37));
 sg13g2_tiehi _24561__38 (.L_HI(net38));
 sg13g2_tiehi _24560__39 (.L_HI(net39));
 sg13g2_tiehi _24559__40 (.L_HI(net40));
 sg13g2_tiehi _24558__41 (.L_HI(net41));
 sg13g2_tiehi _24557__42 (.L_HI(net42));
 sg13g2_tiehi _24556__43 (.L_HI(net43));
 sg13g2_tiehi _24555__44 (.L_HI(net44));
 sg13g2_tiehi _24554__45 (.L_HI(net45));
 sg13g2_tiehi _24553__46 (.L_HI(net46));
 sg13g2_tiehi _24552__47 (.L_HI(net47));
 sg13g2_tiehi _25972__48 (.L_HI(net48));
 sg13g2_tiehi _23331__49 (.L_HI(net49));
 sg13g2_tiehi _25971__50 (.L_HI(net50));
 sg13g2_tiehi _25970__51 (.L_HI(net51));
 sg13g2_tiehi _25969__52 (.L_HI(net52));
 sg13g2_tiehi _25968__53 (.L_HI(net53));
 sg13g2_tiehi _25967__54 (.L_HI(net54));
 sg13g2_tiehi _25966__55 (.L_HI(net55));
 sg13g2_tiehi _25965__56 (.L_HI(net56));
 sg13g2_tiehi _23475__57 (.L_HI(net57));
 sg13g2_tiehi _25964__58 (.L_HI(net58));
 sg13g2_tiehi _25963__59 (.L_HI(net59));
 sg13g2_tiehi _25962__60 (.L_HI(net60));
 sg13g2_tiehi _25961__61 (.L_HI(net61));
 sg13g2_tiehi _25960__62 (.L_HI(net62));
 sg13g2_tiehi _25959__63 (.L_HI(net63));
 sg13g2_tiehi _25958__64 (.L_HI(net64));
 sg13g2_tiehi _25957__65 (.L_HI(net65));
 sg13g2_tiehi _25956__66 (.L_HI(net66));
 sg13g2_tiehi _25955__67 (.L_HI(net67));
 sg13g2_tiehi _25954__68 (.L_HI(net68));
 sg13g2_tiehi _25953__69 (.L_HI(net69));
 sg13g2_tiehi _25952__70 (.L_HI(net70));
 sg13g2_tiehi _25951__71 (.L_HI(net71));
 sg13g2_tiehi _25950__72 (.L_HI(net72));
 sg13g2_tiehi _25949__73 (.L_HI(net73));
 sg13g2_tiehi _25948__74 (.L_HI(net74));
 sg13g2_tiehi _25947__75 (.L_HI(net75));
 sg13g2_tiehi _25946__76 (.L_HI(net76));
 sg13g2_tiehi _25945__77 (.L_HI(net77));
 sg13g2_tiehi _25944__78 (.L_HI(net78));
 sg13g2_tiehi _25943__79 (.L_HI(net79));
 sg13g2_tiehi _25942__80 (.L_HI(net80));
 sg13g2_tiehi _25941__81 (.L_HI(net81));
 sg13g2_tiehi _25940__82 (.L_HI(net82));
 sg13g2_tiehi _25939__83 (.L_HI(net83));
 sg13g2_tiehi _25938__84 (.L_HI(net84));
 sg13g2_tiehi _25937__85 (.L_HI(net85));
 sg13g2_tiehi _25936__86 (.L_HI(net86));
 sg13g2_tiehi _25935__87 (.L_HI(net87));
 sg13g2_tiehi _25934__88 (.L_HI(net88));
 sg13g2_tiehi _25933__89 (.L_HI(net89));
 sg13g2_tiehi _25932__90 (.L_HI(net90));
 sg13g2_tiehi _25931__91 (.L_HI(net91));
 sg13g2_tiehi _25930__92 (.L_HI(net92));
 sg13g2_tiehi _25929__93 (.L_HI(net93));
 sg13g2_tiehi _25928__94 (.L_HI(net94));
 sg13g2_tiehi _25927__95 (.L_HI(net95));
 sg13g2_tiehi _25926__96 (.L_HI(net96));
 sg13g2_tiehi _25925__97 (.L_HI(net97));
 sg13g2_tiehi _25924__98 (.L_HI(net98));
 sg13g2_tiehi _25923__99 (.L_HI(net99));
 sg13g2_tiehi _25922__100 (.L_HI(net100));
 sg13g2_tiehi _25921__101 (.L_HI(net101));
 sg13g2_tiehi _25920__102 (.L_HI(net102));
 sg13g2_tiehi _25919__103 (.L_HI(net103));
 sg13g2_tiehi _25918__104 (.L_HI(net104));
 sg13g2_tiehi _25917__105 (.L_HI(net105));
 sg13g2_tiehi _25916__106 (.L_HI(net106));
 sg13g2_tiehi _25915__107 (.L_HI(net107));
 sg13g2_tiehi _25914__108 (.L_HI(net108));
 sg13g2_tiehi _25913__109 (.L_HI(net109));
 sg13g2_tiehi _25912__110 (.L_HI(net110));
 sg13g2_tiehi _24217__111 (.L_HI(net111));
 sg13g2_tiehi _24216__112 (.L_HI(net112));
 sg13g2_tiehi _24215__113 (.L_HI(net113));
 sg13g2_tiehi _24214__114 (.L_HI(net114));
 sg13g2_tiehi _24213__115 (.L_HI(net115));
 sg13g2_tiehi _24212__116 (.L_HI(net116));
 sg13g2_tiehi _24211__117 (.L_HI(net117));
 sg13g2_tiehi _24210__118 (.L_HI(net118));
 sg13g2_tiehi _24209__119 (.L_HI(net119));
 sg13g2_tiehi _24208__120 (.L_HI(net120));
 sg13g2_tiehi _24207__121 (.L_HI(net121));
 sg13g2_tiehi _24206__122 (.L_HI(net122));
 sg13g2_tiehi _24205__123 (.L_HI(net123));
 sg13g2_tiehi _23807__124 (.L_HI(net124));
 sg13g2_tiehi _24204__125 (.L_HI(net125));
 sg13g2_tiehi _24203__126 (.L_HI(net126));
 sg13g2_tiehi _24202__127 (.L_HI(net127));
 sg13g2_tiehi _24201__128 (.L_HI(net128));
 sg13g2_tiehi _24200__129 (.L_HI(net129));
 sg13g2_tiehi _24199__130 (.L_HI(net130));
 sg13g2_tiehi _24198__131 (.L_HI(net131));
 sg13g2_tiehi _24197__132 (.L_HI(net132));
 sg13g2_tiehi _24196__133 (.L_HI(net133));
 sg13g2_tiehi _24195__134 (.L_HI(net134));
 sg13g2_tiehi _24194__135 (.L_HI(net135));
 sg13g2_tiehi _24193__136 (.L_HI(net136));
 sg13g2_tiehi _24192__137 (.L_HI(net137));
 sg13g2_tiehi _24191__138 (.L_HI(net138));
 sg13g2_tiehi _24190__139 (.L_HI(net139));
 sg13g2_tiehi _24189__140 (.L_HI(net140));
 sg13g2_tiehi _24188__141 (.L_HI(net141));
 sg13g2_tiehi _24187__142 (.L_HI(net142));
 sg13g2_tiehi _24186__143 (.L_HI(net143));
 sg13g2_tiehi _24185__144 (.L_HI(net144));
 sg13g2_tiehi _24184__145 (.L_HI(net145));
 sg13g2_tiehi _24183__146 (.L_HI(net146));
 sg13g2_tiehi _24182__147 (.L_HI(net147));
 sg13g2_tiehi _24181__148 (.L_HI(net148));
 sg13g2_tiehi _24180__149 (.L_HI(net149));
 sg13g2_tiehi _24179__150 (.L_HI(net150));
 sg13g2_tiehi _24178__151 (.L_HI(net151));
 sg13g2_tiehi _24177__152 (.L_HI(net152));
 sg13g2_tiehi _24176__153 (.L_HI(net153));
 sg13g2_tiehi _24175__154 (.L_HI(net154));
 sg13g2_tiehi _24174__155 (.L_HI(net155));
 sg13g2_tiehi _24173__156 (.L_HI(net156));
 sg13g2_tiehi _24172__157 (.L_HI(net157));
 sg13g2_tiehi _24171__158 (.L_HI(net158));
 sg13g2_tiehi _24170__159 (.L_HI(net159));
 sg13g2_tiehi _24169__160 (.L_HI(net160));
 sg13g2_tiehi _24168__161 (.L_HI(net161));
 sg13g2_tiehi _24167__162 (.L_HI(net162));
 sg13g2_tiehi _24166__163 (.L_HI(net163));
 sg13g2_tiehi _24165__164 (.L_HI(net164));
 sg13g2_tiehi _24164__165 (.L_HI(net165));
 sg13g2_tiehi _24163__166 (.L_HI(net166));
 sg13g2_tiehi _24162__167 (.L_HI(net167));
 sg13g2_tiehi _24161__168 (.L_HI(net168));
 sg13g2_tiehi _24160__169 (.L_HI(net169));
 sg13g2_tiehi _24159__170 (.L_HI(net170));
 sg13g2_tiehi _24158__171 (.L_HI(net171));
 sg13g2_tiehi _24157__172 (.L_HI(net172));
 sg13g2_tiehi _24156__173 (.L_HI(net173));
 sg13g2_tiehi _24155__174 (.L_HI(net174));
 sg13g2_tiehi _24154__175 (.L_HI(net175));
 sg13g2_tiehi _24153__176 (.L_HI(net176));
 sg13g2_tiehi _24152__177 (.L_HI(net177));
 sg13g2_tiehi _24151__178 (.L_HI(net178));
 sg13g2_tiehi _24150__179 (.L_HI(net179));
 sg13g2_tiehi _24149__180 (.L_HI(net180));
 sg13g2_tiehi _24148__181 (.L_HI(net181));
 sg13g2_tiehi _24147__182 (.L_HI(net182));
 sg13g2_tiehi _24146__183 (.L_HI(net183));
 sg13g2_tiehi _24145__184 (.L_HI(net184));
 sg13g2_tiehi _24144__185 (.L_HI(net185));
 sg13g2_tiehi _24143__186 (.L_HI(net186));
 sg13g2_tiehi _24142__187 (.L_HI(net187));
 sg13g2_tiehi _24141__188 (.L_HI(net188));
 sg13g2_tiehi _24140__189 (.L_HI(net189));
 sg13g2_tiehi _24139__190 (.L_HI(net190));
 sg13g2_tiehi _24138__191 (.L_HI(net191));
 sg13g2_tiehi _23889__192 (.L_HI(net192));
 sg13g2_tiehi _24137__193 (.L_HI(net193));
 sg13g2_tiehi _24136__194 (.L_HI(net194));
 sg13g2_tiehi _24135__195 (.L_HI(net195));
 sg13g2_tiehi _24134__196 (.L_HI(net196));
 sg13g2_tiehi _24133__197 (.L_HI(net197));
 sg13g2_tiehi _24132__198 (.L_HI(net198));
 sg13g2_tiehi _24131__199 (.L_HI(net199));
 sg13g2_tiehi _24130__200 (.L_HI(net200));
 sg13g2_tiehi _24129__201 (.L_HI(net201));
 sg13g2_tiehi _24128__202 (.L_HI(net202));
 sg13g2_tiehi _24127__203 (.L_HI(net203));
 sg13g2_tiehi _24126__204 (.L_HI(net204));
 sg13g2_tiehi _24125__205 (.L_HI(net205));
 sg13g2_tiehi _24124__206 (.L_HI(net206));
 sg13g2_tiehi _24123__207 (.L_HI(net207));
 sg13g2_tiehi _24122__208 (.L_HI(net208));
 sg13g2_tiehi _24121__209 (.L_HI(net209));
 sg13g2_tiehi _24120__210 (.L_HI(net210));
 sg13g2_tiehi _24119__211 (.L_HI(net211));
 sg13g2_tiehi _24118__212 (.L_HI(net212));
 sg13g2_tiehi _24117__213 (.L_HI(net213));
 sg13g2_tiehi _24116__214 (.L_HI(net214));
 sg13g2_tiehi _24115__215 (.L_HI(net215));
 sg13g2_tiehi _24114__216 (.L_HI(net216));
 sg13g2_tiehi _24113__217 (.L_HI(net217));
 sg13g2_tiehi _24112__218 (.L_HI(net218));
 sg13g2_tiehi _24111__219 (.L_HI(net219));
 sg13g2_tiehi _24110__220 (.L_HI(net220));
 sg13g2_tiehi _24109__221 (.L_HI(net221));
 sg13g2_tiehi _24108__222 (.L_HI(net222));
 sg13g2_tiehi _24107__223 (.L_HI(net223));
 sg13g2_tiehi _24106__224 (.L_HI(net224));
 sg13g2_tiehi _24105__225 (.L_HI(net225));
 sg13g2_tiehi _24104__226 (.L_HI(net226));
 sg13g2_tiehi _24103__227 (.L_HI(net227));
 sg13g2_tiehi _24102__228 (.L_HI(net228));
 sg13g2_tiehi _24101__229 (.L_HI(net229));
 sg13g2_tiehi _24100__230 (.L_HI(net230));
 sg13g2_tiehi _24099__231 (.L_HI(net231));
 sg13g2_tiehi _24098__232 (.L_HI(net232));
 sg13g2_tiehi _24097__233 (.L_HI(net233));
 sg13g2_tiehi _24096__234 (.L_HI(net234));
 sg13g2_tiehi _24095__235 (.L_HI(net235));
 sg13g2_tiehi _24094__236 (.L_HI(net236));
 sg13g2_tiehi _24093__237 (.L_HI(net237));
 sg13g2_tiehi _24092__238 (.L_HI(net238));
 sg13g2_tiehi _24091__239 (.L_HI(net239));
 sg13g2_tiehi _24090__240 (.L_HI(net240));
 sg13g2_tiehi _24084__241 (.L_HI(net241));
 sg13g2_tiehi _24083__242 (.L_HI(net242));
 sg13g2_tiehi _24082__243 (.L_HI(net243));
 sg13g2_tiehi _24081__244 (.L_HI(net244));
 sg13g2_tiehi _24080__245 (.L_HI(net245));
 sg13g2_tiehi _24079__246 (.L_HI(net246));
 sg13g2_tiehi _24078__247 (.L_HI(net247));
 sg13g2_tiehi _24077__248 (.L_HI(net248));
 sg13g2_tiehi _24076__249 (.L_HI(net249));
 sg13g2_tiehi _24075__250 (.L_HI(net250));
 sg13g2_tiehi _24074__251 (.L_HI(net251));
 sg13g2_tiehi _24073__252 (.L_HI(net252));
 sg13g2_tiehi _24072__253 (.L_HI(net253));
 sg13g2_tiehi _24071__254 (.L_HI(net254));
 sg13g2_tiehi _24070__255 (.L_HI(net255));
 sg13g2_tiehi _24069__256 (.L_HI(net256));
 sg13g2_tiehi _24068__257 (.L_HI(net257));
 sg13g2_tiehi _24067__258 (.L_HI(net258));
 sg13g2_tiehi _24066__259 (.L_HI(net259));
 sg13g2_tiehi _24065__260 (.L_HI(net260));
 sg13g2_tiehi _24064__261 (.L_HI(net261));
 sg13g2_tiehi _24063__262 (.L_HI(net262));
 sg13g2_tiehi _24062__263 (.L_HI(net263));
 sg13g2_tiehi _24061__264 (.L_HI(net264));
 sg13g2_tiehi _24060__265 (.L_HI(net265));
 sg13g2_tiehi _24059__266 (.L_HI(net266));
 sg13g2_tiehi _24058__267 (.L_HI(net267));
 sg13g2_tiehi _24057__268 (.L_HI(net268));
 sg13g2_tiehi _24056__269 (.L_HI(net269));
 sg13g2_tiehi _24055__270 (.L_HI(net270));
 sg13g2_tiehi _24054__271 (.L_HI(net271));
 sg13g2_tiehi _24053__272 (.L_HI(net272));
 sg13g2_tiehi _24052__273 (.L_HI(net273));
 sg13g2_tiehi _24051__274 (.L_HI(net274));
 sg13g2_tiehi _24050__275 (.L_HI(net275));
 sg13g2_tiehi _24049__276 (.L_HI(net276));
 sg13g2_tiehi _24048__277 (.L_HI(net277));
 sg13g2_tiehi _24047__278 (.L_HI(net278));
 sg13g2_tiehi _24046__279 (.L_HI(net279));
 sg13g2_tiehi _24045__280 (.L_HI(net280));
 sg13g2_tiehi _24044__281 (.L_HI(net281));
 sg13g2_tiehi _24043__282 (.L_HI(net282));
 sg13g2_tiehi _24042__283 (.L_HI(net283));
 sg13g2_tiehi _24041__284 (.L_HI(net284));
 sg13g2_tiehi _24040__285 (.L_HI(net285));
 sg13g2_tiehi _24039__286 (.L_HI(net286));
 sg13g2_tiehi _24038__287 (.L_HI(net287));
 sg13g2_tiehi _24037__288 (.L_HI(net288));
 sg13g2_tiehi _24036__289 (.L_HI(net289));
 sg13g2_tiehi _24035__290 (.L_HI(net290));
 sg13g2_tiehi _24034__291 (.L_HI(net291));
 sg13g2_tiehi _24033__292 (.L_HI(net292));
 sg13g2_tiehi _24032__293 (.L_HI(net293));
 sg13g2_tiehi _24031__294 (.L_HI(net294));
 sg13g2_tiehi _24030__295 (.L_HI(net295));
 sg13g2_tiehi _24029__296 (.L_HI(net296));
 sg13g2_tiehi _24028__297 (.L_HI(net297));
 sg13g2_tiehi _24027__298 (.L_HI(net298));
 sg13g2_tiehi _24026__299 (.L_HI(net299));
 sg13g2_tiehi _24025__300 (.L_HI(net300));
 sg13g2_tiehi _24024__301 (.L_HI(net301));
 sg13g2_tiehi _24023__302 (.L_HI(net302));
 sg13g2_tiehi _24022__303 (.L_HI(net303));
 sg13g2_tiehi _24021__304 (.L_HI(net304));
 sg13g2_tiehi _24020__305 (.L_HI(net305));
 sg13g2_tiehi _24019__306 (.L_HI(net306));
 sg13g2_tiehi _24018__307 (.L_HI(net307));
 sg13g2_tiehi _24017__308 (.L_HI(net308));
 sg13g2_tiehi _24016__309 (.L_HI(net309));
 sg13g2_tiehi _24015__310 (.L_HI(net310));
 sg13g2_tiehi _24014__311 (.L_HI(net311));
 sg13g2_tiehi _24013__312 (.L_HI(net312));
 sg13g2_tiehi _24012__313 (.L_HI(net313));
 sg13g2_tiehi _24011__314 (.L_HI(net314));
 sg13g2_tiehi _24010__315 (.L_HI(net315));
 sg13g2_tiehi _24009__316 (.L_HI(net316));
 sg13g2_tiehi _24008__317 (.L_HI(net317));
 sg13g2_tiehi _24007__318 (.L_HI(net318));
 sg13g2_tiehi _24006__319 (.L_HI(net319));
 sg13g2_tiehi _24005__320 (.L_HI(net320));
 sg13g2_tiehi _24004__321 (.L_HI(net321));
 sg13g2_tiehi _24003__322 (.L_HI(net322));
 sg13g2_tiehi _24002__323 (.L_HI(net323));
 sg13g2_tiehi _24001__324 (.L_HI(net324));
 sg13g2_tiehi _24000__325 (.L_HI(net325));
 sg13g2_tiehi _23999__326 (.L_HI(net326));
 sg13g2_tiehi _23998__327 (.L_HI(net327));
 sg13g2_tiehi _23997__328 (.L_HI(net328));
 sg13g2_tiehi _23996__329 (.L_HI(net329));
 sg13g2_tiehi _23995__330 (.L_HI(net330));
 sg13g2_tiehi _23994__331 (.L_HI(net331));
 sg13g2_tiehi _23993__332 (.L_HI(net332));
 sg13g2_tiehi _23992__333 (.L_HI(net333));
 sg13g2_tiehi _23991__334 (.L_HI(net334));
 sg13g2_tiehi _23990__335 (.L_HI(net335));
 sg13g2_tiehi _23989__336 (.L_HI(net336));
 sg13g2_tiehi _23988__337 (.L_HI(net337));
 sg13g2_tiehi _23987__338 (.L_HI(net338));
 sg13g2_tiehi _23986__339 (.L_HI(net339));
 sg13g2_tiehi _23985__340 (.L_HI(net340));
 sg13g2_tiehi _23984__341 (.L_HI(net341));
 sg13g2_tiehi _23983__342 (.L_HI(net342));
 sg13g2_tiehi _23982__343 (.L_HI(net343));
 sg13g2_tiehi _23981__344 (.L_HI(net344));
 sg13g2_tiehi _23980__345 (.L_HI(net345));
 sg13g2_tiehi _23979__346 (.L_HI(net346));
 sg13g2_tiehi _23978__347 (.L_HI(net347));
 sg13g2_tiehi _23977__348 (.L_HI(net348));
 sg13g2_tiehi _23976__349 (.L_HI(net349));
 sg13g2_tiehi _23975__350 (.L_HI(net350));
 sg13g2_tiehi _23974__351 (.L_HI(net351));
 sg13g2_tiehi _23973__352 (.L_HI(net352));
 sg13g2_tiehi _23972__353 (.L_HI(net353));
 sg13g2_tiehi _23971__354 (.L_HI(net354));
 sg13g2_tiehi _23970__355 (.L_HI(net355));
 sg13g2_tiehi _23969__356 (.L_HI(net356));
 sg13g2_tiehi _23968__357 (.L_HI(net357));
 sg13g2_tiehi _23967__358 (.L_HI(net358));
 sg13g2_tiehi _23966__359 (.L_HI(net359));
 sg13g2_tiehi _23965__360 (.L_HI(net360));
 sg13g2_tiehi _23964__361 (.L_HI(net361));
 sg13g2_tiehi _23963__362 (.L_HI(net362));
 sg13g2_tiehi _23962__363 (.L_HI(net363));
 sg13g2_tiehi _23961__364 (.L_HI(net364));
 sg13g2_tiehi _23960__365 (.L_HI(net365));
 sg13g2_tiehi _23959__366 (.L_HI(net366));
 sg13g2_tiehi _23958__367 (.L_HI(net367));
 sg13g2_tiehi _23957__368 (.L_HI(net368));
 sg13g2_tiehi _23956__369 (.L_HI(net369));
 sg13g2_tiehi _23955__370 (.L_HI(net370));
 sg13g2_tiehi _23954__371 (.L_HI(net371));
 sg13g2_tiehi _23953__372 (.L_HI(net372));
 sg13g2_tiehi _23952__373 (.L_HI(net373));
 sg13g2_tiehi _23951__374 (.L_HI(net374));
 sg13g2_tiehi _23950__375 (.L_HI(net375));
 sg13g2_tiehi _23949__376 (.L_HI(net376));
 sg13g2_tiehi _23948__377 (.L_HI(net377));
 sg13g2_tiehi _23947__378 (.L_HI(net378));
 sg13g2_tiehi _23946__379 (.L_HI(net379));
 sg13g2_tiehi _23945__380 (.L_HI(net380));
 sg13g2_tiehi _23944__381 (.L_HI(net381));
 sg13g2_tiehi _23943__382 (.L_HI(net382));
 sg13g2_tiehi _23942__383 (.L_HI(net383));
 sg13g2_tiehi _24085__384 (.L_HI(net384));
 sg13g2_tiehi _23941__385 (.L_HI(net385));
 sg13g2_tiehi _23940__386 (.L_HI(net386));
 sg13g2_tiehi _23939__387 (.L_HI(net387));
 sg13g2_tiehi _23938__388 (.L_HI(net388));
 sg13g2_tiehi _23937__389 (.L_HI(net389));
 sg13g2_tiehi _23936__390 (.L_HI(net390));
 sg13g2_tiehi _23935__391 (.L_HI(net391));
 sg13g2_tiehi _23934__392 (.L_HI(net392));
 sg13g2_tiehi _23933__393 (.L_HI(net393));
 sg13g2_tiehi _23932__394 (.L_HI(net394));
 sg13g2_tiehi _23931__395 (.L_HI(net395));
 sg13g2_tiehi _23930__396 (.L_HI(net396));
 sg13g2_tiehi _23929__397 (.L_HI(net397));
 sg13g2_tiehi _23928__398 (.L_HI(net398));
 sg13g2_tiehi _23927__399 (.L_HI(net399));
 sg13g2_tiehi _23926__400 (.L_HI(net400));
 sg13g2_tiehi _23925__401 (.L_HI(net401));
 sg13g2_tiehi _23924__402 (.L_HI(net402));
 sg13g2_tiehi _23923__403 (.L_HI(net403));
 sg13g2_tiehi _23922__404 (.L_HI(net404));
 sg13g2_tiehi _23921__405 (.L_HI(net405));
 sg13g2_tiehi _23920__406 (.L_HI(net406));
 sg13g2_tiehi _23919__407 (.L_HI(net407));
 sg13g2_tiehi _23918__408 (.L_HI(net408));
 sg13g2_tiehi _23917__409 (.L_HI(net409));
 sg13g2_tiehi _23916__410 (.L_HI(net410));
 sg13g2_tiehi _23915__411 (.L_HI(net411));
 sg13g2_tiehi _23914__412 (.L_HI(net412));
 sg13g2_tiehi _23913__413 (.L_HI(net413));
 sg13g2_tiehi _23912__414 (.L_HI(net414));
 sg13g2_tiehi _23911__415 (.L_HI(net415));
 sg13g2_tiehi _23910__416 (.L_HI(net416));
 sg13g2_tiehi _23909__417 (.L_HI(net417));
 sg13g2_tiehi _23908__418 (.L_HI(net418));
 sg13g2_tiehi _23907__419 (.L_HI(net419));
 sg13g2_tiehi _23906__420 (.L_HI(net420));
 sg13g2_tiehi _23905__421 (.L_HI(net421));
 sg13g2_tiehi _23904__422 (.L_HI(net422));
 sg13g2_tiehi _23903__423 (.L_HI(net423));
 sg13g2_tiehi _23902__424 (.L_HI(net424));
 sg13g2_tiehi _23901__425 (.L_HI(net425));
 sg13g2_tiehi _23900__426 (.L_HI(net426));
 sg13g2_tiehi _23899__427 (.L_HI(net427));
 sg13g2_tiehi _23898__428 (.L_HI(net428));
 sg13g2_tiehi _23897__429 (.L_HI(net429));
 sg13g2_tiehi _23896__430 (.L_HI(net430));
 sg13g2_tiehi _23895__431 (.L_HI(net431));
 sg13g2_tiehi _23894__432 (.L_HI(net432));
 sg13g2_tiehi _23888__433 (.L_HI(net433));
 sg13g2_tiehi _23887__434 (.L_HI(net434));
 sg13g2_tiehi _23886__435 (.L_HI(net435));
 sg13g2_tiehi _23885__436 (.L_HI(net436));
 sg13g2_tiehi _23884__437 (.L_HI(net437));
 sg13g2_tiehi _23883__438 (.L_HI(net438));
 sg13g2_tiehi _23882__439 (.L_HI(net439));
 sg13g2_tiehi _23881__440 (.L_HI(net440));
 sg13g2_tiehi _23880__441 (.L_HI(net441));
 sg13g2_tiehi _23879__442 (.L_HI(net442));
 sg13g2_tiehi _23878__443 (.L_HI(net443));
 sg13g2_tiehi _23877__444 (.L_HI(net444));
 sg13g2_tiehi _23876__445 (.L_HI(net445));
 sg13g2_tiehi _23875__446 (.L_HI(net446));
 sg13g2_tiehi _23874__447 (.L_HI(net447));
 sg13g2_tiehi _23873__448 (.L_HI(net448));
 sg13g2_tiehi _23872__449 (.L_HI(net449));
 sg13g2_tiehi _23871__450 (.L_HI(net450));
 sg13g2_tiehi _23870__451 (.L_HI(net451));
 sg13g2_tiehi _23869__452 (.L_HI(net452));
 sg13g2_tiehi _23868__453 (.L_HI(net453));
 sg13g2_tiehi _23867__454 (.L_HI(net454));
 sg13g2_tiehi _23866__455 (.L_HI(net455));
 sg13g2_tiehi _23865__456 (.L_HI(net456));
 sg13g2_tiehi _23864__457 (.L_HI(net457));
 sg13g2_tiehi _23863__458 (.L_HI(net458));
 sg13g2_tiehi _23862__459 (.L_HI(net459));
 sg13g2_tiehi _23861__460 (.L_HI(net460));
 sg13g2_tiehi _23860__461 (.L_HI(net461));
 sg13g2_tiehi _23859__462 (.L_HI(net462));
 sg13g2_tiehi _23858__463 (.L_HI(net463));
 sg13g2_tiehi _23857__464 (.L_HI(net464));
 sg13g2_tiehi _23856__465 (.L_HI(net465));
 sg13g2_tiehi _23855__466 (.L_HI(net466));
 sg13g2_tiehi _23854__467 (.L_HI(net467));
 sg13g2_tiehi _23853__468 (.L_HI(net468));
 sg13g2_tiehi _23852__469 (.L_HI(net469));
 sg13g2_tiehi _23851__470 (.L_HI(net470));
 sg13g2_tiehi _23850__471 (.L_HI(net471));
 sg13g2_tiehi _23849__472 (.L_HI(net472));
 sg13g2_tiehi _23848__473 (.L_HI(net473));
 sg13g2_tiehi _23847__474 (.L_HI(net474));
 sg13g2_tiehi _23846__475 (.L_HI(net475));
 sg13g2_tiehi _23845__476 (.L_HI(net476));
 sg13g2_tiehi _23844__477 (.L_HI(net477));
 sg13g2_tiehi _23843__478 (.L_HI(net478));
 sg13g2_tiehi _23842__479 (.L_HI(net479));
 sg13g2_tiehi _23841__480 (.L_HI(net480));
 sg13g2_tiehi _23840__481 (.L_HI(net481));
 sg13g2_tiehi _23839__482 (.L_HI(net482));
 sg13g2_tiehi _23838__483 (.L_HI(net483));
 sg13g2_tiehi _23837__484 (.L_HI(net484));
 sg13g2_tiehi _23836__485 (.L_HI(net485));
 sg13g2_tiehi _23835__486 (.L_HI(net486));
 sg13g2_tiehi _23834__487 (.L_HI(net487));
 sg13g2_tiehi _23833__488 (.L_HI(net488));
 sg13g2_tiehi _23832__489 (.L_HI(net489));
 sg13g2_tiehi _23831__490 (.L_HI(net490));
 sg13g2_tiehi _23830__491 (.L_HI(net491));
 sg13g2_tiehi _23829__492 (.L_HI(net492));
 sg13g2_tiehi _23828__493 (.L_HI(net493));
 sg13g2_tiehi _23827__494 (.L_HI(net494));
 sg13g2_tiehi _23826__495 (.L_HI(net495));
 sg13g2_tiehi _23806__496 (.L_HI(net496));
 sg13g2_tiehi _23805__497 (.L_HI(net497));
 sg13g2_tiehi _23804__498 (.L_HI(net498));
 sg13g2_tiehi _23803__499 (.L_HI(net499));
 sg13g2_tiehi _23802__500 (.L_HI(net500));
 sg13g2_tiehi _23801__501 (.L_HI(net501));
 sg13g2_tiehi _23800__502 (.L_HI(net502));
 sg13g2_tiehi _23799__503 (.L_HI(net503));
 sg13g2_tiehi _23798__504 (.L_HI(net504));
 sg13g2_tiehi _23797__505 (.L_HI(net505));
 sg13g2_tiehi _23796__506 (.L_HI(net506));
 sg13g2_tiehi _23795__507 (.L_HI(net507));
 sg13g2_tiehi _23794__508 (.L_HI(net508));
 sg13g2_tiehi _23793__509 (.L_HI(net509));
 sg13g2_tiehi _23792__510 (.L_HI(net510));
 sg13g2_tiehi _23791__511 (.L_HI(net511));
 sg13g2_tiehi _23790__512 (.L_HI(net512));
 sg13g2_tiehi _23789__513 (.L_HI(net513));
 sg13g2_tiehi _23788__514 (.L_HI(net514));
 sg13g2_tiehi _23787__515 (.L_HI(net515));
 sg13g2_tiehi _23786__516 (.L_HI(net516));
 sg13g2_tiehi _23785__517 (.L_HI(net517));
 sg13g2_tiehi _23784__518 (.L_HI(net518));
 sg13g2_tiehi _23783__519 (.L_HI(net519));
 sg13g2_tiehi _23782__520 (.L_HI(net520));
 sg13g2_tiehi _23781__521 (.L_HI(net521));
 sg13g2_tiehi _23780__522 (.L_HI(net522));
 sg13g2_tiehi _23779__523 (.L_HI(net523));
 sg13g2_tiehi _23778__524 (.L_HI(net524));
 sg13g2_tiehi _23777__525 (.L_HI(net525));
 sg13g2_tiehi _23776__526 (.L_HI(net526));
 sg13g2_tiehi _23775__527 (.L_HI(net527));
 sg13g2_tiehi _23774__528 (.L_HI(net528));
 sg13g2_tiehi _23773__529 (.L_HI(net529));
 sg13g2_tiehi _23772__530 (.L_HI(net530));
 sg13g2_tiehi _23771__531 (.L_HI(net531));
 sg13g2_tiehi _23770__532 (.L_HI(net532));
 sg13g2_tiehi _23769__533 (.L_HI(net533));
 sg13g2_tiehi _23768__534 (.L_HI(net534));
 sg13g2_tiehi _23767__535 (.L_HI(net535));
 sg13g2_tiehi _23766__536 (.L_HI(net536));
 sg13g2_tiehi _23765__537 (.L_HI(net537));
 sg13g2_tiehi _23764__538 (.L_HI(net538));
 sg13g2_tiehi _23763__539 (.L_HI(net539));
 sg13g2_tiehi _23762__540 (.L_HI(net540));
 sg13g2_tiehi _23761__541 (.L_HI(net541));
 sg13g2_tiehi _23760__542 (.L_HI(net542));
 sg13g2_tiehi _23759__543 (.L_HI(net543));
 sg13g2_tiehi _23758__544 (.L_HI(net544));
 sg13g2_tiehi _23757__545 (.L_HI(net545));
 sg13g2_tiehi _23756__546 (.L_HI(net546));
 sg13g2_tiehi _23755__547 (.L_HI(net547));
 sg13g2_tiehi _23754__548 (.L_HI(net548));
 sg13g2_tiehi _23753__549 (.L_HI(net549));
 sg13g2_tiehi _23752__550 (.L_HI(net550));
 sg13g2_tiehi _23751__551 (.L_HI(net551));
 sg13g2_tiehi _23750__552 (.L_HI(net552));
 sg13g2_tiehi _23749__553 (.L_HI(net553));
 sg13g2_tiehi _23748__554 (.L_HI(net554));
 sg13g2_tiehi _23747__555 (.L_HI(net555));
 sg13g2_tiehi _23746__556 (.L_HI(net556));
 sg13g2_tiehi _23745__557 (.L_HI(net557));
 sg13g2_tiehi _23744__558 (.L_HI(net558));
 sg13g2_tiehi _23743__559 (.L_HI(net559));
 sg13g2_tiehi _23742__560 (.L_HI(net560));
 sg13g2_tiehi _23741__561 (.L_HI(net561));
 sg13g2_tiehi _23740__562 (.L_HI(net562));
 sg13g2_tiehi _23739__563 (.L_HI(net563));
 sg13g2_tiehi _23738__564 (.L_HI(net564));
 sg13g2_tiehi _23737__565 (.L_HI(net565));
 sg13g2_tiehi _23736__566 (.L_HI(net566));
 sg13g2_tiehi _23735__567 (.L_HI(net567));
 sg13g2_tiehi _23734__568 (.L_HI(net568));
 sg13g2_tiehi _23733__569 (.L_HI(net569));
 sg13g2_tiehi _23732__570 (.L_HI(net570));
 sg13g2_tiehi _23731__571 (.L_HI(net571));
 sg13g2_tiehi _23730__572 (.L_HI(net572));
 sg13g2_tiehi _23729__573 (.L_HI(net573));
 sg13g2_tiehi _23728__574 (.L_HI(net574));
 sg13g2_tiehi _23727__575 (.L_HI(net575));
 sg13g2_tiehi _23726__576 (.L_HI(net576));
 sg13g2_tiehi _23725__577 (.L_HI(net577));
 sg13g2_tiehi _23724__578 (.L_HI(net578));
 sg13g2_tiehi _23723__579 (.L_HI(net579));
 sg13g2_tiehi _23722__580 (.L_HI(net580));
 sg13g2_tiehi _23721__581 (.L_HI(net581));
 sg13g2_tiehi _23720__582 (.L_HI(net582));
 sg13g2_tiehi _23719__583 (.L_HI(net583));
 sg13g2_tiehi _23718__584 (.L_HI(net584));
 sg13g2_tiehi _23717__585 (.L_HI(net585));
 sg13g2_tiehi _23716__586 (.L_HI(net586));
 sg13g2_tiehi _23715__587 (.L_HI(net587));
 sg13g2_tiehi _23714__588 (.L_HI(net588));
 sg13g2_tiehi _23713__589 (.L_HI(net589));
 sg13g2_tiehi _23712__590 (.L_HI(net590));
 sg13g2_tiehi _23605__591 (.L_HI(net591));
 sg13g2_tiehi _23604__592 (.L_HI(net592));
 sg13g2_tiehi _23603__593 (.L_HI(net593));
 sg13g2_tiehi _23602__594 (.L_HI(net594));
 sg13g2_tiehi _23601__595 (.L_HI(net595));
 sg13g2_tiehi _23600__596 (.L_HI(net596));
 sg13g2_tiehi _23599__597 (.L_HI(net597));
 sg13g2_tiehi _23598__598 (.L_HI(net598));
 sg13g2_tiehi _23597__599 (.L_HI(net599));
 sg13g2_tiehi _23596__600 (.L_HI(net600));
 sg13g2_tiehi _23595__601 (.L_HI(net601));
 sg13g2_tiehi _23594__602 (.L_HI(net602));
 sg13g2_tiehi _23593__603 (.L_HI(net603));
 sg13g2_tiehi _23592__604 (.L_HI(net604));
 sg13g2_tiehi _23591__605 (.L_HI(net605));
 sg13g2_tiehi _23590__606 (.L_HI(net606));
 sg13g2_tiehi _23589__607 (.L_HI(net607));
 sg13g2_tiehi _23588__608 (.L_HI(net608));
 sg13g2_tiehi _23587__609 (.L_HI(net609));
 sg13g2_tiehi _23586__610 (.L_HI(net610));
 sg13g2_tiehi _23585__611 (.L_HI(net611));
 sg13g2_tiehi _23584__612 (.L_HI(net612));
 sg13g2_tiehi _23583__613 (.L_HI(net613));
 sg13g2_tiehi _23582__614 (.L_HI(net614));
 sg13g2_tiehi _23581__615 (.L_HI(net615));
 sg13g2_tiehi _23580__616 (.L_HI(net616));
 sg13g2_tiehi _23579__617 (.L_HI(net617));
 sg13g2_tiehi _23578__618 (.L_HI(net618));
 sg13g2_tiehi _23577__619 (.L_HI(net619));
 sg13g2_tiehi _23576__620 (.L_HI(net620));
 sg13g2_tiehi _23575__621 (.L_HI(net621));
 sg13g2_tiehi _23574__622 (.L_HI(net622));
 sg13g2_tiehi _24439__623 (.L_HI(net623));
 sg13g2_tiehi _24440__624 (.L_HI(net624));
 sg13g2_tiehi _24441__625 (.L_HI(net625));
 sg13g2_tiehi _25911__626 (.L_HI(net626));
 sg13g2_tiehi _25910__627 (.L_HI(net627));
 sg13g2_tiehi _23474__628 (.L_HI(net628));
 sg13g2_tiehi _23473__629 (.L_HI(net629));
 sg13g2_tiehi _23472__630 (.L_HI(net630));
 sg13g2_tiehi _23471__631 (.L_HI(net631));
 sg13g2_tiehi _23470__632 (.L_HI(net632));
 sg13g2_tiehi _23469__633 (.L_HI(net633));
 sg13g2_tiehi _23468__634 (.L_HI(net634));
 sg13g2_tiehi _23467__635 (.L_HI(net635));
 sg13g2_tiehi _23466__636 (.L_HI(net636));
 sg13g2_tiehi _23465__637 (.L_HI(net637));
 sg13g2_tiehi _23464__638 (.L_HI(net638));
 sg13g2_tiehi _23463__639 (.L_HI(net639));
 sg13g2_tiehi _23462__640 (.L_HI(net640));
 sg13g2_tiehi _23461__641 (.L_HI(net641));
 sg13g2_tiehi _23460__642 (.L_HI(net642));
 sg13g2_tiehi _23459__643 (.L_HI(net643));
 sg13g2_tiehi _23458__644 (.L_HI(net644));
 sg13g2_tiehi _23457__645 (.L_HI(net645));
 sg13g2_tiehi _23456__646 (.L_HI(net646));
 sg13g2_tiehi _23455__647 (.L_HI(net647));
 sg13g2_tiehi _23454__648 (.L_HI(net648));
 sg13g2_tiehi _23453__649 (.L_HI(net649));
 sg13g2_tiehi _23452__650 (.L_HI(net650));
 sg13g2_tiehi _23451__651 (.L_HI(net651));
 sg13g2_tiehi _23450__652 (.L_HI(net652));
 sg13g2_tiehi _23449__653 (.L_HI(net653));
 sg13g2_tiehi _23448__654 (.L_HI(net654));
 sg13g2_tiehi _23447__655 (.L_HI(net655));
 sg13g2_tiehi _23446__656 (.L_HI(net656));
 sg13g2_tiehi _23445__657 (.L_HI(net657));
 sg13g2_tiehi _23444__658 (.L_HI(net658));
 sg13g2_tiehi _23370__659 (.L_HI(net659));
 sg13g2_tiehi _23369__660 (.L_HI(net660));
 sg13g2_tiehi _23368__661 (.L_HI(net661));
 sg13g2_tiehi _23367__662 (.L_HI(net662));
 sg13g2_tiehi _23366__663 (.L_HI(net663));
 sg13g2_tiehi _23365__664 (.L_HI(net664));
 sg13g2_tiehi _23364__665 (.L_HI(net665));
 sg13g2_tiehi _23363__666 (.L_HI(net666));
 sg13g2_tiehi _23362__667 (.L_HI(net667));
 sg13g2_tiehi _23361__668 (.L_HI(net668));
 sg13g2_tiehi _23360__669 (.L_HI(net669));
 sg13g2_tiehi _23359__670 (.L_HI(net670));
 sg13g2_tiehi _23358__671 (.L_HI(net671));
 sg13g2_tiehi _23357__672 (.L_HI(net672));
 sg13g2_tiehi _23356__673 (.L_HI(net673));
 sg13g2_tiehi _23355__674 (.L_HI(net674));
 sg13g2_tiehi _23354__675 (.L_HI(net675));
 sg13g2_tiehi _23353__676 (.L_HI(net676));
 sg13g2_tiehi _23352__677 (.L_HI(net677));
 sg13g2_tiehi _23351__678 (.L_HI(net678));
 sg13g2_tiehi _23350__679 (.L_HI(net679));
 sg13g2_tiehi _23349__680 (.L_HI(net680));
 sg13g2_tiehi _23348__681 (.L_HI(net681));
 sg13g2_tiehi _23347__682 (.L_HI(net682));
 sg13g2_tiehi _23346__683 (.L_HI(net683));
 sg13g2_tiehi _23345__684 (.L_HI(net684));
 sg13g2_tiehi _23344__685 (.L_HI(net685));
 sg13g2_tiehi _23343__686 (.L_HI(net686));
 sg13g2_tiehi _23342__687 (.L_HI(net687));
 sg13g2_tiehi _23341__688 (.L_HI(net688));
 sg13g2_tiehi _23340__689 (.L_HI(net689));
 sg13g2_tiehi _23339__690 (.L_HI(net690));
 sg13g2_tiehi _23338__691 (.L_HI(net691));
 sg13g2_tiehi _23337__692 (.L_HI(net692));
 sg13g2_tiehi _23336__693 (.L_HI(net693));
 sg13g2_tiehi _23335__694 (.L_HI(net694));
 sg13g2_tiehi _23334__695 (.L_HI(net695));
 sg13g2_tiehi _23333__696 (.L_HI(net696));
 sg13g2_tiehi _23332__697 (.L_HI(net697));
 sg13g2_tiehi _25909__698 (.L_HI(net698));
 sg13g2_tiehi _24583__699 (.L_HI(net699));
 sg13g2_tiehi _25908__700 (.L_HI(net700));
 sg13g2_tiehi _25907__701 (.L_HI(net701));
 sg13g2_tiehi _25906__702 (.L_HI(net702));
 sg13g2_tiehi _25905__703 (.L_HI(net703));
 sg13g2_tiehi _25904__704 (.L_HI(net704));
 sg13g2_tiehi _25903__705 (.L_HI(net705));
 sg13g2_tiehi _25902__706 (.L_HI(net706));
 sg13g2_tiehi _25901__707 (.L_HI(net707));
 sg13g2_tiehi _25900__708 (.L_HI(net708));
 sg13g2_tiehi _25899__709 (.L_HI(net709));
 sg13g2_tiehi _25898__710 (.L_HI(net710));
 sg13g2_tiehi _25897__711 (.L_HI(net711));
 sg13g2_tiehi _25896__712 (.L_HI(net712));
 sg13g2_tiehi _25895__713 (.L_HI(net713));
 sg13g2_tiehi _25894__714 (.L_HI(net714));
 sg13g2_tiehi _25893__715 (.L_HI(net715));
 sg13g2_tiehi _25892__716 (.L_HI(net716));
 sg13g2_tiehi _25891__717 (.L_HI(net717));
 sg13g2_tiehi _25890__718 (.L_HI(net718));
 sg13g2_tiehi _25889__719 (.L_HI(net719));
 sg13g2_tiehi _25888__720 (.L_HI(net720));
 sg13g2_tiehi _25887__721 (.L_HI(net721));
 sg13g2_tiehi _25875__722 (.L_HI(net722));
 sg13g2_tiehi _25874__723 (.L_HI(net723));
 sg13g2_tiehi _25873__724 (.L_HI(net724));
 sg13g2_tiehi _25872__725 (.L_HI(net725));
 sg13g2_tiehi _25871__726 (.L_HI(net726));
 sg13g2_tiehi _25870__727 (.L_HI(net727));
 sg13g2_tiehi _25869__728 (.L_HI(net728));
 sg13g2_tiehi _25868__729 (.L_HI(net729));
 sg13g2_tiehi _25867__730 (.L_HI(net730));
 sg13g2_tiehi _25866__731 (.L_HI(net731));
 sg13g2_tiehi _25865__732 (.L_HI(net732));
 sg13g2_tiehi _25864__733 (.L_HI(net733));
 sg13g2_tiehi _25863__734 (.L_HI(net734));
 sg13g2_tiehi _25862__735 (.L_HI(net735));
 sg13g2_tiehi _25861__736 (.L_HI(net736));
 sg13g2_tiehi _25860__737 (.L_HI(net737));
 sg13g2_tiehi _25859__738 (.L_HI(net738));
 sg13g2_tiehi _25858__739 (.L_HI(net739));
 sg13g2_tiehi _25857__740 (.L_HI(net740));
 sg13g2_tiehi _25856__741 (.L_HI(net741));
 sg13g2_tiehi _25855__742 (.L_HI(net742));
 sg13g2_tiehi _25854__743 (.L_HI(net743));
 sg13g2_tiehi _25853__744 (.L_HI(net744));
 sg13g2_tiehi _25852__745 (.L_HI(net745));
 sg13g2_tiehi _25851__746 (.L_HI(net746));
 sg13g2_tiehi _25850__747 (.L_HI(net747));
 sg13g2_tiehi _25849__748 (.L_HI(net748));
 sg13g2_tiehi _25848__749 (.L_HI(net749));
 sg13g2_tiehi _25847__750 (.L_HI(net750));
 sg13g2_tiehi _25846__751 (.L_HI(net751));
 sg13g2_tiehi _25845__752 (.L_HI(net752));
 sg13g2_tiehi _25844__753 (.L_HI(net753));
 sg13g2_tiehi _25843__754 (.L_HI(net754));
 sg13g2_tiehi _25842__755 (.L_HI(net755));
 sg13g2_tiehi _25841__756 (.L_HI(net756));
 sg13g2_tiehi _25840__757 (.L_HI(net757));
 sg13g2_tiehi _25839__758 (.L_HI(net758));
 sg13g2_tiehi _25838__759 (.L_HI(net759));
 sg13g2_tiehi _25837__760 (.L_HI(net760));
 sg13g2_tiehi _25836__761 (.L_HI(net761));
 sg13g2_tiehi _25835__762 (.L_HI(net762));
 sg13g2_tiehi _25834__763 (.L_HI(net763));
 sg13g2_tiehi _25833__764 (.L_HI(net764));
 sg13g2_tiehi _25832__765 (.L_HI(net765));
 sg13g2_tiehi _25831__766 (.L_HI(net766));
 sg13g2_tiehi _25830__767 (.L_HI(net767));
 sg13g2_tiehi _25829__768 (.L_HI(net768));
 sg13g2_tiehi _25828__769 (.L_HI(net769));
 sg13g2_tiehi _25827__770 (.L_HI(net770));
 sg13g2_tiehi _25826__771 (.L_HI(net771));
 sg13g2_tiehi _25825__772 (.L_HI(net772));
 sg13g2_tiehi _25824__773 (.L_HI(net773));
 sg13g2_tiehi _25823__774 (.L_HI(net774));
 sg13g2_tiehi _25822__775 (.L_HI(net775));
 sg13g2_tiehi _25821__776 (.L_HI(net776));
 sg13g2_tiehi _25820__777 (.L_HI(net777));
 sg13g2_tiehi _25819__778 (.L_HI(net778));
 sg13g2_tiehi _25818__779 (.L_HI(net779));
 sg13g2_tiehi _25817__780 (.L_HI(net780));
 sg13g2_tiehi _25816__781 (.L_HI(net781));
 sg13g2_tiehi _25815__782 (.L_HI(net782));
 sg13g2_tiehi _25814__783 (.L_HI(net783));
 sg13g2_tiehi _25813__784 (.L_HI(net784));
 sg13g2_tiehi _25812__785 (.L_HI(net785));
 sg13g2_tiehi _25811__786 (.L_HI(net786));
 sg13g2_tiehi _25810__787 (.L_HI(net787));
 sg13g2_tiehi _25809__788 (.L_HI(net788));
 sg13g2_tiehi _25808__789 (.L_HI(net789));
 sg13g2_tiehi _25807__790 (.L_HI(net790));
 sg13g2_tiehi _25806__791 (.L_HI(net791));
 sg13g2_tiehi _25805__792 (.L_HI(net792));
 sg13g2_tiehi _25804__793 (.L_HI(net793));
 sg13g2_tiehi _25803__794 (.L_HI(net794));
 sg13g2_tiehi _25802__795 (.L_HI(net795));
 sg13g2_tiehi _25801__796 (.L_HI(net796));
 sg13g2_tiehi _25800__797 (.L_HI(net797));
 sg13g2_tiehi _25799__798 (.L_HI(net798));
 sg13g2_tiehi _25798__799 (.L_HI(net799));
 sg13g2_tiehi _25797__800 (.L_HI(net800));
 sg13g2_tiehi _25796__801 (.L_HI(net801));
 sg13g2_tiehi _25795__802 (.L_HI(net802));
 sg13g2_tiehi _25794__803 (.L_HI(net803));
 sg13g2_tiehi _25793__804 (.L_HI(net804));
 sg13g2_tiehi _25792__805 (.L_HI(net805));
 sg13g2_tiehi _25791__806 (.L_HI(net806));
 sg13g2_tiehi _25790__807 (.L_HI(net807));
 sg13g2_tiehi _25789__808 (.L_HI(net808));
 sg13g2_tiehi _25788__809 (.L_HI(net809));
 sg13g2_tiehi _25787__810 (.L_HI(net810));
 sg13g2_tiehi _25783__811 (.L_HI(net811));
 sg13g2_tiehi _25782__812 (.L_HI(net812));
 sg13g2_tiehi _25781__813 (.L_HI(net813));
 sg13g2_tiehi _25780__814 (.L_HI(net814));
 sg13g2_tiehi _25779__815 (.L_HI(net815));
 sg13g2_tiehi _25778__816 (.L_HI(net816));
 sg13g2_tiehi _25777__817 (.L_HI(net817));
 sg13g2_tiehi _25776__818 (.L_HI(net818));
 sg13g2_tiehi _25775__819 (.L_HI(net819));
 sg13g2_tiehi _25774__820 (.L_HI(net820));
 sg13g2_tiehi _25773__821 (.L_HI(net821));
 sg13g2_tiehi _25772__822 (.L_HI(net822));
 sg13g2_tiehi _25771__823 (.L_HI(net823));
 sg13g2_tiehi _25770__824 (.L_HI(net824));
 sg13g2_tiehi _25769__825 (.L_HI(net825));
 sg13g2_tiehi _25768__826 (.L_HI(net826));
 sg13g2_tiehi _25767__827 (.L_HI(net827));
 sg13g2_tiehi _25766__828 (.L_HI(net828));
 sg13g2_tiehi _25765__829 (.L_HI(net829));
 sg13g2_tiehi _25764__830 (.L_HI(net830));
 sg13g2_tiehi _25763__831 (.L_HI(net831));
 sg13g2_tiehi _25762__832 (.L_HI(net832));
 sg13g2_tiehi _25761__833 (.L_HI(net833));
 sg13g2_tiehi _25760__834 (.L_HI(net834));
 sg13g2_tiehi _25759__835 (.L_HI(net835));
 sg13g2_tiehi _25758__836 (.L_HI(net836));
 sg13g2_tiehi _25757__837 (.L_HI(net837));
 sg13g2_tiehi _25756__838 (.L_HI(net838));
 sg13g2_tiehi _25755__839 (.L_HI(net839));
 sg13g2_tiehi _25754__840 (.L_HI(net840));
 sg13g2_tiehi _25753__841 (.L_HI(net841));
 sg13g2_tiehi _25752__842 (.L_HI(net842));
 sg13g2_tiehi _25751__843 (.L_HI(net843));
 sg13g2_tiehi _25750__844 (.L_HI(net844));
 sg13g2_tiehi _25749__845 (.L_HI(net845));
 sg13g2_tiehi _25748__846 (.L_HI(net846));
 sg13g2_tiehi _25747__847 (.L_HI(net847));
 sg13g2_tiehi _25746__848 (.L_HI(net848));
 sg13g2_tiehi _25745__849 (.L_HI(net849));
 sg13g2_tiehi _25744__850 (.L_HI(net850));
 sg13g2_tiehi _25743__851 (.L_HI(net851));
 sg13g2_tiehi _25742__852 (.L_HI(net852));
 sg13g2_tiehi _25741__853 (.L_HI(net853));
 sg13g2_tiehi _25740__854 (.L_HI(net854));
 sg13g2_tiehi _25739__855 (.L_HI(net855));
 sg13g2_tiehi _25738__856 (.L_HI(net856));
 sg13g2_tiehi _25737__857 (.L_HI(net857));
 sg13g2_tiehi _25736__858 (.L_HI(net858));
 sg13g2_tiehi _25735__859 (.L_HI(net859));
 sg13g2_tiehi _25734__860 (.L_HI(net860));
 sg13g2_tiehi _25733__861 (.L_HI(net861));
 sg13g2_tiehi _25732__862 (.L_HI(net862));
 sg13g2_tiehi _25731__863 (.L_HI(net863));
 sg13g2_tiehi _25730__864 (.L_HI(net864));
 sg13g2_tiehi _25729__865 (.L_HI(net865));
 sg13g2_tiehi _25728__866 (.L_HI(net866));
 sg13g2_tiehi _25727__867 (.L_HI(net867));
 sg13g2_tiehi _25726__868 (.L_HI(net868));
 sg13g2_tiehi _25725__869 (.L_HI(net869));
 sg13g2_tiehi _25724__870 (.L_HI(net870));
 sg13g2_tiehi _25723__871 (.L_HI(net871));
 sg13g2_tiehi _25722__872 (.L_HI(net872));
 sg13g2_tiehi _25721__873 (.L_HI(net873));
 sg13g2_tiehi _25720__874 (.L_HI(net874));
 sg13g2_tiehi _25716__875 (.L_HI(net875));
 sg13g2_tiehi _25715__876 (.L_HI(net876));
 sg13g2_tiehi _25714__877 (.L_HI(net877));
 sg13g2_tiehi _25713__878 (.L_HI(net878));
 sg13g2_tiehi _25712__879 (.L_HI(net879));
 sg13g2_tiehi _25711__880 (.L_HI(net880));
 sg13g2_tiehi _25710__881 (.L_HI(net881));
 sg13g2_tiehi _25709__882 (.L_HI(net882));
 sg13g2_tiehi _25708__883 (.L_HI(net883));
 sg13g2_tiehi _25707__884 (.L_HI(net884));
 sg13g2_tiehi _25706__885 (.L_HI(net885));
 sg13g2_tiehi _25705__886 (.L_HI(net886));
 sg13g2_tiehi _25704__887 (.L_HI(net887));
 sg13g2_tiehi _25703__888 (.L_HI(net888));
 sg13g2_tiehi _25702__889 (.L_HI(net889));
 sg13g2_tiehi _25701__890 (.L_HI(net890));
 sg13g2_tiehi _25700__891 (.L_HI(net891));
 sg13g2_tiehi _25699__892 (.L_HI(net892));
 sg13g2_tiehi _25698__893 (.L_HI(net893));
 sg13g2_tiehi _25697__894 (.L_HI(net894));
 sg13g2_tiehi _25696__895 (.L_HI(net895));
 sg13g2_tiehi _25695__896 (.L_HI(net896));
 sg13g2_tiehi _25694__897 (.L_HI(net897));
 sg13g2_tiehi _25693__898 (.L_HI(net898));
 sg13g2_tiehi _25692__899 (.L_HI(net899));
 sg13g2_tiehi _25691__900 (.L_HI(net900));
 sg13g2_tiehi _25690__901 (.L_HI(net901));
 sg13g2_tiehi _25689__902 (.L_HI(net902));
 sg13g2_tiehi _25688__903 (.L_HI(net903));
 sg13g2_tiehi _25687__904 (.L_HI(net904));
 sg13g2_tiehi _25686__905 (.L_HI(net905));
 sg13g2_tiehi _25685__906 (.L_HI(net906));
 sg13g2_tiehi _25684__907 (.L_HI(net907));
 sg13g2_tiehi _25683__908 (.L_HI(net908));
 sg13g2_tiehi _25682__909 (.L_HI(net909));
 sg13g2_tiehi _25681__910 (.L_HI(net910));
 sg13g2_tiehi _25680__911 (.L_HI(net911));
 sg13g2_tiehi _25679__912 (.L_HI(net912));
 sg13g2_tiehi _25678__913 (.L_HI(net913));
 sg13g2_tiehi _25677__914 (.L_HI(net914));
 sg13g2_tiehi _25676__915 (.L_HI(net915));
 sg13g2_tiehi _25675__916 (.L_HI(net916));
 sg13g2_tiehi _25674__917 (.L_HI(net917));
 sg13g2_tiehi _25673__918 (.L_HI(net918));
 sg13g2_tiehi _25672__919 (.L_HI(net919));
 sg13g2_tiehi _25671__920 (.L_HI(net920));
 sg13g2_tiehi _25670__921 (.L_HI(net921));
 sg13g2_tiehi _25669__922 (.L_HI(net922));
 sg13g2_tiehi _25668__923 (.L_HI(net923));
 sg13g2_tiehi _25667__924 (.L_HI(net924));
 sg13g2_tiehi _25666__925 (.L_HI(net925));
 sg13g2_tiehi _25665__926 (.L_HI(net926));
 sg13g2_tiehi _25664__927 (.L_HI(net927));
 sg13g2_tiehi _25663__928 (.L_HI(net928));
 sg13g2_tiehi _25662__929 (.L_HI(net929));
 sg13g2_tiehi _25661__930 (.L_HI(net930));
 sg13g2_tiehi _25660__931 (.L_HI(net931));
 sg13g2_tiehi _25659__932 (.L_HI(net932));
 sg13g2_tiehi _25658__933 (.L_HI(net933));
 sg13g2_tiehi _25657__934 (.L_HI(net934));
 sg13g2_tiehi _25656__935 (.L_HI(net935));
 sg13g2_tiehi _25655__936 (.L_HI(net936));
 sg13g2_tiehi _25654__937 (.L_HI(net937));
 sg13g2_tiehi _25645__938 (.L_HI(net938));
 sg13g2_tiehi _25644__939 (.L_HI(net939));
 sg13g2_tiehi _25643__940 (.L_HI(net940));
 sg13g2_tiehi _25642__941 (.L_HI(net941));
 sg13g2_tiehi _25641__942 (.L_HI(net942));
 sg13g2_tiehi _25640__943 (.L_HI(net943));
 sg13g2_tiehi _25639__944 (.L_HI(net944));
 sg13g2_tiehi _25638__945 (.L_HI(net945));
 sg13g2_tiehi _25637__946 (.L_HI(net946));
 sg13g2_tiehi _25636__947 (.L_HI(net947));
 sg13g2_tiehi _25635__948 (.L_HI(net948));
 sg13g2_tiehi _25634__949 (.L_HI(net949));
 sg13g2_tiehi _25633__950 (.L_HI(net950));
 sg13g2_tiehi _25632__951 (.L_HI(net951));
 sg13g2_tiehi _25631__952 (.L_HI(net952));
 sg13g2_tiehi _25630__953 (.L_HI(net953));
 sg13g2_tiehi _25629__954 (.L_HI(net954));
 sg13g2_tiehi _25628__955 (.L_HI(net955));
 sg13g2_tiehi _25627__956 (.L_HI(net956));
 sg13g2_tiehi _25626__957 (.L_HI(net957));
 sg13g2_tiehi _25625__958 (.L_HI(net958));
 sg13g2_tiehi _25624__959 (.L_HI(net959));
 sg13g2_tiehi _25623__960 (.L_HI(net960));
 sg13g2_tiehi _25622__961 (.L_HI(net961));
 sg13g2_tiehi _25621__962 (.L_HI(net962));
 sg13g2_tiehi _25620__963 (.L_HI(net963));
 sg13g2_tiehi _25619__964 (.L_HI(net964));
 sg13g2_tiehi _25618__965 (.L_HI(net965));
 sg13g2_tiehi _25617__966 (.L_HI(net966));
 sg13g2_tiehi _25616__967 (.L_HI(net967));
 sg13g2_tiehi _25615__968 (.L_HI(net968));
 sg13g2_tiehi _25614__969 (.L_HI(net969));
 sg13g2_tiehi _25613__970 (.L_HI(net970));
 sg13g2_tiehi _25612__971 (.L_HI(net971));
 sg13g2_tiehi _25611__972 (.L_HI(net972));
 sg13g2_tiehi _25610__973 (.L_HI(net973));
 sg13g2_tiehi _25609__974 (.L_HI(net974));
 sg13g2_tiehi _25608__975 (.L_HI(net975));
 sg13g2_tiehi _25607__976 (.L_HI(net976));
 sg13g2_tiehi _25606__977 (.L_HI(net977));
 sg13g2_tiehi _25605__978 (.L_HI(net978));
 sg13g2_tiehi _25604__979 (.L_HI(net979));
 sg13g2_tiehi _25603__980 (.L_HI(net980));
 sg13g2_tiehi _25602__981 (.L_HI(net981));
 sg13g2_tiehi _25601__982 (.L_HI(net982));
 sg13g2_tiehi _25600__983 (.L_HI(net983));
 sg13g2_tiehi _25599__984 (.L_HI(net984));
 sg13g2_tiehi _25598__985 (.L_HI(net985));
 sg13g2_tiehi _25597__986 (.L_HI(net986));
 sg13g2_tiehi _25596__987 (.L_HI(net987));
 sg13g2_tiehi _25595__988 (.L_HI(net988));
 sg13g2_tiehi _25594__989 (.L_HI(net989));
 sg13g2_tiehi _25593__990 (.L_HI(net990));
 sg13g2_tiehi _25592__991 (.L_HI(net991));
 sg13g2_tiehi _25591__992 (.L_HI(net992));
 sg13g2_tiehi _25590__993 (.L_HI(net993));
 sg13g2_tiehi _25589__994 (.L_HI(net994));
 sg13g2_tiehi _25588__995 (.L_HI(net995));
 sg13g2_tiehi _25587__996 (.L_HI(net996));
 sg13g2_tiehi _25586__997 (.L_HI(net997));
 sg13g2_tiehi _25585__998 (.L_HI(net998));
 sg13g2_tiehi _25584__999 (.L_HI(net999));
 sg13g2_tiehi _25583__1000 (.L_HI(net1000));
 sg13g2_tiehi _25582__1001 (.L_HI(net1001));
 sg13g2_tiehi _25581__1002 (.L_HI(net1002));
 sg13g2_tiehi _24992__1003 (.L_HI(net1003));
 sg13g2_tiehi _25221__1004 (.L_HI(net1004));
 sg13g2_tiehi _25222__1005 (.L_HI(net1005));
 sg13g2_tiehi _25223__1006 (.L_HI(net1006));
 sg13g2_tiehi _25224__1007 (.L_HI(net1007));
 sg13g2_tiehi _25322__1008 (.L_HI(net1008));
 sg13g2_tiehi _25321__1009 (.L_HI(net1009));
 sg13g2_tiehi _25320__1010 (.L_HI(net1010));
 sg13g2_tiehi _25319__1011 (.L_HI(net1011));
 sg13g2_tiehi _25318__1012 (.L_HI(net1012));
 sg13g2_tiehi _25317__1013 (.L_HI(net1013));
 sg13g2_tiehi _25316__1014 (.L_HI(net1014));
 sg13g2_tiehi _25315__1015 (.L_HI(net1015));
 sg13g2_tiehi _25314__1016 (.L_HI(net1016));
 sg13g2_tiehi _25313__1017 (.L_HI(net1017));
 sg13g2_tiehi _25312__1018 (.L_HI(net1018));
 sg13g2_tiehi _25311__1019 (.L_HI(net1019));
 sg13g2_tiehi _25310__1020 (.L_HI(net1020));
 sg13g2_tiehi _25309__1021 (.L_HI(net1021));
 sg13g2_tiehi _25308__1022 (.L_HI(net1022));
 sg13g2_tiehi _25307__1023 (.L_HI(net1023));
 sg13g2_tiehi _25306__1024 (.L_HI(net1024));
 sg13g2_tiehi _25305__1025 (.L_HI(net1025));
 sg13g2_tiehi _25304__1026 (.L_HI(net1026));
 sg13g2_tiehi _25303__1027 (.L_HI(net1027));
 sg13g2_tiehi _25302__1028 (.L_HI(net1028));
 sg13g2_tiehi _25301__1029 (.L_HI(net1029));
 sg13g2_tiehi _25300__1030 (.L_HI(net1030));
 sg13g2_tiehi _25299__1031 (.L_HI(net1031));
 sg13g2_tiehi _25298__1032 (.L_HI(net1032));
 sg13g2_tiehi _25297__1033 (.L_HI(net1033));
 sg13g2_tiehi _25296__1034 (.L_HI(net1034));
 sg13g2_tiehi _25295__1035 (.L_HI(net1035));
 sg13g2_tiehi _25294__1036 (.L_HI(net1036));
 sg13g2_tiehi _25293__1037 (.L_HI(net1037));
 sg13g2_tiehi _25292__1038 (.L_HI(net1038));
 sg13g2_tiehi _25291__1039 (.L_HI(net1039));
 sg13g2_tiehi _25290__1040 (.L_HI(net1040));
 sg13g2_tiehi _25289__1041 (.L_HI(net1041));
 sg13g2_tiehi _25288__1042 (.L_HI(net1042));
 sg13g2_tiehi _25287__1043 (.L_HI(net1043));
 sg13g2_tiehi _25286__1044 (.L_HI(net1044));
 sg13g2_tiehi _25285__1045 (.L_HI(net1045));
 sg13g2_tiehi _25284__1046 (.L_HI(net1046));
 sg13g2_tiehi _25283__1047 (.L_HI(net1047));
 sg13g2_tiehi _25282__1048 (.L_HI(net1048));
 sg13g2_tiehi _25281__1049 (.L_HI(net1049));
 sg13g2_tiehi _25280__1050 (.L_HI(net1050));
 sg13g2_tiehi _25279__1051 (.L_HI(net1051));
 sg13g2_tiehi _25278__1052 (.L_HI(net1052));
 sg13g2_tiehi _25277__1053 (.L_HI(net1053));
 sg13g2_tiehi _25276__1054 (.L_HI(net1054));
 sg13g2_tiehi _25275__1055 (.L_HI(net1055));
 sg13g2_tiehi _25274__1056 (.L_HI(net1056));
 sg13g2_tiehi _25273__1057 (.L_HI(net1057));
 sg13g2_tiehi _25272__1058 (.L_HI(net1058));
 sg13g2_tiehi _25271__1059 (.L_HI(net1059));
 sg13g2_tiehi _25270__1060 (.L_HI(net1060));
 sg13g2_tiehi _25269__1061 (.L_HI(net1061));
 sg13g2_tiehi _25268__1062 (.L_HI(net1062));
 sg13g2_tiehi _25267__1063 (.L_HI(net1063));
 sg13g2_tiehi _25266__1064 (.L_HI(net1064));
 sg13g2_tiehi _25265__1065 (.L_HI(net1065));
 sg13g2_tiehi _25264__1066 (.L_HI(net1066));
 sg13g2_tiehi _25263__1067 (.L_HI(net1067));
 sg13g2_tiehi _25262__1068 (.L_HI(net1068));
 sg13g2_tiehi _25261__1069 (.L_HI(net1069));
 sg13g2_tiehi _25260__1070 (.L_HI(net1070));
 sg13g2_tiehi _25259__1071 (.L_HI(net1071));
 sg13g2_tiehi _25258__1072 (.L_HI(net1072));
 sg13g2_tiehi _25257__1073 (.L_HI(net1073));
 sg13g2_tiehi _25256__1074 (.L_HI(net1074));
 sg13g2_tiehi _25255__1075 (.L_HI(net1075));
 sg13g2_tiehi _25254__1076 (.L_HI(net1076));
 sg13g2_tiehi _25253__1077 (.L_HI(net1077));
 sg13g2_tiehi _25252__1078 (.L_HI(net1078));
 sg13g2_tiehi _25251__1079 (.L_HI(net1079));
 sg13g2_tiehi _25250__1080 (.L_HI(net1080));
 sg13g2_tiehi _25249__1081 (.L_HI(net1081));
 sg13g2_tiehi _25248__1082 (.L_HI(net1082));
 sg13g2_tiehi _25247__1083 (.L_HI(net1083));
 sg13g2_tiehi _25246__1084 (.L_HI(net1084));
 sg13g2_tiehi _25245__1085 (.L_HI(net1085));
 sg13g2_tiehi _25244__1086 (.L_HI(net1086));
 sg13g2_tiehi _25243__1087 (.L_HI(net1087));
 sg13g2_tiehi _25242__1088 (.L_HI(net1088));
 sg13g2_tiehi _25241__1089 (.L_HI(net1089));
 sg13g2_tiehi _25240__1090 (.L_HI(net1090));
 sg13g2_tiehi _25239__1091 (.L_HI(net1091));
 sg13g2_tiehi _25238__1092 (.L_HI(net1092));
 sg13g2_tiehi _25237__1093 (.L_HI(net1093));
 sg13g2_tiehi _25236__1094 (.L_HI(net1094));
 sg13g2_tiehi _25235__1095 (.L_HI(net1095));
 sg13g2_tiehi _25234__1096 (.L_HI(net1096));
 sg13g2_tiehi _25233__1097 (.L_HI(net1097));
 sg13g2_tiehi _25232__1098 (.L_HI(net1098));
 sg13g2_tiehi _25231__1099 (.L_HI(net1099));
 sg13g2_tiehi _25230__1100 (.L_HI(net1100));
 sg13g2_tiehi _25229__1101 (.L_HI(net1101));
 sg13g2_tiehi _25228__1102 (.L_HI(net1102));
 sg13g2_tiehi _25227__1103 (.L_HI(net1103));
 sg13g2_tiehi _25226__1104 (.L_HI(net1104));
 sg13g2_tiehi _25220__1105 (.L_HI(net1105));
 sg13g2_tiehi _25219__1106 (.L_HI(net1106));
 sg13g2_tiehi _25218__1107 (.L_HI(net1107));
 sg13g2_tiehi _25217__1108 (.L_HI(net1108));
 sg13g2_tiehi _25216__1109 (.L_HI(net1109));
 sg13g2_tiehi _25215__1110 (.L_HI(net1110));
 sg13g2_tiehi _25214__1111 (.L_HI(net1111));
 sg13g2_tiehi _25213__1112 (.L_HI(net1112));
 sg13g2_tiehi _25212__1113 (.L_HI(net1113));
 sg13g2_tiehi _25211__1114 (.L_HI(net1114));
 sg13g2_tiehi _25210__1115 (.L_HI(net1115));
 sg13g2_tiehi _25209__1116 (.L_HI(net1116));
 sg13g2_tiehi _25208__1117 (.L_HI(net1117));
 sg13g2_tiehi _25207__1118 (.L_HI(net1118));
 sg13g2_tiehi _25206__1119 (.L_HI(net1119));
 sg13g2_tiehi _25205__1120 (.L_HI(net1120));
 sg13g2_tiehi _25204__1121 (.L_HI(net1121));
 sg13g2_tiehi _25203__1122 (.L_HI(net1122));
 sg13g2_tiehi _25202__1123 (.L_HI(net1123));
 sg13g2_tiehi _25201__1124 (.L_HI(net1124));
 sg13g2_tiehi _25200__1125 (.L_HI(net1125));
 sg13g2_tiehi _25199__1126 (.L_HI(net1126));
 sg13g2_tiehi _25198__1127 (.L_HI(net1127));
 sg13g2_tiehi _25197__1128 (.L_HI(net1128));
 sg13g2_tiehi _25196__1129 (.L_HI(net1129));
 sg13g2_tiehi _25195__1130 (.L_HI(net1130));
 sg13g2_tiehi _25194__1131 (.L_HI(net1131));
 sg13g2_tiehi _25193__1132 (.L_HI(net1132));
 sg13g2_tiehi _25192__1133 (.L_HI(net1133));
 sg13g2_tiehi _25191__1134 (.L_HI(net1134));
 sg13g2_tiehi _25190__1135 (.L_HI(net1135));
 sg13g2_tiehi _25189__1136 (.L_HI(net1136));
 sg13g2_tiehi _25188__1137 (.L_HI(net1137));
 sg13g2_tiehi _25187__1138 (.L_HI(net1138));
 sg13g2_tiehi _25186__1139 (.L_HI(net1139));
 sg13g2_tiehi _25185__1140 (.L_HI(net1140));
 sg13g2_tiehi _25184__1141 (.L_HI(net1141));
 sg13g2_tiehi _25183__1142 (.L_HI(net1142));
 sg13g2_tiehi _25182__1143 (.L_HI(net1143));
 sg13g2_tiehi _25181__1144 (.L_HI(net1144));
 sg13g2_tiehi _25180__1145 (.L_HI(net1145));
 sg13g2_tiehi _25179__1146 (.L_HI(net1146));
 sg13g2_tiehi _25178__1147 (.L_HI(net1147));
 sg13g2_tiehi _25177__1148 (.L_HI(net1148));
 sg13g2_tiehi _25176__1149 (.L_HI(net1149));
 sg13g2_tiehi _25175__1150 (.L_HI(net1150));
 sg13g2_tiehi _25174__1151 (.L_HI(net1151));
 sg13g2_tiehi _25173__1152 (.L_HI(net1152));
 sg13g2_tiehi _25172__1153 (.L_HI(net1153));
 sg13g2_tiehi _25171__1154 (.L_HI(net1154));
 sg13g2_tiehi _25170__1155 (.L_HI(net1155));
 sg13g2_tiehi _25169__1156 (.L_HI(net1156));
 sg13g2_tiehi _25168__1157 (.L_HI(net1157));
 sg13g2_tiehi _25167__1158 (.L_HI(net1158));
 sg13g2_tiehi _25166__1159 (.L_HI(net1159));
 sg13g2_tiehi _25165__1160 (.L_HI(net1160));
 sg13g2_tiehi _25164__1161 (.L_HI(net1161));
 sg13g2_tiehi _25163__1162 (.L_HI(net1162));
 sg13g2_tiehi _25162__1163 (.L_HI(net1163));
 sg13g2_tiehi _25161__1164 (.L_HI(net1164));
 sg13g2_tiehi _25160__1165 (.L_HI(net1165));
 sg13g2_tiehi _25159__1166 (.L_HI(net1166));
 sg13g2_tiehi _25158__1167 (.L_HI(net1167));
 sg13g2_tiehi _25157__1168 (.L_HI(net1168));
 sg13g2_tiehi _25156__1169 (.L_HI(net1169));
 sg13g2_tiehi _25155__1170 (.L_HI(net1170));
 sg13g2_tiehi _25154__1171 (.L_HI(net1171));
 sg13g2_tiehi _25153__1172 (.L_HI(net1172));
 sg13g2_tiehi _25152__1173 (.L_HI(net1173));
 sg13g2_tiehi _25151__1174 (.L_HI(net1174));
 sg13g2_tiehi _25150__1175 (.L_HI(net1175));
 sg13g2_tiehi _25149__1176 (.L_HI(net1176));
 sg13g2_tiehi _25148__1177 (.L_HI(net1177));
 sg13g2_tiehi _25147__1178 (.L_HI(net1178));
 sg13g2_tiehi _25146__1179 (.L_HI(net1179));
 sg13g2_tiehi _25145__1180 (.L_HI(net1180));
 sg13g2_tiehi _25144__1181 (.L_HI(net1181));
 sg13g2_tiehi _25143__1182 (.L_HI(net1182));
 sg13g2_tiehi _25142__1183 (.L_HI(net1183));
 sg13g2_tiehi _25141__1184 (.L_HI(net1184));
 sg13g2_tiehi _25140__1185 (.L_HI(net1185));
 sg13g2_tiehi _25139__1186 (.L_HI(net1186));
 sg13g2_tiehi _25138__1187 (.L_HI(net1187));
 sg13g2_tiehi _25137__1188 (.L_HI(net1188));
 sg13g2_tiehi _25136__1189 (.L_HI(net1189));
 sg13g2_tiehi _25135__1190 (.L_HI(net1190));
 sg13g2_tiehi _25134__1191 (.L_HI(net1191));
 sg13g2_tiehi _25133__1192 (.L_HI(net1192));
 sg13g2_tiehi _25132__1193 (.L_HI(net1193));
 sg13g2_tiehi _25131__1194 (.L_HI(net1194));
 sg13g2_tiehi _25130__1195 (.L_HI(net1195));
 sg13g2_tiehi _25129__1196 (.L_HI(net1196));
 sg13g2_tiehi _25128__1197 (.L_HI(net1197));
 sg13g2_tiehi _25127__1198 (.L_HI(net1198));
 sg13g2_tiehi _25126__1199 (.L_HI(net1199));
 sg13g2_tiehi _25125__1200 (.L_HI(net1200));
 sg13g2_tiehi _25124__1201 (.L_HI(net1201));
 sg13g2_tiehi _25123__1202 (.L_HI(net1202));
 sg13g2_tiehi _25122__1203 (.L_HI(net1203));
 sg13g2_tiehi _25121__1204 (.L_HI(net1204));
 sg13g2_tiehi _25120__1205 (.L_HI(net1205));
 sg13g2_tiehi _25119__1206 (.L_HI(net1206));
 sg13g2_tiehi _25118__1207 (.L_HI(net1207));
 sg13g2_tiehi _25117__1208 (.L_HI(net1208));
 sg13g2_tiehi _25116__1209 (.L_HI(net1209));
 sg13g2_tiehi _25115__1210 (.L_HI(net1210));
 sg13g2_tiehi _25114__1211 (.L_HI(net1211));
 sg13g2_tiehi _25113__1212 (.L_HI(net1212));
 sg13g2_tiehi _25112__1213 (.L_HI(net1213));
 sg13g2_tiehi _25111__1214 (.L_HI(net1214));
 sg13g2_tiehi _25110__1215 (.L_HI(net1215));
 sg13g2_tiehi _25109__1216 (.L_HI(net1216));
 sg13g2_tiehi _25108__1217 (.L_HI(net1217));
 sg13g2_tiehi _25107__1218 (.L_HI(net1218));
 sg13g2_tiehi _25106__1219 (.L_HI(net1219));
 sg13g2_tiehi _25105__1220 (.L_HI(net1220));
 sg13g2_tiehi _25104__1221 (.L_HI(net1221));
 sg13g2_tiehi _25103__1222 (.L_HI(net1222));
 sg13g2_tiehi _25102__1223 (.L_HI(net1223));
 sg13g2_tiehi _25101__1224 (.L_HI(net1224));
 sg13g2_tiehi _25100__1225 (.L_HI(net1225));
 sg13g2_tiehi _25099__1226 (.L_HI(net1226));
 sg13g2_tiehi _25098__1227 (.L_HI(net1227));
 sg13g2_tiehi _25097__1228 (.L_HI(net1228));
 sg13g2_tiehi _25096__1229 (.L_HI(net1229));
 sg13g2_tiehi _25095__1230 (.L_HI(net1230));
 sg13g2_tiehi _25094__1231 (.L_HI(net1231));
 sg13g2_tiehi _25225__1232 (.L_HI(net1232));
 sg13g2_tiehi _25579__1233 (.L_HI(net1233));
 sg13g2_tiehi _24991__1234 (.L_HI(net1234));
 sg13g2_tiehi _24990__1235 (.L_HI(net1235));
 sg13g2_tiehi _24989__1236 (.L_HI(net1236));
 sg13g2_tiehi _24988__1237 (.L_HI(net1237));
 sg13g2_tiehi _24987__1238 (.L_HI(net1238));
 sg13g2_tiehi _24986__1239 (.L_HI(net1239));
 sg13g2_tiehi _24985__1240 (.L_HI(net1240));
 sg13g2_tiehi _24984__1241 (.L_HI(net1241));
 sg13g2_tiehi _24983__1242 (.L_HI(net1242));
 sg13g2_tiehi _24982__1243 (.L_HI(net1243));
 sg13g2_tiehi _24981__1244 (.L_HI(net1244));
 sg13g2_tiehi _24980__1245 (.L_HI(net1245));
 sg13g2_tiehi _24979__1246 (.L_HI(net1246));
 sg13g2_tiehi _24978__1247 (.L_HI(net1247));
 sg13g2_tiehi _24977__1248 (.L_HI(net1248));
 sg13g2_tiehi _24976__1249 (.L_HI(net1249));
 sg13g2_tiehi _24975__1250 (.L_HI(net1250));
 sg13g2_tiehi _24974__1251 (.L_HI(net1251));
 sg13g2_tiehi _24973__1252 (.L_HI(net1252));
 sg13g2_tiehi _24972__1253 (.L_HI(net1253));
 sg13g2_tiehi _24971__1254 (.L_HI(net1254));
 sg13g2_tiehi _24970__1255 (.L_HI(net1255));
 sg13g2_tiehi _24969__1256 (.L_HI(net1256));
 sg13g2_tiehi _24968__1257 (.L_HI(net1257));
 sg13g2_tiehi _24967__1258 (.L_HI(net1258));
 sg13g2_tiehi _24966__1259 (.L_HI(net1259));
 sg13g2_tiehi _24965__1260 (.L_HI(net1260));
 sg13g2_tiehi _24964__1261 (.L_HI(net1261));
 sg13g2_tiehi _24963__1262 (.L_HI(net1262));
 sg13g2_tiehi _24962__1263 (.L_HI(net1263));
 sg13g2_tiehi _24961__1264 (.L_HI(net1264));
 sg13g2_tiehi _24960__1265 (.L_HI(net1265));
 sg13g2_tiehi _24959__1266 (.L_HI(net1266));
 sg13g2_tiehi _24958__1267 (.L_HI(net1267));
 sg13g2_tiehi _24957__1268 (.L_HI(net1268));
 sg13g2_tiehi _24956__1269 (.L_HI(net1269));
 sg13g2_tiehi _24955__1270 (.L_HI(net1270));
 sg13g2_tiehi _24954__1271 (.L_HI(net1271));
 sg13g2_tiehi _24953__1272 (.L_HI(net1272));
 sg13g2_tiehi _24952__1273 (.L_HI(net1273));
 sg13g2_tiehi _24951__1274 (.L_HI(net1274));
 sg13g2_tiehi _24950__1275 (.L_HI(net1275));
 sg13g2_tiehi _24949__1276 (.L_HI(net1276));
 sg13g2_tiehi _24948__1277 (.L_HI(net1277));
 sg13g2_tiehi _24947__1278 (.L_HI(net1278));
 sg13g2_tiehi _24946__1279 (.L_HI(net1279));
 sg13g2_tiehi _24945__1280 (.L_HI(net1280));
 sg13g2_tiehi _24944__1281 (.L_HI(net1281));
 sg13g2_tiehi _24943__1282 (.L_HI(net1282));
 sg13g2_tiehi _24942__1283 (.L_HI(net1283));
 sg13g2_tiehi _24941__1284 (.L_HI(net1284));
 sg13g2_tiehi _24940__1285 (.L_HI(net1285));
 sg13g2_tiehi _24939__1286 (.L_HI(net1286));
 sg13g2_tiehi _24938__1287 (.L_HI(net1287));
 sg13g2_tiehi _24937__1288 (.L_HI(net1288));
 sg13g2_tiehi _24936__1289 (.L_HI(net1289));
 sg13g2_tiehi _24935__1290 (.L_HI(net1290));
 sg13g2_tiehi _24934__1291 (.L_HI(net1291));
 sg13g2_tiehi _24933__1292 (.L_HI(net1292));
 sg13g2_tiehi _24932__1293 (.L_HI(net1293));
 sg13g2_tiehi _24931__1294 (.L_HI(net1294));
 sg13g2_tiehi _24930__1295 (.L_HI(net1295));
 sg13g2_tiehi _24929__1296 (.L_HI(net1296));
 sg13g2_tiehi _25580__1297 (.L_HI(net1297));
 sg13g2_tiehi _25717__1298 (.L_HI(net1298));
 sg13g2_tiehi _25718__1299 (.L_HI(net1299));
 sg13g2_tiehi _25786__1300 (.L_HI(net1300));
 sg13g2_tiehi _25974__1301 (.L_HI(net1301));
 sg13g2_tiehi _24856__1302 (.L_HI(net1302));
 sg13g2_tiehi _24855__1303 (.L_HI(net1303));
 sg13g2_tiehi _24854__1304 (.L_HI(net1304));
 sg13g2_tiehi _24853__1305 (.L_HI(net1305));
 sg13g2_tiehi _24852__1306 (.L_HI(net1306));
 sg13g2_tiehi _24851__1307 (.L_HI(net1307));
 sg13g2_tiehi _24850__1308 (.L_HI(net1308));
 sg13g2_tiehi _24849__1309 (.L_HI(net1309));
 sg13g2_tiehi _25719__1310 (.L_HI(net1310));
 sg13g2_tiehi _25784__1311 (.L_HI(net1311));
 sg13g2_tiehi _25785__1312 (.L_HI(net1312));
 sg13g2_tiehi _25973__1313 (.L_HI(net1313));
 sg13g2_tiehi _24857__1314 (.L_HI(net1314));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_8 _27273_ (.A(\fpga_top.qspi_if.sio_en ),
    .X(uio_oe[0]));
 sg13g2_buf_8 _27274_ (.A(\fpga_top.qspi_if.sio_en ),
    .X(uio_oe[1]));
 sg13g2_buf_8 _27275_ (.A(\fpga_top.qspi_if.sio_en ),
    .X(uio_oe[2]));
 sg13g2_buf_8 _27276_ (.A(\fpga_top.qspi_if.sio_en ),
    .X(uio_oe[3]));
 sg13g2_buf_1 _27277_ (.A(\fpga_top.tx ),
    .X(uo_out[0]));
 sg13g2_buf_8 _27278_ (.A(\fpga_top.qspi_if.sck ),
    .X(uo_out[4]));
 sg13g2_buf_8 fanout4075 (.A(_06496_),
    .X(net4075));
 sg13g2_buf_8 fanout4076 (.A(_06496_),
    .X(net4076));
 sg13g2_buf_8 fanout4077 (.A(net4079),
    .X(net4077));
 sg13g2_buf_8 fanout4078 (.A(net4079),
    .X(net4078));
 sg13g2_buf_8 fanout4079 (.A(_06496_),
    .X(net4079));
 sg13g2_buf_8 fanout4080 (.A(_06495_),
    .X(net4080));
 sg13g2_buf_8 fanout4081 (.A(_06495_),
    .X(net4081));
 sg13g2_buf_8 fanout4082 (.A(net4084),
    .X(net4082));
 sg13g2_buf_8 fanout4083 (.A(net4084),
    .X(net4083));
 sg13g2_buf_8 fanout4084 (.A(_06495_),
    .X(net4084));
 sg13g2_buf_8 fanout4085 (.A(_05326_),
    .X(net4085));
 sg13g2_buf_8 fanout4086 (.A(_05326_),
    .X(net4086));
 sg13g2_buf_8 fanout4087 (.A(net4089),
    .X(net4087));
 sg13g2_buf_8 fanout4088 (.A(net4089),
    .X(net4088));
 sg13g2_buf_8 fanout4089 (.A(_05326_),
    .X(net4089));
 sg13g2_buf_8 fanout4090 (.A(net4091),
    .X(net4090));
 sg13g2_buf_8 fanout4091 (.A(_05325_),
    .X(net4091));
 sg13g2_buf_8 fanout4092 (.A(net4094),
    .X(net4092));
 sg13g2_buf_8 fanout4093 (.A(net4094),
    .X(net4093));
 sg13g2_buf_8 fanout4094 (.A(_05325_),
    .X(net4094));
 sg13g2_buf_8 fanout4095 (.A(_05324_),
    .X(net4095));
 sg13g2_buf_8 fanout4096 (.A(_05324_),
    .X(net4096));
 sg13g2_buf_8 fanout4097 (.A(net4099),
    .X(net4097));
 sg13g2_buf_8 fanout4098 (.A(net4099),
    .X(net4098));
 sg13g2_buf_8 fanout4099 (.A(_05324_),
    .X(net4099));
 sg13g2_buf_8 fanout4100 (.A(_05323_),
    .X(net4100));
 sg13g2_buf_8 fanout4101 (.A(_05323_),
    .X(net4101));
 sg13g2_buf_8 fanout4102 (.A(net4104),
    .X(net4102));
 sg13g2_buf_8 fanout4103 (.A(net4104),
    .X(net4103));
 sg13g2_buf_8 fanout4104 (.A(_05323_),
    .X(net4104));
 sg13g2_buf_8 fanout4105 (.A(net4106),
    .X(net4105));
 sg13g2_buf_8 fanout4106 (.A(_05322_),
    .X(net4106));
 sg13g2_buf_8 fanout4107 (.A(net4109),
    .X(net4107));
 sg13g2_buf_8 fanout4108 (.A(net4109),
    .X(net4108));
 sg13g2_buf_8 fanout4109 (.A(_05322_),
    .X(net4109));
 sg13g2_buf_8 fanout4110 (.A(_05321_),
    .X(net4110));
 sg13g2_buf_8 fanout4111 (.A(_05321_),
    .X(net4111));
 sg13g2_buf_8 fanout4112 (.A(net4114),
    .X(net4112));
 sg13g2_buf_8 fanout4113 (.A(net4114),
    .X(net4113));
 sg13g2_buf_8 fanout4114 (.A(_05321_),
    .X(net4114));
 sg13g2_buf_8 fanout4115 (.A(_05320_),
    .X(net4115));
 sg13g2_buf_8 fanout4116 (.A(_05320_),
    .X(net4116));
 sg13g2_buf_8 fanout4117 (.A(net4119),
    .X(net4117));
 sg13g2_buf_8 fanout4118 (.A(net4119),
    .X(net4118));
 sg13g2_buf_8 fanout4119 (.A(_05320_),
    .X(net4119));
 sg13g2_buf_8 fanout4120 (.A(net4121),
    .X(net4120));
 sg13g2_buf_8 fanout4121 (.A(_05238_),
    .X(net4121));
 sg13g2_buf_8 fanout4122 (.A(net4124),
    .X(net4122));
 sg13g2_buf_8 fanout4123 (.A(net4124),
    .X(net4123));
 sg13g2_buf_8 fanout4124 (.A(_05238_),
    .X(net4124));
 sg13g2_buf_8 fanout4125 (.A(net4126),
    .X(net4125));
 sg13g2_buf_8 fanout4126 (.A(_05237_),
    .X(net4126));
 sg13g2_buf_8 fanout4127 (.A(net4129),
    .X(net4127));
 sg13g2_buf_8 fanout4128 (.A(net4129),
    .X(net4128));
 sg13g2_buf_8 fanout4129 (.A(_05237_),
    .X(net4129));
 sg13g2_buf_8 fanout4130 (.A(net4131),
    .X(net4130));
 sg13g2_buf_8 fanout4131 (.A(_04249_),
    .X(net4131));
 sg13g2_buf_8 fanout4132 (.A(net4134),
    .X(net4132));
 sg13g2_buf_8 fanout4133 (.A(net4134),
    .X(net4133));
 sg13g2_buf_8 fanout4134 (.A(_04249_),
    .X(net4134));
 sg13g2_buf_8 fanout4135 (.A(_03193_),
    .X(net4135));
 sg13g2_buf_8 fanout4136 (.A(_03193_),
    .X(net4136));
 sg13g2_buf_8 fanout4137 (.A(net4139),
    .X(net4137));
 sg13g2_buf_8 fanout4138 (.A(net4139),
    .X(net4138));
 sg13g2_buf_8 fanout4139 (.A(_03193_),
    .X(net4139));
 sg13g2_buf_8 fanout4140 (.A(_03192_),
    .X(net4140));
 sg13g2_buf_8 fanout4141 (.A(_03192_),
    .X(net4141));
 sg13g2_buf_8 fanout4142 (.A(net4144),
    .X(net4142));
 sg13g2_buf_8 fanout4143 (.A(net4144),
    .X(net4143));
 sg13g2_buf_8 fanout4144 (.A(_03192_),
    .X(net4144));
 sg13g2_buf_8 fanout4145 (.A(_03190_),
    .X(net4145));
 sg13g2_buf_8 fanout4146 (.A(_03190_),
    .X(net4146));
 sg13g2_buf_8 fanout4147 (.A(net4149),
    .X(net4147));
 sg13g2_buf_8 fanout4148 (.A(net4149),
    .X(net4148));
 sg13g2_buf_8 fanout4149 (.A(_03190_),
    .X(net4149));
 sg13g2_buf_8 fanout4150 (.A(_03183_),
    .X(net4150));
 sg13g2_buf_8 fanout4151 (.A(_03183_),
    .X(net4151));
 sg13g2_buf_8 fanout4152 (.A(net4154),
    .X(net4152));
 sg13g2_buf_8 fanout4153 (.A(net4154),
    .X(net4153));
 sg13g2_buf_8 fanout4154 (.A(_03183_),
    .X(net4154));
 sg13g2_buf_8 fanout4155 (.A(_03181_),
    .X(net4155));
 sg13g2_buf_8 fanout4156 (.A(_03181_),
    .X(net4156));
 sg13g2_buf_8 fanout4157 (.A(net4159),
    .X(net4157));
 sg13g2_buf_8 fanout4158 (.A(net4159),
    .X(net4158));
 sg13g2_buf_8 fanout4159 (.A(_03181_),
    .X(net4159));
 sg13g2_buf_8 fanout4160 (.A(_03172_),
    .X(net4160));
 sg13g2_buf_8 fanout4161 (.A(_03172_),
    .X(net4161));
 sg13g2_buf_8 fanout4162 (.A(net4164),
    .X(net4162));
 sg13g2_buf_8 fanout4163 (.A(net4164),
    .X(net4163));
 sg13g2_buf_8 fanout4164 (.A(_03172_),
    .X(net4164));
 sg13g2_buf_8 fanout4165 (.A(_03171_),
    .X(net4165));
 sg13g2_buf_8 fanout4166 (.A(_03171_),
    .X(net4166));
 sg13g2_buf_8 fanout4167 (.A(net4169),
    .X(net4167));
 sg13g2_buf_8 fanout4168 (.A(net4169),
    .X(net4168));
 sg13g2_buf_8 fanout4169 (.A(_03171_),
    .X(net4169));
 sg13g2_buf_8 fanout4170 (.A(_03170_),
    .X(net4170));
 sg13g2_buf_8 fanout4171 (.A(_03170_),
    .X(net4171));
 sg13g2_buf_8 fanout4172 (.A(net4174),
    .X(net4172));
 sg13g2_buf_8 fanout4173 (.A(net4174),
    .X(net4173));
 sg13g2_buf_8 fanout4174 (.A(_03170_),
    .X(net4174));
 sg13g2_buf_8 fanout4175 (.A(net4176),
    .X(net4175));
 sg13g2_buf_8 fanout4176 (.A(_02994_),
    .X(net4176));
 sg13g2_buf_8 fanout4177 (.A(net4179),
    .X(net4177));
 sg13g2_buf_8 fanout4178 (.A(net4179),
    .X(net4178));
 sg13g2_buf_8 fanout4179 (.A(_02994_),
    .X(net4179));
 sg13g2_buf_8 fanout4180 (.A(net4181),
    .X(net4180));
 sg13g2_buf_8 fanout4181 (.A(_10583_),
    .X(net4181));
 sg13g2_buf_8 fanout4182 (.A(net4184),
    .X(net4182));
 sg13g2_buf_8 fanout4183 (.A(net4184),
    .X(net4183));
 sg13g2_buf_8 fanout4184 (.A(_10583_),
    .X(net4184));
 sg13g2_buf_8 fanout4185 (.A(net4186),
    .X(net4185));
 sg13g2_buf_8 fanout4186 (.A(_10353_),
    .X(net4186));
 sg13g2_buf_8 fanout4187 (.A(net4189),
    .X(net4187));
 sg13g2_buf_8 fanout4188 (.A(net4189),
    .X(net4188));
 sg13g2_buf_8 fanout4189 (.A(_10353_),
    .X(net4189));
 sg13g2_buf_8 fanout4190 (.A(net4194),
    .X(net4190));
 sg13g2_buf_8 fanout4191 (.A(net4194),
    .X(net4191));
 sg13g2_buf_8 fanout4192 (.A(net4194),
    .X(net4192));
 sg13g2_buf_2 fanout4193 (.A(net4194),
    .X(net4193));
 sg13g2_buf_8 fanout4194 (.A(_10339_),
    .X(net4194));
 sg13g2_buf_8 fanout4195 (.A(net4196),
    .X(net4195));
 sg13g2_buf_8 fanout4196 (.A(net4199),
    .X(net4196));
 sg13g2_buf_8 fanout4197 (.A(net4198),
    .X(net4197));
 sg13g2_buf_8 fanout4198 (.A(net4199),
    .X(net4198));
 sg13g2_buf_8 fanout4199 (.A(_10199_),
    .X(net4199));
 sg13g2_buf_8 fanout4200 (.A(net4201),
    .X(net4200));
 sg13g2_buf_8 fanout4201 (.A(_09806_),
    .X(net4201));
 sg13g2_buf_8 fanout4202 (.A(net4204),
    .X(net4202));
 sg13g2_buf_8 fanout4203 (.A(net4204),
    .X(net4203));
 sg13g2_buf_8 fanout4204 (.A(_09806_),
    .X(net4204));
 sg13g2_buf_8 fanout4205 (.A(_09669_),
    .X(net4205));
 sg13g2_buf_8 fanout4206 (.A(_09669_),
    .X(net4206));
 sg13g2_buf_8 fanout4207 (.A(net4209),
    .X(net4207));
 sg13g2_buf_8 fanout4208 (.A(net4209),
    .X(net4208));
 sg13g2_buf_8 fanout4209 (.A(_09669_),
    .X(net4209));
 sg13g2_buf_8 fanout4210 (.A(_06485_),
    .X(net4210));
 sg13g2_buf_8 fanout4211 (.A(_06485_),
    .X(net4211));
 sg13g2_buf_8 fanout4212 (.A(net4214),
    .X(net4212));
 sg13g2_buf_8 fanout4213 (.A(net4214),
    .X(net4213));
 sg13g2_buf_8 fanout4214 (.A(_06485_),
    .X(net4214));
 sg13g2_buf_8 fanout4215 (.A(net4218),
    .X(net4215));
 sg13g2_buf_8 fanout4216 (.A(net4218),
    .X(net4216));
 sg13g2_buf_1 fanout4217 (.A(net4218),
    .X(net4217));
 sg13g2_buf_8 fanout4218 (.A(_06091_),
    .X(net4218));
 sg13g2_buf_8 fanout4219 (.A(_03189_),
    .X(net4219));
 sg13g2_buf_8 fanout4220 (.A(_03189_),
    .X(net4220));
 sg13g2_buf_8 fanout4221 (.A(net4223),
    .X(net4221));
 sg13g2_buf_8 fanout4222 (.A(net4223),
    .X(net4222));
 sg13g2_buf_8 fanout4223 (.A(_03189_),
    .X(net4223));
 sg13g2_buf_8 fanout4224 (.A(_03188_),
    .X(net4224));
 sg13g2_buf_8 fanout4225 (.A(_03188_),
    .X(net4225));
 sg13g2_buf_8 fanout4226 (.A(net4228),
    .X(net4226));
 sg13g2_buf_8 fanout4227 (.A(net4228),
    .X(net4227));
 sg13g2_buf_8 fanout4228 (.A(_03188_),
    .X(net4228));
 sg13g2_buf_8 fanout4229 (.A(_03187_),
    .X(net4229));
 sg13g2_buf_8 fanout4230 (.A(_03187_),
    .X(net4230));
 sg13g2_buf_8 fanout4231 (.A(net4233),
    .X(net4231));
 sg13g2_buf_8 fanout4232 (.A(net4233),
    .X(net4232));
 sg13g2_buf_8 fanout4233 (.A(_03187_),
    .X(net4233));
 sg13g2_buf_8 fanout4234 (.A(_03186_),
    .X(net4234));
 sg13g2_buf_8 fanout4235 (.A(_03186_),
    .X(net4235));
 sg13g2_buf_8 fanout4236 (.A(net4238),
    .X(net4236));
 sg13g2_buf_8 fanout4237 (.A(net4238),
    .X(net4237));
 sg13g2_buf_8 fanout4238 (.A(_03186_),
    .X(net4238));
 sg13g2_buf_8 fanout4239 (.A(_03184_),
    .X(net4239));
 sg13g2_buf_8 fanout4240 (.A(_03184_),
    .X(net4240));
 sg13g2_buf_8 fanout4241 (.A(net4243),
    .X(net4241));
 sg13g2_buf_8 fanout4242 (.A(net4243),
    .X(net4242));
 sg13g2_buf_8 fanout4243 (.A(_03184_),
    .X(net4243));
 sg13g2_buf_8 fanout4244 (.A(_03182_),
    .X(net4244));
 sg13g2_buf_8 fanout4245 (.A(_03182_),
    .X(net4245));
 sg13g2_buf_8 fanout4246 (.A(net4248),
    .X(net4246));
 sg13g2_buf_8 fanout4247 (.A(net4248),
    .X(net4247));
 sg13g2_buf_8 fanout4248 (.A(_03182_),
    .X(net4248));
 sg13g2_buf_8 fanout4249 (.A(_03180_),
    .X(net4249));
 sg13g2_buf_8 fanout4250 (.A(_03180_),
    .X(net4250));
 sg13g2_buf_8 fanout4251 (.A(net4253),
    .X(net4251));
 sg13g2_buf_8 fanout4252 (.A(net4253),
    .X(net4252));
 sg13g2_buf_8 fanout4253 (.A(_03180_),
    .X(net4253));
 sg13g2_buf_8 fanout4254 (.A(net4256),
    .X(net4254));
 sg13g2_buf_1 fanout4255 (.A(net4256),
    .X(net4255));
 sg13g2_buf_2 fanout4256 (.A(_10517_),
    .X(net4256));
 sg13g2_buf_8 fanout4257 (.A(_10517_),
    .X(net4257));
 sg13g2_buf_8 fanout4258 (.A(_10517_),
    .X(net4258));
 sg13g2_buf_8 fanout4259 (.A(net4261),
    .X(net4259));
 sg13g2_buf_1 fanout4260 (.A(net4261),
    .X(net4260));
 sg13g2_buf_8 fanout4261 (.A(_10504_),
    .X(net4261));
 sg13g2_buf_8 fanout4262 (.A(_10504_),
    .X(net4262));
 sg13g2_buf_8 fanout4263 (.A(_10504_),
    .X(net4263));
 sg13g2_buf_8 fanout4264 (.A(_10490_),
    .X(net4264));
 sg13g2_buf_8 fanout4265 (.A(net4268),
    .X(net4265));
 sg13g2_buf_8 fanout4266 (.A(net4268),
    .X(net4266));
 sg13g2_buf_1 fanout4267 (.A(net4268),
    .X(net4267));
 sg13g2_buf_2 fanout4268 (.A(_10490_),
    .X(net4268));
 sg13g2_buf_8 fanout4269 (.A(net4270),
    .X(net4269));
 sg13g2_buf_8 fanout4270 (.A(net4273),
    .X(net4270));
 sg13g2_buf_8 fanout4271 (.A(net4273),
    .X(net4271));
 sg13g2_buf_8 fanout4272 (.A(net4273),
    .X(net4272));
 sg13g2_buf_8 fanout4273 (.A(_10476_),
    .X(net4273));
 sg13g2_buf_8 fanout4274 (.A(net4275),
    .X(net4274));
 sg13g2_buf_1 fanout4275 (.A(net4276),
    .X(net4275));
 sg13g2_buf_8 fanout4276 (.A(_10462_),
    .X(net4276));
 sg13g2_buf_8 fanout4277 (.A(net4278),
    .X(net4277));
 sg13g2_buf_8 fanout4278 (.A(_10462_),
    .X(net4278));
 sg13g2_buf_8 fanout4279 (.A(net4280),
    .X(net4279));
 sg13g2_buf_8 fanout4280 (.A(net4283),
    .X(net4280));
 sg13g2_buf_8 fanout4281 (.A(net4283),
    .X(net4281));
 sg13g2_buf_2 fanout4282 (.A(net4283),
    .X(net4282));
 sg13g2_buf_8 fanout4283 (.A(_10449_),
    .X(net4283));
 sg13g2_buf_8 fanout4284 (.A(net4286),
    .X(net4284));
 sg13g2_buf_1 fanout4285 (.A(net4286),
    .X(net4285));
 sg13g2_buf_2 fanout4286 (.A(_10434_),
    .X(net4286));
 sg13g2_buf_8 fanout4287 (.A(net4288),
    .X(net4287));
 sg13g2_buf_1 fanout4288 (.A(net4289),
    .X(net4288));
 sg13g2_buf_1 fanout4289 (.A(_10434_),
    .X(net4289));
 sg13g2_buf_8 fanout4290 (.A(net4291),
    .X(net4290));
 sg13g2_buf_2 fanout4291 (.A(net4292),
    .X(net4291));
 sg13g2_buf_1 fanout4292 (.A(_10420_),
    .X(net4292));
 sg13g2_buf_8 fanout4293 (.A(net4295),
    .X(net4293));
 sg13g2_buf_1 fanout4294 (.A(net4295),
    .X(net4294));
 sg13g2_buf_2 fanout4295 (.A(_10420_),
    .X(net4295));
 sg13g2_buf_8 fanout4296 (.A(net4300),
    .X(net4296));
 sg13g2_buf_8 fanout4297 (.A(net4300),
    .X(net4297));
 sg13g2_buf_8 fanout4298 (.A(net4299),
    .X(net4298));
 sg13g2_buf_8 fanout4299 (.A(net4300),
    .X(net4299));
 sg13g2_buf_8 fanout4300 (.A(_10404_),
    .X(net4300));
 sg13g2_buf_8 fanout4301 (.A(net4306),
    .X(net4301));
 sg13g2_buf_1 fanout4302 (.A(net4306),
    .X(net4302));
 sg13g2_buf_8 fanout4303 (.A(net4305),
    .X(net4303));
 sg13g2_buf_1 fanout4304 (.A(net4305),
    .X(net4304));
 sg13g2_buf_8 fanout4305 (.A(net4306),
    .X(net4305));
 sg13g2_buf_8 fanout4306 (.A(_10392_),
    .X(net4306));
 sg13g2_buf_2 fanout4307 (.A(net4309),
    .X(net4307));
 sg13g2_buf_1 fanout4308 (.A(net4309),
    .X(net4308));
 sg13g2_buf_2 fanout4309 (.A(_10379_),
    .X(net4309));
 sg13g2_buf_8 fanout4310 (.A(net4311),
    .X(net4310));
 sg13g2_buf_8 fanout4311 (.A(_10379_),
    .X(net4311));
 sg13g2_buf_8 fanout4312 (.A(net4314),
    .X(net4312));
 sg13g2_buf_1 fanout4313 (.A(net4314),
    .X(net4313));
 sg13g2_buf_8 fanout4314 (.A(_10366_),
    .X(net4314));
 sg13g2_buf_8 fanout4315 (.A(net4317),
    .X(net4315));
 sg13g2_buf_1 fanout4316 (.A(net4317),
    .X(net4316));
 sg13g2_buf_2 fanout4317 (.A(_10366_),
    .X(net4317));
 sg13g2_buf_8 fanout4318 (.A(_10323_),
    .X(net4318));
 sg13g2_buf_1 fanout4319 (.A(_10323_),
    .X(net4319));
 sg13g2_buf_8 fanout4320 (.A(net4322),
    .X(net4320));
 sg13g2_buf_1 fanout4321 (.A(net4322),
    .X(net4321));
 sg13g2_buf_8 fanout4322 (.A(net4323),
    .X(net4322));
 sg13g2_buf_2 fanout4323 (.A(_10323_),
    .X(net4323));
 sg13g2_buf_8 fanout4324 (.A(_10300_),
    .X(net4324));
 sg13g2_buf_2 fanout4325 (.A(_10300_),
    .X(net4325));
 sg13g2_buf_8 fanout4326 (.A(net4328),
    .X(net4326));
 sg13g2_buf_1 fanout4327 (.A(net4328),
    .X(net4327));
 sg13g2_buf_8 fanout4328 (.A(_10300_),
    .X(net4328));
 sg13g2_buf_8 fanout4329 (.A(net4331),
    .X(net4329));
 sg13g2_buf_2 fanout4330 (.A(net4331),
    .X(net4330));
 sg13g2_buf_1 fanout4331 (.A(_10269_),
    .X(net4331));
 sg13g2_buf_8 fanout4332 (.A(net4333),
    .X(net4332));
 sg13g2_buf_8 fanout4333 (.A(_10269_),
    .X(net4333));
 sg13g2_buf_8 fanout4334 (.A(net4335),
    .X(net4334));
 sg13g2_buf_8 fanout4335 (.A(_10235_),
    .X(net4335));
 sg13g2_buf_8 fanout4336 (.A(net4338),
    .X(net4336));
 sg13g2_buf_1 fanout4337 (.A(net4338),
    .X(net4337));
 sg13g2_buf_8 fanout4338 (.A(_10235_),
    .X(net4338));
 sg13g2_buf_8 fanout4339 (.A(net4340),
    .X(net4339));
 sg13g2_buf_8 fanout4340 (.A(net4343),
    .X(net4340));
 sg13g2_buf_8 fanout4341 (.A(net4343),
    .X(net4341));
 sg13g2_buf_8 fanout4342 (.A(net4343),
    .X(net4342));
 sg13g2_buf_8 fanout4343 (.A(_10162_),
    .X(net4343));
 sg13g2_buf_8 fanout4344 (.A(net4346),
    .X(net4344));
 sg13g2_buf_8 fanout4345 (.A(net4346),
    .X(net4345));
 sg13g2_buf_8 fanout4346 (.A(_10123_),
    .X(net4346));
 sg13g2_buf_8 fanout4347 (.A(net4348),
    .X(net4347));
 sg13g2_buf_2 fanout4348 (.A(_10123_),
    .X(net4348));
 sg13g2_buf_8 fanout4349 (.A(net4350),
    .X(net4349));
 sg13g2_buf_1 fanout4350 (.A(net4351),
    .X(net4350));
 sg13g2_buf_2 fanout4351 (.A(_10080_),
    .X(net4351));
 sg13g2_buf_8 fanout4352 (.A(net4354),
    .X(net4352));
 sg13g2_buf_1 fanout4353 (.A(net4354),
    .X(net4353));
 sg13g2_buf_2 fanout4354 (.A(_10080_),
    .X(net4354));
 sg13g2_buf_8 fanout4355 (.A(net4357),
    .X(net4355));
 sg13g2_buf_1 fanout4356 (.A(net4357),
    .X(net4356));
 sg13g2_buf_8 fanout4357 (.A(net4360),
    .X(net4357));
 sg13g2_buf_8 fanout4358 (.A(net4360),
    .X(net4358));
 sg13g2_buf_2 fanout4359 (.A(net4360),
    .X(net4359));
 sg13g2_buf_8 fanout4360 (.A(_10026_),
    .X(net4360));
 sg13g2_buf_2 fanout4361 (.A(net4363),
    .X(net4361));
 sg13g2_buf_1 fanout4362 (.A(net4363),
    .X(net4362));
 sg13g2_buf_1 fanout4363 (.A(_09961_),
    .X(net4363));
 sg13g2_buf_8 fanout4364 (.A(net4365),
    .X(net4364));
 sg13g2_buf_2 fanout4365 (.A(net4366),
    .X(net4365));
 sg13g2_buf_1 fanout4366 (.A(_09961_),
    .X(net4366));
 sg13g2_buf_8 fanout4367 (.A(_09801_),
    .X(net4367));
 sg13g2_buf_2 fanout4368 (.A(_09801_),
    .X(net4368));
 sg13g2_buf_8 fanout4369 (.A(net4371),
    .X(net4369));
 sg13g2_buf_1 fanout4370 (.A(net4371),
    .X(net4370));
 sg13g2_buf_8 fanout4371 (.A(_09801_),
    .X(net4371));
 sg13g2_buf_8 fanout4372 (.A(net4373),
    .X(net4372));
 sg13g2_buf_8 fanout4373 (.A(net4376),
    .X(net4373));
 sg13g2_buf_8 fanout4374 (.A(net4376),
    .X(net4374));
 sg13g2_buf_8 fanout4375 (.A(net4376),
    .X(net4375));
 sg13g2_buf_8 fanout4376 (.A(_09789_),
    .X(net4376));
 sg13g2_buf_8 fanout4377 (.A(net4378),
    .X(net4377));
 sg13g2_buf_8 fanout4378 (.A(net4381),
    .X(net4378));
 sg13g2_buf_8 fanout4379 (.A(net4381),
    .X(net4379));
 sg13g2_buf_8 fanout4380 (.A(net4381),
    .X(net4380));
 sg13g2_buf_8 fanout4381 (.A(_09778_),
    .X(net4381));
 sg13g2_buf_8 fanout4382 (.A(net4387),
    .X(net4382));
 sg13g2_buf_1 fanout4383 (.A(net4387),
    .X(net4383));
 sg13g2_buf_8 fanout4384 (.A(net4386),
    .X(net4384));
 sg13g2_buf_1 fanout4385 (.A(net4386),
    .X(net4385));
 sg13g2_buf_8 fanout4386 (.A(net4387),
    .X(net4386));
 sg13g2_buf_8 fanout4387 (.A(_09767_),
    .X(net4387));
 sg13g2_buf_8 fanout4388 (.A(net4389),
    .X(net4388));
 sg13g2_buf_8 fanout4389 (.A(net4392),
    .X(net4389));
 sg13g2_buf_8 fanout4390 (.A(net4392),
    .X(net4390));
 sg13g2_buf_8 fanout4391 (.A(net4392),
    .X(net4391));
 sg13g2_buf_8 fanout4392 (.A(_09756_),
    .X(net4392));
 sg13g2_buf_8 fanout4393 (.A(net4394),
    .X(net4393));
 sg13g2_buf_1 fanout4394 (.A(_09744_),
    .X(net4394));
 sg13g2_buf_8 fanout4395 (.A(net4397),
    .X(net4395));
 sg13g2_buf_2 fanout4396 (.A(net4397),
    .X(net4396));
 sg13g2_buf_8 fanout4397 (.A(_09744_),
    .X(net4397));
 sg13g2_buf_8 fanout4398 (.A(net4400),
    .X(net4398));
 sg13g2_buf_1 fanout4399 (.A(net4400),
    .X(net4399));
 sg13g2_buf_2 fanout4400 (.A(_09731_),
    .X(net4400));
 sg13g2_buf_8 fanout4401 (.A(_09731_),
    .X(net4401));
 sg13g2_buf_8 fanout4402 (.A(_09731_),
    .X(net4402));
 sg13g2_buf_2 fanout4403 (.A(net4404),
    .X(net4403));
 sg13g2_buf_8 fanout4404 (.A(net4407),
    .X(net4404));
 sg13g2_buf_8 fanout4405 (.A(net4407),
    .X(net4405));
 sg13g2_buf_8 fanout4406 (.A(net4407),
    .X(net4406));
 sg13g2_buf_8 fanout4407 (.A(_09710_),
    .X(net4407));
 sg13g2_buf_8 fanout4408 (.A(_06383_),
    .X(net4408));
 sg13g2_buf_2 fanout4409 (.A(_06383_),
    .X(net4409));
 sg13g2_buf_8 fanout4410 (.A(_06362_),
    .X(net4410));
 sg13g2_buf_8 fanout4411 (.A(_06362_),
    .X(net4411));
 sg13g2_buf_8 fanout4412 (.A(net4413),
    .X(net4412));
 sg13g2_buf_8 fanout4413 (.A(_06355_),
    .X(net4413));
 sg13g2_buf_8 fanout4414 (.A(_06088_),
    .X(net4414));
 sg13g2_buf_8 fanout4415 (.A(_06088_),
    .X(net4415));
 sg13g2_buf_8 fanout4416 (.A(net4417),
    .X(net4416));
 sg13g2_buf_8 fanout4417 (.A(net4418),
    .X(net4417));
 sg13g2_buf_8 fanout4418 (.A(_06088_),
    .X(net4418));
 sg13g2_buf_8 fanout4419 (.A(net4420),
    .X(net4419));
 sg13g2_buf_8 fanout4420 (.A(_03572_),
    .X(net4420));
 sg13g2_buf_8 fanout4421 (.A(_03033_),
    .X(net4421));
 sg13g2_buf_8 fanout4422 (.A(_03033_),
    .X(net4422));
 sg13g2_buf_8 fanout4423 (.A(_06390_),
    .X(net4423));
 sg13g2_buf_8 fanout4424 (.A(_06390_),
    .X(net4424));
 sg13g2_buf_8 fanout4425 (.A(net4426),
    .X(net4425));
 sg13g2_buf_8 fanout4426 (.A(_06369_),
    .X(net4426));
 sg13g2_buf_8 fanout4427 (.A(net4429),
    .X(net4427));
 sg13g2_buf_1 fanout4428 (.A(net4429),
    .X(net4428));
 sg13g2_buf_1 fanout4429 (.A(net4433),
    .X(net4429));
 sg13g2_buf_8 fanout4430 (.A(net4431),
    .X(net4430));
 sg13g2_buf_2 fanout4431 (.A(net4432),
    .X(net4431));
 sg13g2_buf_1 fanout4432 (.A(net4433),
    .X(net4432));
 sg13g2_buf_8 fanout4433 (.A(_03597_),
    .X(net4433));
 sg13g2_buf_2 fanout4434 (.A(net4435),
    .X(net4434));
 sg13g2_buf_8 fanout4435 (.A(_03589_),
    .X(net4435));
 sg13g2_buf_8 fanout4436 (.A(net4438),
    .X(net4436));
 sg13g2_buf_1 fanout4437 (.A(net4438),
    .X(net4437));
 sg13g2_buf_2 fanout4438 (.A(_03581_),
    .X(net4438));
 sg13g2_buf_8 fanout4439 (.A(_03556_),
    .X(net4439));
 sg13g2_buf_8 fanout4440 (.A(_03556_),
    .X(net4440));
 sg13g2_buf_8 fanout4441 (.A(_03539_),
    .X(net4441));
 sg13g2_buf_8 fanout4442 (.A(net4446),
    .X(net4442));
 sg13g2_buf_8 fanout4443 (.A(net4445),
    .X(net4443));
 sg13g2_buf_8 fanout4444 (.A(net4445),
    .X(net4444));
 sg13g2_buf_8 fanout4445 (.A(net4446),
    .X(net4445));
 sg13g2_buf_8 fanout4446 (.A(_03053_),
    .X(net4446));
 sg13g2_buf_8 fanout4447 (.A(_03052_),
    .X(net4447));
 sg13g2_buf_2 fanout4448 (.A(_03052_),
    .X(net4448));
 sg13g2_buf_8 fanout4449 (.A(net4450),
    .X(net4449));
 sg13g2_buf_1 fanout4450 (.A(net4451),
    .X(net4450));
 sg13g2_buf_1 fanout4451 (.A(net4452),
    .X(net4451));
 sg13g2_buf_8 fanout4452 (.A(_03051_),
    .X(net4452));
 sg13g2_buf_8 fanout4453 (.A(net4454),
    .X(net4453));
 sg13g2_buf_8 fanout4454 (.A(net4457),
    .X(net4454));
 sg13g2_buf_8 fanout4455 (.A(net4456),
    .X(net4455));
 sg13g2_buf_8 fanout4456 (.A(net4457),
    .X(net4456));
 sg13g2_buf_8 fanout4457 (.A(_03051_),
    .X(net4457));
 sg13g2_buf_8 fanout4458 (.A(_02998_),
    .X(net4458));
 sg13g2_buf_8 fanout4459 (.A(net4460),
    .X(net4459));
 sg13g2_buf_8 fanout4460 (.A(_02996_),
    .X(net4460));
 sg13g2_buf_8 fanout4461 (.A(_09618_),
    .X(net4461));
 sg13g2_buf_1 fanout4462 (.A(_09618_),
    .X(net4462));
 sg13g2_buf_8 fanout4463 (.A(net4464),
    .X(net4463));
 sg13g2_buf_8 fanout4464 (.A(net4465),
    .X(net4464));
 sg13g2_buf_8 fanout4465 (.A(_06486_),
    .X(net4465));
 sg13g2_buf_8 fanout4466 (.A(_03537_),
    .X(net4466));
 sg13g2_buf_8 fanout4467 (.A(_03049_),
    .X(net4467));
 sg13g2_buf_1 fanout4468 (.A(_03049_),
    .X(net4468));
 sg13g2_buf_8 fanout4469 (.A(_10584_),
    .X(net4469));
 sg13g2_buf_1 fanout4470 (.A(_10584_),
    .X(net4470));
 sg13g2_buf_8 fanout4471 (.A(net4473),
    .X(net4471));
 sg13g2_buf_1 fanout4472 (.A(net4473),
    .X(net4472));
 sg13g2_buf_1 fanout4473 (.A(_10584_),
    .X(net4473));
 sg13g2_buf_8 fanout4474 (.A(net4475),
    .X(net4474));
 sg13g2_buf_8 fanout4475 (.A(net4481),
    .X(net4475));
 sg13g2_buf_8 fanout4476 (.A(net4481),
    .X(net4476));
 sg13g2_buf_1 fanout4477 (.A(net4481),
    .X(net4477));
 sg13g2_buf_8 fanout4478 (.A(net4479),
    .X(net4478));
 sg13g2_buf_8 fanout4479 (.A(net4480),
    .X(net4479));
 sg13g2_buf_8 fanout4480 (.A(net4481),
    .X(net4480));
 sg13g2_buf_8 fanout4481 (.A(_09458_),
    .X(net4481));
 sg13g2_buf_8 fanout4482 (.A(net4484),
    .X(net4482));
 sg13g2_buf_1 fanout4483 (.A(net4484),
    .X(net4483));
 sg13g2_buf_8 fanout4484 (.A(_09457_),
    .X(net4484));
 sg13g2_buf_8 fanout4485 (.A(net4487),
    .X(net4485));
 sg13g2_buf_1 fanout4486 (.A(net4487),
    .X(net4486));
 sg13g2_buf_2 fanout4487 (.A(net4488),
    .X(net4487));
 sg13g2_buf_1 fanout4488 (.A(net4489),
    .X(net4488));
 sg13g2_buf_8 fanout4489 (.A(_06055_),
    .X(net4489));
 sg13g2_buf_8 fanout4490 (.A(net4493),
    .X(net4490));
 sg13g2_buf_8 fanout4491 (.A(net4493),
    .X(net4491));
 sg13g2_buf_1 fanout4492 (.A(net4493),
    .X(net4492));
 sg13g2_buf_2 fanout4493 (.A(_06055_),
    .X(net4493));
 sg13g2_buf_8 fanout4494 (.A(net4496),
    .X(net4494));
 sg13g2_buf_1 fanout4495 (.A(net4496),
    .X(net4495));
 sg13g2_buf_8 fanout4496 (.A(_06055_),
    .X(net4496));
 sg13g2_buf_8 fanout4497 (.A(net4499),
    .X(net4497));
 sg13g2_buf_8 fanout4498 (.A(net4499),
    .X(net4498));
 sg13g2_buf_8 fanout4499 (.A(net4500),
    .X(net4499));
 sg13g2_buf_8 fanout4500 (.A(_04971_),
    .X(net4500));
 sg13g2_buf_8 fanout4501 (.A(net4504),
    .X(net4501));
 sg13g2_buf_8 fanout4502 (.A(net4504),
    .X(net4502));
 sg13g2_buf_8 fanout4503 (.A(net4504),
    .X(net4503));
 sg13g2_buf_8 fanout4504 (.A(_03048_),
    .X(net4504));
 sg13g2_buf_8 fanout4505 (.A(net4506),
    .X(net4505));
 sg13g2_buf_8 fanout4506 (.A(net4516),
    .X(net4506));
 sg13g2_buf_8 fanout4507 (.A(net4509),
    .X(net4507));
 sg13g2_buf_1 fanout4508 (.A(net4509),
    .X(net4508));
 sg13g2_buf_1 fanout4509 (.A(net4516),
    .X(net4509));
 sg13g2_buf_8 fanout4510 (.A(net4511),
    .X(net4510));
 sg13g2_buf_8 fanout4511 (.A(net4516),
    .X(net4511));
 sg13g2_buf_8 fanout4512 (.A(net4515),
    .X(net4512));
 sg13g2_buf_8 fanout4513 (.A(net4515),
    .X(net4513));
 sg13g2_buf_2 fanout4514 (.A(net4515),
    .X(net4514));
 sg13g2_buf_8 fanout4515 (.A(net4516),
    .X(net4515));
 sg13g2_buf_8 fanout4516 (.A(_03046_),
    .X(net4516));
 sg13g2_buf_2 fanout4517 (.A(net4518),
    .X(net4517));
 sg13g2_buf_2 fanout4518 (.A(net4519),
    .X(net4518));
 sg13g2_buf_8 fanout4519 (.A(_02741_),
    .X(net4519));
 sg13g2_buf_8 fanout4520 (.A(net4522),
    .X(net4520));
 sg13g2_buf_1 fanout4521 (.A(net4522),
    .X(net4521));
 sg13g2_buf_8 fanout4522 (.A(net4523),
    .X(net4522));
 sg13g2_buf_8 fanout4523 (.A(_02741_),
    .X(net4523));
 sg13g2_buf_8 fanout4524 (.A(net4525),
    .X(net4524));
 sg13g2_buf_8 fanout4525 (.A(net4526),
    .X(net4525));
 sg13g2_buf_8 fanout4526 (.A(net4527),
    .X(net4526));
 sg13g2_buf_8 fanout4527 (.A(_02741_),
    .X(net4527));
 sg13g2_buf_8 fanout4528 (.A(net4534),
    .X(net4528));
 sg13g2_buf_1 fanout4529 (.A(net4534),
    .X(net4529));
 sg13g2_buf_8 fanout4530 (.A(net4533),
    .X(net4530));
 sg13g2_buf_8 fanout4531 (.A(net4532),
    .X(net4531));
 sg13g2_buf_2 fanout4532 (.A(net4533),
    .X(net4532));
 sg13g2_buf_8 fanout4533 (.A(net4534),
    .X(net4533));
 sg13g2_buf_8 fanout4534 (.A(net4535),
    .X(net4534));
 sg13g2_buf_8 fanout4535 (.A(_09552_),
    .X(net4535));
 sg13g2_buf_8 fanout4536 (.A(net4537),
    .X(net4536));
 sg13g2_buf_1 fanout4537 (.A(net4538),
    .X(net4537));
 sg13g2_buf_1 fanout4538 (.A(net4539),
    .X(net4538));
 sg13g2_buf_8 fanout4539 (.A(net4540),
    .X(net4539));
 sg13g2_buf_8 fanout4540 (.A(_04972_),
    .X(net4540));
 sg13g2_buf_8 fanout4541 (.A(net4543),
    .X(net4541));
 sg13g2_buf_2 fanout4542 (.A(net4543),
    .X(net4542));
 sg13g2_buf_8 fanout4543 (.A(_03201_),
    .X(net4543));
 sg13g2_buf_8 fanout4544 (.A(net4545),
    .X(net4544));
 sg13g2_buf_8 fanout4545 (.A(_03201_),
    .X(net4545));
 sg13g2_buf_8 fanout4546 (.A(net4547),
    .X(net4546));
 sg13g2_buf_8 fanout4547 (.A(net4548),
    .X(net4547));
 sg13g2_buf_8 fanout4548 (.A(_03200_),
    .X(net4548));
 sg13g2_buf_8 fanout4549 (.A(_03200_),
    .X(net4549));
 sg13g2_buf_8 fanout4550 (.A(net4559),
    .X(net4550));
 sg13g2_buf_8 fanout4551 (.A(net4553),
    .X(net4551));
 sg13g2_buf_1 fanout4552 (.A(net4553),
    .X(net4552));
 sg13g2_buf_8 fanout4553 (.A(net4554),
    .X(net4553));
 sg13g2_buf_8 fanout4554 (.A(net4559),
    .X(net4554));
 sg13g2_buf_8 fanout4555 (.A(net4556),
    .X(net4555));
 sg13g2_buf_8 fanout4556 (.A(net4558),
    .X(net4556));
 sg13g2_buf_8 fanout4557 (.A(net4558),
    .X(net4557));
 sg13g2_buf_8 fanout4558 (.A(net4559),
    .X(net4558));
 sg13g2_buf_8 fanout4559 (.A(_09560_),
    .X(net4559));
 sg13g2_buf_8 fanout4560 (.A(_08893_),
    .X(net4560));
 sg13g2_buf_8 fanout4561 (.A(_04965_),
    .X(net4561));
 sg13g2_buf_1 fanout4562 (.A(_04965_),
    .X(net4562));
 sg13g2_buf_8 fanout4563 (.A(net4568),
    .X(net4563));
 sg13g2_buf_2 fanout4564 (.A(net4568),
    .X(net4564));
 sg13g2_buf_8 fanout4565 (.A(net4567),
    .X(net4565));
 sg13g2_buf_2 fanout4566 (.A(net4567),
    .X(net4566));
 sg13g2_buf_2 fanout4567 (.A(net4568),
    .X(net4567));
 sg13g2_buf_1 fanout4568 (.A(net4569),
    .X(net4568));
 sg13g2_buf_8 fanout4569 (.A(_09547_),
    .X(net4569));
 sg13g2_buf_8 fanout4570 (.A(_08849_),
    .X(net4570));
 sg13g2_buf_8 fanout4571 (.A(net4573),
    .X(net4571));
 sg13g2_buf_1 fanout4572 (.A(net4573),
    .X(net4572));
 sg13g2_buf_2 fanout4573 (.A(net4574),
    .X(net4573));
 sg13g2_buf_8 fanout4574 (.A(_04964_),
    .X(net4574));
 sg13g2_buf_8 fanout4575 (.A(net4576),
    .X(net4575));
 sg13g2_buf_8 fanout4576 (.A(net4577),
    .X(net4576));
 sg13g2_buf_1 fanout4577 (.A(net4578),
    .X(net4577));
 sg13g2_buf_1 fanout4578 (.A(net4579),
    .X(net4578));
 sg13g2_buf_1 fanout4579 (.A(_04964_),
    .X(net4579));
 sg13g2_buf_8 fanout4580 (.A(_05546_),
    .X(net4580));
 sg13g2_buf_8 fanout4581 (.A(net4582),
    .X(net4581));
 sg13g2_buf_8 fanout4582 (.A(_03835_),
    .X(net4582));
 sg13g2_buf_8 fanout4583 (.A(net4585),
    .X(net4583));
 sg13g2_buf_1 fanout4584 (.A(net4585),
    .X(net4584));
 sg13g2_buf_8 fanout4585 (.A(net4586),
    .X(net4585));
 sg13g2_buf_8 fanout4586 (.A(_03835_),
    .X(net4586));
 sg13g2_buf_8 fanout4587 (.A(_03834_),
    .X(net4587));
 sg13g2_buf_8 fanout4588 (.A(net4589),
    .X(net4588));
 sg13g2_buf_8 fanout4589 (.A(_03834_),
    .X(net4589));
 sg13g2_buf_8 fanout4590 (.A(_05943_),
    .X(net4590));
 sg13g2_buf_8 fanout4591 (.A(_05938_),
    .X(net4591));
 sg13g2_buf_1 fanout4592 (.A(_05938_),
    .X(net4592));
 sg13g2_buf_8 fanout4593 (.A(net4594),
    .X(net4593));
 sg13g2_buf_8 fanout4594 (.A(_05937_),
    .X(net4594));
 sg13g2_buf_8 fanout4595 (.A(net4596),
    .X(net4595));
 sg13g2_buf_1 fanout4596 (.A(net4597),
    .X(net4596));
 sg13g2_buf_8 fanout4597 (.A(net4598),
    .X(net4597));
 sg13g2_buf_8 fanout4598 (.A(_05937_),
    .X(net4598));
 sg13g2_buf_8 fanout4599 (.A(net4600),
    .X(net4599));
 sg13g2_buf_8 fanout4600 (.A(net4607),
    .X(net4600));
 sg13g2_buf_8 fanout4601 (.A(net4607),
    .X(net4601));
 sg13g2_buf_8 fanout4602 (.A(net4606),
    .X(net4602));
 sg13g2_buf_8 fanout4603 (.A(net4606),
    .X(net4603));
 sg13g2_buf_1 fanout4604 (.A(net4606),
    .X(net4604));
 sg13g2_buf_8 fanout4605 (.A(net4606),
    .X(net4605));
 sg13g2_buf_8 fanout4606 (.A(net4607),
    .X(net4606));
 sg13g2_buf_8 fanout4607 (.A(_05879_),
    .X(net4607));
 sg13g2_buf_8 fanout4608 (.A(_05570_),
    .X(net4608));
 sg13g2_buf_8 fanout4609 (.A(net4610),
    .X(net4609));
 sg13g2_buf_8 fanout4610 (.A(_05570_),
    .X(net4610));
 sg13g2_buf_8 fanout4611 (.A(net4612),
    .X(net4611));
 sg13g2_buf_1 fanout4612 (.A(net4617),
    .X(net4612));
 sg13g2_buf_8 fanout4613 (.A(net4617),
    .X(net4613));
 sg13g2_buf_8 fanout4614 (.A(net4615),
    .X(net4614));
 sg13g2_buf_8 fanout4615 (.A(net4616),
    .X(net4615));
 sg13g2_buf_8 fanout4616 (.A(net4617),
    .X(net4616));
 sg13g2_buf_8 fanout4617 (.A(_05569_),
    .X(net4617));
 sg13g2_buf_8 fanout4618 (.A(net4619),
    .X(net4618));
 sg13g2_buf_8 fanout4619 (.A(_05358_),
    .X(net4619));
 sg13g2_buf_8 fanout4620 (.A(net4621),
    .X(net4620));
 sg13g2_buf_8 fanout4621 (.A(_05358_),
    .X(net4621));
 sg13g2_buf_8 fanout4622 (.A(net4627),
    .X(net4622));
 sg13g2_buf_8 fanout4623 (.A(net4626),
    .X(net4623));
 sg13g2_buf_8 fanout4624 (.A(net4625),
    .X(net4624));
 sg13g2_buf_8 fanout4625 (.A(net4626),
    .X(net4625));
 sg13g2_buf_8 fanout4626 (.A(net4627),
    .X(net4626));
 sg13g2_buf_8 fanout4627 (.A(_05358_),
    .X(net4627));
 sg13g2_buf_8 fanout4628 (.A(net4629),
    .X(net4628));
 sg13g2_buf_8 fanout4629 (.A(_03829_),
    .X(net4629));
 sg13g2_buf_8 fanout4630 (.A(net4631),
    .X(net4630));
 sg13g2_buf_8 fanout4631 (.A(net4632),
    .X(net4631));
 sg13g2_buf_8 fanout4632 (.A(_03829_),
    .X(net4632));
 sg13g2_buf_8 fanout4633 (.A(_05936_),
    .X(net4633));
 sg13g2_buf_8 fanout4634 (.A(_05936_),
    .X(net4634));
 sg13g2_buf_8 fanout4635 (.A(_05883_),
    .X(net4635));
 sg13g2_buf_8 fanout4636 (.A(_05878_),
    .X(net4636));
 sg13g2_buf_8 fanout4637 (.A(_05878_),
    .X(net4637));
 sg13g2_buf_8 fanout4638 (.A(net4639),
    .X(net4638));
 sg13g2_buf_8 fanout4639 (.A(net4641),
    .X(net4639));
 sg13g2_buf_8 fanout4640 (.A(net4641),
    .X(net4640));
 sg13g2_buf_8 fanout4641 (.A(_05577_),
    .X(net4641));
 sg13g2_buf_8 fanout4642 (.A(net4647),
    .X(net4642));
 sg13g2_buf_8 fanout4643 (.A(net4645),
    .X(net4643));
 sg13g2_buf_1 fanout4644 (.A(net4645),
    .X(net4644));
 sg13g2_buf_2 fanout4645 (.A(net4647),
    .X(net4645));
 sg13g2_buf_8 fanout4646 (.A(net4647),
    .X(net4646));
 sg13g2_buf_8 fanout4647 (.A(_05577_),
    .X(net4647));
 sg13g2_buf_8 fanout4648 (.A(net4649),
    .X(net4648));
 sg13g2_buf_8 fanout4649 (.A(net4650),
    .X(net4649));
 sg13g2_buf_8 fanout4650 (.A(net4651),
    .X(net4650));
 sg13g2_buf_8 fanout4651 (.A(_05359_),
    .X(net4651));
 sg13g2_buf_8 fanout4652 (.A(net4657),
    .X(net4652));
 sg13g2_buf_8 fanout4653 (.A(net4657),
    .X(net4653));
 sg13g2_buf_2 fanout4654 (.A(net4656),
    .X(net4654));
 sg13g2_buf_1 fanout4655 (.A(net4656),
    .X(net4655));
 sg13g2_buf_1 fanout4656 (.A(net4657),
    .X(net4656));
 sg13g2_buf_8 fanout4657 (.A(_05359_),
    .X(net4657));
 sg13g2_buf_8 fanout4658 (.A(_03872_),
    .X(net4658));
 sg13g2_buf_8 fanout4659 (.A(_03872_),
    .X(net4659));
 sg13g2_buf_8 fanout4660 (.A(net4661),
    .X(net4660));
 sg13g2_buf_8 fanout4661 (.A(_03865_),
    .X(net4661));
 sg13g2_buf_8 fanout4662 (.A(net4663),
    .X(net4662));
 sg13g2_buf_8 fanout4663 (.A(_03852_),
    .X(net4663));
 sg13g2_buf_8 fanout4664 (.A(_03852_),
    .X(net4664));
 sg13g2_buf_8 fanout4665 (.A(net4666),
    .X(net4665));
 sg13g2_buf_8 fanout4666 (.A(_03850_),
    .X(net4666));
 sg13g2_buf_8 fanout4667 (.A(net4668),
    .X(net4667));
 sg13g2_buf_8 fanout4668 (.A(net4669),
    .X(net4668));
 sg13g2_buf_8 fanout4669 (.A(_03850_),
    .X(net4669));
 sg13g2_buf_8 fanout4670 (.A(_03846_),
    .X(net4670));
 sg13g2_buf_8 fanout4671 (.A(net4673),
    .X(net4671));
 sg13g2_buf_1 fanout4672 (.A(net4673),
    .X(net4672));
 sg13g2_buf_8 fanout4673 (.A(_03845_),
    .X(net4673));
 sg13g2_buf_8 fanout4674 (.A(net4676),
    .X(net4674));
 sg13g2_buf_1 fanout4675 (.A(net4676),
    .X(net4675));
 sg13g2_buf_8 fanout4676 (.A(_03845_),
    .X(net4676));
 sg13g2_buf_8 fanout4677 (.A(net4679),
    .X(net4677));
 sg13g2_buf_1 fanout4678 (.A(net4679),
    .X(net4678));
 sg13g2_buf_8 fanout4679 (.A(net4683),
    .X(net4679));
 sg13g2_buf_8 fanout4680 (.A(net4681),
    .X(net4680));
 sg13g2_buf_8 fanout4681 (.A(net4683),
    .X(net4681));
 sg13g2_buf_8 fanout4682 (.A(net4683),
    .X(net4682));
 sg13g2_buf_8 fanout4683 (.A(_05989_),
    .X(net4683));
 sg13g2_buf_8 fanout4684 (.A(net4685),
    .X(net4684));
 sg13g2_buf_8 fanout4685 (.A(_05987_),
    .X(net4685));
 sg13g2_buf_8 fanout4686 (.A(_03892_),
    .X(net4686));
 sg13g2_buf_8 fanout4687 (.A(net4689),
    .X(net4687));
 sg13g2_buf_1 fanout4688 (.A(net4689),
    .X(net4688));
 sg13g2_buf_8 fanout4689 (.A(_03892_),
    .X(net4689));
 sg13g2_buf_8 fanout4690 (.A(net4691),
    .X(net4690));
 sg13g2_buf_8 fanout4691 (.A(_09295_),
    .X(net4691));
 sg13g2_buf_8 fanout4692 (.A(net4693),
    .X(net4692));
 sg13g2_buf_8 fanout4693 (.A(net4694),
    .X(net4693));
 sg13g2_buf_8 fanout4694 (.A(_03863_),
    .X(net4694));
 sg13g2_buf_8 fanout4695 (.A(_03859_),
    .X(net4695));
 sg13g2_buf_8 fanout4696 (.A(net4698),
    .X(net4696));
 sg13g2_buf_1 fanout4697 (.A(net4698),
    .X(net4697));
 sg13g2_buf_8 fanout4698 (.A(_03858_),
    .X(net4698));
 sg13g2_buf_8 fanout4699 (.A(_03858_),
    .X(net4699));
 sg13g2_buf_8 fanout4700 (.A(net4701),
    .X(net4700));
 sg13g2_buf_1 fanout4701 (.A(net4710),
    .X(net4701));
 sg13g2_buf_8 fanout4702 (.A(net4704),
    .X(net4702));
 sg13g2_buf_1 fanout4703 (.A(net4704),
    .X(net4703));
 sg13g2_buf_8 fanout4704 (.A(net4709),
    .X(net4704));
 sg13g2_buf_8 fanout4705 (.A(net4709),
    .X(net4705));
 sg13g2_buf_1 fanout4706 (.A(net4709),
    .X(net4706));
 sg13g2_buf_8 fanout4707 (.A(net4708),
    .X(net4707));
 sg13g2_buf_8 fanout4708 (.A(net4709),
    .X(net4708));
 sg13g2_buf_8 fanout4709 (.A(net4710),
    .X(net4709));
 sg13g2_buf_8 fanout4710 (.A(_03268_),
    .X(net4710));
 sg13g2_buf_8 fanout4711 (.A(net4712),
    .X(net4711));
 sg13g2_buf_8 fanout4712 (.A(net4713),
    .X(net4712));
 sg13g2_buf_8 fanout4713 (.A(net4718),
    .X(net4713));
 sg13g2_buf_8 fanout4714 (.A(net4715),
    .X(net4714));
 sg13g2_buf_8 fanout4715 (.A(net4718),
    .X(net4715));
 sg13g2_buf_8 fanout4716 (.A(net4717),
    .X(net4716));
 sg13g2_buf_8 fanout4717 (.A(net4718),
    .X(net4717));
 sg13g2_buf_8 fanout4718 (.A(\fpga_top.uart_top.uart_rec_char.word_valid_pre ),
    .X(net4718));
 sg13g2_buf_8 fanout4719 (.A(net4722),
    .X(net4719));
 sg13g2_buf_1 fanout4720 (.A(net4722),
    .X(net4720));
 sg13g2_buf_8 fanout4721 (.A(net4722),
    .X(net4721));
 sg13g2_buf_8 fanout4722 (.A(_04983_),
    .X(net4722));
 sg13g2_buf_8 fanout4723 (.A(net4724),
    .X(net4723));
 sg13g2_buf_8 fanout4724 (.A(_04969_),
    .X(net4724));
 sg13g2_buf_8 fanout4725 (.A(net4726),
    .X(net4725));
 sg13g2_buf_8 fanout4726 (.A(_04968_),
    .X(net4726));
 sg13g2_buf_8 fanout4727 (.A(net4729),
    .X(net4727));
 sg13g2_buf_1 fanout4728 (.A(net4729),
    .X(net4728));
 sg13g2_buf_8 fanout4729 (.A(net4732),
    .X(net4729));
 sg13g2_buf_8 fanout4730 (.A(net4731),
    .X(net4730));
 sg13g2_buf_8 fanout4731 (.A(net4732),
    .X(net4731));
 sg13g2_buf_8 fanout4732 (.A(net4740),
    .X(net4732));
 sg13g2_buf_8 fanout4733 (.A(net4740),
    .X(net4733));
 sg13g2_buf_1 fanout4734 (.A(net4740),
    .X(net4734));
 sg13g2_buf_8 fanout4735 (.A(net4737),
    .X(net4735));
 sg13g2_buf_1 fanout4736 (.A(net4737),
    .X(net4736));
 sg13g2_buf_2 fanout4737 (.A(net4738),
    .X(net4737));
 sg13g2_buf_2 fanout4738 (.A(net4739),
    .X(net4738));
 sg13g2_buf_8 fanout4739 (.A(net4740),
    .X(net4739));
 sg13g2_buf_8 fanout4740 (.A(_04926_),
    .X(net4740));
 sg13g2_buf_8 fanout4741 (.A(net4744),
    .X(net4741));
 sg13g2_buf_8 fanout4742 (.A(net4744),
    .X(net4742));
 sg13g2_buf_1 fanout4743 (.A(net4744),
    .X(net4743));
 sg13g2_buf_8 fanout4744 (.A(_04925_),
    .X(net4744));
 sg13g2_buf_8 fanout4745 (.A(net4746),
    .X(net4745));
 sg13g2_buf_1 fanout4746 (.A(net4747),
    .X(net4746));
 sg13g2_buf_2 fanout4747 (.A(_04424_),
    .X(net4747));
 sg13g2_buf_8 fanout4748 (.A(net4749),
    .X(net4748));
 sg13g2_buf_8 fanout4749 (.A(_04424_),
    .X(net4749));
 sg13g2_buf_8 fanout4750 (.A(net4754),
    .X(net4750));
 sg13g2_buf_1 fanout4751 (.A(net4754),
    .X(net4751));
 sg13g2_buf_8 fanout4752 (.A(net4754),
    .X(net4752));
 sg13g2_buf_8 fanout4753 (.A(net4754),
    .X(net4753));
 sg13g2_buf_8 fanout4754 (.A(net4755),
    .X(net4754));
 sg13g2_buf_8 fanout4755 (.A(_03249_),
    .X(net4755));
 sg13g2_buf_8 fanout4756 (.A(_07687_),
    .X(net4756));
 sg13g2_buf_8 fanout4757 (.A(_05574_),
    .X(net4757));
 sg13g2_buf_1 fanout4758 (.A(_05574_),
    .X(net4758));
 sg13g2_buf_8 fanout4759 (.A(net4760),
    .X(net4759));
 sg13g2_buf_8 fanout4760 (.A(net4761),
    .X(net4760));
 sg13g2_buf_2 fanout4761 (.A(_05574_),
    .X(net4761));
 sg13g2_buf_8 fanout4762 (.A(net4766),
    .X(net4762));
 sg13g2_buf_1 fanout4763 (.A(net4766),
    .X(net4763));
 sg13g2_buf_8 fanout4764 (.A(net4765),
    .X(net4764));
 sg13g2_buf_8 fanout4765 (.A(net4766),
    .X(net4765));
 sg13g2_buf_8 fanout4766 (.A(net4774),
    .X(net4766));
 sg13g2_buf_8 fanout4767 (.A(net4774),
    .X(net4767));
 sg13g2_buf_1 fanout4768 (.A(net4774),
    .X(net4768));
 sg13g2_buf_8 fanout4769 (.A(net4773),
    .X(net4769));
 sg13g2_buf_8 fanout4770 (.A(net4771),
    .X(net4770));
 sg13g2_buf_1 fanout4771 (.A(net4772),
    .X(net4771));
 sg13g2_buf_1 fanout4772 (.A(net4773),
    .X(net4772));
 sg13g2_buf_8 fanout4773 (.A(net4774),
    .X(net4773));
 sg13g2_buf_8 fanout4774 (.A(_05328_),
    .X(net4774));
 sg13g2_buf_8 fanout4775 (.A(_04923_),
    .X(net4775));
 sg13g2_buf_2 fanout4776 (.A(_04923_),
    .X(net4776));
 sg13g2_buf_8 fanout4777 (.A(net4778),
    .X(net4777));
 sg13g2_buf_8 fanout4778 (.A(net4779),
    .X(net4778));
 sg13g2_buf_2 fanout4779 (.A(_04923_),
    .X(net4779));
 sg13g2_buf_8 fanout4780 (.A(net4783),
    .X(net4780));
 sg13g2_buf_8 fanout4781 (.A(net4782),
    .X(net4781));
 sg13g2_buf_8 fanout4782 (.A(net4783),
    .X(net4782));
 sg13g2_buf_2 fanout4783 (.A(_09637_),
    .X(net4783));
 sg13g2_buf_8 fanout4784 (.A(_07629_),
    .X(net4784));
 sg13g2_buf_2 fanout4785 (.A(_07629_),
    .X(net4785));
 sg13g2_buf_8 fanout4786 (.A(_07580_),
    .X(net4786));
 sg13g2_buf_8 fanout4787 (.A(_05370_),
    .X(net4787));
 sg13g2_buf_1 fanout4788 (.A(_05370_),
    .X(net4788));
 sg13g2_buf_8 fanout4789 (.A(net4790),
    .X(net4789));
 sg13g2_buf_8 fanout4790 (.A(net4791),
    .X(net4790));
 sg13g2_buf_8 fanout4791 (.A(_05370_),
    .X(net4791));
 sg13g2_buf_8 fanout4792 (.A(net4793),
    .X(net4792));
 sg13g2_buf_2 fanout4793 (.A(net4794),
    .X(net4793));
 sg13g2_buf_8 fanout4794 (.A(_05351_),
    .X(net4794));
 sg13g2_buf_8 fanout4795 (.A(net4796),
    .X(net4795));
 sg13g2_buf_1 fanout4796 (.A(net4797),
    .X(net4796));
 sg13g2_buf_8 fanout4797 (.A(_05351_),
    .X(net4797));
 sg13g2_buf_8 fanout4798 (.A(_05350_),
    .X(net4798));
 sg13g2_buf_1 fanout4799 (.A(_05350_),
    .X(net4799));
 sg13g2_buf_8 fanout4800 (.A(net4801),
    .X(net4800));
 sg13g2_buf_8 fanout4801 (.A(net4802),
    .X(net4801));
 sg13g2_buf_1 fanout4802 (.A(_05350_),
    .X(net4802));
 sg13g2_buf_8 fanout4803 (.A(net4805),
    .X(net4803));
 sg13g2_buf_1 fanout4804 (.A(net4805),
    .X(net4804));
 sg13g2_buf_1 fanout4805 (.A(_05329_),
    .X(net4805));
 sg13g2_buf_8 fanout4806 (.A(net4807),
    .X(net4806));
 sg13g2_buf_8 fanout4807 (.A(_05329_),
    .X(net4807));
 sg13g2_buf_8 fanout4808 (.A(net4810),
    .X(net4808));
 sg13g2_buf_8 fanout4809 (.A(net4810),
    .X(net4809));
 sg13g2_buf_8 fanout4810 (.A(net4811),
    .X(net4810));
 sg13g2_buf_8 fanout4811 (.A(_04667_),
    .X(net4811));
 sg13g2_buf_8 fanout4812 (.A(net4814),
    .X(net4812));
 sg13g2_buf_1 fanout4813 (.A(net4814),
    .X(net4813));
 sg13g2_buf_8 fanout4814 (.A(net4815),
    .X(net4814));
 sg13g2_buf_8 fanout4815 (.A(_04666_),
    .X(net4815));
 sg13g2_buf_8 fanout4816 (.A(net4817),
    .X(net4816));
 sg13g2_buf_8 fanout4817 (.A(_04508_),
    .X(net4817));
 sg13g2_buf_8 fanout4818 (.A(net4821),
    .X(net4818));
 sg13g2_buf_1 fanout4819 (.A(net4821),
    .X(net4819));
 sg13g2_buf_8 fanout4820 (.A(net4821),
    .X(net4820));
 sg13g2_buf_8 fanout4821 (.A(_04357_),
    .X(net4821));
 sg13g2_buf_8 fanout4822 (.A(net4824),
    .X(net4822));
 sg13g2_buf_1 fanout4823 (.A(net4824),
    .X(net4823));
 sg13g2_buf_1 fanout4824 (.A(net4825),
    .X(net4824));
 sg13g2_buf_2 fanout4825 (.A(net4827),
    .X(net4825));
 sg13g2_buf_8 fanout4826 (.A(net4827),
    .X(net4826));
 sg13g2_buf_8 fanout4827 (.A(_04357_),
    .X(net4827));
 sg13g2_buf_8 fanout4828 (.A(_03833_),
    .X(net4828));
 sg13g2_buf_2 fanout4829 (.A(_03833_),
    .X(net4829));
 sg13g2_buf_8 fanout4830 (.A(_02759_),
    .X(net4830));
 sg13g2_buf_8 fanout4831 (.A(_02759_),
    .X(net4831));
 sg13g2_buf_8 fanout4832 (.A(_02755_),
    .X(net4832));
 sg13g2_buf_8 fanout4833 (.A(_02755_),
    .X(net4833));
 sg13g2_buf_8 fanout4834 (.A(_02752_),
    .X(net4834));
 sg13g2_buf_8 fanout4835 (.A(_02751_),
    .X(net4835));
 sg13g2_buf_8 fanout4836 (.A(_02751_),
    .X(net4836));
 sg13g2_buf_8 fanout4837 (.A(net4840),
    .X(net4837));
 sg13g2_buf_8 fanout4838 (.A(net4840),
    .X(net4838));
 sg13g2_buf_8 fanout4839 (.A(net4840),
    .X(net4839));
 sg13g2_buf_8 fanout4840 (.A(_02747_),
    .X(net4840));
 sg13g2_buf_8 fanout4841 (.A(net4842),
    .X(net4841));
 sg13g2_buf_8 fanout4842 (.A(_10590_),
    .X(net4842));
 sg13g2_buf_8 fanout4843 (.A(net4844),
    .X(net4843));
 sg13g2_buf_8 fanout4844 (.A(_10590_),
    .X(net4844));
 sg13g2_buf_8 fanout4845 (.A(_10530_),
    .X(net4845));
 sg13g2_buf_8 fanout4846 (.A(_10530_),
    .X(net4846));
 sg13g2_buf_8 fanout4847 (.A(net4848),
    .X(net4847));
 sg13g2_buf_8 fanout4848 (.A(_09357_),
    .X(net4848));
 sg13g2_buf_8 fanout4849 (.A(net4851),
    .X(net4849));
 sg13g2_buf_8 fanout4850 (.A(net4851),
    .X(net4850));
 sg13g2_buf_8 fanout4851 (.A(net4852),
    .X(net4851));
 sg13g2_buf_8 fanout4852 (.A(_08914_),
    .X(net4852));
 sg13g2_buf_8 fanout4853 (.A(net4855),
    .X(net4853));
 sg13g2_buf_2 fanout4854 (.A(net4855),
    .X(net4854));
 sg13g2_buf_8 fanout4855 (.A(_07628_),
    .X(net4855));
 sg13g2_buf_8 fanout4856 (.A(net4859),
    .X(net4856));
 sg13g2_buf_8 fanout4857 (.A(net4859),
    .X(net4857));
 sg13g2_buf_8 fanout4858 (.A(net4859),
    .X(net4858));
 sg13g2_buf_8 fanout4859 (.A(net4860),
    .X(net4859));
 sg13g2_buf_8 fanout4860 (.A(_07413_),
    .X(net4860));
 sg13g2_buf_8 fanout4861 (.A(_06279_),
    .X(net4861));
 sg13g2_buf_8 fanout4862 (.A(_06275_),
    .X(net4862));
 sg13g2_buf_8 fanout4863 (.A(net6593),
    .X(net4863));
 sg13g2_buf_8 fanout4864 (.A(net6591),
    .X(net4864));
 sg13g2_buf_8 fanout4865 (.A(_06265_),
    .X(net4865));
 sg13g2_buf_8 fanout4866 (.A(_06263_),
    .X(net4866));
 sg13g2_buf_8 fanout4867 (.A(net4869),
    .X(net4867));
 sg13g2_buf_1 fanout4868 (.A(net4869),
    .X(net4868));
 sg13g2_buf_8 fanout4869 (.A(net4870),
    .X(net4869));
 sg13g2_buf_8 fanout4870 (.A(_05262_),
    .X(net4870));
 sg13g2_buf_8 fanout4871 (.A(net4873),
    .X(net4871));
 sg13g2_buf_8 fanout4872 (.A(net4873),
    .X(net4872));
 sg13g2_buf_8 fanout4873 (.A(_05262_),
    .X(net4873));
 sg13g2_buf_8 fanout4874 (.A(_05262_),
    .X(net4874));
 sg13g2_buf_8 fanout4875 (.A(net4878),
    .X(net4875));
 sg13g2_buf_8 fanout4876 (.A(net4878),
    .X(net4876));
 sg13g2_buf_1 fanout4877 (.A(net4878),
    .X(net4877));
 sg13g2_buf_8 fanout4878 (.A(_04954_),
    .X(net4878));
 sg13g2_buf_8 fanout4879 (.A(_04804_),
    .X(net4879));
 sg13g2_buf_8 fanout4880 (.A(net4881),
    .X(net4880));
 sg13g2_buf_8 fanout4881 (.A(_04665_),
    .X(net4881));
 sg13g2_buf_8 fanout4882 (.A(net4886),
    .X(net4882));
 sg13g2_buf_8 fanout4883 (.A(net4886),
    .X(net4883));
 sg13g2_buf_1 fanout4884 (.A(net4886),
    .X(net4884));
 sg13g2_buf_8 fanout4885 (.A(net4886),
    .X(net4885));
 sg13g2_buf_8 fanout4886 (.A(net4889),
    .X(net4886));
 sg13g2_buf_8 fanout4887 (.A(net4889),
    .X(net4887));
 sg13g2_buf_8 fanout4888 (.A(net4889),
    .X(net4888));
 sg13g2_buf_8 fanout4889 (.A(_04664_),
    .X(net4889));
 sg13g2_buf_8 fanout4890 (.A(net4893),
    .X(net4890));
 sg13g2_buf_1 fanout4891 (.A(net4893),
    .X(net4891));
 sg13g2_buf_8 fanout4892 (.A(net4893),
    .X(net4892));
 sg13g2_buf_2 fanout4893 (.A(_04507_),
    .X(net4893));
 sg13g2_buf_8 fanout4894 (.A(net4895),
    .X(net4894));
 sg13g2_buf_8 fanout4895 (.A(_04503_),
    .X(net4895));
 sg13g2_buf_8 fanout4896 (.A(net4897),
    .X(net4896));
 sg13g2_buf_8 fanout4897 (.A(net4905),
    .X(net4897));
 sg13g2_buf_8 fanout4898 (.A(net4899),
    .X(net4898));
 sg13g2_buf_2 fanout4899 (.A(net4900),
    .X(net4899));
 sg13g2_buf_2 fanout4900 (.A(net4901),
    .X(net4900));
 sg13g2_buf_8 fanout4901 (.A(net4905),
    .X(net4901));
 sg13g2_buf_8 fanout4902 (.A(net4903),
    .X(net4902));
 sg13g2_buf_2 fanout4903 (.A(net4905),
    .X(net4903));
 sg13g2_buf_8 fanout4904 (.A(net4905),
    .X(net4904));
 sg13g2_buf_8 fanout4905 (.A(_04466_),
    .X(net4905));
 sg13g2_buf_8 fanout4906 (.A(net4907),
    .X(net4906));
 sg13g2_buf_8 fanout4907 (.A(_04253_),
    .X(net4907));
 sg13g2_buf_8 fanout4908 (.A(_03788_),
    .X(net4908));
 sg13g2_buf_8 fanout4909 (.A(_03657_),
    .X(net4909));
 sg13g2_buf_2 fanout4910 (.A(_03657_),
    .X(net4910));
 sg13g2_buf_8 fanout4911 (.A(net4913),
    .X(net4911));
 sg13g2_buf_8 fanout4912 (.A(net4913),
    .X(net4912));
 sg13g2_buf_8 fanout4913 (.A(net4915),
    .X(net4913));
 sg13g2_buf_8 fanout4914 (.A(net4915),
    .X(net4914));
 sg13g2_buf_8 fanout4915 (.A(_03202_),
    .X(net4915));
 sg13g2_buf_8 fanout4916 (.A(net4918),
    .X(net4916));
 sg13g2_buf_8 fanout4917 (.A(net4918),
    .X(net4917));
 sg13g2_buf_8 fanout4918 (.A(_10529_),
    .X(net4918));
 sg13g2_buf_8 fanout4919 (.A(net4920),
    .X(net4919));
 sg13g2_buf_8 fanout4920 (.A(_10525_),
    .X(net4920));
 sg13g2_buf_8 fanout4921 (.A(_10525_),
    .X(net4921));
 sg13g2_buf_8 fanout4922 (.A(net4923),
    .X(net4922));
 sg13g2_buf_8 fanout4923 (.A(_09706_),
    .X(net4923));
 sg13g2_buf_8 fanout4924 (.A(net4925),
    .X(net4924));
 sg13g2_buf_8 fanout4925 (.A(_09677_),
    .X(net4925));
 sg13g2_buf_8 fanout4926 (.A(net4927),
    .X(net4926));
 sg13g2_buf_8 fanout4927 (.A(net4938),
    .X(net4927));
 sg13g2_buf_2 fanout4928 (.A(net4929),
    .X(net4928));
 sg13g2_buf_1 fanout4929 (.A(net4935),
    .X(net4929));
 sg13g2_buf_8 fanout4930 (.A(net4935),
    .X(net4930));
 sg13g2_buf_8 fanout4931 (.A(net4935),
    .X(net4931));
 sg13g2_buf_8 fanout4932 (.A(net4933),
    .X(net4932));
 sg13g2_buf_2 fanout4933 (.A(net4934),
    .X(net4933));
 sg13g2_buf_2 fanout4934 (.A(net4935),
    .X(net4934));
 sg13g2_buf_2 fanout4935 (.A(net4938),
    .X(net4935));
 sg13g2_buf_8 fanout4936 (.A(net4937),
    .X(net4936));
 sg13g2_buf_8 fanout4937 (.A(net4938),
    .X(net4937));
 sg13g2_buf_8 fanout4938 (.A(_09652_),
    .X(net4938));
 sg13g2_buf_8 fanout4939 (.A(net4940),
    .X(net4939));
 sg13g2_buf_8 fanout4940 (.A(net4941),
    .X(net4940));
 sg13g2_buf_8 fanout4941 (.A(_09558_),
    .X(net4941));
 sg13g2_buf_8 fanout4942 (.A(net4944),
    .X(net4942));
 sg13g2_buf_1 fanout4943 (.A(net4944),
    .X(net4943));
 sg13g2_buf_8 fanout4944 (.A(_09348_),
    .X(net4944));
 sg13g2_buf_8 fanout4945 (.A(_09347_),
    .X(net4945));
 sg13g2_buf_1 fanout4946 (.A(_09347_),
    .X(net4946));
 sg13g2_buf_8 fanout4947 (.A(net4948),
    .X(net4947));
 sg13g2_buf_8 fanout4948 (.A(net6595),
    .X(net4948));
 sg13g2_buf_8 fanout4949 (.A(_09001_),
    .X(net4949));
 sg13g2_buf_8 fanout4950 (.A(net4953),
    .X(net4950));
 sg13g2_buf_1 fanout4951 (.A(net4952),
    .X(net4951));
 sg13g2_buf_8 fanout4952 (.A(net4953),
    .X(net4952));
 sg13g2_buf_8 fanout4953 (.A(net4954),
    .X(net4953));
 sg13g2_buf_8 fanout4954 (.A(_07414_),
    .X(net4954));
 sg13g2_buf_8 fanout4955 (.A(net4957),
    .X(net4955));
 sg13g2_buf_8 fanout4956 (.A(net4963),
    .X(net4956));
 sg13g2_buf_1 fanout4957 (.A(net4963),
    .X(net4957));
 sg13g2_buf_8 fanout4958 (.A(net4962),
    .X(net4958));
 sg13g2_buf_8 fanout4959 (.A(net4961),
    .X(net4959));
 sg13g2_buf_8 fanout4960 (.A(net4961),
    .X(net4960));
 sg13g2_buf_8 fanout4961 (.A(net4962),
    .X(net4961));
 sg13g2_buf_8 fanout4962 (.A(net4963),
    .X(net4962));
 sg13g2_buf_8 fanout4963 (.A(_07404_),
    .X(net4963));
 sg13g2_buf_8 fanout4964 (.A(net4965),
    .X(net4964));
 sg13g2_buf_8 fanout4965 (.A(_07403_),
    .X(net4965));
 sg13g2_buf_8 fanout4966 (.A(net4968),
    .X(net4966));
 sg13g2_buf_8 fanout4967 (.A(net4968),
    .X(net4967));
 sg13g2_buf_8 fanout4968 (.A(net4974),
    .X(net4968));
 sg13g2_buf_8 fanout4969 (.A(net4973),
    .X(net4969));
 sg13g2_buf_1 fanout4970 (.A(net4973),
    .X(net4970));
 sg13g2_buf_8 fanout4971 (.A(net4973),
    .X(net4971));
 sg13g2_buf_1 fanout4972 (.A(net4973),
    .X(net4972));
 sg13g2_buf_2 fanout4973 (.A(net4974),
    .X(net4973));
 sg13g2_buf_8 fanout4974 (.A(_07403_),
    .X(net4974));
 sg13g2_buf_8 fanout4975 (.A(net4976),
    .X(net4975));
 sg13g2_buf_2 fanout4976 (.A(net4977),
    .X(net4976));
 sg13g2_buf_2 fanout4977 (.A(net4981),
    .X(net4977));
 sg13g2_buf_8 fanout4978 (.A(net4979),
    .X(net4978));
 sg13g2_buf_8 fanout4979 (.A(net4980),
    .X(net4979));
 sg13g2_buf_8 fanout4980 (.A(net4981),
    .X(net4980));
 sg13g2_buf_8 fanout4981 (.A(_07394_),
    .X(net4981));
 sg13g2_buf_8 fanout4982 (.A(net4983),
    .X(net4982));
 sg13g2_buf_8 fanout4983 (.A(net4989),
    .X(net4983));
 sg13g2_buf_8 fanout4984 (.A(net4985),
    .X(net4984));
 sg13g2_buf_8 fanout4985 (.A(net4986),
    .X(net4985));
 sg13g2_buf_8 fanout4986 (.A(net4989),
    .X(net4986));
 sg13g2_buf_8 fanout4987 (.A(net4989),
    .X(net4987));
 sg13g2_buf_8 fanout4988 (.A(net4989),
    .X(net4988));
 sg13g2_buf_8 fanout4989 (.A(_07394_),
    .X(net4989));
 sg13g2_buf_8 fanout4990 (.A(_07389_),
    .X(net4990));
 sg13g2_buf_2 fanout4991 (.A(_07389_),
    .X(net4991));
 sg13g2_buf_8 fanout4992 (.A(net4993),
    .X(net4992));
 sg13g2_buf_8 fanout4993 (.A(net4994),
    .X(net4993));
 sg13g2_buf_8 fanout4994 (.A(_07389_),
    .X(net4994));
 sg13g2_buf_8 fanout4995 (.A(net4996),
    .X(net4995));
 sg13g2_buf_8 fanout4996 (.A(net4997),
    .X(net4996));
 sg13g2_buf_8 fanout4997 (.A(_07388_),
    .X(net4997));
 sg13g2_buf_8 fanout4998 (.A(net5001),
    .X(net4998));
 sg13g2_buf_8 fanout4999 (.A(net5001),
    .X(net4999));
 sg13g2_buf_8 fanout5000 (.A(net5001),
    .X(net5000));
 sg13g2_buf_8 fanout5001 (.A(net5002),
    .X(net5001));
 sg13g2_buf_8 fanout5002 (.A(_07388_),
    .X(net5002));
 sg13g2_buf_8 fanout5003 (.A(net5004),
    .X(net5003));
 sg13g2_buf_8 fanout5004 (.A(net5011),
    .X(net5004));
 sg13g2_buf_8 fanout5005 (.A(net5006),
    .X(net5005));
 sg13g2_buf_8 fanout5006 (.A(net5011),
    .X(net5006));
 sg13g2_buf_8 fanout5007 (.A(net5010),
    .X(net5007));
 sg13g2_buf_8 fanout5008 (.A(net5009),
    .X(net5008));
 sg13g2_buf_8 fanout5009 (.A(net5010),
    .X(net5009));
 sg13g2_buf_8 fanout5010 (.A(net5011),
    .X(net5010));
 sg13g2_buf_8 fanout5011 (.A(_07380_),
    .X(net5011));
 sg13g2_buf_8 fanout5012 (.A(net5020),
    .X(net5012));
 sg13g2_buf_8 fanout5013 (.A(net5014),
    .X(net5013));
 sg13g2_buf_1 fanout5014 (.A(net5019),
    .X(net5014));
 sg13g2_buf_8 fanout5015 (.A(net5016),
    .X(net5015));
 sg13g2_buf_8 fanout5016 (.A(net5019),
    .X(net5016));
 sg13g2_buf_8 fanout5017 (.A(net5019),
    .X(net5017));
 sg13g2_buf_1 fanout5018 (.A(net5019),
    .X(net5018));
 sg13g2_buf_8 fanout5019 (.A(net5020),
    .X(net5019));
 sg13g2_buf_8 fanout5020 (.A(_07379_),
    .X(net5020));
 sg13g2_buf_8 fanout5021 (.A(net5022),
    .X(net5021));
 sg13g2_buf_8 fanout5022 (.A(net5026),
    .X(net5022));
 sg13g2_buf_8 fanout5023 (.A(net5024),
    .X(net5023));
 sg13g2_buf_2 fanout5024 (.A(net5025),
    .X(net5024));
 sg13g2_buf_2 fanout5025 (.A(net5026),
    .X(net5025));
 sg13g2_buf_8 fanout5026 (.A(_05286_),
    .X(net5026));
 sg13g2_buf_8 fanout5027 (.A(net5028),
    .X(net5027));
 sg13g2_buf_1 fanout5028 (.A(net5029),
    .X(net5028));
 sg13g2_buf_8 fanout5029 (.A(_05284_),
    .X(net5029));
 sg13g2_buf_8 fanout5030 (.A(net5031),
    .X(net5030));
 sg13g2_buf_2 fanout5031 (.A(net5032),
    .X(net5031));
 sg13g2_buf_8 fanout5032 (.A(_05284_),
    .X(net5032));
 sg13g2_buf_8 fanout5033 (.A(net5034),
    .X(net5033));
 sg13g2_buf_8 fanout5034 (.A(net5035),
    .X(net5034));
 sg13g2_buf_8 fanout5035 (.A(_04978_),
    .X(net5035));
 sg13g2_buf_2 fanout5036 (.A(net5037),
    .X(net5036));
 sg13g2_buf_8 fanout5037 (.A(net5038),
    .X(net5037));
 sg13g2_buf_1 fanout5038 (.A(net5039),
    .X(net5038));
 sg13g2_buf_2 fanout5039 (.A(net5040),
    .X(net5039));
 sg13g2_buf_8 fanout5040 (.A(_04978_),
    .X(net5040));
 sg13g2_buf_8 fanout5041 (.A(net5042),
    .X(net5041));
 sg13g2_buf_8 fanout5042 (.A(_04977_),
    .X(net5042));
 sg13g2_buf_8 fanout5043 (.A(_04956_),
    .X(net5043));
 sg13g2_buf_8 fanout5044 (.A(net5046),
    .X(net5044));
 sg13g2_buf_8 fanout5045 (.A(net5046),
    .X(net5045));
 sg13g2_buf_8 fanout5046 (.A(_04252_),
    .X(net5046));
 sg13g2_buf_8 fanout5047 (.A(net5050),
    .X(net5047));
 sg13g2_buf_8 fanout5048 (.A(net5050),
    .X(net5048));
 sg13g2_buf_8 fanout5049 (.A(net5050),
    .X(net5049));
 sg13g2_buf_8 fanout5050 (.A(_03830_),
    .X(net5050));
 sg13g2_buf_8 fanout5051 (.A(net5054),
    .X(net5051));
 sg13g2_buf_8 fanout5052 (.A(net5053),
    .X(net5052));
 sg13g2_buf_1 fanout5053 (.A(net5054),
    .X(net5053));
 sg13g2_buf_2 fanout5054 (.A(_03830_),
    .X(net5054));
 sg13g2_buf_8 fanout5055 (.A(net5064),
    .X(net5055));
 sg13g2_buf_8 fanout5056 (.A(net5059),
    .X(net5056));
 sg13g2_buf_8 fanout5057 (.A(net5058),
    .X(net5057));
 sg13g2_buf_8 fanout5058 (.A(net5059),
    .X(net5058));
 sg13g2_buf_8 fanout5059 (.A(net5060),
    .X(net5059));
 sg13g2_buf_2 fanout5060 (.A(net5064),
    .X(net5060));
 sg13g2_buf_8 fanout5061 (.A(net5063),
    .X(net5061));
 sg13g2_buf_8 fanout5062 (.A(net5063),
    .X(net5062));
 sg13g2_buf_8 fanout5063 (.A(net5064),
    .X(net5063));
 sg13g2_buf_8 fanout5064 (.A(_03830_),
    .X(net5064));
 sg13g2_buf_8 fanout5065 (.A(_03785_),
    .X(net5065));
 sg13g2_buf_2 fanout5066 (.A(_03785_),
    .X(net5066));
 sg13g2_buf_8 fanout5067 (.A(_10541_),
    .X(net5067));
 sg13g2_buf_8 fanout5068 (.A(_09723_),
    .X(net5068));
 sg13g2_buf_8 fanout5069 (.A(_09294_),
    .X(net5069));
 sg13g2_buf_8 fanout5070 (.A(_09293_),
    .X(net5070));
 sg13g2_buf_1 fanout5071 (.A(_09293_),
    .X(net5071));
 sg13g2_buf_8 fanout5072 (.A(net5073),
    .X(net5072));
 sg13g2_buf_8 fanout5073 (.A(_09293_),
    .X(net5073));
 sg13g2_buf_8 fanout5074 (.A(_09004_),
    .X(net5074));
 sg13g2_buf_8 fanout5075 (.A(net5076),
    .X(net5075));
 sg13g2_buf_8 fanout5076 (.A(net1622),
    .X(net5076));
 sg13g2_buf_8 fanout5077 (.A(net5079),
    .X(net5077));
 sg13g2_buf_8 fanout5078 (.A(net5079),
    .X(net5078));
 sg13g2_buf_8 fanout5079 (.A(net5080),
    .X(net5079));
 sg13g2_buf_8 fanout5080 (.A(_08875_),
    .X(net5080));
 sg13g2_buf_8 fanout5081 (.A(net5082),
    .X(net5081));
 sg13g2_buf_8 fanout5082 (.A(net5083),
    .X(net5082));
 sg13g2_buf_2 fanout5083 (.A(net5084),
    .X(net5083));
 sg13g2_buf_8 fanout5084 (.A(net5091),
    .X(net5084));
 sg13g2_buf_8 fanout5085 (.A(net5086),
    .X(net5085));
 sg13g2_buf_8 fanout5086 (.A(net5088),
    .X(net5086));
 sg13g2_buf_8 fanout5087 (.A(net5088),
    .X(net5087));
 sg13g2_buf_8 fanout5088 (.A(net5091),
    .X(net5088));
 sg13g2_buf_8 fanout5089 (.A(net5091),
    .X(net5089));
 sg13g2_buf_1 fanout5090 (.A(net5091),
    .X(net5090));
 sg13g2_buf_8 fanout5091 (.A(_08875_),
    .X(net5091));
 sg13g2_buf_8 fanout5092 (.A(net5094),
    .X(net5092));
 sg13g2_buf_8 fanout5093 (.A(net5094),
    .X(net5093));
 sg13g2_buf_2 fanout5094 (.A(net5097),
    .X(net5094));
 sg13g2_buf_8 fanout5095 (.A(net5097),
    .X(net5095));
 sg13g2_buf_1 fanout5096 (.A(net5097),
    .X(net5096));
 sg13g2_buf_8 fanout5097 (.A(net5098),
    .X(net5097));
 sg13g2_buf_8 fanout5098 (.A(_08729_),
    .X(net5098));
 sg13g2_buf_8 fanout5099 (.A(net5100),
    .X(net5099));
 sg13g2_buf_8 fanout5100 (.A(_07613_),
    .X(net5100));
 sg13g2_buf_8 fanout5101 (.A(net5102),
    .X(net5101));
 sg13g2_buf_2 fanout5102 (.A(net5103),
    .X(net5102));
 sg13g2_buf_1 fanout5103 (.A(_07613_),
    .X(net5103));
 sg13g2_buf_8 fanout5104 (.A(net5105),
    .X(net5104));
 sg13g2_buf_8 fanout5105 (.A(net5106),
    .X(net5105));
 sg13g2_buf_8 fanout5106 (.A(_07314_),
    .X(net5106));
 sg13g2_buf_8 fanout5107 (.A(net5110),
    .X(net5107));
 sg13g2_buf_8 fanout5108 (.A(net5110),
    .X(net5108));
 sg13g2_buf_8 fanout5109 (.A(net5110),
    .X(net5109));
 sg13g2_buf_8 fanout5110 (.A(_07313_),
    .X(net5110));
 sg13g2_buf_8 fanout5111 (.A(_07310_),
    .X(net5111));
 sg13g2_buf_8 fanout5112 (.A(net5113),
    .X(net5112));
 sg13g2_buf_8 fanout5113 (.A(_07310_),
    .X(net5113));
 sg13g2_buf_8 fanout5114 (.A(_07306_),
    .X(net5114));
 sg13g2_buf_8 fanout5115 (.A(net5116),
    .X(net5115));
 sg13g2_buf_8 fanout5116 (.A(_07306_),
    .X(net5116));
 sg13g2_buf_8 fanout5117 (.A(net5120),
    .X(net5117));
 sg13g2_buf_8 fanout5118 (.A(net5119),
    .X(net5118));
 sg13g2_buf_8 fanout5119 (.A(net5120),
    .X(net5119));
 sg13g2_buf_8 fanout5120 (.A(_04993_),
    .X(net5120));
 sg13g2_buf_8 fanout5121 (.A(_04990_),
    .X(net5121));
 sg13g2_buf_8 fanout5122 (.A(net5124),
    .X(net5122));
 sg13g2_buf_8 fanout5123 (.A(net5124),
    .X(net5123));
 sg13g2_buf_8 fanout5124 (.A(_04250_),
    .X(net5124));
 sg13g2_buf_8 fanout5125 (.A(net5126),
    .X(net5125));
 sg13g2_buf_8 fanout5126 (.A(_04250_),
    .X(net5126));
 sg13g2_buf_2 fanout5127 (.A(net5128),
    .X(net5127));
 sg13g2_buf_1 fanout5128 (.A(_04250_),
    .X(net5128));
 sg13g2_buf_8 fanout5129 (.A(_03839_),
    .X(net5129));
 sg13g2_buf_2 fanout5130 (.A(_03839_),
    .X(net5130));
 sg13g2_buf_8 fanout5131 (.A(net5133),
    .X(net5131));
 sg13g2_buf_2 fanout5132 (.A(net5133),
    .X(net5132));
 sg13g2_buf_8 fanout5133 (.A(_03839_),
    .X(net5133));
 sg13g2_buf_8 fanout5134 (.A(net5135),
    .X(net5134));
 sg13g2_buf_8 fanout5135 (.A(net5136),
    .X(net5135));
 sg13g2_buf_2 fanout5136 (.A(net5137),
    .X(net5136));
 sg13g2_buf_8 fanout5137 (.A(net5138),
    .X(net5137));
 sg13g2_buf_8 fanout5138 (.A(_03831_),
    .X(net5138));
 sg13g2_buf_8 fanout5139 (.A(net5145),
    .X(net5139));
 sg13g2_buf_1 fanout5140 (.A(net5145),
    .X(net5140));
 sg13g2_buf_8 fanout5141 (.A(net5144),
    .X(net5141));
 sg13g2_buf_8 fanout5142 (.A(net5143),
    .X(net5142));
 sg13g2_buf_8 fanout5143 (.A(net5144),
    .X(net5143));
 sg13g2_buf_8 fanout5144 (.A(net5145),
    .X(net5144));
 sg13g2_buf_8 fanout5145 (.A(_03831_),
    .X(net5145));
 sg13g2_buf_8 fanout5146 (.A(_03653_),
    .X(net5146));
 sg13g2_buf_8 fanout5147 (.A(net5148),
    .X(net5147));
 sg13g2_buf_8 fanout5148 (.A(net5150),
    .X(net5148));
 sg13g2_buf_8 fanout5149 (.A(net5150),
    .X(net5149));
 sg13g2_buf_2 fanout5150 (.A(net5151),
    .X(net5150));
 sg13g2_buf_8 fanout5151 (.A(_10627_),
    .X(net5151));
 sg13g2_buf_8 fanout5152 (.A(net5156),
    .X(net5152));
 sg13g2_buf_1 fanout5153 (.A(net5156),
    .X(net5153));
 sg13g2_buf_8 fanout5154 (.A(net5156),
    .X(net5154));
 sg13g2_buf_1 fanout5155 (.A(net5156),
    .X(net5155));
 sg13g2_buf_2 fanout5156 (.A(net5157),
    .X(net5156));
 sg13g2_buf_8 fanout5157 (.A(_10625_),
    .X(net5157));
 sg13g2_buf_8 fanout5158 (.A(net5160),
    .X(net5158));
 sg13g2_buf_8 fanout5159 (.A(net5160),
    .X(net5159));
 sg13g2_buf_8 fanout5160 (.A(_09564_),
    .X(net5160));
 sg13g2_buf_8 fanout5161 (.A(net5163),
    .X(net5161));
 sg13g2_buf_1 fanout5162 (.A(net5163),
    .X(net5162));
 sg13g2_buf_8 fanout5163 (.A(_09550_),
    .X(net5163));
 sg13g2_buf_8 fanout5164 (.A(net5165),
    .X(net5164));
 sg13g2_buf_8 fanout5165 (.A(net5168),
    .X(net5165));
 sg13g2_buf_2 fanout5166 (.A(net5167),
    .X(net5166));
 sg13g2_buf_8 fanout5167 (.A(net5168),
    .X(net5167));
 sg13g2_buf_8 fanout5168 (.A(_09549_),
    .X(net5168));
 sg13g2_buf_8 fanout5169 (.A(net5170),
    .X(net5169));
 sg13g2_buf_8 fanout5170 (.A(net5171),
    .X(net5170));
 sg13g2_buf_8 fanout5171 (.A(net5172),
    .X(net5171));
 sg13g2_buf_1 fanout5172 (.A(net5173),
    .X(net5172));
 sg13g2_buf_8 fanout5173 (.A(_09300_),
    .X(net5173));
 sg13g2_buf_8 fanout5174 (.A(net5176),
    .X(net5174));
 sg13g2_buf_1 fanout5175 (.A(net5176),
    .X(net5175));
 sg13g2_buf_2 fanout5176 (.A(_08730_),
    .X(net5176));
 sg13g2_buf_8 fanout5177 (.A(net5179),
    .X(net5177));
 sg13g2_buf_1 fanout5178 (.A(net5179),
    .X(net5178));
 sg13g2_buf_8 fanout5179 (.A(_07649_),
    .X(net5179));
 sg13g2_buf_8 fanout5180 (.A(net5182),
    .X(net5180));
 sg13g2_buf_8 fanout5181 (.A(net5182),
    .X(net5181));
 sg13g2_buf_8 fanout5182 (.A(_07649_),
    .X(net5182));
 sg13g2_buf_8 fanout5183 (.A(net5184),
    .X(net5183));
 sg13g2_buf_8 fanout5184 (.A(_07615_),
    .X(net5184));
 sg13g2_buf_8 fanout5185 (.A(net5186),
    .X(net5185));
 sg13g2_buf_8 fanout5186 (.A(_07615_),
    .X(net5186));
 sg13g2_buf_8 fanout5187 (.A(net5189),
    .X(net5187));
 sg13g2_buf_8 fanout5188 (.A(net5189),
    .X(net5188));
 sg13g2_buf_8 fanout5189 (.A(_07612_),
    .X(net5189));
 sg13g2_buf_8 fanout5190 (.A(_07604_),
    .X(net5190));
 sg13g2_buf_8 fanout5191 (.A(net5192),
    .X(net5191));
 sg13g2_buf_8 fanout5192 (.A(net5193),
    .X(net5192));
 sg13g2_buf_8 fanout5193 (.A(_07578_),
    .X(net5193));
 sg13g2_buf_8 fanout5194 (.A(net5195),
    .X(net5194));
 sg13g2_buf_8 fanout5195 (.A(_07578_),
    .X(net5195));
 sg13g2_buf_8 fanout5196 (.A(net5197),
    .X(net5196));
 sg13g2_buf_8 fanout5197 (.A(_07573_),
    .X(net5197));
 sg13g2_buf_8 fanout5198 (.A(net5199),
    .X(net5198));
 sg13g2_buf_8 fanout5199 (.A(net5200),
    .X(net5199));
 sg13g2_buf_2 fanout5200 (.A(net5201),
    .X(net5200));
 sg13g2_buf_1 fanout5201 (.A(_07572_),
    .X(net5201));
 sg13g2_buf_8 fanout5202 (.A(net5204),
    .X(net5202));
 sg13g2_buf_2 fanout5203 (.A(net5204),
    .X(net5203));
 sg13g2_buf_8 fanout5204 (.A(_07572_),
    .X(net5204));
 sg13g2_buf_8 fanout5205 (.A(_07309_),
    .X(net5205));
 sg13g2_buf_8 fanout5206 (.A(_07305_),
    .X(net5206));
 sg13g2_buf_8 fanout5207 (.A(_07304_),
    .X(net5207));
 sg13g2_buf_8 fanout5208 (.A(net5209),
    .X(net5208));
 sg13g2_buf_2 fanout5209 (.A(_07291_),
    .X(net5209));
 sg13g2_buf_2 fanout5210 (.A(net5211),
    .X(net5210));
 sg13g2_buf_1 fanout5211 (.A(net5212),
    .X(net5211));
 sg13g2_buf_8 fanout5212 (.A(net5213),
    .X(net5212));
 sg13g2_buf_8 fanout5213 (.A(_07082_),
    .X(net5213));
 sg13g2_buf_8 fanout5214 (.A(net5216),
    .X(net5214));
 sg13g2_buf_8 fanout5215 (.A(net5216),
    .X(net5215));
 sg13g2_buf_8 fanout5216 (.A(_07082_),
    .X(net5216));
 sg13g2_buf_8 fanout5217 (.A(net5218),
    .X(net5217));
 sg13g2_buf_8 fanout5218 (.A(net5219),
    .X(net5218));
 sg13g2_buf_8 fanout5219 (.A(_07081_),
    .X(net5219));
 sg13g2_buf_8 fanout5220 (.A(_07034_),
    .X(net5220));
 sg13g2_buf_8 fanout5221 (.A(net5224),
    .X(net5221));
 sg13g2_buf_8 fanout5222 (.A(net5224),
    .X(net5222));
 sg13g2_buf_8 fanout5223 (.A(net5224),
    .X(net5223));
 sg13g2_buf_8 fanout5224 (.A(_07033_),
    .X(net5224));
 sg13g2_buf_8 fanout5225 (.A(_07033_),
    .X(net5225));
 sg13g2_buf_8 fanout5226 (.A(_07033_),
    .X(net5226));
 sg13g2_buf_8 fanout5227 (.A(net5228),
    .X(net5227));
 sg13g2_buf_8 fanout5228 (.A(_06996_),
    .X(net5228));
 sg13g2_buf_8 fanout5229 (.A(_06992_),
    .X(net5229));
 sg13g2_buf_2 fanout5230 (.A(net5231),
    .X(net5230));
 sg13g2_buf_2 fanout5231 (.A(net5233),
    .X(net5231));
 sg13g2_buf_8 fanout5232 (.A(net5233),
    .X(net5232));
 sg13g2_buf_1 fanout5233 (.A(net5234),
    .X(net5233));
 sg13g2_buf_8 fanout5234 (.A(net5235),
    .X(net5234));
 sg13g2_buf_8 fanout5235 (.A(_06991_),
    .X(net5235));
 sg13g2_buf_8 fanout5236 (.A(net5237),
    .X(net5236));
 sg13g2_buf_8 fanout5237 (.A(_06476_),
    .X(net5237));
 sg13g2_buf_8 fanout5238 (.A(net5239),
    .X(net5238));
 sg13g2_buf_8 fanout5239 (.A(_06467_),
    .X(net5239));
 sg13g2_buf_8 fanout5240 (.A(net5241),
    .X(net5240));
 sg13g2_buf_8 fanout5241 (.A(_06458_),
    .X(net5241));
 sg13g2_buf_8 fanout5242 (.A(net5243),
    .X(net5242));
 sg13g2_buf_8 fanout5243 (.A(_06449_),
    .X(net5243));
 sg13g2_buf_8 fanout5244 (.A(net5246),
    .X(net5244));
 sg13g2_buf_1 fanout5245 (.A(net5246),
    .X(net5245));
 sg13g2_buf_8 fanout5246 (.A(_06440_),
    .X(net5246));
 sg13g2_buf_8 fanout5247 (.A(net5249),
    .X(net5247));
 sg13g2_buf_1 fanout5248 (.A(net5249),
    .X(net5248));
 sg13g2_buf_8 fanout5249 (.A(_06431_),
    .X(net5249));
 sg13g2_buf_8 fanout5250 (.A(net5251),
    .X(net5250));
 sg13g2_buf_8 fanout5251 (.A(net5252),
    .X(net5251));
 sg13g2_buf_8 fanout5252 (.A(_06422_),
    .X(net5252));
 sg13g2_buf_8 fanout5253 (.A(net5254),
    .X(net5253));
 sg13g2_buf_8 fanout5254 (.A(net5256),
    .X(net5254));
 sg13g2_buf_8 fanout5255 (.A(net5256),
    .X(net5255));
 sg13g2_buf_8 fanout5256 (.A(_04924_),
    .X(net5256));
 sg13g2_buf_8 fanout5257 (.A(net5258),
    .X(net5257));
 sg13g2_buf_8 fanout5258 (.A(_04499_),
    .X(net5258));
 sg13g2_buf_8 fanout5259 (.A(net5260),
    .X(net5259));
 sg13g2_buf_2 fanout5260 (.A(net5261),
    .X(net5260));
 sg13g2_buf_1 fanout5261 (.A(_04499_),
    .X(net5261));
 sg13g2_buf_8 fanout5262 (.A(net5263),
    .X(net5262));
 sg13g2_buf_8 fanout5263 (.A(net5265),
    .X(net5263));
 sg13g2_buf_8 fanout5264 (.A(net5265),
    .X(net5264));
 sg13g2_buf_8 fanout5265 (.A(_04498_),
    .X(net5265));
 sg13g2_buf_8 fanout5266 (.A(net5267),
    .X(net5266));
 sg13g2_buf_8 fanout5267 (.A(_04498_),
    .X(net5267));
 sg13g2_buf_8 fanout5268 (.A(net5269),
    .X(net5268));
 sg13g2_buf_8 fanout5269 (.A(net5270),
    .X(net5269));
 sg13g2_buf_8 fanout5270 (.A(_10581_),
    .X(net5270));
 sg13g2_buf_8 fanout5271 (.A(net5273),
    .X(net5271));
 sg13g2_buf_8 fanout5272 (.A(net5273),
    .X(net5272));
 sg13g2_buf_8 fanout5273 (.A(_09454_),
    .X(net5273));
 sg13g2_buf_1 fanout5274 (.A(_09454_),
    .X(net5274));
 sg13g2_buf_8 fanout5275 (.A(net5276),
    .X(net5275));
 sg13g2_buf_8 fanout5276 (.A(net5277),
    .X(net5276));
 sg13g2_buf_8 fanout5277 (.A(_09454_),
    .X(net5277));
 sg13g2_buf_8 fanout5278 (.A(_09453_),
    .X(net5278));
 sg13g2_buf_2 fanout5279 (.A(_09453_),
    .X(net5279));
 sg13g2_buf_2 fanout5280 (.A(net5281),
    .X(net5280));
 sg13g2_buf_2 fanout5281 (.A(_09394_),
    .X(net5281));
 sg13g2_buf_8 fanout5282 (.A(_09336_),
    .X(net5282));
 sg13g2_buf_1 fanout5283 (.A(_09336_),
    .X(net5283));
 sg13g2_buf_8 fanout5284 (.A(_09336_),
    .X(net5284));
 sg13g2_buf_8 fanout5285 (.A(net6574),
    .X(net5285));
 sg13g2_buf_8 fanout5286 (.A(_07650_),
    .X(net5286));
 sg13g2_buf_1 fanout5287 (.A(_07650_),
    .X(net5287));
 sg13g2_buf_8 fanout5288 (.A(_07608_),
    .X(net5288));
 sg13g2_buf_8 fanout5289 (.A(net5290),
    .X(net5289));
 sg13g2_buf_8 fanout5290 (.A(net5291),
    .X(net5290));
 sg13g2_buf_8 fanout5291 (.A(net5292),
    .X(net5291));
 sg13g2_buf_8 fanout5292 (.A(_07577_),
    .X(net5292));
 sg13g2_buf_8 fanout5293 (.A(_07577_),
    .X(net5293));
 sg13g2_buf_8 fanout5294 (.A(_07298_),
    .X(net5294));
 sg13g2_buf_8 fanout5295 (.A(_07080_),
    .X(net5295));
 sg13g2_buf_1 fanout5296 (.A(_07080_),
    .X(net5296));
 sg13g2_buf_8 fanout5297 (.A(net5298),
    .X(net5297));
 sg13g2_buf_8 fanout5298 (.A(net5300),
    .X(net5298));
 sg13g2_buf_8 fanout5299 (.A(net5300),
    .X(net5299));
 sg13g2_buf_8 fanout5300 (.A(_07042_),
    .X(net5300));
 sg13g2_buf_8 fanout5301 (.A(net5303),
    .X(net5301));
 sg13g2_buf_8 fanout5302 (.A(net5303),
    .X(net5302));
 sg13g2_buf_8 fanout5303 (.A(_07041_),
    .X(net5303));
 sg13g2_buf_8 fanout5304 (.A(net5306),
    .X(net5304));
 sg13g2_buf_8 fanout5305 (.A(net5306),
    .X(net5305));
 sg13g2_buf_8 fanout5306 (.A(_07041_),
    .X(net5306));
 sg13g2_buf_8 fanout5307 (.A(net5308),
    .X(net5307));
 sg13g2_buf_8 fanout5308 (.A(net5309),
    .X(net5308));
 sg13g2_buf_8 fanout5309 (.A(_07032_),
    .X(net5309));
 sg13g2_buf_8 fanout5310 (.A(net5312),
    .X(net5310));
 sg13g2_buf_8 fanout5311 (.A(net5312),
    .X(net5311));
 sg13g2_buf_8 fanout5312 (.A(net5313),
    .X(net5312));
 sg13g2_buf_8 fanout5313 (.A(net5314),
    .X(net5313));
 sg13g2_buf_8 fanout5314 (.A(_07032_),
    .X(net5314));
 sg13g2_buf_8 fanout5315 (.A(_04974_),
    .X(net5315));
 sg13g2_buf_8 fanout5316 (.A(net5317),
    .X(net5316));
 sg13g2_buf_8 fanout5317 (.A(net5318),
    .X(net5317));
 sg13g2_buf_8 fanout5318 (.A(_04497_),
    .X(net5318));
 sg13g2_buf_8 fanout5319 (.A(net5323),
    .X(net5319));
 sg13g2_buf_2 fanout5320 (.A(net5321),
    .X(net5320));
 sg13g2_buf_1 fanout5321 (.A(net5322),
    .X(net5321));
 sg13g2_buf_2 fanout5322 (.A(net5323),
    .X(net5322));
 sg13g2_buf_1 fanout5323 (.A(net5324),
    .X(net5323));
 sg13g2_buf_8 fanout5324 (.A(_04496_),
    .X(net5324));
 sg13g2_buf_8 fanout5325 (.A(net5326),
    .X(net5325));
 sg13g2_buf_8 fanout5326 (.A(_04496_),
    .X(net5326));
 sg13g2_buf_8 fanout5327 (.A(_02737_),
    .X(net5327));
 sg13g2_buf_2 fanout5328 (.A(_02737_),
    .X(net5328));
 sg13g2_buf_8 fanout5329 (.A(_09702_),
    .X(net5329));
 sg13g2_buf_8 fanout5330 (.A(net5331),
    .X(net5330));
 sg13g2_buf_8 fanout5331 (.A(_09125_),
    .X(net5331));
 sg13g2_buf_8 fanout5332 (.A(net5335),
    .X(net5332));
 sg13g2_buf_8 fanout5333 (.A(net5334),
    .X(net5333));
 sg13g2_buf_8 fanout5334 (.A(net5335),
    .X(net5334));
 sg13g2_buf_8 fanout5335 (.A(_09117_),
    .X(net5335));
 sg13g2_buf_8 fanout5336 (.A(net5337),
    .X(net5336));
 sg13g2_buf_8 fanout5337 (.A(net5338),
    .X(net5337));
 sg13g2_buf_8 fanout5338 (.A(net1391),
    .X(net5338));
 sg13g2_buf_8 fanout5339 (.A(_08852_),
    .X(net5339));
 sg13g2_buf_8 fanout5340 (.A(_08742_),
    .X(net5340));
 sg13g2_buf_8 fanout5341 (.A(_08741_),
    .X(net5341));
 sg13g2_buf_8 fanout5342 (.A(net5343),
    .X(net5342));
 sg13g2_buf_8 fanout5343 (.A(_07302_),
    .X(net5343));
 sg13g2_buf_8 fanout5344 (.A(_07030_),
    .X(net5344));
 sg13g2_buf_8 fanout5345 (.A(net5346),
    .X(net5345));
 sg13g2_buf_8 fanout5346 (.A(_06935_),
    .X(net5346));
 sg13g2_buf_2 fanout5347 (.A(net5348),
    .X(net5347));
 sg13g2_buf_8 fanout5348 (.A(_06934_),
    .X(net5348));
 sg13g2_buf_8 fanout5349 (.A(_06933_),
    .X(net5349));
 sg13g2_buf_8 fanout5350 (.A(net5351),
    .X(net5350));
 sg13g2_buf_8 fanout5351 (.A(net5352),
    .X(net5351));
 sg13g2_buf_8 fanout5352 (.A(_06932_),
    .X(net5352));
 sg13g2_buf_8 fanout5353 (.A(net5354),
    .X(net5353));
 sg13g2_buf_8 fanout5354 (.A(net5355),
    .X(net5354));
 sg13g2_buf_8 fanout5355 (.A(_06931_),
    .X(net5355));
 sg13g2_buf_8 fanout5356 (.A(_06870_),
    .X(net5356));
 sg13g2_buf_1 fanout5357 (.A(_06870_),
    .X(net5357));
 sg13g2_buf_8 fanout5358 (.A(_06864_),
    .X(net5358));
 sg13g2_buf_8 fanout5359 (.A(_06864_),
    .X(net5359));
 sg13g2_buf_8 fanout5360 (.A(net5361),
    .X(net5360));
 sg13g2_buf_8 fanout5361 (.A(_06864_),
    .X(net5361));
 sg13g2_buf_8 fanout5362 (.A(net5364),
    .X(net5362));
 sg13g2_buf_8 fanout5363 (.A(net5364),
    .X(net5363));
 sg13g2_buf_8 fanout5364 (.A(net5367),
    .X(net5364));
 sg13g2_buf_8 fanout5365 (.A(net5366),
    .X(net5365));
 sg13g2_buf_8 fanout5366 (.A(net5367),
    .X(net5366));
 sg13g2_buf_8 fanout5367 (.A(_06863_),
    .X(net5367));
 sg13g2_buf_8 fanout5368 (.A(net5372),
    .X(net5368));
 sg13g2_buf_8 fanout5369 (.A(net5371),
    .X(net5369));
 sg13g2_buf_8 fanout5370 (.A(net5371),
    .X(net5370));
 sg13g2_buf_8 fanout5371 (.A(net5372),
    .X(net5371));
 sg13g2_buf_8 fanout5372 (.A(_06863_),
    .X(net5372));
 sg13g2_buf_8 fanout5373 (.A(_06797_),
    .X(net5373));
 sg13g2_buf_8 fanout5374 (.A(_06795_),
    .X(net5374));
 sg13g2_buf_8 fanout5375 (.A(_06794_),
    .X(net5375));
 sg13g2_buf_8 fanout5376 (.A(_06794_),
    .X(net5376));
 sg13g2_buf_8 fanout5377 (.A(net5378),
    .X(net5377));
 sg13g2_buf_8 fanout5378 (.A(_06662_),
    .X(net5378));
 sg13g2_buf_8 fanout5379 (.A(_06553_),
    .X(net5379));
 sg13g2_buf_8 fanout5380 (.A(_06553_),
    .X(net5380));
 sg13g2_buf_8 fanout5381 (.A(net5382),
    .X(net5381));
 sg13g2_buf_8 fanout5382 (.A(net5385),
    .X(net5382));
 sg13g2_buf_8 fanout5383 (.A(net5384),
    .X(net5383));
 sg13g2_buf_2 fanout5384 (.A(net5385),
    .X(net5384));
 sg13g2_buf_8 fanout5385 (.A(_06551_),
    .X(net5385));
 sg13g2_buf_8 fanout5386 (.A(_06547_),
    .X(net5386));
 sg13g2_buf_8 fanout5387 (.A(_00007_),
    .X(net5387));
 sg13g2_buf_8 fanout5388 (.A(net5389),
    .X(net5388));
 sg13g2_buf_8 fanout5389 (.A(net5390),
    .X(net5389));
 sg13g2_buf_8 fanout5390 (.A(_00006_),
    .X(net5390));
 sg13g2_buf_8 fanout5391 (.A(_00006_),
    .X(net5391));
 sg13g2_buf_8 fanout5392 (.A(net5394),
    .X(net5392));
 sg13g2_buf_8 fanout5393 (.A(net5394),
    .X(net5393));
 sg13g2_buf_8 fanout5394 (.A(net5398),
    .X(net5394));
 sg13g2_buf_8 fanout5395 (.A(net5398),
    .X(net5395));
 sg13g2_buf_8 fanout5396 (.A(net5397),
    .X(net5396));
 sg13g2_buf_8 fanout5397 (.A(net5398),
    .X(net5397));
 sg13g2_buf_8 fanout5398 (.A(_00005_),
    .X(net5398));
 sg13g2_buf_8 fanout5399 (.A(net5401),
    .X(net5399));
 sg13g2_buf_1 fanout5400 (.A(net5401),
    .X(net5400));
 sg13g2_buf_8 fanout5401 (.A(_00010_),
    .X(net5401));
 sg13g2_buf_8 fanout5402 (.A(net5403),
    .X(net5402));
 sg13g2_buf_8 fanout5403 (.A(_00009_),
    .X(net5403));
 sg13g2_buf_8 fanout5404 (.A(net5405),
    .X(net5404));
 sg13g2_buf_8 fanout5405 (.A(_00008_),
    .X(net5405));
 sg13g2_buf_8 fanout5406 (.A(net5407),
    .X(net5406));
 sg13g2_buf_8 fanout5407 (.A(_00013_),
    .X(net5407));
 sg13g2_buf_8 fanout5408 (.A(net5410),
    .X(net5408));
 sg13g2_buf_1 fanout5409 (.A(net5410),
    .X(net5409));
 sg13g2_buf_8 fanout5410 (.A(_00012_),
    .X(net5410));
 sg13g2_buf_8 fanout5411 (.A(_00012_),
    .X(net5411));
 sg13g2_buf_1 fanout5412 (.A(_00012_),
    .X(net5412));
 sg13g2_buf_8 fanout5413 (.A(net5416),
    .X(net5413));
 sg13g2_buf_8 fanout5414 (.A(net5416),
    .X(net5414));
 sg13g2_buf_8 fanout5415 (.A(net5416),
    .X(net5415));
 sg13g2_buf_8 fanout5416 (.A(_00011_),
    .X(net5416));
 sg13g2_buf_8 fanout5417 (.A(net5418),
    .X(net5417));
 sg13g2_buf_8 fanout5418 (.A(net5421),
    .X(net5418));
 sg13g2_buf_8 fanout5419 (.A(net5421),
    .X(net5419));
 sg13g2_buf_1 fanout5420 (.A(net5421),
    .X(net5420));
 sg13g2_buf_2 fanout5421 (.A(_00011_),
    .X(net5421));
 sg13g2_buf_8 fanout5422 (.A(\fpga_top.uart_top.uart_send_char.send_cntr[3] ),
    .X(net5422));
 sg13g2_buf_8 fanout5423 (.A(net6507),
    .X(net5423));
 sg13g2_buf_8 fanout5424 (.A(net5425),
    .X(net5424));
 sg13g2_buf_8 fanout5425 (.A(net6584),
    .X(net5425));
 sg13g2_buf_8 fanout5426 (.A(net6280),
    .X(net5426));
 sg13g2_buf_8 fanout5427 (.A(net6280),
    .X(net5427));
 sg13g2_buf_2 fanout5428 (.A(net5433),
    .X(net5428));
 sg13g2_buf_2 fanout5429 (.A(net5433),
    .X(net5429));
 sg13g2_buf_1 fanout5430 (.A(net5433),
    .X(net5430));
 sg13g2_buf_2 fanout5431 (.A(net5432),
    .X(net5431));
 sg13g2_buf_1 fanout5432 (.A(net5433),
    .X(net5432));
 sg13g2_buf_1 fanout5433 (.A(net5437),
    .X(net5433));
 sg13g2_buf_8 fanout5434 (.A(net5437),
    .X(net5434));
 sg13g2_buf_8 fanout5435 (.A(net5436),
    .X(net5435));
 sg13g2_buf_8 fanout5436 (.A(net5437),
    .X(net5436));
 sg13g2_buf_8 fanout5437 (.A(\fpga_top.cpu_top.data_rw_mem.dma_io_ren_wb ),
    .X(net5437));
 sg13g2_buf_8 fanout5438 (.A(net5439),
    .X(net5438));
 sg13g2_buf_2 fanout5439 (.A(net5440),
    .X(net5439));
 sg13g2_buf_2 fanout5440 (.A(net6482),
    .X(net5440));
 sg13g2_buf_8 fanout5441 (.A(net5445),
    .X(net5441));
 sg13g2_buf_8 fanout5442 (.A(net5445),
    .X(net5442));
 sg13g2_buf_8 fanout5443 (.A(net5445),
    .X(net5443));
 sg13g2_buf_1 fanout5444 (.A(net5445),
    .X(net5444));
 sg13g2_buf_8 fanout5445 (.A(_00004_),
    .X(net5445));
 sg13g2_buf_8 fanout5446 (.A(net5451),
    .X(net5446));
 sg13g2_buf_8 fanout5447 (.A(net5451),
    .X(net5447));
 sg13g2_buf_8 fanout5448 (.A(net5450),
    .X(net5448));
 sg13g2_buf_8 fanout5449 (.A(net5451),
    .X(net5449));
 sg13g2_buf_8 fanout5450 (.A(net5451),
    .X(net5450));
 sg13g2_buf_8 fanout5451 (.A(_00004_),
    .X(net5451));
 sg13g2_buf_8 fanout5452 (.A(net5456),
    .X(net5452));
 sg13g2_buf_8 fanout5453 (.A(net5456),
    .X(net5453));
 sg13g2_buf_8 fanout5454 (.A(net5456),
    .X(net5454));
 sg13g2_buf_8 fanout5455 (.A(net5456),
    .X(net5455));
 sg13g2_buf_8 fanout5456 (.A(_00003_),
    .X(net5456));
 sg13g2_buf_8 fanout5457 (.A(net5462),
    .X(net5457));
 sg13g2_buf_8 fanout5458 (.A(net5461),
    .X(net5458));
 sg13g2_buf_8 fanout5459 (.A(net5460),
    .X(net5459));
 sg13g2_buf_8 fanout5460 (.A(net5461),
    .X(net5460));
 sg13g2_buf_8 fanout5461 (.A(net5462),
    .X(net5461));
 sg13g2_buf_8 fanout5462 (.A(_00003_),
    .X(net5462));
 sg13g2_buf_8 fanout5463 (.A(net5464),
    .X(net5463));
 sg13g2_buf_8 fanout5464 (.A(net5468),
    .X(net5464));
 sg13g2_buf_8 fanout5465 (.A(net5466),
    .X(net5465));
 sg13g2_buf_8 fanout5466 (.A(net5468),
    .X(net5466));
 sg13g2_buf_2 fanout5467 (.A(net5468),
    .X(net5467));
 sg13g2_buf_8 fanout5468 (.A(net5478),
    .X(net5468));
 sg13g2_buf_8 fanout5469 (.A(net5478),
    .X(net5469));
 sg13g2_buf_8 fanout5470 (.A(net5471),
    .X(net5470));
 sg13g2_buf_8 fanout5471 (.A(net5477),
    .X(net5471));
 sg13g2_buf_8 fanout5472 (.A(net5476),
    .X(net5472));
 sg13g2_buf_1 fanout5473 (.A(net5476),
    .X(net5473));
 sg13g2_buf_8 fanout5474 (.A(net5476),
    .X(net5474));
 sg13g2_buf_8 fanout5475 (.A(net5476),
    .X(net5475));
 sg13g2_buf_8 fanout5476 (.A(net5477),
    .X(net5476));
 sg13g2_buf_8 fanout5477 (.A(net5478),
    .X(net5477));
 sg13g2_buf_8 fanout5478 (.A(_00002_),
    .X(net5478));
 sg13g2_buf_8 fanout5479 (.A(net5482),
    .X(net5479));
 sg13g2_buf_8 fanout5480 (.A(net5481),
    .X(net5480));
 sg13g2_buf_8 fanout5481 (.A(net5482),
    .X(net5481));
 sg13g2_buf_8 fanout5482 (.A(net5488),
    .X(net5482));
 sg13g2_buf_8 fanout5483 (.A(net5485),
    .X(net5483));
 sg13g2_buf_8 fanout5484 (.A(net5485),
    .X(net5484));
 sg13g2_buf_8 fanout5485 (.A(net5488),
    .X(net5485));
 sg13g2_buf_8 fanout5486 (.A(net5488),
    .X(net5486));
 sg13g2_buf_8 fanout5487 (.A(net5488),
    .X(net5487));
 sg13g2_buf_8 fanout5488 (.A(net5523),
    .X(net5488));
 sg13g2_buf_8 fanout5489 (.A(net5490),
    .X(net5489));
 sg13g2_buf_8 fanout5490 (.A(net5493),
    .X(net5490));
 sg13g2_buf_8 fanout5491 (.A(net5493),
    .X(net5491));
 sg13g2_buf_8 fanout5492 (.A(net5493),
    .X(net5492));
 sg13g2_buf_8 fanout5493 (.A(net5523),
    .X(net5493));
 sg13g2_buf_8 fanout5494 (.A(net5496),
    .X(net5494));
 sg13g2_buf_8 fanout5495 (.A(net5499),
    .X(net5495));
 sg13g2_buf_8 fanout5496 (.A(net5499),
    .X(net5496));
 sg13g2_buf_8 fanout5497 (.A(net5499),
    .X(net5497));
 sg13g2_buf_8 fanout5498 (.A(net5499),
    .X(net5498));
 sg13g2_buf_8 fanout5499 (.A(net5523),
    .X(net5499));
 sg13g2_buf_8 fanout5500 (.A(net5511),
    .X(net5500));
 sg13g2_buf_8 fanout5501 (.A(net5511),
    .X(net5501));
 sg13g2_buf_8 fanout5502 (.A(net5504),
    .X(net5502));
 sg13g2_buf_8 fanout5503 (.A(net5504),
    .X(net5503));
 sg13g2_buf_8 fanout5504 (.A(net5511),
    .X(net5504));
 sg13g2_buf_8 fanout5505 (.A(net5510),
    .X(net5505));
 sg13g2_buf_8 fanout5506 (.A(net5510),
    .X(net5506));
 sg13g2_buf_8 fanout5507 (.A(net5509),
    .X(net5507));
 sg13g2_buf_8 fanout5508 (.A(net5510),
    .X(net5508));
 sg13g2_buf_8 fanout5509 (.A(net5510),
    .X(net5509));
 sg13g2_buf_8 fanout5510 (.A(net5511),
    .X(net5510));
 sg13g2_buf_8 fanout5511 (.A(net5523),
    .X(net5511));
 sg13g2_buf_8 fanout5512 (.A(net5516),
    .X(net5512));
 sg13g2_buf_2 fanout5513 (.A(net5516),
    .X(net5513));
 sg13g2_buf_8 fanout5514 (.A(net5515),
    .X(net5514));
 sg13g2_buf_8 fanout5515 (.A(net5516),
    .X(net5515));
 sg13g2_buf_8 fanout5516 (.A(net5523),
    .X(net5516));
 sg13g2_buf_8 fanout5517 (.A(net5519),
    .X(net5517));
 sg13g2_buf_8 fanout5518 (.A(net5519),
    .X(net5518));
 sg13g2_buf_8 fanout5519 (.A(net5522),
    .X(net5519));
 sg13g2_buf_8 fanout5520 (.A(net5521),
    .X(net5520));
 sg13g2_buf_8 fanout5521 (.A(net5522),
    .X(net5521));
 sg13g2_buf_8 fanout5522 (.A(net5523),
    .X(net5522));
 sg13g2_buf_8 fanout5523 (.A(_00001_),
    .X(net5523));
 sg13g2_buf_8 fanout5524 (.A(net5527),
    .X(net5524));
 sg13g2_buf_8 fanout5525 (.A(net5526),
    .X(net5525));
 sg13g2_buf_8 fanout5526 (.A(net5527),
    .X(net5526));
 sg13g2_buf_8 fanout5527 (.A(net5533),
    .X(net5527));
 sg13g2_buf_8 fanout5528 (.A(net5530),
    .X(net5528));
 sg13g2_buf_8 fanout5529 (.A(net5530),
    .X(net5529));
 sg13g2_buf_8 fanout5530 (.A(net5533),
    .X(net5530));
 sg13g2_buf_8 fanout5531 (.A(net5533),
    .X(net5531));
 sg13g2_buf_8 fanout5532 (.A(net5533),
    .X(net5532));
 sg13g2_buf_8 fanout5533 (.A(net5568),
    .X(net5533));
 sg13g2_buf_8 fanout5534 (.A(net5535),
    .X(net5534));
 sg13g2_buf_8 fanout5535 (.A(net5538),
    .X(net5535));
 sg13g2_buf_8 fanout5536 (.A(net5538),
    .X(net5536));
 sg13g2_buf_8 fanout5537 (.A(net5538),
    .X(net5537));
 sg13g2_buf_8 fanout5538 (.A(net5568),
    .X(net5538));
 sg13g2_buf_8 fanout5539 (.A(net5541),
    .X(net5539));
 sg13g2_buf_8 fanout5540 (.A(net5544),
    .X(net5540));
 sg13g2_buf_8 fanout5541 (.A(net5544),
    .X(net5541));
 sg13g2_buf_8 fanout5542 (.A(net5544),
    .X(net5542));
 sg13g2_buf_8 fanout5543 (.A(net5544),
    .X(net5543));
 sg13g2_buf_8 fanout5544 (.A(net5568),
    .X(net5544));
 sg13g2_buf_8 fanout5545 (.A(net5556),
    .X(net5545));
 sg13g2_buf_8 fanout5546 (.A(net5556),
    .X(net5546));
 sg13g2_buf_8 fanout5547 (.A(net5549),
    .X(net5547));
 sg13g2_buf_8 fanout5548 (.A(net5549),
    .X(net5548));
 sg13g2_buf_8 fanout5549 (.A(net5556),
    .X(net5549));
 sg13g2_buf_8 fanout5550 (.A(net5555),
    .X(net5550));
 sg13g2_buf_8 fanout5551 (.A(net5555),
    .X(net5551));
 sg13g2_buf_8 fanout5552 (.A(net5554),
    .X(net5552));
 sg13g2_buf_8 fanout5553 (.A(net5555),
    .X(net5553));
 sg13g2_buf_8 fanout5554 (.A(net5555),
    .X(net5554));
 sg13g2_buf_8 fanout5555 (.A(net5556),
    .X(net5555));
 sg13g2_buf_8 fanout5556 (.A(net5568),
    .X(net5556));
 sg13g2_buf_8 fanout5557 (.A(net5561),
    .X(net5557));
 sg13g2_buf_8 fanout5558 (.A(net5561),
    .X(net5558));
 sg13g2_buf_8 fanout5559 (.A(net5560),
    .X(net5559));
 sg13g2_buf_8 fanout5560 (.A(net5561),
    .X(net5560));
 sg13g2_buf_8 fanout5561 (.A(net5568),
    .X(net5561));
 sg13g2_buf_8 fanout5562 (.A(net5564),
    .X(net5562));
 sg13g2_buf_8 fanout5563 (.A(net5564),
    .X(net5563));
 sg13g2_buf_8 fanout5564 (.A(net5567),
    .X(net5564));
 sg13g2_buf_8 fanout5565 (.A(net5566),
    .X(net5565));
 sg13g2_buf_8 fanout5566 (.A(net5567),
    .X(net5566));
 sg13g2_buf_8 fanout5567 (.A(net5568),
    .X(net5567));
 sg13g2_buf_8 fanout5568 (.A(_00000_),
    .X(net5568));
 sg13g2_buf_8 fanout5569 (.A(net6438),
    .X(net5569));
 sg13g2_buf_8 fanout5570 (.A(net6568),
    .X(net5570));
 sg13g2_buf_8 fanout5571 (.A(net6555),
    .X(net5571));
 sg13g2_buf_8 fanout5572 (.A(net5573),
    .X(net5572));
 sg13g2_buf_8 fanout5573 (.A(net6340),
    .X(net5573));
 sg13g2_buf_8 fanout5574 (.A(net5575),
    .X(net5574));
 sg13g2_buf_2 fanout5575 (.A(net5576),
    .X(net5575));
 sg13g2_buf_8 fanout5576 (.A(net5577),
    .X(net5576));
 sg13g2_buf_8 fanout5577 (.A(net6456),
    .X(net5577));
 sg13g2_buf_8 fanout5578 (.A(net5579),
    .X(net5578));
 sg13g2_buf_8 fanout5579 (.A(net5580),
    .X(net5579));
 sg13g2_buf_8 fanout5580 (.A(\fpga_top.cpu_top.alu_code[2] ),
    .X(net5580));
 sg13g2_buf_8 fanout5581 (.A(net6463),
    .X(net5581));
 sg13g2_buf_8 fanout5582 (.A(\fpga_top.cpu_top.alu_code[1] ),
    .X(net5582));
 sg13g2_buf_8 fanout5583 (.A(net5584),
    .X(net5583));
 sg13g2_buf_8 fanout5584 (.A(net6331),
    .X(net5584));
 sg13g2_buf_8 fanout5585 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[2] ),
    .X(net5585));
 sg13g2_buf_1 fanout5586 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[2] ),
    .X(net5586));
 sg13g2_buf_8 fanout5587 (.A(net5589),
    .X(net5587));
 sg13g2_buf_2 fanout5588 (.A(net5589),
    .X(net5588));
 sg13g2_buf_8 fanout5589 (.A(net6475),
    .X(net5589));
 sg13g2_buf_8 fanout5590 (.A(net6559),
    .X(net5590));
 sg13g2_buf_8 fanout5591 (.A(\fpga_top.bus_gather.i_read_adr[22] ),
    .X(net5591));
 sg13g2_buf_1 fanout5592 (.A(net6583),
    .X(net5592));
 sg13g2_buf_8 fanout5593 (.A(\fpga_top.bus_gather.i_read_adr[16] ),
    .X(net5593));
 sg13g2_buf_1 fanout5594 (.A(net6552),
    .X(net5594));
 sg13g2_buf_8 fanout5595 (.A(\fpga_top.bus_gather.i_read_adr[8] ),
    .X(net5595));
 sg13g2_buf_8 fanout5596 (.A(net6540),
    .X(net5596));
 sg13g2_buf_8 fanout5597 (.A(net6498),
    .X(net5597));
 sg13g2_buf_1 fanout5598 (.A(\fpga_top.bus_gather.i_read_adr[4] ),
    .X(net5598));
 sg13g2_buf_8 fanout5599 (.A(net5601),
    .X(net5599));
 sg13g2_buf_1 fanout5600 (.A(net5601),
    .X(net5600));
 sg13g2_buf_8 fanout5601 (.A(net5602),
    .X(net5601));
 sg13g2_buf_8 fanout5602 (.A(net5603),
    .X(net5602));
 sg13g2_buf_8 fanout5603 (.A(net5604),
    .X(net5603));
 sg13g2_buf_8 fanout5604 (.A(net3940),
    .X(net5604));
 sg13g2_buf_8 fanout5605 (.A(net3168),
    .X(net5605));
 sg13g2_buf_8 fanout5606 (.A(net3488),
    .X(net5606));
 sg13g2_buf_8 fanout5607 (.A(net3659),
    .X(net5607));
 sg13g2_buf_8 fanout5608 (.A(\fpga_top.uart_top.uart_if.byte_data[4] ),
    .X(net5608));
 sg13g2_buf_8 fanout5609 (.A(net6408),
    .X(net5609));
 sg13g2_buf_8 fanout5610 (.A(net6521),
    .X(net5610));
 sg13g2_buf_8 fanout5611 (.A(net6404),
    .X(net5611));
 sg13g2_buf_8 fanout5612 (.A(net6419),
    .X(net5612));
 sg13g2_buf_8 fanout5613 (.A(net6554),
    .X(net5613));
 sg13g2_buf_8 fanout5614 (.A(net6527),
    .X(net5614));
 sg13g2_buf_8 fanout5615 (.A(net3851),
    .X(net5615));
 sg13g2_buf_8 fanout5616 (.A(net6396),
    .X(net5616));
 sg13g2_buf_8 fanout5617 (.A(net5621),
    .X(net5617));
 sg13g2_buf_8 fanout5618 (.A(net5619),
    .X(net5618));
 sg13g2_buf_1 fanout5619 (.A(net5620),
    .X(net5619));
 sg13g2_buf_1 fanout5620 (.A(net5621),
    .X(net5620));
 sg13g2_buf_2 fanout5621 (.A(net5623),
    .X(net5621));
 sg13g2_buf_8 fanout5622 (.A(net5623),
    .X(net5622));
 sg13g2_buf_8 fanout5623 (.A(net5624),
    .X(net5623));
 sg13g2_buf_8 fanout5624 (.A(net6378),
    .X(net5624));
 sg13g2_buf_2 fanout5625 (.A(net5626),
    .X(net5625));
 sg13g2_buf_8 fanout5626 (.A(\fpga_top.uart_top.uart_rec_char.pdata[3] ),
    .X(net5626));
 sg13g2_buf_2 fanout5627 (.A(net2232),
    .X(net5627));
 sg13g2_buf_8 fanout5628 (.A(\fpga_top.uart_top.uart_rec_char.pdata[1] ),
    .X(net5628));
 sg13g2_buf_8 fanout5629 (.A(net6338),
    .X(net5629));
 sg13g2_buf_8 fanout5630 (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[1] ),
    .X(net5630));
 sg13g2_buf_1 fanout5631 (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[1] ),
    .X(net5631));
 sg13g2_buf_8 fanout5632 (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[0] ),
    .X(net5632));
 sg13g2_buf_8 fanout5633 (.A(net5634),
    .X(net5633));
 sg13g2_buf_8 fanout5634 (.A(net6525),
    .X(net5634));
 sg13g2_buf_8 fanout5635 (.A(net2558),
    .X(net5635));
 sg13g2_buf_1 fanout5636 (.A(\fpga_top.cpu_start_adr[30] ),
    .X(net5636));
 sg13g2_buf_8 fanout5637 (.A(net3635),
    .X(net5637));
 sg13g2_buf_8 fanout5638 (.A(net2054),
    .X(net5638));
 sg13g2_buf_2 fanout5639 (.A(\fpga_top.cpu_start_adr[28] ),
    .X(net5639));
 sg13g2_buf_8 fanout5640 (.A(net3920),
    .X(net5640));
 sg13g2_buf_8 fanout5641 (.A(net3920),
    .X(net5641));
 sg13g2_buf_8 fanout5642 (.A(\fpga_top.cpu_start_adr[23] ),
    .X(net5642));
 sg13g2_buf_8 fanout5643 (.A(\fpga_top.cpu_start_adr[22] ),
    .X(net5643));
 sg13g2_buf_8 fanout5644 (.A(net3952),
    .X(net5644));
 sg13g2_buf_8 fanout5645 (.A(net3952),
    .X(net5645));
 sg13g2_buf_8 fanout5646 (.A(\fpga_top.cpu_start_adr[20] ),
    .X(net5646));
 sg13g2_buf_8 fanout5647 (.A(\fpga_top.cpu_start_adr[18] ),
    .X(net5647));
 sg13g2_buf_8 fanout5648 (.A(\fpga_top.cpu_start_adr[17] ),
    .X(net5648));
 sg13g2_buf_8 fanout5649 (.A(\fpga_top.cpu_start_adr[16] ),
    .X(net5649));
 sg13g2_buf_8 fanout5650 (.A(\fpga_top.cpu_start_adr[14] ),
    .X(net5650));
 sg13g2_buf_8 fanout5651 (.A(net2190),
    .X(net5651));
 sg13g2_buf_8 fanout5652 (.A(\fpga_top.cpu_start_adr[10] ),
    .X(net5652));
 sg13g2_buf_8 fanout5653 (.A(net6432),
    .X(net5653));
 sg13g2_buf_8 fanout5654 (.A(net3778),
    .X(net5654));
 sg13g2_buf_8 fanout5655 (.A(\fpga_top.cpu_start_adr[8] ),
    .X(net5655));
 sg13g2_buf_8 fanout5656 (.A(net3719),
    .X(net5656));
 sg13g2_buf_2 fanout5657 (.A(net3719),
    .X(net5657));
 sg13g2_buf_8 fanout5658 (.A(net6098),
    .X(net5658));
 sg13g2_buf_8 fanout5659 (.A(net6098),
    .X(net5659));
 sg13g2_buf_8 fanout5660 (.A(\fpga_top.cpu_start_adr[4] ),
    .X(net5660));
 sg13g2_buf_8 fanout5661 (.A(\fpga_top.cpu_start_adr[4] ),
    .X(net5661));
 sg13g2_buf_8 fanout5662 (.A(net6472),
    .X(net5662));
 sg13g2_buf_8 fanout5663 (.A(\fpga_top.cpu_start_adr[3] ),
    .X(net5663));
 sg13g2_buf_8 fanout5664 (.A(net6582),
    .X(net5664));
 sg13g2_buf_8 fanout5665 (.A(net6575),
    .X(net5665));
 sg13g2_buf_8 fanout5666 (.A(\fpga_top.io_uart_out.rout_en ),
    .X(net5666));
 sg13g2_buf_2 fanout5667 (.A(net6388),
    .X(net5667));
 sg13g2_buf_8 fanout5668 (.A(net6324),
    .X(net5668));
 sg13g2_buf_8 fanout5669 (.A(net5670),
    .X(net5669));
 sg13g2_buf_8 fanout5670 (.A(\fpga_top.uart_top.uart_if.rx_fifo.radr[2] ),
    .X(net5670));
 sg13g2_buf_8 fanout5671 (.A(net5674),
    .X(net5671));
 sg13g2_buf_1 fanout5672 (.A(net5674),
    .X(net5672));
 sg13g2_buf_8 fanout5673 (.A(net5674),
    .X(net5673));
 sg13g2_buf_8 fanout5674 (.A(\fpga_top.uart_top.uart_if.rx_fifo.radr[1] ),
    .X(net5674));
 sg13g2_buf_8 fanout5675 (.A(net5676),
    .X(net5675));
 sg13g2_buf_8 fanout5676 (.A(net5679),
    .X(net5676));
 sg13g2_buf_8 fanout5677 (.A(net5678),
    .X(net5677));
 sg13g2_buf_8 fanout5678 (.A(net5679),
    .X(net5678));
 sg13g2_buf_8 fanout5679 (.A(\fpga_top.uart_top.uart_if.rx_fifo.radr[0] ),
    .X(net5679));
 sg13g2_buf_8 fanout5680 (.A(net6466),
    .X(net5680));
 sg13g2_buf_8 fanout5681 (.A(net6464),
    .X(net5681));
 sg13g2_buf_8 fanout5682 (.A(net6545),
    .X(net5682));
 sg13g2_buf_8 fanout5683 (.A(net6361),
    .X(net5683));
 sg13g2_buf_8 fanout5684 (.A(\fpga_top.qspi_if.rdwrch[5] ),
    .X(net5684));
 sg13g2_buf_1 fanout5685 (.A(\fpga_top.qspi_if.rdwrch[5] ),
    .X(net5685));
 sg13g2_buf_8 fanout5686 (.A(net5688),
    .X(net5686));
 sg13g2_buf_8 fanout5687 (.A(net5688),
    .X(net5687));
 sg13g2_buf_2 fanout5688 (.A(net6385),
    .X(net5688));
 sg13g2_buf_8 fanout5689 (.A(net5690),
    .X(net5689));
 sg13g2_buf_8 fanout5690 (.A(\fpga_top.qspi_if.re_qspi_latency_dly[8] ),
    .X(net5690));
 sg13g2_buf_8 fanout5691 (.A(\fpga_top.qspi_if.re_qspi_latency_dly[6] ),
    .X(net5691));
 sg13g2_buf_8 fanout5692 (.A(\fpga_top.qspi_if.re_qspi_latency_dly[4] ),
    .X(net5692));
 sg13g2_buf_8 fanout5693 (.A(\fpga_top.qspi_if.re_qspi_latency_dly[4] ),
    .X(net5693));
 sg13g2_buf_8 fanout5694 (.A(net5695),
    .X(net5694));
 sg13g2_buf_8 fanout5695 (.A(net5697),
    .X(net5695));
 sg13g2_buf_8 fanout5696 (.A(net5697),
    .X(net5696));
 sg13g2_buf_8 fanout5697 (.A(\fpga_top.qspi_if.re_qspi_latency_dly[3] ),
    .X(net5697));
 sg13g2_buf_8 fanout5698 (.A(\fpga_top.qspi_if.re_qspi_latency_dly[2] ),
    .X(net5698));
 sg13g2_buf_8 fanout5699 (.A(net5709),
    .X(net5699));
 sg13g2_buf_8 fanout5700 (.A(net5701),
    .X(net5700));
 sg13g2_buf_8 fanout5701 (.A(net5709),
    .X(net5701));
 sg13g2_buf_8 fanout5702 (.A(net5708),
    .X(net5702));
 sg13g2_buf_2 fanout5703 (.A(net5704),
    .X(net5703));
 sg13g2_buf_1 fanout5704 (.A(net5705),
    .X(net5704));
 sg13g2_buf_1 fanout5705 (.A(net5706),
    .X(net5705));
 sg13g2_buf_1 fanout5706 (.A(net5707),
    .X(net5706));
 sg13g2_buf_8 fanout5707 (.A(net5708),
    .X(net5707));
 sg13g2_buf_2 fanout5708 (.A(net5709),
    .X(net5708));
 sg13g2_buf_8 fanout5709 (.A(\fpga_top.qspi_if.word_w ),
    .X(net5709));
 sg13g2_buf_8 fanout5710 (.A(\fpga_top.io_led.re_gpio_value_dly[0] ),
    .X(net5710));
 sg13g2_buf_8 fanout5711 (.A(net5712),
    .X(net5711));
 sg13g2_buf_1 fanout5712 (.A(net5713),
    .X(net5712));
 sg13g2_buf_1 fanout5713 (.A(\fpga_top.io_uart_out.uart_io_we ),
    .X(net5713));
 sg13g2_buf_8 fanout5714 (.A(net5716),
    .X(net5714));
 sg13g2_buf_2 fanout5715 (.A(net5716),
    .X(net5715));
 sg13g2_buf_8 fanout5716 (.A(\fpga_top.io_uart_out.re_uart_rdflg_dly[2] ),
    .X(net5716));
 sg13g2_buf_8 fanout5717 (.A(\fpga_top.io_uart_out.re_uart_rdflg_dly[0] ),
    .X(net5717));
 sg13g2_buf_8 fanout5718 (.A(net5719),
    .X(net5718));
 sg13g2_buf_8 fanout5719 (.A(net5721),
    .X(net5719));
 sg13g2_buf_8 fanout5720 (.A(net5721),
    .X(net5720));
 sg13g2_buf_8 fanout5721 (.A(\fpga_top.io_frc.re_frc_dly[3] ),
    .X(net5721));
 sg13g2_buf_8 fanout5722 (.A(net5724),
    .X(net5722));
 sg13g2_buf_1 fanout5723 (.A(net5724),
    .X(net5723));
 sg13g2_buf_8 fanout5724 (.A(net5731),
    .X(net5724));
 sg13g2_buf_2 fanout5725 (.A(net5730),
    .X(net5725));
 sg13g2_buf_1 fanout5726 (.A(net5730),
    .X(net5726));
 sg13g2_buf_8 fanout5727 (.A(net5729),
    .X(net5727));
 sg13g2_buf_1 fanout5728 (.A(net5729),
    .X(net5728));
 sg13g2_buf_8 fanout5729 (.A(net5730),
    .X(net5729));
 sg13g2_buf_8 fanout5730 (.A(net5731),
    .X(net5730));
 sg13g2_buf_8 fanout5731 (.A(\fpga_top.io_frc.re_frc_dly[2] ),
    .X(net5731));
 sg13g2_buf_2 fanout5732 (.A(net5733),
    .X(net5732));
 sg13g2_buf_2 fanout5733 (.A(net5734),
    .X(net5733));
 sg13g2_buf_2 fanout5734 (.A(\fpga_top.io_frc.re_frc_dly[1] ),
    .X(net5734));
 sg13g2_buf_2 fanout5735 (.A(net5736),
    .X(net5735));
 sg13g2_buf_1 fanout5736 (.A(net5737),
    .X(net5736));
 sg13g2_buf_2 fanout5737 (.A(net5742),
    .X(net5737));
 sg13g2_buf_8 fanout5738 (.A(net5740),
    .X(net5738));
 sg13g2_buf_1 fanout5739 (.A(net5740),
    .X(net5739));
 sg13g2_buf_8 fanout5740 (.A(net5741),
    .X(net5740));
 sg13g2_buf_2 fanout5741 (.A(net5742),
    .X(net5741));
 sg13g2_buf_2 fanout5742 (.A(\fpga_top.io_frc.re_frc_dly[1] ),
    .X(net5742));
 sg13g2_buf_2 fanout5743 (.A(net5744),
    .X(net5743));
 sg13g2_buf_1 fanout5744 (.A(net5745),
    .X(net5744));
 sg13g2_buf_8 fanout5745 (.A(net5753),
    .X(net5745));
 sg13g2_buf_8 fanout5746 (.A(net5747),
    .X(net5746));
 sg13g2_buf_2 fanout5747 (.A(net5748),
    .X(net5747));
 sg13g2_buf_1 fanout5748 (.A(net5753),
    .X(net5748));
 sg13g2_buf_2 fanout5749 (.A(net5750),
    .X(net5749));
 sg13g2_buf_8 fanout5750 (.A(net5751),
    .X(net5750));
 sg13g2_buf_1 fanout5751 (.A(net5752),
    .X(net5751));
 sg13g2_buf_1 fanout5752 (.A(net5753),
    .X(net5752));
 sg13g2_buf_8 fanout5753 (.A(\fpga_top.io_frc.re_frc_dly[0] ),
    .X(net5753));
 sg13g2_buf_8 fanout5754 (.A(net5755),
    .X(net5754));
 sg13g2_buf_8 fanout5755 (.A(net6389),
    .X(net5755));
 sg13g2_buf_8 fanout5756 (.A(net6495),
    .X(net5756));
 sg13g2_buf_8 fanout5757 (.A(net5758),
    .X(net5757));
 sg13g2_buf_8 fanout5758 (.A(net5759),
    .X(net5758));
 sg13g2_buf_8 fanout5759 (.A(net6377),
    .X(net5759));
 sg13g2_buf_8 fanout5760 (.A(net6478),
    .X(net5760));
 sg13g2_buf_8 fanout5761 (.A(net5763),
    .X(net5761));
 sg13g2_buf_1 fanout5762 (.A(net5763),
    .X(net5762));
 sg13g2_buf_8 fanout5763 (.A(net6382),
    .X(net5763));
 sg13g2_buf_8 fanout5764 (.A(net5765),
    .X(net5764));
 sg13g2_buf_8 fanout5765 (.A(net6452),
    .X(net5765));
 sg13g2_buf_8 fanout5766 (.A(net5767),
    .X(net5766));
 sg13g2_buf_2 fanout5767 (.A(net5768),
    .X(net5767));
 sg13g2_buf_8 fanout5768 (.A(net6334),
    .X(net5768));
 sg13g2_buf_8 fanout5769 (.A(net5770),
    .X(net5769));
 sg13g2_buf_8 fanout5770 (.A(net6585),
    .X(net5770));
 sg13g2_buf_8 fanout5771 (.A(net5773),
    .X(net5771));
 sg13g2_buf_1 fanout5772 (.A(net5773),
    .X(net5772));
 sg13g2_buf_2 fanout5773 (.A(net6567),
    .X(net5773));
 sg13g2_buf_8 fanout5774 (.A(net6477),
    .X(net5774));
 sg13g2_buf_8 fanout5775 (.A(net5776),
    .X(net5775));
 sg13g2_buf_8 fanout5776 (.A(net6381),
    .X(net5776));
 sg13g2_buf_8 fanout5777 (.A(net6532),
    .X(net5777));
 sg13g2_buf_8 fanout5778 (.A(net5779),
    .X(net5778));
 sg13g2_buf_8 fanout5779 (.A(net5780),
    .X(net5779));
 sg13g2_buf_8 fanout5780 (.A(net6333),
    .X(net5780));
 sg13g2_buf_8 fanout5781 (.A(net5782),
    .X(net5781));
 sg13g2_buf_8 fanout5782 (.A(net6523),
    .X(net5782));
 sg13g2_buf_8 fanout5783 (.A(net5784),
    .X(net5783));
 sg13g2_buf_8 fanout5784 (.A(net5785),
    .X(net5784));
 sg13g2_buf_8 fanout5785 (.A(net6383),
    .X(net5785));
 sg13g2_buf_8 fanout5786 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[16] ),
    .X(net5786));
 sg13g2_buf_8 fanout5787 (.A(net5788),
    .X(net5787));
 sg13g2_buf_8 fanout5788 (.A(net5789),
    .X(net5788));
 sg13g2_buf_8 fanout5789 (.A(net6368),
    .X(net5789));
 sg13g2_buf_8 fanout5790 (.A(net6511),
    .X(net5790));
 sg13g2_buf_8 fanout5791 (.A(net5792),
    .X(net5791));
 sg13g2_buf_8 fanout5792 (.A(net5793),
    .X(net5792));
 sg13g2_buf_1 fanout5793 (.A(net6444),
    .X(net5793));
 sg13g2_buf_8 fanout5794 (.A(net5795),
    .X(net5794));
 sg13g2_buf_8 fanout5795 (.A(net5796),
    .X(net5795));
 sg13g2_buf_1 fanout5796 (.A(net6462),
    .X(net5796));
 sg13g2_buf_8 fanout5797 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[11] ),
    .X(net5797));
 sg13g2_buf_8 fanout5798 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[10] ),
    .X(net5798));
 sg13g2_buf_1 fanout5799 (.A(net6531),
    .X(net5799));
 sg13g2_buf_8 fanout5800 (.A(net5801),
    .X(net5800));
 sg13g2_buf_8 fanout5801 (.A(net5802),
    .X(net5801));
 sg13g2_buf_8 fanout5802 (.A(net6384),
    .X(net5802));
 sg13g2_buf_8 fanout5803 (.A(net5804),
    .X(net5803));
 sg13g2_buf_8 fanout5804 (.A(net6372),
    .X(net5804));
 sg13g2_buf_8 fanout5805 (.A(net5806),
    .X(net5805));
 sg13g2_buf_8 fanout5806 (.A(net6563),
    .X(net5806));
 sg13g2_buf_8 fanout5807 (.A(net5809),
    .X(net5807));
 sg13g2_buf_8 fanout5808 (.A(net5809),
    .X(net5808));
 sg13g2_buf_8 fanout5809 (.A(net6399),
    .X(net5809));
 sg13g2_buf_8 fanout5810 (.A(net5812),
    .X(net5810));
 sg13g2_buf_1 fanout5811 (.A(net5812),
    .X(net5811));
 sg13g2_buf_8 fanout5812 (.A(net6395),
    .X(net5812));
 sg13g2_buf_8 fanout5813 (.A(net5814),
    .X(net5813));
 sg13g2_buf_8 fanout5814 (.A(net5815),
    .X(net5814));
 sg13g2_buf_8 fanout5815 (.A(net6356),
    .X(net5815));
 sg13g2_buf_8 fanout5816 (.A(net5817),
    .X(net5816));
 sg13g2_buf_8 fanout5817 (.A(net5818),
    .X(net5817));
 sg13g2_buf_8 fanout5818 (.A(net6362),
    .X(net5818));
 sg13g2_buf_8 fanout5819 (.A(net5821),
    .X(net5819));
 sg13g2_buf_2 fanout5820 (.A(net5821),
    .X(net5820));
 sg13g2_buf_8 fanout5821 (.A(net6561),
    .X(net5821));
 sg13g2_buf_8 fanout5822 (.A(net5823),
    .X(net5822));
 sg13g2_buf_1 fanout5823 (.A(net5824),
    .X(net5823));
 sg13g2_buf_8 fanout5824 (.A(net6344),
    .X(net5824));
 sg13g2_buf_8 fanout5825 (.A(net6512),
    .X(net5825));
 sg13g2_buf_8 fanout5826 (.A(net6484),
    .X(net5826));
 sg13g2_buf_8 fanout5827 (.A(net5829),
    .X(net5827));
 sg13g2_buf_1 fanout5828 (.A(net5829),
    .X(net5828));
 sg13g2_buf_8 fanout5829 (.A(net5830),
    .X(net5829));
 sg13g2_buf_8 fanout5830 (.A(net6417),
    .X(net5830));
 sg13g2_buf_8 fanout5831 (.A(net5833),
    .X(net5831));
 sg13g2_buf_8 fanout5832 (.A(net5833),
    .X(net5832));
 sg13g2_buf_8 fanout5833 (.A(\fpga_top.io_spi_lite.miso_fifo.rnext ),
    .X(net5833));
 sg13g2_buf_8 fanout5834 (.A(\fpga_top.io_spi_lite.re_spi_value_dly[1] ),
    .X(net5834));
 sg13g2_buf_2 fanout5835 (.A(\fpga_top.io_spi_lite.re_spi_value_dly[1] ),
    .X(net5835));
 sg13g2_buf_8 fanout5836 (.A(net5837),
    .X(net5836));
 sg13g2_buf_8 fanout5837 (.A(\fpga_top.io_spi_lite.re_spi_value_dly[0] ),
    .X(net5837));
 sg13g2_buf_8 fanout5838 (.A(\fpga_top.io_spi_lite.re_spi_value_dly[0] ),
    .X(net5838));
 sg13g2_buf_8 fanout5839 (.A(net5858),
    .X(net5839));
 sg13g2_buf_8 fanout5840 (.A(net5842),
    .X(net5840));
 sg13g2_buf_8 fanout5841 (.A(net5842),
    .X(net5841));
 sg13g2_buf_8 fanout5842 (.A(net5843),
    .X(net5842));
 sg13g2_buf_8 fanout5843 (.A(net5857),
    .X(net5843));
 sg13g2_buf_8 fanout5844 (.A(net5845),
    .X(net5844));
 sg13g2_buf_8 fanout5845 (.A(net5846),
    .X(net5845));
 sg13g2_buf_8 fanout5846 (.A(net5857),
    .X(net5846));
 sg13g2_buf_8 fanout5847 (.A(net5850),
    .X(net5847));
 sg13g2_buf_8 fanout5848 (.A(net5850),
    .X(net5848));
 sg13g2_buf_8 fanout5849 (.A(net5850),
    .X(net5849));
 sg13g2_buf_8 fanout5850 (.A(net5856),
    .X(net5850));
 sg13g2_buf_8 fanout5851 (.A(net5853),
    .X(net5851));
 sg13g2_buf_8 fanout5852 (.A(net5853),
    .X(net5852));
 sg13g2_buf_8 fanout5853 (.A(net5856),
    .X(net5853));
 sg13g2_buf_8 fanout5854 (.A(net5856),
    .X(net5854));
 sg13g2_buf_8 fanout5855 (.A(net5856),
    .X(net5855));
 sg13g2_buf_8 fanout5856 (.A(net5857),
    .X(net5856));
 sg13g2_buf_8 fanout5857 (.A(net5858),
    .X(net5857));
 sg13g2_buf_8 fanout5858 (.A(net5959),
    .X(net5858));
 sg13g2_buf_8 fanout5859 (.A(net5863),
    .X(net5859));
 sg13g2_buf_8 fanout5860 (.A(net5862),
    .X(net5860));
 sg13g2_buf_1 fanout5861 (.A(net5862),
    .X(net5861));
 sg13g2_buf_8 fanout5862 (.A(net5863),
    .X(net5862));
 sg13g2_buf_8 fanout5863 (.A(net5871),
    .X(net5863));
 sg13g2_buf_8 fanout5864 (.A(net5865),
    .X(net5864));
 sg13g2_buf_8 fanout5865 (.A(net5866),
    .X(net5865));
 sg13g2_buf_8 fanout5866 (.A(net5867),
    .X(net5866));
 sg13g2_buf_8 fanout5867 (.A(net5871),
    .X(net5867));
 sg13g2_buf_8 fanout5868 (.A(net5870),
    .X(net5868));
 sg13g2_buf_8 fanout5869 (.A(net5871),
    .X(net5869));
 sg13g2_buf_8 fanout5870 (.A(net5871),
    .X(net5870));
 sg13g2_buf_8 fanout5871 (.A(net5959),
    .X(net5871));
 sg13g2_buf_8 fanout5872 (.A(net5874),
    .X(net5872));
 sg13g2_buf_8 fanout5873 (.A(net5874),
    .X(net5873));
 sg13g2_buf_8 fanout5874 (.A(net5876),
    .X(net5874));
 sg13g2_buf_8 fanout5875 (.A(net5876),
    .X(net5875));
 sg13g2_buf_8 fanout5876 (.A(net5886),
    .X(net5876));
 sg13g2_buf_8 fanout5877 (.A(net5880),
    .X(net5877));
 sg13g2_buf_8 fanout5878 (.A(net5880),
    .X(net5878));
 sg13g2_buf_2 fanout5879 (.A(net5880),
    .X(net5879));
 sg13g2_buf_8 fanout5880 (.A(net5886),
    .X(net5880));
 sg13g2_buf_8 fanout5881 (.A(net5886),
    .X(net5881));
 sg13g2_buf_8 fanout5882 (.A(net5883),
    .X(net5882));
 sg13g2_buf_2 fanout5883 (.A(net5886),
    .X(net5883));
 sg13g2_buf_8 fanout5884 (.A(net5886),
    .X(net5884));
 sg13g2_buf_8 fanout5885 (.A(net5886),
    .X(net5885));
 sg13g2_buf_8 fanout5886 (.A(net5959),
    .X(net5886));
 sg13g2_buf_8 fanout5887 (.A(net5891),
    .X(net5887));
 sg13g2_buf_8 fanout5888 (.A(net5890),
    .X(net5888));
 sg13g2_buf_8 fanout5889 (.A(net5890),
    .X(net5889));
 sg13g2_buf_8 fanout5890 (.A(net5891),
    .X(net5890));
 sg13g2_buf_8 fanout5891 (.A(net5897),
    .X(net5891));
 sg13g2_buf_8 fanout5892 (.A(net5893),
    .X(net5892));
 sg13g2_buf_8 fanout5893 (.A(net5894),
    .X(net5893));
 sg13g2_buf_8 fanout5894 (.A(net5897),
    .X(net5894));
 sg13g2_buf_8 fanout5895 (.A(net5896),
    .X(net5895));
 sg13g2_buf_8 fanout5896 (.A(net5897),
    .X(net5896));
 sg13g2_buf_8 fanout5897 (.A(net5958),
    .X(net5897));
 sg13g2_buf_8 fanout5898 (.A(net5899),
    .X(net5898));
 sg13g2_buf_8 fanout5899 (.A(net5904),
    .X(net5899));
 sg13g2_buf_8 fanout5900 (.A(net5901),
    .X(net5900));
 sg13g2_buf_8 fanout5901 (.A(net5903),
    .X(net5901));
 sg13g2_buf_8 fanout5902 (.A(net5903),
    .X(net5902));
 sg13g2_buf_8 fanout5903 (.A(net5904),
    .X(net5903));
 sg13g2_buf_8 fanout5904 (.A(net5958),
    .X(net5904));
 sg13g2_buf_8 fanout5905 (.A(net5906),
    .X(net5905));
 sg13g2_buf_8 fanout5906 (.A(net5914),
    .X(net5906));
 sg13g2_buf_8 fanout5907 (.A(net5908),
    .X(net5907));
 sg13g2_buf_8 fanout5908 (.A(net5914),
    .X(net5908));
 sg13g2_buf_8 fanout5909 (.A(net5910),
    .X(net5909));
 sg13g2_buf_8 fanout5910 (.A(net5913),
    .X(net5910));
 sg13g2_buf_8 fanout5911 (.A(net5913),
    .X(net5911));
 sg13g2_buf_8 fanout5912 (.A(net5913),
    .X(net5912));
 sg13g2_buf_8 fanout5913 (.A(net5914),
    .X(net5913));
 sg13g2_buf_8 fanout5914 (.A(net5921),
    .X(net5914));
 sg13g2_buf_8 fanout5915 (.A(net5918),
    .X(net5915));
 sg13g2_buf_8 fanout5916 (.A(net5917),
    .X(net5916));
 sg13g2_buf_8 fanout5917 (.A(net5918),
    .X(net5917));
 sg13g2_buf_8 fanout5918 (.A(net5921),
    .X(net5918));
 sg13g2_buf_8 fanout5919 (.A(net5921),
    .X(net5919));
 sg13g2_buf_8 fanout5920 (.A(net5921),
    .X(net5920));
 sg13g2_buf_8 fanout5921 (.A(net5958),
    .X(net5921));
 sg13g2_buf_8 fanout5922 (.A(net5925),
    .X(net5922));
 sg13g2_buf_2 fanout5923 (.A(net5925),
    .X(net5923));
 sg13g2_buf_8 fanout5924 (.A(net5925),
    .X(net5924));
 sg13g2_buf_8 fanout5925 (.A(net5932),
    .X(net5925));
 sg13g2_buf_8 fanout5926 (.A(net5932),
    .X(net5926));
 sg13g2_buf_8 fanout5927 (.A(net5932),
    .X(net5927));
 sg13g2_buf_8 fanout5928 (.A(net5929),
    .X(net5928));
 sg13g2_buf_8 fanout5929 (.A(net5932),
    .X(net5929));
 sg13g2_buf_8 fanout5930 (.A(net5932),
    .X(net5930));
 sg13g2_buf_8 fanout5931 (.A(net5932),
    .X(net5931));
 sg13g2_buf_8 fanout5932 (.A(net5957),
    .X(net5932));
 sg13g2_buf_8 fanout5933 (.A(net5934),
    .X(net5933));
 sg13g2_buf_8 fanout5934 (.A(net5941),
    .X(net5934));
 sg13g2_buf_8 fanout5935 (.A(net5941),
    .X(net5935));
 sg13g2_buf_8 fanout5936 (.A(net5941),
    .X(net5936));
 sg13g2_buf_8 fanout5937 (.A(net5938),
    .X(net5937));
 sg13g2_buf_8 fanout5938 (.A(net5941),
    .X(net5938));
 sg13g2_buf_8 fanout5939 (.A(net5940),
    .X(net5939));
 sg13g2_buf_8 fanout5940 (.A(net5941),
    .X(net5940));
 sg13g2_buf_8 fanout5941 (.A(net5957),
    .X(net5941));
 sg13g2_buf_8 fanout5942 (.A(net5945),
    .X(net5942));
 sg13g2_buf_8 fanout5943 (.A(net5945),
    .X(net5943));
 sg13g2_buf_8 fanout5944 (.A(net5945),
    .X(net5944));
 sg13g2_buf_8 fanout5945 (.A(net5957),
    .X(net5945));
 sg13g2_buf_8 fanout5946 (.A(net5949),
    .X(net5946));
 sg13g2_buf_8 fanout5947 (.A(net5949),
    .X(net5947));
 sg13g2_buf_8 fanout5948 (.A(net5949),
    .X(net5948));
 sg13g2_buf_8 fanout5949 (.A(net5957),
    .X(net5949));
 sg13g2_buf_8 fanout5950 (.A(net5956),
    .X(net5950));
 sg13g2_buf_2 fanout5951 (.A(net5956),
    .X(net5951));
 sg13g2_buf_8 fanout5952 (.A(net5956),
    .X(net5952));
 sg13g2_buf_8 fanout5953 (.A(net5956),
    .X(net5953));
 sg13g2_buf_8 fanout5954 (.A(net5955),
    .X(net5954));
 sg13g2_buf_8 fanout5955 (.A(net5956),
    .X(net5955));
 sg13g2_buf_8 fanout5956 (.A(net5957),
    .X(net5956));
 sg13g2_buf_8 fanout5957 (.A(net5958),
    .X(net5957));
 sg13g2_buf_8 fanout5958 (.A(net5959),
    .X(net5958));
 sg13g2_buf_8 fanout5959 (.A(net6078),
    .X(net5959));
 sg13g2_buf_8 fanout5960 (.A(net5962),
    .X(net5960));
 sg13g2_buf_8 fanout5961 (.A(net5962),
    .X(net5961));
 sg13g2_buf_8 fanout5962 (.A(net5970),
    .X(net5962));
 sg13g2_buf_8 fanout5963 (.A(net5970),
    .X(net5963));
 sg13g2_buf_8 fanout5964 (.A(net5970),
    .X(net5964));
 sg13g2_buf_8 fanout5965 (.A(net5970),
    .X(net5965));
 sg13g2_buf_2 fanout5966 (.A(net5967),
    .X(net5966));
 sg13g2_buf_8 fanout5967 (.A(net5970),
    .X(net5967));
 sg13g2_buf_8 fanout5968 (.A(net5969),
    .X(net5968));
 sg13g2_buf_2 fanout5969 (.A(net5970),
    .X(net5969));
 sg13g2_buf_8 fanout5970 (.A(net6031),
    .X(net5970));
 sg13g2_buf_8 fanout5971 (.A(net5972),
    .X(net5971));
 sg13g2_buf_8 fanout5972 (.A(net5977),
    .X(net5972));
 sg13g2_buf_8 fanout5973 (.A(net5977),
    .X(net5973));
 sg13g2_buf_8 fanout5974 (.A(net5977),
    .X(net5974));
 sg13g2_buf_8 fanout5975 (.A(net5977),
    .X(net5975));
 sg13g2_buf_8 fanout5976 (.A(net5977),
    .X(net5976));
 sg13g2_buf_8 fanout5977 (.A(net6031),
    .X(net5977));
 sg13g2_buf_8 fanout5978 (.A(net5980),
    .X(net5978));
 sg13g2_buf_2 fanout5979 (.A(net5980),
    .X(net5979));
 sg13g2_buf_8 fanout5980 (.A(net5983),
    .X(net5980));
 sg13g2_buf_8 fanout5981 (.A(net5983),
    .X(net5981));
 sg13g2_buf_8 fanout5982 (.A(net5983),
    .X(net5982));
 sg13g2_buf_8 fanout5983 (.A(net5996),
    .X(net5983));
 sg13g2_buf_8 fanout5984 (.A(net5986),
    .X(net5984));
 sg13g2_buf_8 fanout5985 (.A(net5986),
    .X(net5985));
 sg13g2_buf_8 fanout5986 (.A(net5988),
    .X(net5986));
 sg13g2_buf_8 fanout5987 (.A(net5988),
    .X(net5987));
 sg13g2_buf_8 fanout5988 (.A(net5996),
    .X(net5988));
 sg13g2_buf_8 fanout5989 (.A(net5992),
    .X(net5989));
 sg13g2_buf_1 fanout5990 (.A(net5992),
    .X(net5990));
 sg13g2_buf_8 fanout5991 (.A(net5992),
    .X(net5991));
 sg13g2_buf_8 fanout5992 (.A(net5996),
    .X(net5992));
 sg13g2_buf_8 fanout5993 (.A(net5994),
    .X(net5993));
 sg13g2_buf_8 fanout5994 (.A(net5996),
    .X(net5994));
 sg13g2_buf_8 fanout5995 (.A(net5996),
    .X(net5995));
 sg13g2_buf_8 fanout5996 (.A(net6031),
    .X(net5996));
 sg13g2_buf_8 fanout5997 (.A(net6004),
    .X(net5997));
 sg13g2_buf_1 fanout5998 (.A(net6004),
    .X(net5998));
 sg13g2_buf_8 fanout5999 (.A(net6000),
    .X(net5999));
 sg13g2_buf_8 fanout6000 (.A(net6004),
    .X(net6000));
 sg13g2_buf_8 fanout6001 (.A(net6003),
    .X(net6001));
 sg13g2_buf_8 fanout6002 (.A(net6003),
    .X(net6002));
 sg13g2_buf_8 fanout6003 (.A(net6004),
    .X(net6003));
 sg13g2_buf_8 fanout6004 (.A(net6031),
    .X(net6004));
 sg13g2_buf_8 fanout6005 (.A(net6009),
    .X(net6005));
 sg13g2_buf_8 fanout6006 (.A(net6009),
    .X(net6006));
 sg13g2_buf_8 fanout6007 (.A(net6009),
    .X(net6007));
 sg13g2_buf_8 fanout6008 (.A(net6009),
    .X(net6008));
 sg13g2_buf_8 fanout6009 (.A(net6013),
    .X(net6009));
 sg13g2_buf_8 fanout6010 (.A(net6011),
    .X(net6010));
 sg13g2_buf_8 fanout6011 (.A(net6013),
    .X(net6011));
 sg13g2_buf_8 fanout6012 (.A(net6013),
    .X(net6012));
 sg13g2_buf_8 fanout6013 (.A(net6031),
    .X(net6013));
 sg13g2_buf_8 fanout6014 (.A(net6015),
    .X(net6014));
 sg13g2_buf_8 fanout6015 (.A(net6030),
    .X(net6015));
 sg13g2_buf_8 fanout6016 (.A(net6018),
    .X(net6016));
 sg13g2_buf_8 fanout6017 (.A(net6030),
    .X(net6017));
 sg13g2_buf_8 fanout6018 (.A(net6030),
    .X(net6018));
 sg13g2_buf_8 fanout6019 (.A(net6022),
    .X(net6019));
 sg13g2_buf_8 fanout6020 (.A(net6022),
    .X(net6020));
 sg13g2_buf_2 fanout6021 (.A(net6022),
    .X(net6021));
 sg13g2_buf_8 fanout6022 (.A(net6029),
    .X(net6022));
 sg13g2_buf_8 fanout6023 (.A(net6024),
    .X(net6023));
 sg13g2_buf_8 fanout6024 (.A(net6029),
    .X(net6024));
 sg13g2_buf_8 fanout6025 (.A(net6029),
    .X(net6025));
 sg13g2_buf_8 fanout6026 (.A(net6028),
    .X(net6026));
 sg13g2_buf_8 fanout6027 (.A(net6028),
    .X(net6027));
 sg13g2_buf_8 fanout6028 (.A(net6029),
    .X(net6028));
 sg13g2_buf_8 fanout6029 (.A(net6030),
    .X(net6029));
 sg13g2_buf_8 fanout6030 (.A(net6031),
    .X(net6030));
 sg13g2_buf_8 fanout6031 (.A(net6078),
    .X(net6031));
 sg13g2_buf_8 fanout6032 (.A(net6035),
    .X(net6032));
 sg13g2_buf_8 fanout6033 (.A(net6035),
    .X(net6033));
 sg13g2_buf_8 fanout6034 (.A(net6035),
    .X(net6034));
 sg13g2_buf_8 fanout6035 (.A(net6064),
    .X(net6035));
 sg13g2_buf_8 fanout6036 (.A(net6037),
    .X(net6036));
 sg13g2_buf_8 fanout6037 (.A(net6040),
    .X(net6037));
 sg13g2_buf_8 fanout6038 (.A(net6040),
    .X(net6038));
 sg13g2_buf_8 fanout6039 (.A(net6040),
    .X(net6039));
 sg13g2_buf_8 fanout6040 (.A(net6064),
    .X(net6040));
 sg13g2_buf_8 fanout6041 (.A(net6044),
    .X(net6041));
 sg13g2_buf_8 fanout6042 (.A(net6044),
    .X(net6042));
 sg13g2_buf_8 fanout6043 (.A(net6044),
    .X(net6043));
 sg13g2_buf_8 fanout6044 (.A(net6064),
    .X(net6044));
 sg13g2_buf_8 fanout6045 (.A(net6047),
    .X(net6045));
 sg13g2_buf_1 fanout6046 (.A(net6047),
    .X(net6046));
 sg13g2_buf_8 fanout6047 (.A(net6056),
    .X(net6047));
 sg13g2_buf_8 fanout6048 (.A(net6056),
    .X(net6048));
 sg13g2_buf_8 fanout6049 (.A(net6056),
    .X(net6049));
 sg13g2_buf_8 fanout6050 (.A(net6052),
    .X(net6050));
 sg13g2_buf_8 fanout6051 (.A(net6052),
    .X(net6051));
 sg13g2_buf_8 fanout6052 (.A(net6055),
    .X(net6052));
 sg13g2_buf_8 fanout6053 (.A(net6054),
    .X(net6053));
 sg13g2_buf_8 fanout6054 (.A(net6055),
    .X(net6054));
 sg13g2_buf_8 fanout6055 (.A(net6056),
    .X(net6055));
 sg13g2_buf_8 fanout6056 (.A(net6063),
    .X(net6056));
 sg13g2_buf_8 fanout6057 (.A(net6063),
    .X(net6057));
 sg13g2_buf_1 fanout6058 (.A(net6063),
    .X(net6058));
 sg13g2_buf_8 fanout6059 (.A(net6061),
    .X(net6059));
 sg13g2_buf_8 fanout6060 (.A(net6061),
    .X(net6060));
 sg13g2_buf_8 fanout6061 (.A(net6062),
    .X(net6061));
 sg13g2_buf_8 fanout6062 (.A(net6063),
    .X(net6062));
 sg13g2_buf_8 fanout6063 (.A(net6064),
    .X(net6063));
 sg13g2_buf_8 fanout6064 (.A(net6078),
    .X(net6064));
 sg13g2_buf_8 fanout6065 (.A(net6069),
    .X(net6065));
 sg13g2_buf_8 fanout6066 (.A(net6068),
    .X(net6066));
 sg13g2_buf_8 fanout6067 (.A(net6068),
    .X(net6067));
 sg13g2_buf_8 fanout6068 (.A(net6069),
    .X(net6068));
 sg13g2_buf_8 fanout6069 (.A(net6077),
    .X(net6069));
 sg13g2_buf_8 fanout6070 (.A(net6071),
    .X(net6070));
 sg13g2_buf_8 fanout6071 (.A(net6072),
    .X(net6071));
 sg13g2_buf_8 fanout6072 (.A(net6076),
    .X(net6072));
 sg13g2_buf_8 fanout6073 (.A(net6075),
    .X(net6073));
 sg13g2_buf_8 fanout6074 (.A(net6075),
    .X(net6074));
 sg13g2_buf_8 fanout6075 (.A(net6076),
    .X(net6075));
 sg13g2_buf_8 fanout6076 (.A(net6077),
    .X(net6076));
 sg13g2_buf_8 fanout6077 (.A(net6078),
    .X(net6077));
 sg13g2_buf_8 fanout6078 (.A(rst_n),
    .X(net6078));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_2 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_2 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_2 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tiehi _24582__17 (.L_HI(net17));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_8 clkbuf_leaf_313_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_8 clkbuf_leaf_314_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_314_clk));
 sg13g2_buf_8 clkbuf_leaf_315_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_315_clk));
 sg13g2_buf_8 clkbuf_leaf_316_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_316_clk));
 sg13g2_buf_8 clkbuf_leaf_317_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_317_clk));
 sg13g2_buf_8 clkbuf_leaf_318_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_318_clk));
 sg13g2_buf_8 clkbuf_leaf_319_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_319_clk));
 sg13g2_buf_8 clkbuf_leaf_320_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_320_clk));
 sg13g2_buf_8 clkbuf_leaf_321_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_321_clk));
 sg13g2_buf_8 clkbuf_leaf_322_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_322_clk));
 sg13g2_buf_8 clkbuf_leaf_323_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_323_clk));
 sg13g2_buf_8 clkbuf_leaf_324_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_324_clk));
 sg13g2_buf_8 clkbuf_leaf_325_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_325_clk));
 sg13g2_buf_8 clkbuf_leaf_326_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_326_clk));
 sg13g2_buf_8 clkbuf_leaf_327_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_327_clk));
 sg13g2_buf_8 clkbuf_leaf_328_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_328_clk));
 sg13g2_buf_8 clkbuf_leaf_329_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_329_clk));
 sg13g2_buf_8 clkbuf_leaf_330_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_330_clk));
 sg13g2_buf_8 clkbuf_leaf_331_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_331_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sg13g2_buf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sg13g2_buf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sg13g2_buf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sg13g2_buf_8 clkbuf_5_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0_0_clk));
 sg13g2_buf_8 clkbuf_5_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1_0_clk));
 sg13g2_buf_8 clkbuf_5_2_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2_0_clk));
 sg13g2_buf_8 clkbuf_5_3_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3_0_clk));
 sg13g2_buf_8 clkbuf_5_4_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4_0_clk));
 sg13g2_buf_8 clkbuf_5_5_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5_0_clk));
 sg13g2_buf_8 clkbuf_5_6_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6_0_clk));
 sg13g2_buf_8 clkbuf_5_7_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7_0_clk));
 sg13g2_buf_8 clkbuf_5_8_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8_0_clk));
 sg13g2_buf_8 clkbuf_5_9_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9_0_clk));
 sg13g2_buf_8 clkbuf_5_10_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10_0_clk));
 sg13g2_buf_8 clkbuf_5_11_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11_0_clk));
 sg13g2_buf_8 clkbuf_5_12_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12_0_clk));
 sg13g2_buf_8 clkbuf_5_13_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13_0_clk));
 sg13g2_buf_8 clkbuf_5_14_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14_0_clk));
 sg13g2_buf_8 clkbuf_5_15_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15_0_clk));
 sg13g2_buf_8 clkbuf_5_16_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16_0_clk));
 sg13g2_buf_8 clkbuf_5_17_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17_0_clk));
 sg13g2_buf_8 clkbuf_5_18_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18_0_clk));
 sg13g2_buf_8 clkbuf_5_19_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19_0_clk));
 sg13g2_buf_8 clkbuf_5_20_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20_0_clk));
 sg13g2_buf_8 clkbuf_5_21_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21_0_clk));
 sg13g2_buf_8 clkbuf_5_22_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22_0_clk));
 sg13g2_buf_8 clkbuf_5_23_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23_0_clk));
 sg13g2_buf_8 clkbuf_5_24_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24_0_clk));
 sg13g2_buf_8 clkbuf_5_25_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25_0_clk));
 sg13g2_buf_8 clkbuf_5_26_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26_0_clk));
 sg13g2_buf_8 clkbuf_5_27_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27_0_clk));
 sg13g2_buf_8 clkbuf_5_28_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28_0_clk));
 sg13g2_buf_8 clkbuf_5_29_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29_0_clk));
 sg13g2_buf_8 clkbuf_5_30_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30_0_clk));
 sg13g2_buf_8 clkbuf_5_31_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31_0_clk));
 sg13g2_buf_8 clkbuf_6_0__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_8 clkbuf_6_1__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkbuf_6_2__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_8 clkbuf_6_3__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkbuf_6_4__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_8 clkbuf_6_5__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkbuf_6_6__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_8 clkbuf_6_7__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkbuf_6_8__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_8 clkbuf_6_9__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkbuf_6_10__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_8 clkbuf_6_11__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkbuf_6_12__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_8 clkbuf_6_13__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkbuf_6_14__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_8 clkbuf_6_15__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkbuf_6_16__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_8 clkbuf_6_17__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkbuf_6_18__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_8 clkbuf_6_19__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkbuf_6_20__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_8 clkbuf_6_21__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkbuf_6_22__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_8 clkbuf_6_23__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkbuf_6_24__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_8 clkbuf_6_25__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkbuf_6_26__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_8 clkbuf_6_27__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkbuf_6_28__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_8 clkbuf_6_29__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkbuf_6_30__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_8 clkbuf_6_31__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkbuf_6_32__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_8 clkbuf_6_33__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkbuf_6_34__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_8 clkbuf_6_35__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkbuf_6_36__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_8 clkbuf_6_37__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkbuf_6_38__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_8 clkbuf_6_39__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkbuf_6_40__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_8 clkbuf_6_41__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkbuf_6_42__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_8 clkbuf_6_43__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkbuf_6_44__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_8 clkbuf_6_45__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkbuf_6_46__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_8 clkbuf_6_47__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkbuf_6_48__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_8 clkbuf_6_49__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkbuf_6_50__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_8 clkbuf_6_51__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkbuf_6_52__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_8 clkbuf_6_53__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkbuf_6_54__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_8 clkbuf_6_55__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkbuf_6_56__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_8 clkbuf_6_57__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_8 clkbuf_6_58__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_8 clkbuf_6_59__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkbuf_6_60__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_8 clkbuf_6_61__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_8 clkbuf_6_62__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_8 clkbuf_6_63__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_6_57__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_331_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_125_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_129_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_198_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_leaf_133_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_244_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\fpga_top.qspi_if.sio_in_mt1[0] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold2 (.A(\fpga_top.qspi_if.sio_in_mt0[1] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold3 (.A(\fpga_top.qspi_if.sio_out_dly[0] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold4 (.A(\fpga_top.io_led.gpi_init_lat1[2] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold5 (.A(\fpga_top.qspi_if.sio_in_mt0[2] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold6 (.A(\fpga_top.interrupter.int0_1lat ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold7 (.A(\fpga_top.qspi_if.sio_out_enbl_dly ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold8 (.A(\fpga_top.io_led.gpi_init_lat1[5] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold9 (.A(\fpga_top.qspi_if.sio_in_mt1[1] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold10 (.A(\fpga_top.io_spi_lite.sel_mosi[2] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold11 (.A(\fpga_top.qspi_if.sio_out_dly[1] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold12 (.A(\fpga_top.uart_top.uart_rec_char.g_crlf_dly2 ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold13 (.A(\fpga_top.io_led.gpi_init_lat1[4] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold14 (.A(\fpga_top.qspi_if.sio_in_mt0[0] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold15 (.A(\fpga_top.uart_top.uart_rec_char.g_crlf_dly ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold16 (.A(\fpga_top.io_led.gpio_in_lat1[1] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold17 (.A(\fpga_top.qspi_if.sio_out_dly[3] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold18 (.A(\fpga_top.io_led.gpi_init_lat1[1] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold19 (.A(\fpga_top.io_led.gpio_in_lat1[3] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold20 (.A(\fpga_top.io_led.gpio_in_lat1[0] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold21 (.A(\fpga_top.qspi_if.sio_out_dly[2] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold22 (.A(\fpga_top.io_spi_lite.sel_sck[6] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold23 (.A(\fpga_top.io_led.gpi_init_lat1[3] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold24 (.A(\fpga_top.io_led.gpio_in_lat1[2] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold25 (.A(\fpga_top.qspi_if.sio_in_mt0[3] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold26 (.A(\fpga_top.io_spi_lite.sel_cs[4] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold27 (.A(\fpga_top.io_spi_lite.sel_cs[6] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold28 (.A(\fpga_top.io_spi_lite.sel_mosi[4] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold29 (.A(\fpga_top.io_spi_lite.sel_mosi[6] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold30 (.A(\fpga_top.io_spi_lite.sel_cs[3] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold31 (.A(\fpga_top.io_spi_lite.miso_lat[5] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold32 (.A(\fpga_top.io_led.gpi_init_lat1[0] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold33 (.A(\fpga_top.io_spi_lite.sel_cs[2] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold34 (.A(\fpga_top.io_spi_lite.sel_mosi[1] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold35 (.A(\fpga_top.io_spi_lite.sel_sck[1] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold36 (.A(\fpga_top.io_spi_lite.sel_mosi[5] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold37 (.A(\fpga_top.io_spi_lite.sel_sck[3] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold38 (.A(\fpga_top.io_spi_lite.sel_sck[4] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold39 (.A(\fpga_top.io_spi_lite.sel_cs[1] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold40 (.A(\fpga_top.io_spi_lite.sel_sck[2] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold41 (.A(\fpga_top.io_spi_lite.sel_sck[5] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold42 (.A(\fpga_top.io_spi_lite.miso_lat[6] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold43 (.A(\fpga_top.io_spi_lite.miso_lat[2] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold44 (.A(\fpga_top.io_spi_lite.miso_lat[4] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold45 (.A(\fpga_top.io_spi_lite.sel_cs[5] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold46 (.A(\fpga_top.io_spi_lite.miso_lat[3] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold47 (.A(\fpga_top.qspi_if.sio_in_mt1[2] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold48 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_radr[2] ),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold49 (.A(\fpga_top.io_spi_lite.sel_mosi[3] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold50 (.A(\fpga_top.uart_top.rx_fifo_rcntr[2] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold51 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_radr[1] ),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold52 (.A(\fpga_top.qspi_if.sio_in_mt1[3] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold53 (.A(\fpga_top.uart_top.rx_fifo_rcntr[1] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold54 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_radr[0] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold55 (.A(\fpga_top.io_spi_lite.org_sck ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold56 (.A(\fpga_top.uart_top.rx_fifo_rcntr[0] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold57 (.A(\fpga_top.io_led.gpi_init_lat2[0] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold58 (.A(_00119_),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold59 (.A(\fpga_top.interrupter.int0_2lat ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold60 (.A(_00126_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold61 (.A(\fpga_top.qspi_if.dbg_2div_cew_pre ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold62 (.A(\fpga_top.interrupter.g_interrupt_dly ),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold63 (.A(_01510_),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold64 (.A(\fpga_top.uart_top.uart_logics.write_stat ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold65 (.A(_00084_),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold66 (.A(\fpga_top.cpu_top.inst_mem_read.imr_stat ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold67 (.A(\fpga_top.io_frc.frc_cntr_val_rst_lat ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold68 (.A(_00328_),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold69 (.A(_00116_),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold70 (.A(_00088_),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold71 (.A(\fpga_top.uart_top.uart_if.tx_out_data[1] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold72 (.A(_01131_),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold73 (.A(\fpga_top.io_uart_out.re_uart_rdflg_dly[3] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold74 (.A(_00382_),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold75 (.A(_00120_),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold76 (.A(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[1] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold77 (.A(_08873_),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold78 (.A(\fpga_top.uart_top.uart_if.tx_out_cntr[3] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold79 (.A(_09519_),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold80 (.A(_00117_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold81 (.A(_00118_),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold82 (.A(\fpga_top.uart_top.uart_rec_char.data_cntr[3] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold83 (.A(_01301_),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold84 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][2] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold85 (.A(_02343_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold86 (.A(\fpga_top.qspi_if.qspi_state[7] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold87 (.A(_00145_),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold88 (.A(\fpga_top.qspi_if.word_data[31] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold89 (.A(_00988_),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold90 (.A(\fpga_top.io_spi_lite.sck_div[0] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold91 (.A(\fpga_top.io_uart_out.rx_write_error ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold92 (.A(_03036_),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold93 (.A(\fpga_top.io_spi_lite.miso_bit_cntr[2] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold94 (.A(_10570_),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold95 (.A(_00207_),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold96 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[30] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold97 (.A(\fpga_top.uart_top.uart_if.tx_out_data[7] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold98 (.A(_01138_),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold99 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][4] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold100 (.A(_02345_),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold101 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[7] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold102 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[16] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold103 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[10] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold104 (.A(_01457_),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold105 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][5] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold106 (.A(_06359_),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold107 (.A(_02282_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold108 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][6] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold109 (.A(_02347_),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold110 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[22] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold111 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][0] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold112 (.A(_02309_),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold113 (.A(\fpga_top.io_spi_lite.miso_bit_cntr[1] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold114 (.A(_10568_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold115 (.A(_00206_),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold116 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[26] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold117 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][0] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold118 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[12] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold119 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[7] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold120 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][5] ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold121 (.A(_02346_),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold122 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[17] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold123 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[16] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold124 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[31] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold125 (.A(_01478_),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold126 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[17] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold127 (.A(_01464_),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold128 (.A(\fpga_top.qspi_if.word_data[30] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold129 (.A(_00987_),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold130 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[25] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold131 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sie ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold132 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[15] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold133 (.A(_01462_),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold134 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][7] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold135 (.A(_02284_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold136 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[9] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold137 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[1] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold138 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[31] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold139 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][1] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold140 (.A(_02310_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold141 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[3] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold142 (.A(_01582_),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold143 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[28] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold144 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][7] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold145 (.A(_02316_),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold146 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][6] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold147 (.A(_02283_),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold148 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[17] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold149 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[28] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold150 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[19] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold151 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[9] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold152 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[28] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold153 (.A(\fpga_top.cpu_top.data_rw_mem.unsigned_bit_dly ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold154 (.A(_05341_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold155 (.A(_01901_),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold156 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][5] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold157 (.A(_02314_),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold158 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][2] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold159 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[27] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold160 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[15] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold161 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[6] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold162 (.A(_01453_),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold163 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[9] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold164 (.A(_01456_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold165 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[14] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold166 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][6] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold167 (.A(_02315_),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold168 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[30] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold169 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][3] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold170 (.A(_02344_),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold171 (.A(\fpga_top.qspi_if.sck_cntr[0] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold172 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[5] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold173 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][0] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold174 (.A(_02277_),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold175 (.A(\fpga_top.qspi_if.read_cntr[3] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold176 (.A(_01018_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold177 (.A(\fpga_top.uart_top.uart_if.tx_out_data[3] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold178 (.A(_01134_),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold179 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][7] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold180 (.A(_02348_),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold181 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[13] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold182 (.A(_01460_),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold183 (.A(\fpga_top.qspi_if.word_data[28] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold184 (.A(_00985_),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold185 (.A(_00107_),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold186 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[11] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold187 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[27] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold188 (.A(_02037_),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold189 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[13] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold190 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[3] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold191 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[3] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold192 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[21] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold193 (.A(_01468_),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold194 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[24] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold195 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[11] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold196 (.A(_01458_),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold197 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[3] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold198 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[20] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold199 (.A(_01467_),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold200 (.A(\fpga_top.uart_top.uart_if.tx_out_data[5] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold201 (.A(_01136_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold202 (.A(_00095_),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold203 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[16] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold204 (.A(_02026_),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold205 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[0] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold206 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[5] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold207 (.A(_01452_),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold208 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][2] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold209 (.A(_02311_),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold210 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[18] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold211 (.A(_01465_),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold212 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][1] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold213 (.A(_02342_),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold214 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[5] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold215 (.A(_01584_),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold216 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[2] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold217 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[12] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold218 (.A(_01459_),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold219 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[10] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold220 (.A(\fpga_top.qspi_if.qspi_state[1] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold221 (.A(_00016_),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold222 (.A(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[0] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold223 (.A(_01123_),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold224 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[4] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold225 (.A(_00089_),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold226 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[14] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold227 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[7] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold228 (.A(_01454_),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold229 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[1] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold230 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[18] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold231 (.A(_00087_),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold232 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[24] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold233 (.A(_01471_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold234 (.A(\fpga_top.uart_top.uart_rec_char.data_word[8] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold235 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[14] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold236 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[14] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold237 (.A(_01461_),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold238 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[9] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold239 (.A(_01986_),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold240 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[1] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold241 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[23] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold242 (.A(_01470_),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold243 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][1] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold244 (.A(_06357_),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold245 (.A(_02278_),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold246 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[27] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold247 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[11] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold248 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[5] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold249 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[16] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold250 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[7][0] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold251 (.A(_02341_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold252 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[6] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold253 (.A(_01912_),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold254 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[2] ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold255 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[1] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold256 (.A(_01907_),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold257 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[6] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold258 (.A(\fpga_top.io_spi_lite.mosi_fifo.radr[2] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold259 (.A(\fpga_top.io_spi_lite.mosi_fifo.radr_early[2] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold260 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[3] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold261 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[2] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold262 (.A(\fpga_top.uart_top.uart_if.tx_out_data[6] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold263 (.A(_01137_),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold264 (.A(\fpga_top.uart_top.uart_rec_char.data_word[22] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold265 (.A(_01261_),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold266 (.A(\fpga_top.io_spi_lite.mosi_pp_cntr[2] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00203_),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold268 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[19] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold269 (.A(_01466_),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold270 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[7] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold271 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[9] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold272 (.A(_02019_),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold273 (.A(\fpga_top.io_spi_lite.mosi_fifo.radr[1] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold274 (.A(_08976_),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold275 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[17] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold276 (.A(_02027_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold277 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[27] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold278 (.A(_01474_),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold279 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[20] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold280 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[29] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold281 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[30] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold282 (.A(\fpga_top.uart_top.uart_if.tx_out_data[9] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold283 (.A(\fpga_top.qspi_if.adr_rw[0] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold284 (.A(\fpga_top.uart_top.uart_rec_char.data_word[27] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold285 (.A(_04462_),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold286 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[26] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold287 (.A(_01473_),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold288 (.A(\fpga_top.uart_top.uart_if.rx_state[1] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold289 (.A(\fpga_top.uart_top.uart_if.next_rx_state[3] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold290 (.A(\fpga_top.uart_top.uart_if.tx_out_data[8] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold291 (.A(_01139_),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold292 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[19] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold293 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][1] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold294 (.A(_06451_),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold295 (.A(_02374_),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold296 (.A(\fpga_top.qspi_if.word_data[17] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold297 (.A(_00974_),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold298 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[16] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold299 (.A(_01993_),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold300 (.A(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[0] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold301 (.A(\fpga_top.qspi_if.word_data[29] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold302 (.A(_00986_),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold303 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][0] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold304 (.A(_06477_),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold305 (.A(_02397_),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold306 (.A(_00115_),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold307 (.A(\fpga_top.io_spi_lite.spi_sck_div[7] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold308 (.A(_08950_),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold309 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[7] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold310 (.A(_01147_),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold311 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[23] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold312 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[4] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold313 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][5] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold314 (.A(_02354_),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold315 (.A(\fpga_top.qspi_if.sio_in_sync[2] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold316 (.A(_00959_),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold317 (.A(\fpga_top.uart_top.uart_if.tx_out_data[2] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold318 (.A(_01132_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold319 (.A(\fpga_top.qspi_if.adr_rw[1] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold320 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][7] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold321 (.A(_02396_),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold322 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][3] ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold323 (.A(_06444_),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold324 (.A(_02368_),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold325 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[11] ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold326 (.A(_01590_),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold327 (.A(\fpga_top.uart_top.uart_logics.cmd_read_adr[32] ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold328 (.A(_01431_),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold329 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[6] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold330 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][7] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold331 (.A(_02404_),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold332 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[14] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold333 (.A(\fpga_top.uart_top.uart_rec_char.data_word[15] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold334 (.A(_01254_),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold335 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][5] ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold336 (.A(_02370_),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold337 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[15] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold338 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][7] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold339 (.A(_06389_),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold340 (.A(_02324_),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold341 (.A(\fpga_top.io_spi_lite.miso_bit_cntr[0] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold342 (.A(_00205_),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold343 (.A(\fpga_top.qspi_if.word_data[20] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold344 (.A(_00977_),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold345 (.A(\fpga_top.uart_top.uart_rec_char.data_word[9] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold346 (.A(\fpga_top.qspi_if.word_data[21] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold347 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[13] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold348 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][0] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold349 (.A(_06459_),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold350 (.A(_02381_),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold351 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][4] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold352 (.A(_02353_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold353 (.A(\fpga_top.qspi_if.wdata[9] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold354 (.A(_00932_),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold355 (.A(\fpga_top.qspi_if.word_data[22] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold356 (.A(_00979_),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold357 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][7] ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold358 (.A(_02372_),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold359 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][3] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold360 (.A(_06453_),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold361 (.A(_02376_),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold362 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[30] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold363 (.A(_01477_),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold364 (.A(\fpga_top.uart_top.uart_rec_char.data_word[24] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold365 (.A(_04459_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold366 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[29] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold367 (.A(\fpga_top.io_spi_lite.mosi_pp_cntr[3] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold368 (.A(_00204_),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold369 (.A(\fpga_top.qspi_if.word_data[27] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold370 (.A(_00984_),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold371 (.A(_00122_),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold372 (.A(\fpga_top.io_uart_out.rx_data_latch[0] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold373 (.A(_00383_),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold374 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[30] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold375 (.A(_01366_),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold376 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][5] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold377 (.A(_02394_),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold378 (.A(\fpga_top.uart_top.uart_rec_char.data_word[13] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold379 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][1] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold380 (.A(_03697_),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold381 (.A(_03702_),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold382 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][1] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold383 (.A(_06478_),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold384 (.A(_02398_),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold385 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[3] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold386 (.A(_01450_),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold387 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][6] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold388 (.A(_02387_),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold389 (.A(\fpga_top.io_spi_lite.bit_sel_org[0] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold390 (.A(_00208_),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold391 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mcause[1] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold392 (.A(_01939_),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold393 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[18] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold394 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][3] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold395 (.A(_06462_),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold396 (.A(_02384_),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold397 (.A(\fpga_top.io_uart_out.rx_data_latch[7] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold398 (.A(_00390_),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold399 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][5] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold400 (.A(_02402_),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold401 (.A(\fpga_top.qspi_if.word_data[26] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold402 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[9] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold403 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[26] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold404 (.A(\fpga_top.qspi_if.word_data[13] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold405 (.A(_00970_),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold406 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][1] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold407 (.A(_06460_),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold408 (.A(_02382_),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold409 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][2] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold410 (.A(\fpga_top.uart_top.uart_rec_char.data_word[11] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold411 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][1] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold412 (.A(_06469_),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold413 (.A(_02390_),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold414 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][0] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold415 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][0] ),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold416 (.A(_06450_),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold417 (.A(_02373_),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold418 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][0] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold419 (.A(\fpga_top.qspi_if.rdcmd1[2] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold420 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][6] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold421 (.A(_02371_),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold422 (.A(\fpga_top.uart_top.uart_rec_char.data_word[6] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold423 (.A(\fpga_top.uart_top.uart_rec_char.data_word[16] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold424 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][3] ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold425 (.A(_02192_),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold426 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mcause[5] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold427 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[11] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold428 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[22] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold429 (.A(_01601_),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold430 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][1] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold431 (.A(_06364_),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold432 (.A(_02286_),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold433 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][1] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold434 (.A(_06385_),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold435 (.A(_02318_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold436 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][6] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold437 (.A(_02403_),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold438 (.A(\fpga_top.cpu_top.csr_mepc_ex[3] ),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold439 (.A(_01946_),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold440 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][2] ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold441 (.A(_02351_),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold442 (.A(\fpga_top.io_spi_lite.mosi_pp_cntr[1] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold443 (.A(_00202_),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold444 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][3] ),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold445 (.A(_06480_),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold446 (.A(_02400_),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold447 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][7] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold448 (.A(_02380_),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold449 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][2] ),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold450 (.A(_02399_),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold451 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][2] ),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold452 (.A(_06386_),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold453 (.A(_02319_),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold454 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[23] ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold455 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][5] ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold456 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][4] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold457 (.A(_02361_),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold458 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[8] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold459 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][7] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold460 (.A(_02388_),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold461 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][2] ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold462 (.A(_02383_),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold463 (.A(\fpga_top.io_spi_lite.spi_mode[1] ),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold464 (.A(_09646_),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold465 (.A(\fpga_top.uart_top.uart_rec_char.data_word[14] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold466 (.A(_01253_),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold467 (.A(\fpga_top.interrupter.int_enable_int0 ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold468 (.A(\fpga_top.qspi_if.wdata[6] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold469 (.A(_00929_),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold470 (.A(\fpga_top.qspi_if.word_data[18] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold471 (.A(_00975_),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold472 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[11] ),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold473 (.A(_01151_),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold474 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[31] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold475 (.A(_01937_),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold476 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][6] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold477 (.A(_02379_),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold478 (.A(\fpga_top.cpu_top.csr_mepc_ex[29] ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold479 (.A(_01972_),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold480 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[12] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold481 (.A(_01591_),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold482 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[12] ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold483 (.A(_01152_),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold484 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][5] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold485 (.A(_06387_),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold486 (.A(_02322_),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold487 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[21] ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold488 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[16] ),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold489 (.A(_01352_),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold490 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][2] ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold491 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][7] ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold492 (.A(_02364_),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold493 (.A(\fpga_top.qspi_if.inner_state[0] ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold494 (.A(\fpga_top.qspi_if.inner_machine$func$/home/runner/work/ttihp-26a-risc-v-wg-swc1/ttihp-26a-risc-v-wg-swc1/src/qspi_if.v:768$329.$result[1] ),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold495 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][1] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold496 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[2] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold497 (.A(_01449_),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold498 (.A(\fpga_top.uart_top.uart_rec_char.data_word[18] ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold499 (.A(_01257_),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold500 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][2] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold501 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][6] ),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold502 (.A(_02395_),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold503 (.A(\fpga_top.cpu_top.csr_mepc_ex[15] ),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold504 (.A(_01958_),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold505 (.A(\fpga_top.cpu_top.csr_mepc_ex[11] ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold506 (.A(_01954_),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold507 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][0] ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold508 (.A(_06268_),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold509 (.A(_02165_),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold510 (.A(\fpga_top.uart_top.uart_rec_char.data_word[26] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold511 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][1] ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold512 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[30] ),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold513 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][6] ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold514 (.A(_06388_),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold515 (.A(_02323_),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold516 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][1] ),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold517 (.A(_02174_),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold518 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[20] ),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold519 (.A(_01599_),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold520 (.A(\fpga_top.interrupter.int_enable_rx ),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold521 (.A(\fpga_top.uart_top.uart_rec_char.data_word[20] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold522 (.A(_01259_),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold523 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][0] ),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold524 (.A(\fpga_top.qspi_if.wdata[8] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold525 (.A(_00931_),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold526 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[0][4] ),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold527 (.A(_06481_),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold528 (.A(_02401_),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold529 (.A(\fpga_top.cpu_top.pc_stage.cmd_ebreak_pc_pre ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold530 (.A(_05235_),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold531 (.A(_01514_),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold532 (.A(\fpga_top.qspi_if.word_data[19] ),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold533 (.A(_00976_),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold534 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][3] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold535 (.A(_06471_),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold536 (.A(_02392_),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold537 (.A(\fpga_top.uart_top.uart_logics.status_dump[1] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold538 (.A(\fpga_top.uart_top.uart_logics.rdata_snd_wait ),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold539 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][3] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold540 (.A(_02176_),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold541 (.A(\fpga_top.uart_top.uart_rec_char.data_word[2] ),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold542 (.A(_01241_),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold543 (.A(\fpga_top.cpu_top.csr_msie ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold544 (.A(\fpga_top.qspi_if.word_data[25] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold545 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[10] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold546 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[26] ),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold547 (.A(\fpga_top.io_spi_lite.miso_fifo.radr[0] ),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold548 (.A(\fpga_top.io_spi_lite.miso_fifo.radr_early[0] ),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold549 (.A(\fpga_top.qspi_if.word_data[10] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold550 (.A(_00967_),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold551 (.A(\fpga_top.uart_top.uart_rec_char.data_word[1] ),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold552 (.A(_01303_),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold553 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[24] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold554 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][0] ),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold555 (.A(_06280_),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold556 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][7] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold557 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][5] ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold558 (.A(_02386_),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold559 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[22] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold560 (.A(_01358_),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold561 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][1] ),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold562 (.A(_06442_),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold563 (.A(_02366_),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold564 (.A(\fpga_top.cpu_top.csr_mepc_ex[4] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold565 (.A(_01947_),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold566 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][0] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold567 (.A(_06274_),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold568 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][6] ),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold569 (.A(_02355_),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold570 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][6] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold571 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][6] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold572 (.A(_02363_),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold573 (.A(\fpga_top.uart_top.uart_rec_char.data_word[25] ),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold574 (.A(_04460_),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold575 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][5] ),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold576 (.A(_06366_),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold577 (.A(_02290_),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold578 (.A(\fpga_top.io_spi_lite.mosi_fifo.radr[0] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold579 (.A(\fpga_top.io_spi_lite.mosi_fifo.radr_early[0] ),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold580 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][3] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold581 (.A(_06435_),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold582 (.A(_02360_),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold583 (.A(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[3] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold584 (.A(_01116_),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold585 (.A(\fpga_top.io_spi_lite.sck_div[2] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold586 (.A(_08952_),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold587 (.A(_00030_),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold588 (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[0] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold589 (.A(_00068_),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold590 (.A(\fpga_top.qspi_if.wdata[7] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold591 (.A(_00930_),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold592 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][1] ),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold593 (.A(_06371_),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold594 (.A(_02294_),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold595 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[1] ),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold596 (.A(\fpga_top.qspi_if.word_data[15] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold597 (.A(_00972_),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold598 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][7] ),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold599 (.A(_02356_),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold600 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[19] ),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold601 (.A(\fpga_top.io_spi_lite.bit_sel_org[2] ),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold602 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][0] ),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold603 (.A(_02365_),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold604 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[6] ),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold605 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[11] ),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold606 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][0] ),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold607 (.A(_06384_),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold608 (.A(_02317_),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold609 (.A(\fpga_top.cpu_top.csr_mepc_ex[5] ),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold610 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[28] ),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold611 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][0] ),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold612 (.A(_02349_),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold613 (.A(\fpga_top.qspi_if.word_data[24] ),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold614 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][7] ),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold615 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[8] ),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold616 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[15] ),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold617 (.A(\fpga_top.uart_top.uart_rec_char.data_word[5] ),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold618 (.A(\fpga_top.uart_top.uart_logics.data_0[8] ),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold619 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[29] ),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold620 (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[15] ),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold621 (.A(_09393_),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold622 (.A(_00074_),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold623 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[6] ),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold624 (.A(\fpga_top.cpu_top.pc_stage.cmd_ecall_pc_pre ),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold625 (.A(_05318_),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold626 (.A(_01675_),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold627 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[28] ),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold628 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[23] ),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold629 (.A(_02033_),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold630 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[25] ),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold631 (.A(_01472_),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold632 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[8] ),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold633 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[8] ),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold634 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[19] ),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold635 (.A(_01355_),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold636 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[15] ),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold637 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[2] ),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold638 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][2] ),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold639 (.A(_02375_),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold640 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[8] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold641 (.A(_01344_),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold642 (.A(\fpga_top.uart_top.uart_if.tx_out_data[4] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold643 (.A(_01135_),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold644 (.A(\fpga_top.io_frc.frc_cntr_val[47] ),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold645 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[3] ),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold646 (.A(_01269_),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold647 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][0] ),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold648 (.A(_06468_),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold649 (.A(_02389_),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold650 (.A(\fpga_top.cpu_top.csr_mepc_ex[2] ),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold651 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][1] ),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold652 (.A(_06433_),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold653 (.A(_02358_),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold654 (.A(\fpga_top.uart_top.uart_logics.data_0[22] ),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold655 (.A(_01390_),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold656 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[7] ),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold657 (.A(_01273_),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold658 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[29] ),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold659 (.A(\fpga_top.io_uart_out.uart_term[1] ),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold660 (.A(_00075_),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold661 (.A(\fpga_top.io_spi_lite.bit_sel_org[1] ),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold662 (.A(_10574_),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold663 (.A(_00209_),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold664 (.A(\fpga_top.uart_top.uart_logics.data_0[4] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold665 (.A(\fpga_top.cpu_top.csr_mepc_ex[14] ),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold666 (.A(_01957_),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold667 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[31] ),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold668 (.A(_01297_),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold669 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[23] ),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold670 (.A(_01163_),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold671 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[18] ),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold672 (.A(\fpga_top.uart_top.uart_logics.data_0[16] ),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold673 (.A(_01384_),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold674 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[10] ),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold675 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[22] ),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold676 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[2] ),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold677 (.A(\fpga_top.io_spi_lite.miso_fifo.radr[2] ),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold678 (.A(\fpga_top.io_spi_lite.miso_fifo.radr_early[2] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold679 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mcause[4] ),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold680 (.A(\fpga_top.io_frc.frc_cmp_val[11] ),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold681 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[27] ),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold682 (.A(\fpga_top.cpu_top.csr_mepc_ex[25] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold683 (.A(_01968_),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold684 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[24] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold685 (.A(\fpga_top.qspi_if.word_data[11] ),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold686 (.A(_00968_),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold687 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[27] ),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold688 (.A(_02069_),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold689 (.A(\fpga_top.qspi_if.sck_cntr[6] ),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold690 (.A(_09263_),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold691 (.A(_00048_),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold692 (.A(\fpga_top.qspi_if.word_data[16] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold693 (.A(_00973_),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold694 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[24] ),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold695 (.A(_01290_),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold696 (.A(\fpga_top.cpu_top.csr_mepc_ex[31] ),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold697 (.A(_01974_),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold698 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][4] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold699 (.A(_02369_),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold700 (.A(\fpga_top.uart_top.uart_rec_char.data_word[10] ),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold701 (.A(_01249_),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold702 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][4] ),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold703 (.A(_06454_),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold704 (.A(_02377_),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold705 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[15] ),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold706 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][0] ),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold707 (.A(_06269_),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold708 (.A(_02173_),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold709 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[13] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold710 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[28] ),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold711 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][0] ),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold712 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[18] ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold713 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[29] ),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold714 (.A(_01476_),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold715 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][6] ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold716 (.A(_06367_),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold717 (.A(_02291_),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold718 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[30] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold719 (.A(_01609_),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold720 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][2] ),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold721 (.A(_02391_),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold722 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[3][5] ),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold723 (.A(_02378_),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold724 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[23] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold725 (.A(_02000_),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold726 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[21] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold727 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[20] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold728 (.A(\fpga_top.qspi_if.word_data[23] ),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold729 (.A(\fpga_top.uart_top.uart_logics.data_0[23] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold730 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][3] ),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold731 (.A(_06426_),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold732 (.A(_02352_),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold733 (.A(\fpga_top.io_spi_lite.spi_sck_div[9] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold734 (.A(\fpga_top.cpu_top.csr_mepc_ex[28] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold735 (.A(_01971_),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold736 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[13] ),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold737 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][5] ),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold738 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][5] ),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold739 (.A(_02362_),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold740 (.A(\fpga_top.cpu_start_adr[28] ),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold741 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[25] ),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold742 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][0] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold743 (.A(_06363_),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold744 (.A(_02285_),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold745 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[6][1] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold746 (.A(_06424_),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold747 (.A(_02350_),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold748 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[1] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold749 (.A(_00378_),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold750 (.A(\fpga_top.uart_top.uart_logics.data_0[24] ),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold751 (.A(_01392_),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold752 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mpie ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold753 (.A(_01905_),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold754 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[12] ),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold755 (.A(\fpga_top.uart_top.uart_rec_char.bpoint_en ),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold756 (.A(_01267_),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold757 (.A(\fpga_top.uart_top.uart_rec_char.data_word[12] ),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold758 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][5] ),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold759 (.A(_02194_),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold760 (.A(\fpga_top.io_frc.frc_cntr_val[41] ),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold761 (.A(_02121_),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold762 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[5] ),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold763 (.A(\fpga_top.io_frc.frc_cmp_val[7] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold764 (.A(\fpga_top.io_frc.frc_cntr_val[46] ),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold765 (.A(_02126_),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold766 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtval[0] ),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold767 (.A(_01906_),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold768 (.A(\fpga_top.uart_top.uart_logics.data_0[30] ),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold769 (.A(_01398_),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold770 (.A(\fpga_top.cpu_top.csr_mepc_ex[12] ),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold771 (.A(\fpga_top.uart_top.uart_rec_char.data_word[4] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold772 (.A(_04439_),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold773 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[19] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold774 (.A(_01285_),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold775 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[14] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold776 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[22] ),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold777 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[12] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold778 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[21] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold779 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][2] ),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold780 (.A(_02359_),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold781 (.A(\fpga_top.qspi_if.word_data[5] ),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold782 (.A(_00962_),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold783 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[21] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold784 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[24] ),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold785 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[6] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold786 (.A(_01272_),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold787 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[2] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold788 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[26] ),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold789 (.A(\fpga_top.cpu_top.csr_mepc_ex[13] ),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold790 (.A(\fpga_top.cpu_top.csr_mepc_ex[7] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold791 (.A(_00123_),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold792 (.A(\fpga_top.io_frc.frc_cmp_val[15] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold793 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][5] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold794 (.A(_02234_),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold795 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[17] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold796 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[10] ),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold797 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[17] ),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold798 (.A(_01994_),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold799 (.A(\fpga_top.io_uart_out.uart_term[3] ),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold800 (.A(_00077_),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold801 (.A(\fpga_top.qspi_if.wdata[11] ),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold802 (.A(_00934_),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold803 (.A(\fpga_top.uart_top.uart_rec_char.data_word[21] ),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold804 (.A(_01260_),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold805 (.A(\fpga_top.io_led.led_value[1] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold806 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][0] ),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold807 (.A(_02229_),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold808 (.A(\fpga_top.cpu_top.csr_mepc_ex[9] ),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold809 (.A(\fpga_top.io_uart_out.uart_term[2] ),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold810 (.A(_00076_),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold811 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[29] ),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold812 (.A(\fpga_top.qspi_if.sck_div[5] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold813 (.A(\fpga_top.cpu_top.csr_mepc_ex[8] ),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold814 (.A(_01951_),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold815 (.A(\fpga_top.uart_top.uart_rec_char.data_word[7] ),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold816 (.A(\fpga_top.io_frc.frc_cntr_val[63] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold817 (.A(_02143_),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold818 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[26] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold819 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][6] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold820 (.A(_02235_),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold821 (.A(\fpga_top.uart_top.uart_logics.data_0[28] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold822 (.A(_01396_),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold823 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[2] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold824 (.A(\fpga_top.io_frc.frc_cntr_val[52] ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold825 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[15] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold826 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][20] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold827 (.A(\fpga_top.uart_top.uart_rec_char.data_cntr[2] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold828 (.A(_01300_),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold829 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[14] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold830 (.A(_01280_),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold831 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][6] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold832 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][19] ),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold833 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[0] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold834 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][4] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold835 (.A(_02233_),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold836 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[4][2] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold837 (.A(_02367_),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold838 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][0] ),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold839 (.A(_02205_),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold840 (.A(\fpga_top.cpu_top.csr_mepc_ex[27] ),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold841 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][5] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold842 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][7] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold843 (.A(_06368_),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold844 (.A(_02292_),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold845 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][2] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold846 (.A(\fpga_top.bus_gather.d_write_data[5] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold847 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][19] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold848 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][10] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold849 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][4] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold850 (.A(_02257_),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold851 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][7] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold852 (.A(_02212_),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold853 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][6] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold854 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][23] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold855 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][12] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold856 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[15] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold857 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][30] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold858 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][14] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold859 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][8] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold860 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][5] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold861 (.A(_02274_),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold862 (.A(\fpga_top.uart_top.uart_if.rx_fifo_dcntr[2] ),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold863 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][4] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold864 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][13] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold865 (.A(\fpga_top.uart_top.uart_logics.data_0[2] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold866 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][11] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold867 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][15] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold868 (.A(\fpga_top.io_frc.frc_cntr_val[33] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold869 (.A(_02113_),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold870 (.A(\fpga_top.cpu_top.execution.csr_array.csr_spie ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold871 (.A(\fpga_top.uart_top.uart_logics.data_0[26] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold872 (.A(_01394_),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold873 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][5] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold874 (.A(_02210_),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold875 (.A(\fpga_top.io_frc.frc_cmp_val[32] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold876 (.A(\fpga_top.cpu_start_adr[11] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold877 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][7] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold878 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[1][4] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold879 (.A(_06472_),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold880 (.A(_02393_),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold881 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][0] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold882 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][28] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold883 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[10] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold884 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][1] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold885 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][26] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold886 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][6] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold887 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[1] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold888 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][2] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold889 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][2] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold890 (.A(_02231_),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold891 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][4] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold892 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][16] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold893 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][21] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold894 (.A(\fpga_top.io_frc.frc_cntr_val[58] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold895 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][29] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold896 (.A(\fpga_top.cpu_top.csr_mepc_ex[20] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold897 (.A(_01963_),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold898 (.A(\fpga_top.io_frc.frc_cntr_val[36] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold899 (.A(_02116_),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold900 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[21] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold901 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][9] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold902 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][26] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold903 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][9] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold904 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][2] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold905 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][26] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold906 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][30] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold907 (.A(\fpga_top.cpu_start_adr[31] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold908 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][9] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold909 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][26] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold910 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][0] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold911 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][10] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold912 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][4] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold913 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][30] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold914 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][2] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold915 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][3] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold916 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[9] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold917 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][5] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold918 (.A(\fpga_top.uart_top.uart_rec_char.pdata[2] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold919 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][3] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold920 (.A(_02256_),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold921 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][7] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold922 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][21] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold923 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][16] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold924 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][15] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold925 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][30] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold926 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][20] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold927 (.A(\fpga_top.qspi_if.word_data[9] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold928 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][28] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold929 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][0] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold930 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][30] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold931 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][27] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold932 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][4] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold933 (.A(_02289_),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold934 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][5] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold935 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][3] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold936 (.A(_02232_),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold937 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][23] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold938 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][19] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold939 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][2] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold940 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][4] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold941 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][10] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold942 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][23] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold943 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][30] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold944 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][30] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold945 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][6] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold946 (.A(_02211_),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold947 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][1] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold948 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][4] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold949 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][6] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold950 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][29] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold951 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][11] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold952 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][29] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold953 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][7] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold954 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[25] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold955 (.A(_01361_),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold956 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][6] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold957 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][29] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold958 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][16] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold959 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][14] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold960 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][7] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold961 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][28] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold962 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][11] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold963 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][27] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold964 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[6] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold965 (.A(_01342_),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold966 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][1] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold967 (.A(_02230_),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold968 (.A(\fpga_top.uart_top.uart_rec_char.data_word[3] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold969 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][26] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold970 (.A(\fpga_top.cpu_top.csr_mepc_ex[10] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold971 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][5] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold972 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][1] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold973 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][1] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold974 (.A(_02206_),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold975 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][30] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold976 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][11] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold977 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][3] ),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold978 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][12] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold979 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][22] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold980 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][5] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold981 (.A(_02250_),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold982 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][4] ),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold983 (.A(_02321_),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold984 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][4] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold985 (.A(_02153_),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold986 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][12] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold987 (.A(\fpga_top.cpu_top.data_rw_mem.req_hw_dly ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold988 (.A(_06051_),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold989 (.A(_02076_),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold990 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][21] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold991 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][6] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold992 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][5] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold993 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][15] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold994 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][4] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold995 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][30] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold996 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][2] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold997 (.A(\fpga_top.cpu_top.csr_mepc_ex[6] ),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold998 (.A(\fpga_top.cpu_top.csr_mepc_ex[26] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold999 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][2] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][30] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][26] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][29] ),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][27] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][23] ),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][7] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][2] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][25] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][18] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][31] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][13] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][12] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][21] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[26] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_01362_),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\fpga_top.cpu_top.csr_mepc_ex[24] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][19] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][16] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][22] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][5] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][5] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][11] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][16] ),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][9] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][2] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold1025 (.A(_02271_),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][1] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][23] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][7] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[10] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][14] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][28] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][11] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\fpga_top.io_frc.frc_cmp_val[24] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][18] ),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][30] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][5] ),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][2] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_06365_),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold1039 (.A(_02287_),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][25] ),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][28] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][12] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\fpga_top.qspi_if.rdwrch[5] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][15] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][25] ),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][4] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold1047 (.A(_02209_),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][7] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][7] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][1] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][0] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][16] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][30] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][27] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][25] ),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][25] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][23] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][3] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\fpga_top.io_uart_out.uart_term[5] ),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold1060 (.A(_00079_),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][11] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][15] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][21] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][11] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][5] ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][17] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][6] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][25] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][24] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][27] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][24] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][24] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][22] ),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][9] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][11] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][22] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][10] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][13] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[6][3] ),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][16] ),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][9] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][12] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][8] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\fpga_top.qspi_if.rwait_cntr[3] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold1085 (.A(_01022_),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][6] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][25] ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][27] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][18] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][22] ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][30] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][3] ),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][0] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][10] ),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][9] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][1] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][14] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][1] ),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][18] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[11] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][5] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][23] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][8] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][14] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[18] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold1106 (.A(_01354_),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][0] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][15] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][2] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][17] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][19] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][15] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][7] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold1114 (.A(_02188_),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][31] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][3] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold1117 (.A(_02208_),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[29] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][25] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][1] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][13] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][29] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][0] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][26] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][15] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][19] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][30] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][10] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][30] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][19] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][25] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][20] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][25] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][26] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][26] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][1] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold1137 (.A(_02262_),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][4] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold1139 (.A(_02161_),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][31] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][24] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][2] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold1143 (.A(_02263_),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][31] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][28] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][8] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][14] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][26] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][24] ),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][5] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][5] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][25] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][22] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][15] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][18] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][27] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][2] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][22] ),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][13] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][1] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][3] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][30] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][0] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[5][0] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold1165 (.A(_02357_),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][1] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][4] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][21] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][29] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][13] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][29] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][16] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][23] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][20] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\fpga_top.cpu_top.csr_mepc_ex[18] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][2] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][2] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][17] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][3] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][17] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][25] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][5] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][13] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][11] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][10] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[31] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][17] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][25] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][31] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][5] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][20] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][16] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\fpga_top.uart_top.uart_logics.data_0[21] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][4] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][10] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][13] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][17] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][20] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][24] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][19] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][15] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][29] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][21] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][9] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][6] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[7][2] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold1207 (.A(_02207_),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][12] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][0] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram[2][4] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold1211 (.A(_06463_),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold1212 (.A(_02385_),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][8] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][11] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][27] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][6] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold1217 (.A(_02251_),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][27] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][1] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][1] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][21] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][7] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold1223 (.A(_02228_),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][12] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][12] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][26] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\fpga_top.bus_gather.i_read_adr[8] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold1228 (.A(_01486_),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][0] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][13] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][27] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][7] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold1233 (.A(_02252_),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][30] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][24] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][4] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold1237 (.A(_02241_),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\fpga_top.uart_top.uart_logics.data_0[25] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold1239 (.A(_01393_),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][16] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][31] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][26] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][8] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\fpga_top.cpu_start_adr[30] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[14] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold1246 (.A(_01350_),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][22] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\fpga_top.uart_top.uart_logics.data_0[20] ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold1249 (.A(_01388_),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][14] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][11] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][0] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold1253 (.A(_02269_),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][6] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][4] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][30] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][16] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][10] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[5][7] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold1260 (.A(_02236_),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][7] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][20] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][1] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][9] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][7] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold1266 (.A(_02260_),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][11] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][23] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][29] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][26] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][10] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][20] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][9] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][17] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][31] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][5] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold1277 (.A(_02242_),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][3] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][21] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[0] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][0] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][3] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][27] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][21] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][9] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][13] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][3] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][22] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][14] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][8] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][18] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][0] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][26] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][7] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][12] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][20] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][27] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][0] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][3] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][28] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][29] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][4] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][3] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][8] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][4] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][18] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][10] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][16] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][27] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][24] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[26] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][2] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold1313 (.A(_02247_),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][3] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][4] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[30] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][7] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][4] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][9] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][5] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][9] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][23] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][31] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][14] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][26] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][1] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][24] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][11] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][12] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][27] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][29] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][6] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][19] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][1] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][15] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][28] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][14] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][19] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][21] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][8] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][13] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][1] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][24] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][5] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][23] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][7] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][16] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][17] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][21] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][5] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][3] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][4] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][0] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold1354 (.A(_02221_),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][10] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][17] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][7] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][14] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][20] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][10] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][5] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][1] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][10] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][6] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][6] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][12] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][6] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][14] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][7] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][4] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][31] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][26] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][0] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][8] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][5] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][19] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][14] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][7] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][31] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][19] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][28] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][0] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold1383 (.A(_02237_),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][15] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][2] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][20] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][22] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][14] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][2] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][24] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[25] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][11] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][16] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][22] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][11] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][21] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][10] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][23] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][4] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][12] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][27] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][4] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][21] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][3] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][8] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[18] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_01284_),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][7] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][18] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\fpga_top.io_uart_out.rout[0] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold1411 (.A(_04463_),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold1412 (.A(_01330_),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][0] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][31] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][23] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][0] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][19] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][15] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][31] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][17] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][13] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][10] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][8] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][23] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][21] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][2] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold1427 (.A(_02239_),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][3] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][17] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][24] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][26] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][2] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][13] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][0] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][21] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][26] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][20] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[7] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][9] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][20] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][4] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold1442 (.A(_02249_),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][27] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][30] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[9] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold1446 (.A(_01345_),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][25] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][3] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][0] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][23] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][14] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][12] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][24] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[8] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold1455 (.A(_01274_),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][25] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][3] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][28] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][19] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][2] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold1461 (.A(_02223_),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][20] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\fpga_top.cpu_top.execution.csr_array.csr_spp ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][17] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][24] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][27] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][7] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][7] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][31] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][29] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][11] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][28] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][6] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][7] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\fpga_top.cpu_top.csr_mepc_ex[23] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\fpga_top.uart_top.uart_rec_char.data_cntr[1] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold1477 (.A(_01299_),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][26] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[8] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][22] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][2] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\fpga_top.qspi_if.wdata[2] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold1483 (.A(_00925_),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][25] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][31] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][3] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold1487 (.A(_02264_),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][5] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][17] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][1] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold1491 (.A(_02222_),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][30] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][13] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][8] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][7] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][25] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][24] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][26] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][12] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][6] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][31] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][28] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][7] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][6] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][6] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold1506 (.A(_02243_),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][18] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][22] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][5] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][7] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\fpga_top.uart_top.uart_logics.data_0[10] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][2] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][8] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][23] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][18] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][5] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][24] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][30] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][13] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][16] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\fpga_top.interrupter.int_status_rx ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold1522 (.A(_00292_),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][22] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][13] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][4] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][4] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][0] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][12] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][1] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][7] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][0] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][25] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][4] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][9] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][0] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][3] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][7] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\fpga_top.io_uart_out.rout[2] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold1539 (.A(_04464_),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold1540 (.A(_01332_),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][27] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\fpga_top.io_frc.frc_cmp_val[44] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][23] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][6] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][16] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][4] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][14] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][12] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][18] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][4] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][31] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[13] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][30] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][30] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\fpga_top.io_frc.frc_cmp_val[52] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][3] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][2] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][12] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][29] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][8] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[22] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold1562 (.A(_01288_),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][6] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][15] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][29] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][1] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][3] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][10] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][20] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][5] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][17] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][5] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][3] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][9] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][10] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][9] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[25] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold1578 (.A(_01291_),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[4] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][21] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][2] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[17] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][25] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][28] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][21] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][15] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][18] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][16] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][12] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][10] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][5] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold1592 (.A(_02226_),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][29] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][16] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][17] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][11] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][7] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][9] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold1599 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][18] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][2] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][17] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][7] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][13] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][1] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold1605 (.A(_02270_),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][9] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][27] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][3] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][2] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][4] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold1611 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][27] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][8] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][7] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][29] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][26] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][7] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][0] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][21] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][0] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][2] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][5] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\fpga_top.cpu_top.csr_mepc_ex[30] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][3] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\fpga_top.bus_gather.d_write_data[10] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][21] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][3] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[3][4] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][26] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][11] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mscrach[18] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][3] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold1632 (.A(_02248_),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][23] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][4] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][4] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][5] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][4] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold1638 (.A(_02169_),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][9] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][6] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][6] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][20] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\fpga_top.io_frc.frc_cmp_val[43] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][31] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][26] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][26] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][3] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold1648 (.A(_02240_),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][16] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][5] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][5] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][3] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][4] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][12] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][3] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[27] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\fpga_top.uart_top.uart_logics.data_0[13] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][19] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][24] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][8] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][1] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold1662 (.A(_02238_),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][25] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][2] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][31] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][18] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][18] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][1] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[1][7] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold1670 (.A(_02196_),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[2][3] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][2] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][2] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][30] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][1] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][9] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][6] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][9] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[23] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold1680 (.A(_01289_),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][19] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][26] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][26] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][22] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][8] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][10] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][3] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][3] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][13] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][21] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][24] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][1] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][14] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][27] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][13] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][0] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][16] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold1698 (.A(_00101_),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][12] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][23] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][31] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][6] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][5] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold1704 (.A(_02258_),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][20] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][2] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold1707 (.A(_00104_),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][6] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][8] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][6] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][12] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\fpga_top.io_spi_lite.spi_sck_div[8] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[3] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_01339_),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][17] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][19] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][17] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[0] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][2] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][16] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][18] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][25] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][29] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][6] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][24] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][4] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold1727 (.A(_02273_),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][30] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][21] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][16] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][15] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][24] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][27] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][10] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][12] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][17] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][2] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][3] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][18] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][21] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][28] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[19] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][22] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][27] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][19] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][16] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][4] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][31] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][23] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][12] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][23] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][15] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][15] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][24] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][27] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][2] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold1757 (.A(_02255_),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][13] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][9] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][24] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][4] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][10] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][6] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][31] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\fpga_top.qspi_if.qspi_state[9] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold1766 (.A(_02079_),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][22] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][5] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][7] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][10] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[25] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][11] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][5] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][27] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][12] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][5] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][20] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][23] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][25] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][16] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[3][5] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][25] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][14] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[19] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][22] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][13] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][3] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][10] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][24] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][28] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][27] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][8] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][1] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][20] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[31] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][20] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][0] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][0] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\fpga_top.io_frc.frc_cntr_val[43] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold1800 (.A(_02123_),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][10] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][8] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][23] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][10] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][2] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\fpga_top.io_uart_out.uart_io_char[6] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][22] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][17] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][8] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][12] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\fpga_top.io_frc.frc_cntr_val[34] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold1812 (.A(_02114_),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][18] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][2] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][14] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][8] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][21] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][28] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][28] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[6][1] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[2] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][19] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][21] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[5] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold1825 (.A(_01341_),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][16] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][1] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\fpga_top.io_uart_out.uart_term[6] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold1829 (.A(_00080_),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\fpga_top.io_uart_out.uart_io_char[2] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][3] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][9] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\fpga_top.qspi_if.sck_div[2] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][6] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][5] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][23] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][9] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][14] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\fpga_top.io_led.led_value[0] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][15] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[4] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold1842 (.A(_01583_),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\fpga_top.io_frc.frc_cmp_val[59] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][25] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][19] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][22] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][7] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[4][7] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold1849 (.A(_02244_),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][20] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][31] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][3] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][25] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\fpga_top.uart_top.uart_if.byte_data[7] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][29] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][6] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\fpga_top.io_uart_out.uart_io_char[5] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][7] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\fpga_top.qspi_if.adr_rw[12] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold1860 (.A(_01001_),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][22] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\fpga_top.io_frc.frc_cmp_val[18] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][14] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][3] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold1865 (.A(_02168_),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][24] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\fpga_top.io_spi_lite.spi_mode[2] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][19] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][7] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][29] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][29] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][19] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][6] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][2] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][0] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][21] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][4] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][13] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][3] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][6] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][6] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold1882 (.A(_02227_),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[20] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[11] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][20] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][9] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\fpga_top.io_spi_lite.mosi_pp_cntr[0] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][12] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\fpga_top.io_uart_out.uart_io_char[0] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold1890 (.A(_00111_),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][22] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\fpga_top.uart_top.uart_rec_char.data_word[17] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\fpga_top.qspi_if.word_data[14] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][20] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][28] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][0] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][13] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][2] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][26] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][15] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][7] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][15] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][24] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][19] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][20] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[5][3] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][17] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][28] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][1] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][13] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\fpga_top.uart_top.uart_logics.data_0[3] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][28] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][22] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][10] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][4] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][22] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][31] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][18] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][15] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\fpga_top.io_frc.frc_cmp_val[47] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][31] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][9] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][8] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][23] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][11] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][6] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][17] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][31] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][23] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][28] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][14] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][14] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][30] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][25] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][11] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][28] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[7][4] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold1938 (.A(_02281_),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][31] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][1] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][21] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][13] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][14] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][12] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][17] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][19] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][17] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][26] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][23] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][6] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold1951 (.A(_02259_),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][11] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][7] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][20] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\fpga_top.io_frc.frc_cmp_val[23] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][24] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][29] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][15] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][4] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][19] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][6] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][27] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][14] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][19] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][18] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][14] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][1] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold1968 (.A(_02254_),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][19] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][15] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][18] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][25] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][6] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\fpga_top.qspi_if.word_data[4] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold1975 (.A(_00961_),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][28] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][7] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][5] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][4] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][4] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][27] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][19] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\fpga_top.io_frc.frc_cmp_val[49] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[0] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][31] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][30] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][11] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][2] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\fpga_top.bus_gather.d_write_data[1] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][26] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\fpga_top.io_uart_out.uart_term[9] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold1992 (.A(_00083_),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][3] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][3] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold1995 (.A(_02272_),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][4] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold1997 (.A(_02265_),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[8] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][31] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][22] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\fpga_top.uart_top.uart_logics.trash_cond_dly ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold2002 (.A(_01440_),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][28] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[1][4] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][9] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][27] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][3] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][30] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[5][1] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][6] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][4] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\fpga_top.qspi_if.dbg_2div_wirte_half_end ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold2013 (.A(_00019_),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][4] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][0] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][15] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][17] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][9] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][3] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][31] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][31] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\fpga_top.uart_top.uart_logics.data_0[17] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\fpga_top.cpu_top.csr_mepc_ex[22] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold2024 (.A(_01965_),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][0] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][18] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][29] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][29] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][3] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold2030 (.A(_02224_),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][16] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][11] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\fpga_top.qspi_if.wredge[2] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\fpga_top.cpu_top.csr_mepc_ex[16] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold2035 (.A(_01959_),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][28] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[16] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold2038 (.A(_01282_),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][24] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][29] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][24] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[2] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold2043 (.A(_06279_),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][6] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][3] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][30] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][22] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\fpga_top.io_frc.frc_cmp_val[8] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[4][3] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\fpga_top.io_frc.frc_cmp_val[25] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold2051 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][28] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][26] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[4] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold2054 (.A(_01451_),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold2055 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][17] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][0] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][15] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][7] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][7] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[24][14] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][29] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][22] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][20] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][7] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold2065 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][10] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][2] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][30] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\fpga_top.io_uart_out.uart_io_char[7] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][29] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][31] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[31] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold2072 (.A(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[2] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold2073 (.A(_01125_),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\fpga_top.io_frc.frc_cntr_val[59] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][13] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\fpga_top.io_frc.frc_cmp_val[53] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][12] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][6] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][15] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][0] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\fpga_top.cpu_top.br_ofs[1] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][10] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][16] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][25] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold2085 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][6] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][28] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][30] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][6] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][5] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][3] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][7] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][2] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\fpga_top.io_frc.frc_cntr_val[62] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold2094 (.A(_02142_),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold2095 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][25] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][1] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][21] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][18] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][12] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\fpga_top.cpu_top.pc_stage.frc_cntr_val_leq_latch ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold2101 (.A(_05233_),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][19] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold2103 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][20] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][5] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\fpga_top.io_frc.frc_cmp_val[60] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][24] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\fpga_top.io_frc.frc_cmp_val[34] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][25] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][5] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold2110 (.A(\fpga_top.uart_top.uart_rec_char.data_word[23] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold2111 (.A(_04458_),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][29] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][24] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][19] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold2115 (.A(\fpga_top.qspi_if.sck_div[7] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][1] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][27] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][0] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold2119 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[24] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold2120 (.A(_01360_),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold2121 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][25] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\fpga_top.io_frc.frc_cmp_val[63] ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][23] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[17] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][23] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][13] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[12] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold2128 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][15] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\fpga_top.uart_top.uart_if.tx_out_cntr[2] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold2130 (.A(_03679_),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold2131 (.A(_01130_),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][14] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[6][4] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold2134 (.A(_02225_),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\fpga_top.io_frc.frc_cntr_val[38] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold2136 (.A(_02118_),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][12] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][24] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][21] ),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\fpga_top.io_frc.frc_cmp_val[0] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][1] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold2142 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][13] ),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][29] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[12][6] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][18] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold2146 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][13] ),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][10] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold2148 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][4] ),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[8][17] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold2150 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][15] ),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][26] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold2152 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][11] ),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][1] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\fpga_top.io_frc.frc_cmp_val[20] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][28] ),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold2156 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][29] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][13] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold2158 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][29] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][8] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][23] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][20] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][1] ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][13] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][19] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[4][22] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\fpga_top.uart_top.uart_logics.data_0[31] ),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold2167 (.A(_01399_),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][23] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold2169 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][21] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][5] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][28] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold2172 (.A(_00100_),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][18] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\fpga_top.uart_top.uart_if.byte_data[6] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mcause[3] ),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold2176 (.A(_01941_),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][20] ),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\fpga_top.qspi_if.wrcmd1[7] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mcause[0] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold2180 (.A(_01938_),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][27] ),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold2182 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][1] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[20] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][0] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold2185 (.A(_02261_),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold2186 (.A(_00090_),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[20][8] ),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\fpga_top.io_spi_lite.spi_mode[9] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][11] ),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][28] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\fpga_top.bus_gather.d_write_data[15] ),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold2192 (.A(\fpga_top.io_frc.frc_cmp_val[12] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][5] ),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold2194 (.A(_02266_),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold2195 (.A(\fpga_top.io_spi_lite.miso_byte_org[4] ),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold2196 (.A(_10549_),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][20] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\fpga_top.io_frc.frc_cmp_val[14] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\fpga_top.uart_top.uart_rec_char.data_cntr[0] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold2200 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][17] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][18] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][4] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold2203 (.A(_00109_),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][8] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][28] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold2206 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][5] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[0][11] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][1] ),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][2] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\fpga_top.qspi_if.rst_cntr[1] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold2211 (.A(_03633_),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold2212 (.A(_01104_),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold2213 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][22] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\fpga_top.io_frc.frc_cmp_val[55] ),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][22] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold2216 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][19] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][22] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][16] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][18] ),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][18] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][18] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][13] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold2223 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[7] ),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold2224 (.A(_01343_),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][29] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\fpga_top.io_frc.frc_cmp_val[22] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold2227 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][4] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][9] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][21] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[4][1] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold2231 (.A(_02166_),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][24] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][11] ),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[23] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][17] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[2][23] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][5] ),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold2238 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][2] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][6] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][14] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[1][6] ),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][0] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold2243 (.A(_02245_),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\fpga_top.cpu_top.csr_mepc_ex[19] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][14] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[0] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][11] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][18] ),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[6][30] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][8] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][16] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][7] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[28] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][9] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[13][17] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][12] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\fpga_top.bus_gather.d_write_data[3] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[2] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][7] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold2260 (.A(\fpga_top.io_spi_lite.miso_byte_org[3] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold2261 (.A(_10548_),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[17][1] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[29][4] ),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold2264 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][1] ),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][0] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\fpga_top.io_frc.frc_cmp_val[48] ),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[13] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold2268 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][15] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[0] ),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold2270 (.A(_01579_),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[3][1] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold2272 (.A(_02246_),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold2273 (.A(\fpga_top.io_frc.frc_cmp_val[62] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[14][16] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\fpga_top.qspi_if.rst_cntr[3] ),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold2276 (.A(_03638_),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][21] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold2278 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[25][5] ),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\fpga_top.uart_top.uart_logics.data_0[11] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold2280 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[1][8] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\fpga_top.io_uart_out.rx_data_latch[6] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold2282 (.A(_00389_),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold2283 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][8] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mcause[6] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold2285 (.A(_01944_),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\fpga_top.qspi_if.rdedge[0] ),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold2287 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][2] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][3] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold2289 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[21][8] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[27][4] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold2291 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][15] ),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\fpga_top.io_uart_out.uart_term[7] ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold2293 (.A(_00081_),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold2294 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][25] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold2295 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][20] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold2296 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][11] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][2] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[25] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[22][10] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\fpga_top.qspi_if.sck_div[6] ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold2301 (.A(\fpga_top.io_frc.frc_cntr_val[61] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][17] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][1] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold2304 (.A(\fpga_top.io_frc.frc_cntr_val[44] ),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold2305 (.A(_02124_),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[31][18] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold2307 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[2][0] ),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold2308 (.A(_02253_),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\fpga_top.io_uart_out.rout[4] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold2310 (.A(_04465_),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold2311 (.A(_01334_),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[26][16] ),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\fpga_top.io_uart_out.rx_disable_echoback_value ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[10][16] ),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold2315 (.A(\fpga_top.uart_top.uart_rec_char.data_word[19] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold2316 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[28][6] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][7] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold2318 (.A(_02276_),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\fpga_top.bus_gather.d_write_data[4] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold2320 (.A(\fpga_top.io_frc.frc_cmp_val[6] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold2321 (.A(\fpga_top.cpu_start_adr[29] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[5][20] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][14] ),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\fpga_top.uart_top.uart_logics.data_0[1] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram[0][3] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][15] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold2327 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[16] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold2328 (.A(\fpga_top.io_frc.frc_cmp_val[31] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold2329 (.A(_00105_),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold2330 (.A(_00102_),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\fpga_top.io_frc.frc_cntr_val[50] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\fpga_top.io_frc.frc_cmp_val[5] ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold2333 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[28] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold2334 (.A(_01475_),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[28] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold2336 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[15][14] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold2337 (.A(\fpga_top.io_spi_lite.miso_byte_org[2] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold2338 (.A(_10547_),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold2339 (.A(_00108_),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold2340 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[30][8] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][31] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][18] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[10] ),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold2344 (.A(\fpga_top.io_frc.frc_cmp_val[46] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\fpga_top.uart_top.uart_if.byte_data[5] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold2346 (.A(_01436_),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold2347 (.A(\fpga_top.qspi_if.rdwrch[2] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[23][9] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[11][28] ),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\fpga_top.uart_top.uart_if.tx_state[0] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold2351 (.A(_09516_),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\fpga_top.qspi_if.sck_div[1] ),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\fpga_top.io_frc.frc_cmp_val[40] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold2354 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[16][26] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\fpga_top.io_frc.frc_cmp_val[61] ),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold2356 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram[0][6] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold2357 (.A(_02275_),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\fpga_top.io_frc.frc_cmp_val[9] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold2359 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[9][6] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\fpga_top.cpu_top.execution.csr_array.csr_sscrach[31] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[6] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold2362 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[12] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold2363 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[3][17] ),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold2364 (.A(_00096_),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold2365 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[7][2] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\fpga_top.uart_top.uart_logics.data_0[7] ),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold2367 (.A(\fpga_top.dbg_bpoint_en[0] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold2368 (.A(_00123_),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold2369 (.A(_00098_),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold2370 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][27] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\fpga_top.io_frc.frc_cmp_val[51] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\fpga_top.io_frc.frc_cmp_val[56] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold2373 (.A(\fpga_top.uart_top.uart_logics.data_0[12] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[21] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold2375 (.A(_01357_),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold2376 (.A(\fpga_top.qspi_if.dbg_reg_2div_cec_read ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[2] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\fpga_top.io_spi_lite.miso_byte_org[5] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold2379 (.A(_10550_),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold2380 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[0][3] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold2381 (.A(\fpga_top.bus_gather.d_write_data[0] ),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold2382 (.A(_05285_),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold2383 (.A(_00114_),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold2384 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[7][10] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold2385 (.A(\fpga_top.io_frc.frc_cmp_val[41] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold2386 (.A(\fpga_top.qspi_if.read_latency_0[3] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\fpga_top.qspi_if.wrcmd1[2] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold2388 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][11] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\fpga_top.qspi_if.wrcmd0[0] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold2390 (.A(\fpga_top.io_frc.frc_cmp_val[45] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[19][0] ),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold2392 (.A(\fpga_top.cpu_top.csr_mepc_ex[17] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold2393 (.A(\fpga_top.uart_top.uart_logics.data_0[18] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold2394 (.A(\fpga_top.qspi_if.rdwrch[3] ),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold2395 (.A(\fpga_top.io_frc.frc_cntr_val[42] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold2396 (.A(_02122_),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\fpga_top.io_frc.frc_cmp_val[54] ),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\fpga_top.qspi_if.wrcmd0[7] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\fpga_top.io_spi_lite.miso_byte_org[1] ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold2400 (.A(_10546_),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold2401 (.A(_00097_),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\fpga_top.io_frc.frc_cmp_val[2] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold2403 (.A(\fpga_top.io_frc.frc_cmp_val[39] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\fpga_top.uart_top.uart_logics.data_0[9] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold2405 (.A(\fpga_top.cpu_start_adr[7] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\fpga_top.uart_top.uart_logics.data_0[15] ),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold2407 (.A(\fpga_top.io_frc.frc_cntr_val[53] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold2408 (.A(_06196_),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold2409 (.A(\fpga_top.cpu_top.execution.csr_array.csr_rd_data[1] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold2410 (.A(\fpga_top.qspi_if.wrcmd0[1] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\fpga_top.io_spi_lite.sck_div[7] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold2412 (.A(_08962_),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold2413 (.A(_00035_),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold2414 (.A(\fpga_top.qspi_if.word_data[12] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold2415 (.A(_00969_),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold2416 (.A(\fpga_top.uart_top.uart_if.tx_state[1] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold2417 (.A(_09335_),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold2418 (.A(_01129_),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold2419 (.A(\fpga_top.io_spi_lite.miso_byte_org[0] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold2420 (.A(_10545_),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold2421 (.A(\fpga_top.io_uart_out.rx_data_latch[5] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold2422 (.A(_00388_),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold2423 (.A(\fpga_top.qspi_if.sio_in_sync[0] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold2424 (.A(_00957_),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold2425 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[30] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold2426 (.A(_02072_),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold2427 (.A(\fpga_top.io_frc.frc_cmp_val[57] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold2428 (.A(\fpga_top.qspi_if.read_latency_0[2] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold2429 (.A(\fpga_top.qspi_if.sio_in_sync[3] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold2430 (.A(_00960_),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold2431 (.A(\fpga_top.io_frc.frc_cntr_val[13] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold2432 (.A(_00409_),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold2433 (.A(\fpga_top.io_frc.frc_cntr_val[32] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold2434 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[29] ),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold2435 (.A(\fpga_top.cpu_top.csr_mepc_ex[21] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold2436 (.A(\fpga_top.qspi_if.read_latency_0[1] ),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold2437 (.A(\fpga_top.qspi_if.wrcmd1[1] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold2438 (.A(\fpga_top.cpu_top.register_file.rf_1r1w.ram[18][22] ),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold2439 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[16] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold2440 (.A(_01463_),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold2441 (.A(\fpga_top.io_frc.frc_cmp_val[38] ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold2442 (.A(\fpga_top.io_frc.frc_cntr_val[20] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold2443 (.A(_00416_),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold2444 (.A(\fpga_top.io_frc.frc_cmp_val[1] ),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold2445 (.A(\fpga_top.io_frc.frc_cmp_val[28] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold2446 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram[2][2] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold2447 (.A(_02183_),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold2448 (.A(\fpga_top.qspi_if.qspi_state[8] ),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold2449 (.A(_00023_),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold2450 (.A(\fpga_top.qspi_if.wrcmd0[6] ),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold2451 (.A(\fpga_top.qspi_if.sio_in_sync[1] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold2452 (.A(_00958_),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold2453 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[22] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold2454 (.A(\fpga_top.io_frc.frc_cmp_val[33] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold2455 (.A(\fpga_top.io_frc.frc_cmp_val[16] ),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold2456 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mpp[0] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold2457 (.A(\fpga_top.uart_top.uart_logics.data_0[29] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold2458 (.A(\fpga_top.qspi_if.rdwrch[0] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold2459 (.A(\fpga_top.qspi_if.dbg_reg_2div_cec_write ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold2460 (.A(\fpga_top.io_frc.frc_cntr_val[49] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold2461 (.A(_02129_),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold2462 (.A(\fpga_top.qspi_if.sck_cntr[4] ),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold2463 (.A(_09261_),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold2464 (.A(\fpga_top.cpu_start_adr[8] ),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold2465 (.A(\fpga_top.cpu_top.execution.csr_array.pc_excep2[22] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold2466 (.A(_01469_),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold2467 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mcause[2] ),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold2468 (.A(_01940_),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold2469 (.A(\fpga_top.uart_top.uart_if.sample_cntr[1] ),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold2470 (.A(_09302_),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold2471 (.A(\fpga_top.qspi_if.rdcmd1[7] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold2472 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[5] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold2473 (.A(\fpga_top.io_frc.frc_cmp_val[26] ),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold2474 (.A(\fpga_top.qspi_if.rst_cntr[2] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold2475 (.A(_01105_),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold2476 (.A(\fpga_top.qspi_if.word_data[7] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold2477 (.A(_00964_),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold2478 (.A(\fpga_top.io_spi_lite.spi_sck_div[0] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold2479 (.A(\fpga_top.qspi_if.read_latency_1[3] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold2480 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[20] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold2481 (.A(\fpga_top.qspi_if.wrcmd1[6] ),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold2482 (.A(\fpga_top.qspi_if.wrcmd0[2] ),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold2483 (.A(\fpga_top.io_spi_lite.sck_div[1] ),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold2484 (.A(\fpga_top.uart_top.uart_rec_char.data_word[0] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold2485 (.A(_01239_),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold2486 (.A(\fpga_top.io_frc.frc_cmp_val[17] ),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold2487 (.A(_00103_),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold2488 (.A(_00110_),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold2489 (.A(\fpga_top.io_frc.frc_cntr_val[19] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold2490 (.A(_00415_),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold2491 (.A(\fpga_top.io_uart_out.uart_io_char[1] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold2492 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[6] ),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold2493 (.A(\fpga_top.dbg_bpoint_en[2] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold2494 (.A(\fpga_top.io_frc.frc_cmp_val[50] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold2495 (.A(\fpga_top.io_uart_out.rx_data_latch[2] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold2496 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[20] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold2497 (.A(\fpga_top.uart_top.uart_logics.data_0[6] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold2498 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[24] ),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold2499 (.A(\fpga_top.qspi_if.rdwrch[1] ),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold2500 (.A(\fpga_top.io_frc.frc_cmp_val[19] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold2501 (.A(\fpga_top.io_uart_out.rx_data_latch[3] ),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold2502 (.A(_00386_),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold2503 (.A(\fpga_top.io_frc.frc_cmp_val[13] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold2504 (.A(\fpga_top.qspi_if.read_latency_1[1] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold2505 (.A(\fpga_top.qspi_if.read_latency_1[2] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold2506 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[13] ),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold2507 (.A(\fpga_top.io_frc.frc_cntr_val[40] ),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold2508 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[4] ),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold2509 (.A(_01340_),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold2510 (.A(\fpga_top.io_frc.frc_cntr_val[21] ),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold2511 (.A(_00106_),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold2512 (.A(\fpga_top.io_frc.frc_cmp_val[37] ),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold2513 (.A(\fpga_top.io_spi_lite.spi_state[1] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold2514 (.A(_00192_),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold2515 (.A(\fpga_top.io_spi_lite.spi_mode[6] ),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold2516 (.A(_00099_),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold2517 (.A(\fpga_top.io_led.led_value[2] ),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold2518 (.A(\fpga_top.qspi_if.read_latency_1[0] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold2519 (.A(\fpga_top.uart_top.uart_logics.cmd_read_end[27] ),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold2520 (.A(_01363_),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold2521 (.A(\fpga_top.io_frc.frc_cntr_val[54] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold2522 (.A(\fpga_top.io_frc.frc_cmp_val[27] ),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold2523 (.A(\fpga_top.qspi_if.word_data[8] ),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold2524 (.A(\fpga_top.io_uart_out.uart_term[0] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold2525 (.A(\fpga_top.dbg_bpoint_en[1] ),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold2526 (.A(\fpga_top.qspi_if.rdcmd0[2] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold2527 (.A(\fpga_top.io_spi_lite.miso_byte_org[6] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold2528 (.A(_10551_),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold2529 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[24] ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold2530 (.A(_02066_),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold2531 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mstatush[25] ),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold2532 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[7] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold2533 (.A(\fpga_top.io_spi_lite.spi_sck_div[5] ),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold2534 (.A(\fpga_top.io_frc.frc_cmp_val[3] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold2535 (.A(_00094_),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold2536 (.A(\fpga_top.io_frc.frc_cmp_val[29] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold2537 (.A(\fpga_top.bus_gather.u_read_adr[3] ),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold2538 (.A(_01402_),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold2539 (.A(\fpga_top.qspi_if.sck_div[8] ),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold2540 (.A(\fpga_top.io_uart_out.uart_io_char[3] ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold2541 (.A(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[1] ),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold2542 (.A(\fpga_top.uart_top.uart_logics.data_0[19] ),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold2543 (.A(\fpga_top.qspi_if.sck_div[3] ),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold2544 (.A(\fpga_top.io_frc.frc_cmp_val[10] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold2545 (.A(\fpga_top.qspi_if.sck_cntr[7] ),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold2546 (.A(_09265_),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold2547 (.A(\fpga_top.io_frc.frc_cmp_val[58] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold2548 (.A(\fpga_top.io_frc.frc_cntr_val[27] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold2549 (.A(_00423_),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold2550 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[0] ),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold2551 (.A(_09641_),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold2552 (.A(_00026_),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold2553 (.A(\fpga_top.uart_top.uart_if.sample_cntr[15] ),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold2554 (.A(_09333_),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold2555 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[11] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold2556 (.A(\fpga_top.qspi_if.rst_cntr[0] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold2557 (.A(\fpga_top.io_spi_lite.sck_div[4] ),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold2558 (.A(_08956_),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold2559 (.A(_00032_),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold2560 (.A(\fpga_top.io_spi_lite.sck_div[5] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold2561 (.A(_08958_),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold2562 (.A(\fpga_top.qspi_if.wdata[31] ),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold2563 (.A(_00954_),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold2564 (.A(\fpga_top.io_spi_lite.sck_div[6] ),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold2565 (.A(\fpga_top.qspi_if.word_data[6] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold2566 (.A(_00963_),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold2567 (.A(\fpga_top.io_uart_out.uart_io_char[4] ),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold2568 (.A(\fpga_top.io_frc.frc_cmp_val[21] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold2569 (.A(\fpga_top.io_uart_out.rx_data_latch[1] ),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold2570 (.A(_00384_),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold2571 (.A(\fpga_top.uart_top.uart_rec_char.pdata[0] ),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold2572 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[20] ),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold2573 (.A(_02062_),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold2574 (.A(\fpga_top.qspi_if.read_latency_2[0] ),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold2575 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[1] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold2576 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[8] ),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold2577 (.A(\fpga_top.qspi_if.rdcmd1[4] ),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold2578 (.A(\fpga_top.io_spi_lite.spi_mode[8] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold2579 (.A(\fpga_top.io_spi_lite.sck_div[8] ),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold2580 (.A(\fpga_top.cpu_top.register_file.rfr_state[0] ),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold2581 (.A(_09444_),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold2582 (.A(\fpga_top.cpu_top.register_file.next_rfr_state[2] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold2583 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[0] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold2584 (.A(\fpga_top.qspi_if.qspi_state[6] ),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold2585 (.A(_08933_),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold2586 (.A(_00018_),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold2587 (.A(\fpga_top.bus_gather.u_read_adr[23] ),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold2588 (.A(\fpga_top.io_frc.frc_cntr_val[15] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold2589 (.A(_00411_),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold2590 (.A(\fpga_top.io_frc.frc_cntr_val[39] ),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold2591 (.A(_00113_),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold2592 (.A(\fpga_top.qspi_if.sck_div[4] ),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold2593 (.A(\fpga_top.io_spi_lite.spi_sck_div[6] ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold2594 (.A(\fpga_top.io_spi_lite.spi_sck_div[2] ),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold2595 (.A(\fpga_top.bus_gather.u_read_adr[28] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold2596 (.A(\fpga_top.qspi_if.rdcmd0[4] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold2597 (.A(\fpga_top.qspi_if.read_cntr[1] ),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold2598 (.A(_01016_),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold2599 (.A(\fpga_top.qspi_if.read_latency_0[0] ),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold2600 (.A(\fpga_top.io_uart_out.rout[1] ),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold2601 (.A(_01331_),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold2602 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[26] ),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold2603 (.A(\fpga_top.qspi_if.read_latency_2[3] ),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold2604 (.A(\fpga_top.uart_top.uart_rec_char.pdata[3] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold2605 (.A(_01333_),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold2606 (.A(\fpga_top.cpu_start_adr[27] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold2607 (.A(\fpga_top.io_spi_lite.spi_sck_div[1] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold2608 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[1] ),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold2609 (.A(\fpga_top.io_frc.frc_cntr_val[60] ),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold2610 (.A(_02140_),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold2611 (.A(\fpga_top.io_uart_out.rx_data_latch[4] ),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold2612 (.A(\fpga_top.qspi_if.qspi_state[2] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold2613 (.A(_09097_),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold2614 (.A(\fpga_top.uart_top.uart_if.rx_state[2] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold2615 (.A(_09522_),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold2616 (.A(\fpga_top.io_frc.frc_cntr_val[2] ),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold2617 (.A(\fpga_top.io_spi_lite.spi_sck_div[4] ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold2618 (.A(\fpga_top.uart_top.uart_if.sample_cntr[0] ),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold2619 (.A(\fpga_top.qspi_if.wrcmd1[0] ),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold2620 (.A(\fpga_top.cpu_top.data_rw_mem.data_state[2] ),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold2621 (.A(\fpga_top.cpu_top.data_rw_mem.next_data_state[2] ),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold2622 (.A(_00112_),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold2623 (.A(\fpga_top.cpu_top.csr_wadr_mon[5] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold2624 (.A(\fpga_top.cpu_top.br_ofs[3] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold2625 (.A(\fpga_top.cpu_top.br_ofs[4] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold2626 (.A(_00127_),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold2627 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[17] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold2628 (.A(_02059_),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold2629 (.A(\fpga_top.io_frc.frc_cmp_val[30] ),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold2630 (.A(\fpga_top.qspi_if.read_cntr[0] ),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold2631 (.A(\fpga_top.bus_gather.u_read_adr[27] ),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold2632 (.A(\fpga_top.uart_top.uart_if.tx_out_cntr[2] ),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold2633 (.A(\fpga_top.qspi_if.read_latency_2[2] ),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold2634 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[18] ),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold2635 (.A(\fpga_top.io_frc.frc_cntr_val[18] ),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold2636 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[13] ),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold2637 (.A(_02055_),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold2638 (.A(\fpga_top.cpu_start_adr[21] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold2639 (.A(\fpga_top.qspi_if.sck_cntr[1] ),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold2640 (.A(\fpga_top.bus_gather.u_read_adr[26] ),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold2641 (.A(_01425_),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold2642 (.A(\fpga_top.qspi_if.sck_cntr[8] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold2643 (.A(_09267_),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold2644 (.A(\fpga_top.io_uart_out.rout[3] ),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold2645 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[4] ),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold2646 (.A(_01270_),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold2647 (.A(\fpga_top.qspi_if.read_latency_2[1] ),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold2648 (.A(\fpga_top.qspi_if.wdata[21] ),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold2649 (.A(_00944_),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold2650 (.A(\fpga_top.io_frc.frc_cmp_val[36] ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold2651 (.A(\fpga_top.io_uart_out.uart_term[8] ),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold2652 (.A(_00082_),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold2653 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[27] ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold2654 (.A(\fpga_top.interrupter.int0_3lat ),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold2655 (.A(_02732_),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold2656 (.A(_00291_),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold2657 (.A(\fpga_top.io_frc.frc_cntr_val[35] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold2658 (.A(_02115_),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold2659 (.A(\fpga_top.io_uart_out.uart_term[4] ),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold2660 (.A(_00061_),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold2661 (.A(_00125_),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold2662 (.A(_08924_),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold2663 (.A(_00021_),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold2664 (.A(\fpga_top.qspi_if.qspi_state[11] ),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold2665 (.A(_08871_),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold2666 (.A(\fpga_top.io_frc.frc_cmp_val[4] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold2667 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[30] ),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold2668 (.A(_01232_),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold2669 (.A(\fpga_top.qspi_if.wdata[27] ),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold2670 (.A(_00950_),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold2671 (.A(\fpga_top.uart_top.uart_rec_char.pdata[5] ),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold2672 (.A(_01335_),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold2673 (.A(\fpga_top.io_spi_lite.spi_sck_div[3] ),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold2674 (.A(\fpga_top.io_uart_out.uart_term[10] ),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold2675 (.A(_00069_),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold2676 (.A(\fpga_top.qspi_if.wdata[22] ),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold2677 (.A(_03231_),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold2678 (.A(_00945_),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold2679 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[4] ),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold2680 (.A(\fpga_top.uart_top.uart_if.sample_cntr[8] ),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold2681 (.A(_09317_),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold2682 (.A(_09318_),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold2683 (.A(_00066_),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold2684 (.A(\fpga_top.uart_top.uart_logics.rdata_snd_wait_dly ),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold2685 (.A(_02147_),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold2686 (.A(\fpga_top.qspi_if.sck_cntr[5] ),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold2687 (.A(\fpga_top.io_spi_lite.sck_div[3] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold2688 (.A(\fpga_top.io_uart_out.rout[5] ),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold2689 (.A(_02218_),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold2690 (.A(\fpga_top.io_frc.frc_cntr_val[37] ),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold2691 (.A(\fpga_top.io_frc.frc_cntr_val[24] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold2692 (.A(_00420_),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold2693 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[27] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold2694 (.A(_01229_),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold2695 (.A(\fpga_top.io_frc.frc_cntr_val[45] ),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold2696 (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[4] ),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold2697 (.A(_09366_),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold2698 (.A(\fpga_top.io_led.dbg_smpl_trgsig ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold2699 (.A(_00391_),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold2700 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[9] ),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold2701 (.A(_02051_),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold2702 (.A(\fpga_top.io_frc.frc_cntr_val[10] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold2703 (.A(_00406_),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold2704 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[16] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold2705 (.A(_02058_),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold2706 (.A(\fpga_top.uart_top.uart_rec_char.pdata[6] ),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold2707 (.A(_01336_),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold2708 (.A(\fpga_top.io_uart_out.uart_term[12] ),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold2709 (.A(_00071_),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold2710 (.A(\fpga_top.io_frc.frc_cmp_val[35] ),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold2711 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[21] ),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold2712 (.A(\fpga_top.uart_top.uart_if.sample_cntr[4] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold2713 (.A(_09309_),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold2714 (.A(\fpga_top.io_frc.frc_cntr_val[9] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold2715 (.A(_00405_),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold2716 (.A(\fpga_top.qspi_if.wdata[19] ),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold2717 (.A(_03228_),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold2718 (.A(_00942_),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold2719 (.A(\fpga_top.uart_top.uart_rec_char.pdata[7] ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold2720 (.A(_01337_),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold2721 (.A(\fpga_top.cpu_top.csr_wadr_mon[10] ),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold2722 (.A(_04291_),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold2723 (.A(_01214_),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold2724 (.A(\fpga_top.bus_gather.d_write_data[20] ),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold2725 (.A(\fpga_top.io_frc.frc_cntr_val[16] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold2726 (.A(\fpga_top.io_frc.frc_cntr_val[26] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold2727 (.A(_00422_),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold2728 (.A(\fpga_top.cpu_top.br_ofs[11] ),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold2729 (.A(\fpga_top.io_uart_out.uart_term[13] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold2730 (.A(_00072_),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold2731 (.A(\fpga_top.uart_top.uart_rec_char.bpoint[5] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold2732 (.A(_01271_),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold2733 (.A(\fpga_top.io_frc.frc_cntr_val[48] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold2734 (.A(\fpga_top.io_frc.frc_cntr_val[57] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold2735 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[26] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold2736 (.A(_01228_),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold2737 (.A(\fpga_top.io_frc.frc_cntr_val[14] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold2738 (.A(\fpga_top.io_frc.frc_cntr_val[11] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold2739 (.A(\fpga_top.qspi_if.wdata[4] ),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold2740 (.A(_03208_),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold2741 (.A(\fpga_top.io_frc.frc_cntr_val[30] ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold2742 (.A(\fpga_top.qspi_if.sck_div[9] ),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold2743 (.A(\fpga_top.cpu_top.pc_stage.pc_int_ecall_syn_state ),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold2744 (.A(\fpga_top.qspi_if.wdata[23] ),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold2745 (.A(_03232_),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold2746 (.A(_00946_),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold2747 (.A(\fpga_top.io_frc.frc_cntr_val[6] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold2748 (.A(\fpga_top.qspi_if.wdata[26] ),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold2749 (.A(_03235_),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold2750 (.A(_00949_),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold2751 (.A(\fpga_top.io_frc.frc_cntr_val[51] ),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold2752 (.A(_06186_),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold2753 (.A(\fpga_top.qspi_if.read_cntr[2] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold2754 (.A(_03508_),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold2755 (.A(\fpga_top.uart_top.uart_logics.data_0[0] ),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold2756 (.A(\fpga_top.qspi_if.wdata[28] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold2757 (.A(_00951_),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold2758 (.A(\fpga_top.io_frc.frc_cntr_val[22] ),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold2759 (.A(\fpga_top.bus_gather.d_write_data[28] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold2760 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[29] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold2761 (.A(_01231_),
    .X(net6079));
 sg13g2_dlygate4sd3_1 hold2762 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[3] ),
    .X(net6080));
 sg13g2_dlygate4sd3_1 hold2763 (.A(_02045_),
    .X(net6081));
 sg13g2_dlygate4sd3_1 hold2764 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[23] ),
    .X(net6082));
 sg13g2_dlygate4sd3_1 hold2765 (.A(_01225_),
    .X(net6083));
 sg13g2_dlygate4sd3_1 hold2766 (.A(\fpga_top.io_spi_lite.sck_div[9] ),
    .X(net6084));
 sg13g2_dlygate4sd3_1 hold2767 (.A(\fpga_top.io_spi_lite.spi_mode[12] ),
    .X(net6085));
 sg13g2_dlygate4sd3_1 hold2768 (.A(\fpga_top.io_frc.frc_cntr_val[31] ),
    .X(net6086));
 sg13g2_dlygate4sd3_1 hold2769 (.A(_00427_),
    .X(net6087));
 sg13g2_dlygate4sd3_1 hold2770 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[15] ),
    .X(net6088));
 sg13g2_dlygate4sd3_1 hold2771 (.A(\fpga_top.io_spi_lite.spi_mode[0] ),
    .X(net6089));
 sg13g2_dlygate4sd3_1 hold2772 (.A(\fpga_top.cpu_top.br_ofs[2] ),
    .X(net6090));
 sg13g2_dlygate4sd3_1 hold2773 (.A(\fpga_top.uart_top.uart_rec_char.bpoint_ld ),
    .X(net6091));
 sg13g2_dlygate4sd3_1 hold2774 (.A(_04358_),
    .X(net6092));
 sg13g2_dlygate4sd3_1 hold2775 (.A(\fpga_top.cpu_top.csr_uimm[1] ),
    .X(net6093));
 sg13g2_dlygate4sd3_1 hold2776 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[18] ),
    .X(net6094));
 sg13g2_dlygate4sd3_1 hold2777 (.A(_04313_),
    .X(net6095));
 sg13g2_dlygate4sd3_1 hold2778 (.A(_01220_),
    .X(net6096));
 sg13g2_dlygate4sd3_1 hold2779 (.A(\fpga_top.uart_top.uart_logics.data_0[27] ),
    .X(net6097));
 sg13g2_dlygate4sd3_1 hold2780 (.A(\fpga_top.cpu_start_adr[5] ),
    .X(net6098));
 sg13g2_dlygate4sd3_1 hold2781 (.A(\fpga_top.qspi_if.rdedge[2] ),
    .X(net6099));
 sg13g2_dlygate4sd3_1 hold2782 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[12] ),
    .X(net6100));
 sg13g2_dlygate4sd3_1 hold2783 (.A(\fpga_top.io_frc.frc_cmp_val[42] ),
    .X(net6101));
 sg13g2_dlygate4sd3_1 hold2784 (.A(\fpga_top.io_frc.frc_cntr_val[56] ),
    .X(net6102));
 sg13g2_dlygate4sd3_1 hold2785 (.A(\fpga_top.qspi_if.wdata[24] ),
    .X(net6103));
 sg13g2_dlygate4sd3_1 hold2786 (.A(_03233_),
    .X(net6104));
 sg13g2_dlygate4sd3_1 hold2787 (.A(_00947_),
    .X(net6105));
 sg13g2_dlygate4sd3_1 hold2788 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[22] ),
    .X(net6106));
 sg13g2_dlygate4sd3_1 hold2789 (.A(_02064_),
    .X(net6107));
 sg13g2_dlygate4sd3_1 hold2790 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[22] ),
    .X(net6108));
 sg13g2_dlygate4sd3_1 hold2791 (.A(_04325_),
    .X(net6109));
 sg13g2_dlygate4sd3_1 hold2792 (.A(_01224_),
    .X(net6110));
 sg13g2_dlygate4sd3_1 hold2793 (.A(\fpga_top.io_uart_out.uart_term[14] ),
    .X(net6111));
 sg13g2_dlygate4sd3_1 hold2794 (.A(_00073_),
    .X(net6112));
 sg13g2_dlygate4sd3_1 hold2795 (.A(\fpga_top.qspi_if.wdata[30] ),
    .X(net6113));
 sg13g2_dlygate4sd3_1 hold2796 (.A(_00953_),
    .X(net6114));
 sg13g2_dlygate4sd3_1 hold2797 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[21] ),
    .X(net6115));
 sg13g2_dlygate4sd3_1 hold2798 (.A(_01223_),
    .X(net6116));
 sg13g2_dlygate4sd3_1 hold2799 (.A(\fpga_top.uart_top.uart_if.tx_fifo_dcntr[3] ),
    .X(net6117));
 sg13g2_dlygate4sd3_1 hold2800 (.A(_03653_),
    .X(net6118));
 sg13g2_dlygate4sd3_1 hold2801 (.A(\fpga_top.bus_gather.u_read_adr[9] ),
    .X(net6119));
 sg13g2_dlygate4sd3_1 hold2802 (.A(_04693_),
    .X(net6120));
 sg13g2_dlygate4sd3_1 hold2803 (.A(_01408_),
    .X(net6121));
 sg13g2_dlygate4sd3_1 hold2804 (.A(\fpga_top.uart_top.uart_if.sample_cntr[6] ),
    .X(net6122));
 sg13g2_dlygate4sd3_1 hold2805 (.A(_09313_),
    .X(net6123));
 sg13g2_dlygate4sd3_1 hold2806 (.A(\fpga_top.bus_gather.d_write_data[9] ),
    .X(net6124));
 sg13g2_dlygate4sd3_1 hold2807 (.A(\fpga_top.bus_gather.d_write_data[16] ),
    .X(net6125));
 sg13g2_dlygate4sd3_1 hold2808 (.A(\fpga_top.qspi_if.wdata[18] ),
    .X(net6126));
 sg13g2_dlygate4sd3_1 hold2809 (.A(_03227_),
    .X(net6127));
 sg13g2_dlygate4sd3_1 hold2810 (.A(_00941_),
    .X(net6128));
 sg13g2_dlygate4sd3_1 hold2811 (.A(\fpga_top.io_frc.frc_cntr_val[8] ),
    .X(net6129));
 sg13g2_dlygate4sd3_1 hold2812 (.A(\fpga_top.qspi_if.adr_rw[13] ),
    .X(net6130));
 sg13g2_dlygate4sd3_1 hold2813 (.A(_01002_),
    .X(net6131));
 sg13g2_dlygate4sd3_1 hold2814 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[29] ),
    .X(net6132));
 sg13g2_dlygate4sd3_1 hold2815 (.A(\fpga_top.io_frc.frc_cntr_val[55] ),
    .X(net6133));
 sg13g2_dlygate4sd3_1 hold2816 (.A(\fpga_top.qspi_if.wdata[1] ),
    .X(net6134));
 sg13g2_dlygate4sd3_1 hold2817 (.A(_03204_),
    .X(net6135));
 sg13g2_dlygate4sd3_1 hold2818 (.A(\fpga_top.io_frc.frc_cntr_val[29] ),
    .X(net6136));
 sg13g2_dlygate4sd3_1 hold2819 (.A(_00425_),
    .X(net6137));
 sg13g2_dlygate4sd3_1 hold2820 (.A(\fpga_top.qspi_if.wdata[15] ),
    .X(net6138));
 sg13g2_dlygate4sd3_1 hold2821 (.A(_03224_),
    .X(net6139));
 sg13g2_dlygate4sd3_1 hold2822 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[19] ),
    .X(net6140));
 sg13g2_dlygate4sd3_1 hold2823 (.A(_04316_),
    .X(net6141));
 sg13g2_dlygate4sd3_1 hold2824 (.A(_01221_),
    .X(net6142));
 sg13g2_dlygate4sd3_1 hold2825 (.A(\fpga_top.io_frc.frc_cntr_val[0] ),
    .X(net6143));
 sg13g2_dlygate4sd3_1 hold2826 (.A(\fpga_top.qspi_if.wdata[25] ),
    .X(net6144));
 sg13g2_dlygate4sd3_1 hold2827 (.A(_03234_),
    .X(net6145));
 sg13g2_dlygate4sd3_1 hold2828 (.A(_00948_),
    .X(net6146));
 sg13g2_dlygate4sd3_1 hold2829 (.A(\fpga_top.io_uart_out.uart_term[15] ),
    .X(net6147));
 sg13g2_dlygate4sd3_1 hold2830 (.A(_00057_),
    .X(net6148));
 sg13g2_dlygate4sd3_1 hold2831 (.A(\fpga_top.bus_gather.u_read_adr[7] ),
    .X(net6149));
 sg13g2_dlygate4sd3_1 hold2832 (.A(_01406_),
    .X(net6150));
 sg13g2_dlygate4sd3_1 hold2833 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[16] ),
    .X(net6151));
 sg13g2_dlygate4sd3_1 hold2834 (.A(_01218_),
    .X(net6152));
 sg13g2_dlygate4sd3_1 hold2835 (.A(\fpga_top.qspi_if.qspi_state[4] ),
    .X(net6153));
 sg13g2_dlygate4sd3_1 hold2836 (.A(_08917_),
    .X(net6154));
 sg13g2_dlygate4sd3_1 hold2837 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[31] ),
    .X(net6155));
 sg13g2_dlygate4sd3_1 hold2838 (.A(\fpga_top.bus_gather.d_write_data[19] ),
    .X(net6156));
 sg13g2_dlygate4sd3_1 hold2839 (.A(\fpga_top.qspi_if.adr_ofs[1] ),
    .X(net6157));
 sg13g2_dlygate4sd3_1 hold2840 (.A(_03627_),
    .X(net6158));
 sg13g2_dlygate4sd3_1 hold2841 (.A(_01101_),
    .X(net6159));
 sg13g2_dlygate4sd3_1 hold2842 (.A(\fpga_top.qspi_if.wdata[3] ),
    .X(net6160));
 sg13g2_dlygate4sd3_1 hold2843 (.A(_03207_),
    .X(net6161));
 sg13g2_dlygate4sd3_1 hold2844 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[24] ),
    .X(net6162));
 sg13g2_dlygate4sd3_1 hold2845 (.A(_04332_),
    .X(net6163));
 sg13g2_dlygate4sd3_1 hold2846 (.A(_01226_),
    .X(net6164));
 sg13g2_dlygate4sd3_1 hold2847 (.A(\fpga_top.io_frc.frc_cntr_val[23] ),
    .X(net6165));
 sg13g2_dlygate4sd3_1 hold2848 (.A(\fpga_top.uart_top.uart_if.tx_cycle_cntr[11] ),
    .X(net6166));
 sg13g2_dlygate4sd3_1 hold2849 (.A(_09382_),
    .X(net6167));
 sg13g2_dlygate4sd3_1 hold2850 (.A(_00070_),
    .X(net6168));
 sg13g2_dlygate4sd3_1 hold2851 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[17] ),
    .X(net6169));
 sg13g2_dlygate4sd3_1 hold2852 (.A(_01219_),
    .X(net6170));
 sg13g2_dlygate4sd3_1 hold2853 (.A(\fpga_top.uart_top.uart_if.sample_cntr[13] ),
    .X(net6171));
 sg13g2_dlygate4sd3_1 hold2854 (.A(_09328_),
    .X(net6172));
 sg13g2_dlygate4sd3_1 hold2855 (.A(_09329_),
    .X(net6173));
 sg13g2_dlygate4sd3_1 hold2856 (.A(\fpga_top.io_uart_out.uart_term[11] ),
    .X(net6174));
 sg13g2_dlygate4sd3_1 hold2857 (.A(_09325_),
    .X(net6175));
 sg13g2_dlygate4sd3_1 hold2858 (.A(_00054_),
    .X(net6176));
 sg13g2_dlygate4sd3_1 hold2859 (.A(\fpga_top.qspi_if.wdata[29] ),
    .X(net6177));
 sg13g2_dlygate4sd3_1 hold2860 (.A(_00952_),
    .X(net6178));
 sg13g2_dlygate4sd3_1 hold2861 (.A(\fpga_top.io_frc.frc_cntr_val[3] ),
    .X(net6179));
 sg13g2_dlygate4sd3_1 hold2862 (.A(_00399_),
    .X(net6180));
 sg13g2_dlygate4sd3_1 hold2863 (.A(\fpga_top.io_frc.frc_cntr_val[25] ),
    .X(net6181));
 sg13g2_dlygate4sd3_1 hold2864 (.A(_00421_),
    .X(net6182));
 sg13g2_dlygate4sd3_1 hold2865 (.A(\fpga_top.qspi_if.wdata[14] ),
    .X(net6183));
 sg13g2_dlygate4sd3_1 hold2866 (.A(_03223_),
    .X(net6184));
 sg13g2_dlygate4sd3_1 hold2867 (.A(_00937_),
    .X(net6185));
 sg13g2_dlygate4sd3_1 hold2868 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[20] ),
    .X(net6186));
 sg13g2_dlygate4sd3_1 hold2869 (.A(\fpga_top.qspi_if.wdata[20] ),
    .X(net6187));
 sg13g2_dlygate4sd3_1 hold2870 (.A(\fpga_top.uart_top.uart_if.rx_state[0] ),
    .X(net6188));
 sg13g2_dlygate4sd3_1 hold2871 (.A(_09524_),
    .X(net6189));
 sg13g2_dlygate4sd3_1 hold2872 (.A(\fpga_top.uart_top.uart_if.next_rx_state[0] ),
    .X(net6190));
 sg13g2_dlygate4sd3_1 hold2873 (.A(\fpga_top.qspi_if.wdata[10] ),
    .X(net6191));
 sg13g2_dlygate4sd3_1 hold2874 (.A(\fpga_top.io_spi_lite.spi_state[0] ),
    .X(net6192));
 sg13g2_dlygate4sd3_1 hold2875 (.A(_00191_),
    .X(net6193));
 sg13g2_dlygate4sd3_1 hold2876 (.A(\fpga_top.qspi_if.dbg_2div_read_half_end ),
    .X(net6194));
 sg13g2_dlygate4sd3_1 hold2877 (.A(\fpga_top.qspi_if.wdata_ofs[1] ),
    .X(net6195));
 sg13g2_dlygate4sd3_1 hold2878 (.A(_03569_),
    .X(net6196));
 sg13g2_dlygate4sd3_1 hold2879 (.A(\fpga_top.io_frc.frc_cntr_val[7] ),
    .X(net6197));
 sg13g2_dlygate4sd3_1 hold2880 (.A(_00403_),
    .X(net6198));
 sg13g2_dlygate4sd3_1 hold2881 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[14] ),
    .X(net6199));
 sg13g2_dlygate4sd3_1 hold2882 (.A(_02056_),
    .X(net6200));
 sg13g2_dlygate4sd3_1 hold2883 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[23] ),
    .X(net6201));
 sg13g2_dlygate4sd3_1 hold2884 (.A(_02065_),
    .X(net6202));
 sg13g2_dlygate4sd3_1 hold2885 (.A(\fpga_top.io_frc.frc_cntrl_val ),
    .X(net6203));
 sg13g2_dlygate4sd3_1 hold2886 (.A(\fpga_top.bus_gather.d_write_data[22] ),
    .X(net6204));
 sg13g2_dlygate4sd3_1 hold2887 (.A(\fpga_top.qspi_if.sck_cntr[9] ),
    .X(net6205));
 sg13g2_dlygate4sd3_1 hold2888 (.A(\fpga_top.uart_top.uart_if.sample_cntr[10] ),
    .X(net6206));
 sg13g2_dlygate4sd3_1 hold2889 (.A(_09322_),
    .X(net6207));
 sg13g2_dlygate4sd3_1 hold2890 (.A(_09323_),
    .X(net6208));
 sg13g2_dlygate4sd3_1 hold2891 (.A(_00053_),
    .X(net6209));
 sg13g2_dlygate4sd3_1 hold2892 (.A(\fpga_top.qspi_if.dbg_2div_trt ),
    .X(net6210));
 sg13g2_dlygate4sd3_1 hold2893 (.A(\fpga_top.cpu_top.csr_uimm[2] ),
    .X(net6211));
 sg13g2_dlygate4sd3_1 hold2894 (.A(\fpga_top.cpu_top.csr_mtie ),
    .X(net6212));
 sg13g2_dlygate4sd3_1 hold2895 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[25] ),
    .X(net6213));
 sg13g2_dlygate4sd3_1 hold2896 (.A(\fpga_top.bus_gather.u_read_adr[11] ),
    .X(net6214));
 sg13g2_dlygate4sd3_1 hold2897 (.A(_04703_),
    .X(net6215));
 sg13g2_dlygate4sd3_1 hold2898 (.A(\fpga_top.uart_top.uart_if.sample_cntr[5] ),
    .X(net6216));
 sg13g2_dlygate4sd3_1 hold2899 (.A(\fpga_top.cpu_top.csr_uimm[0] ),
    .X(net6217));
 sg13g2_dlygate4sd3_1 hold2900 (.A(\fpga_top.bus_gather.d_write_data[2] ),
    .X(net6218));
 sg13g2_dlygate4sd3_1 hold2901 (.A(\fpga_top.cpu_top.register_file.rfr_state[2] ),
    .X(net6219));
 sg13g2_dlygate4sd3_1 hold2902 (.A(_09442_),
    .X(net6220));
 sg13g2_dlygate4sd3_1 hold2903 (.A(\fpga_top.cpu_top.register_file.next_rfr_state[0] ),
    .X(net6221));
 sg13g2_dlygate4sd3_1 hold2904 (.A(\fpga_top.qspi_if.wdata[17] ),
    .X(net6222));
 sg13g2_dlygate4sd3_1 hold2905 (.A(_00940_),
    .X(net6223));
 sg13g2_dlygate4sd3_1 hold2906 (.A(\fpga_top.bus_gather.u_read_adr[15] ),
    .X(net6224));
 sg13g2_dlygate4sd3_1 hold2907 (.A(_04714_),
    .X(net6225));
 sg13g2_dlygate4sd3_1 hold2908 (.A(_01414_),
    .X(net6226));
 sg13g2_dlygate4sd3_1 hold2909 (.A(\fpga_top.qspi_if.wdata[0] ),
    .X(net6227));
 sg13g2_dlygate4sd3_1 hold2910 (.A(_03203_),
    .X(net6228));
 sg13g2_dlygate4sd3_1 hold2911 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[10] ),
    .X(net6229));
 sg13g2_dlygate4sd3_1 hold2912 (.A(\fpga_top.qspi_if.wdata[5] ),
    .X(net6230));
 sg13g2_dlygate4sd3_1 hold2913 (.A(\fpga_top.bus_gather.u_read_adr[16] ),
    .X(net6231));
 sg13g2_dlygate4sd3_1 hold2914 (.A(_01415_),
    .X(net6232));
 sg13g2_dlygate4sd3_1 hold2915 (.A(\fpga_top.bus_gather.u_read_adr[22] ),
    .X(net6233));
 sg13g2_dlygate4sd3_1 hold2916 (.A(_01421_),
    .X(net6234));
 sg13g2_dlygate4sd3_1 hold2917 (.A(\fpga_top.qspi_if.wdata[13] ),
    .X(net6235));
 sg13g2_dlygate4sd3_1 hold2918 (.A(_03222_),
    .X(net6236));
 sg13g2_dlygate4sd3_1 hold2919 (.A(_00936_),
    .X(net6237));
 sg13g2_dlygate4sd3_1 hold2920 (.A(\fpga_top.cpu_top.csr_wadr_mon[9] ),
    .X(net6238));
 sg13g2_dlygate4sd3_1 hold2921 (.A(\fpga_top.bus_gather.u_read_adr[25] ),
    .X(net6239));
 sg13g2_dlygate4sd3_1 hold2922 (.A(_01424_),
    .X(net6240));
 sg13g2_dlygate4sd3_1 hold2923 (.A(\fpga_top.uart_top.uart_if.sample_cntr[7] ),
    .X(net6241));
 sg13g2_dlygate4sd3_1 hold2924 (.A(\fpga_top.bus_gather.d_write_data[7] ),
    .X(net6242));
 sg13g2_dlygate4sd3_1 hold2925 (.A(\fpga_top.qspi_if.wdata[12] ),
    .X(net6243));
 sg13g2_dlygate4sd3_1 hold2926 (.A(_03221_),
    .X(net6244));
 sg13g2_dlygate4sd3_1 hold2927 (.A(_00935_),
    .X(net6245));
 sg13g2_dlygate4sd3_1 hold2928 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[28] ),
    .X(net6246));
 sg13g2_dlygate4sd3_1 hold2929 (.A(\fpga_top.qspi_if.rwait_cntr[0] ),
    .X(net6247));
 sg13g2_dlygate4sd3_1 hold2930 (.A(\fpga_top.qspi_if.adr_rw[3] ),
    .X(net6248));
 sg13g2_dlygate4sd3_1 hold2931 (.A(_00992_),
    .X(net6249));
 sg13g2_dlygate4sd3_1 hold2932 (.A(\fpga_top.io_frc.frc_cntr_val[12] ),
    .X(net6250));
 sg13g2_dlygate4sd3_1 hold2933 (.A(\fpga_top.qspi_if.wdata[16] ),
    .X(net6251));
 sg13g2_dlygate4sd3_1 hold2934 (.A(_03225_),
    .X(net6252));
 sg13g2_dlygate4sd3_1 hold2935 (.A(\fpga_top.qspi_if.adr_rw[9] ),
    .X(net6253));
 sg13g2_dlygate4sd3_1 hold2936 (.A(_00998_),
    .X(net6254));
 sg13g2_dlygate4sd3_1 hold2937 (.A(\fpga_top.bus_gather.u_read_adr[17] ),
    .X(net6255));
 sg13g2_dlygate4sd3_1 hold2938 (.A(_01416_),
    .X(net6256));
 sg13g2_dlygate4sd3_1 hold2939 (.A(\fpga_top.bus_gather.u_read_adr[14] ),
    .X(net6257));
 sg13g2_dlygate4sd3_1 hold2940 (.A(_01413_),
    .X(net6258));
 sg13g2_dlygate4sd3_1 hold2941 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mpp[1] ),
    .X(net6259));
 sg13g2_dlygate4sd3_1 hold2942 (.A(_05877_),
    .X(net6260));
 sg13g2_dlygate4sd3_1 hold2943 (.A(\fpga_top.qspi_if.adr_rw[16] ),
    .X(net6261));
 sg13g2_dlygate4sd3_1 hold2944 (.A(\fpga_top.qspi_if.word_adr[25] ),
    .X(net6262));
 sg13g2_dlygate4sd3_1 hold2945 (.A(_00132_),
    .X(net6263));
 sg13g2_dlygate4sd3_1 hold2946 (.A(\fpga_top.bus_gather.u_read_adr[19] ),
    .X(net6264));
 sg13g2_dlygate4sd3_1 hold2947 (.A(_01418_),
    .X(net6265));
 sg13g2_dlygate4sd3_1 hold2948 (.A(\fpga_top.uart_top.uart_if.sample_cntr[2] ),
    .X(net6266));
 sg13g2_dlygate4sd3_1 hold2949 (.A(\fpga_top.qspi_if.adr_rw[7] ),
    .X(net6267));
 sg13g2_dlygate4sd3_1 hold2950 (.A(_00996_),
    .X(net6268));
 sg13g2_dlygate4sd3_1 hold2951 (.A(\fpga_top.bus_gather.d_write_data[31] ),
    .X(net6269));
 sg13g2_dlygate4sd3_1 hold2952 (.A(\fpga_top.bus_gather.d_write_data[26] ),
    .X(net6270));
 sg13g2_dlygate4sd3_1 hold2953 (.A(\fpga_top.qspi_if.adr_rw[14] ),
    .X(net6271));
 sg13g2_dlygate4sd3_1 hold2954 (.A(_01003_),
    .X(net6272));
 sg13g2_dlygate4sd3_1 hold2955 (.A(\fpga_top.io_frc.frc_cntr_val[17] ),
    .X(net6273));
 sg13g2_dlygate4sd3_1 hold2956 (.A(\fpga_top.cpu_top.csr_wadr_mon[11] ),
    .X(net6274));
 sg13g2_dlygate4sd3_1 hold2957 (.A(_01216_),
    .X(net6275));
 sg13g2_dlygate4sd3_1 hold2958 (.A(\fpga_top.bus_gather.d_write_data[17] ),
    .X(net6276));
 sg13g2_dlygate4sd3_1 hold2959 (.A(\fpga_top.qspi_if.adr_rw[4] ),
    .X(net6277));
 sg13g2_dlygate4sd3_1 hold2960 (.A(_00993_),
    .X(net6278));
 sg13g2_dlygate4sd3_1 hold2961 (.A(\fpga_top.uart_top.uart_logics.data_0[14] ),
    .X(net6279));
 sg13g2_dlygate4sd3_1 hold2962 (.A(\fpga_top.cpu_run_state ),
    .X(net6280));
 sg13g2_dlygate4sd3_1 hold2963 (.A(_06053_),
    .X(net6281));
 sg13g2_dlygate4sd3_1 hold2964 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[3] ),
    .X(net6282));
 sg13g2_dlygate4sd3_1 hold2965 (.A(\fpga_top.uart_top.uart_if.tx_out_cntr[0] ),
    .X(net6283));
 sg13g2_dlygate4sd3_1 hold2966 (.A(_03673_),
    .X(net6284));
 sg13g2_dlygate4sd3_1 hold2967 (.A(\fpga_top.bus_gather.d_write_data[8] ),
    .X(net6285));
 sg13g2_dlygate4sd3_1 hold2968 (.A(\fpga_top.bus_gather.u_read_adr[13] ),
    .X(net6286));
 sg13g2_dlygate4sd3_1 hold2969 (.A(_01412_),
    .X(net6287));
 sg13g2_dlygate4sd3_1 hold2970 (.A(\fpga_top.io_spi_lite.spi_mode[11] ),
    .X(net6288));
 sg13g2_dlygate4sd3_1 hold2971 (.A(\fpga_top.bus_gather.u_read_adr[18] ),
    .X(net6289));
 sg13g2_dlygate4sd3_1 hold2972 (.A(_01417_),
    .X(net6290));
 sg13g2_dlygate4sd3_1 hold2973 (.A(\fpga_top.bus_gather.u_read_adr[20] ),
    .X(net6291));
 sg13g2_dlygate4sd3_1 hold2974 (.A(_01419_),
    .X(net6292));
 sg13g2_dlygate4sd3_1 hold2975 (.A(\fpga_top.bus_gather.d_write_data[11] ),
    .X(net6293));
 sg13g2_dlygate4sd3_1 hold2976 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[21] ),
    .X(net6294));
 sg13g2_dlygate4sd3_1 hold2977 (.A(\fpga_top.qspi_if.adr_rw[2] ),
    .X(net6295));
 sg13g2_dlygate4sd3_1 hold2978 (.A(_00991_),
    .X(net6296));
 sg13g2_dlygate4sd3_1 hold2979 (.A(\fpga_top.uart_top.uart_send_char.send_cntr[2] ),
    .X(net6297));
 sg13g2_dlygate4sd3_1 hold2980 (.A(_02146_),
    .X(net6298));
 sg13g2_dlygate4sd3_1 hold2981 (.A(\fpga_top.uart_top.uart_if.sample_cntr[9] ),
    .X(net6299));
 sg13g2_dlygate4sd3_1 hold2982 (.A(_09320_),
    .X(net6300));
 sg13g2_dlygate4sd3_1 hold2983 (.A(\fpga_top.bus_gather.u_read_adr[12] ),
    .X(net6301));
 sg13g2_dlygate4sd3_1 hold2984 (.A(uio_out[5]),
    .X(net6302));
 sg13g2_dlygate4sd3_1 hold2985 (.A(\fpga_top.bus_gather.u_read_adr[5] ),
    .X(net6303));
 sg13g2_dlygate4sd3_1 hold2986 (.A(_04680_),
    .X(net6304));
 sg13g2_dlygate4sd3_1 hold2987 (.A(uio_out[4]),
    .X(net6305));
 sg13g2_dlygate4sd3_1 hold2988 (.A(\fpga_top.qspi_if.inner_state[1] ),
    .X(net6306));
 sg13g2_dlygate4sd3_1 hold2989 (.A(\fpga_top.cpu_top.cpu_state_machine.cpu_state[2] ),
    .X(net6307));
 sg13g2_dlygate4sd3_1 hold2990 (.A(_09459_),
    .X(net6308));
 sg13g2_dlygate4sd3_1 hold2991 (.A(_00024_),
    .X(net6309));
 sg13g2_dlygate4sd3_1 hold2992 (.A(\fpga_top.io_uart_out.rout[7] ),
    .X(net6310));
 sg13g2_dlygate4sd3_1 hold2993 (.A(\fpga_top.io_uart_out.rout[6] ),
    .X(net6311));
 sg13g2_dlygate4sd3_1 hold2994 (.A(\fpga_top.io_spi_lite.spi_mode[10] ),
    .X(net6312));
 sg13g2_dlygate4sd3_1 hold2995 (.A(uio_oe[5]),
    .X(net6313));
 sg13g2_dlygate4sd3_1 hold2996 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[5] ),
    .X(net6314));
 sg13g2_dlygate4sd3_1 hold2997 (.A(\fpga_top.bus_gather.u_read_adr[6] ),
    .X(net6315));
 sg13g2_dlygate4sd3_1 hold2998 (.A(_01405_),
    .X(net6316));
 sg13g2_dlygate4sd3_1 hold2999 (.A(\fpga_top.bus_gather.u_read_adr[29] ),
    .X(net6317));
 sg13g2_dlygate4sd3_1 hold3000 (.A(\fpga_top.uart_top.uart_send_char.send_cntr[4] ),
    .X(net6318));
 sg13g2_dlygate4sd3_1 hold3001 (.A(\fpga_top.bus_gather.u_read_adr[24] ),
    .X(net6319));
 sg13g2_dlygate4sd3_1 hold3002 (.A(_01423_),
    .X(net6320));
 sg13g2_dlygate4sd3_1 hold3003 (.A(\fpga_top.io_frc.frc_cntr_val[4] ),
    .X(net6321));
 sg13g2_dlygate4sd3_1 hold3004 (.A(_00400_),
    .X(net6322));
 sg13g2_dlygate4sd3_1 hold3005 (.A(\fpga_top.qspi_if.wredge[0] ),
    .X(net6323));
 sg13g2_dlygate4sd3_1 hold3006 (.A(\fpga_top.uart_top.uart_if.rx_fifo.ram_wadr[2] ),
    .X(net6324));
 sg13g2_dlygate4sd3_1 hold3007 (.A(uio_out[6]),
    .X(net6325));
 sg13g2_dlygate4sd3_1 hold3008 (.A(\fpga_top.bus_gather.d_write_data[29] ),
    .X(net6326));
 sg13g2_dlygate4sd3_1 hold3009 (.A(\fpga_top.qspi_if.word_hw ),
    .X(net6327));
 sg13g2_dlygate4sd3_1 hold3010 (.A(_00956_),
    .X(net6328));
 sg13g2_dlygate4sd3_1 hold3011 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[19] ),
    .X(net6329));
 sg13g2_dlygate4sd3_1 hold3012 (.A(\fpga_top.io_frc.frc_cntr_val[5] ),
    .X(net6330));
 sg13g2_dlygate4sd3_1 hold3013 (.A(\fpga_top.cpu_top.alu_code[0] ),
    .X(net6331));
 sg13g2_dlygate4sd3_1 hold3014 (.A(\fpga_top.io_spi_lite.spi_mode[5] ),
    .X(net6332));
 sg13g2_dlygate4sd3_1 hold3015 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[19] ),
    .X(net6333));
 sg13g2_dlygate4sd3_1 hold3016 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[25] ),
    .X(net6334));
 sg13g2_dlygate4sd3_1 hold3017 (.A(\fpga_top.io_frc.frc_cntr_val[1] ),
    .X(net6335));
 sg13g2_dlygate4sd3_1 hold3018 (.A(\fpga_top.bus_gather.d_write_data[6] ),
    .X(net6336));
 sg13g2_dlygate4sd3_1 hold3019 (.A(\fpga_top.bus_gather.d_write_data[18] ),
    .X(net6337));
 sg13g2_dlygate4sd3_1 hold3020 (.A(\fpga_top.qspi_if.qspi_state[10] ),
    .X(net6338));
 sg13g2_dlygate4sd3_1 hold3021 (.A(\fpga_top.qspi_if.sio_out_pre[1] ),
    .X(net6339));
 sg13g2_dlygate4sd3_1 hold3022 (.A(\fpga_top.cpu_top.alui_shamt[0] ),
    .X(net6340));
 sg13g2_dlygate4sd3_1 hold3023 (.A(\fpga_top.bus_gather.u_read_adr[10] ),
    .X(net6341));
 sg13g2_dlygate4sd3_1 hold3024 (.A(_01409_),
    .X(net6342));
 sg13g2_dlygate4sd3_1 hold3025 (.A(\fpga_top.cpu_top.register_file.rfr_state[2] ),
    .X(net6343));
 sg13g2_dlygate4sd3_1 hold3026 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[1] ),
    .X(net6344));
 sg13g2_dlygate4sd3_1 hold3027 (.A(\fpga_top.bus_gather.d_write_data[13] ),
    .X(net6345));
 sg13g2_dlygate4sd3_1 hold3028 (.A(\fpga_top.cpu_top.register_file.rfr_state[1] ),
    .X(net6346));
 sg13g2_dlygate4sd3_1 hold3029 (.A(\fpga_top.io_frc.frc_cntr_val[28] ),
    .X(net6347));
 sg13g2_dlygate4sd3_1 hold3030 (.A(\fpga_top.uart_top.uart_if.tx_out_cntr[1] ),
    .X(net6348));
 sg13g2_dlygate4sd3_1 hold3031 (.A(_03676_),
    .X(net6349));
 sg13g2_dlygate4sd3_1 hold3032 (.A(\fpga_top.uart_top.uart_if.rx_state[3] ),
    .X(net6350));
 sg13g2_dlygate4sd3_1 hold3033 (.A(\fpga_top.qspi_if.rwait_cntr[1] ),
    .X(net6351));
 sg13g2_dlygate4sd3_1 hold3034 (.A(\fpga_top.bus_gather.d_write_data[23] ),
    .X(net6352));
 sg13g2_dlygate4sd3_1 hold3035 (.A(\fpga_top.cpu_top.csr_rmie ),
    .X(net6353));
 sg13g2_dlygate4sd3_1 hold3036 (.A(_00027_),
    .X(net6354));
 sg13g2_dlygate4sd3_1 hold3037 (.A(\fpga_top.qspi_if.sck_cntr[2] ),
    .X(net6355));
 sg13g2_dlygate4sd3_1 hold3038 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[4] ),
    .X(net6356));
 sg13g2_dlygate4sd3_1 hold3039 (.A(\fpga_top.uart_top.uart_if.sample_cntr[12] ),
    .X(net6357));
 sg13g2_dlygate4sd3_1 hold3040 (.A(_09326_),
    .X(net6358));
 sg13g2_dlygate4sd3_1 hold3041 (.A(\fpga_top.io_spi_lite.spi_mode[4] ),
    .X(net6359));
 sg13g2_dlygate4sd3_1 hold3042 (.A(uio_oe[6]),
    .X(net6360));
 sg13g2_dlygate4sd3_1 hold3043 (.A(\fpga_top.qspi_if.wdata_ofs[0] ),
    .X(net6361));
 sg13g2_dlygate4sd3_1 hold3044 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[3] ),
    .X(net6362));
 sg13g2_dlygate4sd3_1 hold3045 (.A(\fpga_top.bus_gather.d_write_data[12] ),
    .X(net6363));
 sg13g2_dlygate4sd3_1 hold3046 (.A(\fpga_top.bus_gather.u_read_adr[8] ),
    .X(net6364));
 sg13g2_dlygate4sd3_1 hold3047 (.A(\fpga_top.dma_io_wadr_u[15] ),
    .X(net6365));
 sg13g2_dlygate4sd3_1 hold3048 (.A(_04301_),
    .X(net6366));
 sg13g2_dlygate4sd3_1 hold3049 (.A(_01217_),
    .X(net6367));
 sg13g2_dlygate4sd3_1 hold3050 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[15] ),
    .X(net6368));
 sg13g2_dlygate4sd3_1 hold3051 (.A(\fpga_top.cmd_ld_ma ),
    .X(net6369));
 sg13g2_dlygate4sd3_1 hold3052 (.A(\fpga_top.cpu_top.csr_wadr_mon[4] ),
    .X(net6370));
 sg13g2_dlygate4sd3_1 hold3053 (.A(_01208_),
    .X(net6371));
 sg13g2_dlygate4sd3_1 hold3054 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[8] ),
    .X(net6372));
 sg13g2_dlygate4sd3_1 hold3055 (.A(uio_oe[4]),
    .X(net6373));
 sg13g2_dlygate4sd3_1 hold3056 (.A(\fpga_top.cpu_top.csr_wadr_mon[7] ),
    .X(net6374));
 sg13g2_dlygate4sd3_1 hold3057 (.A(\fpga_top.cpu_top.csr_uimm[4] ),
    .X(net6375));
 sg13g2_dlygate4sd3_1 hold3058 (.A(\fpga_top.bus_gather.d_write_data[25] ),
    .X(net6376));
 sg13g2_dlygate4sd3_1 hold3059 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[29] ),
    .X(net6377));
 sg13g2_dlygate4sd3_1 hold3060 (.A(\fpga_top.uart_top.trush_running ),
    .X(net6378));
 sg13g2_dlygate4sd3_1 hold3061 (.A(_04662_),
    .X(net6379));
 sg13g2_dlygate4sd3_1 hold3062 (.A(_01400_),
    .X(net6380));
 sg13g2_dlygate4sd3_1 hold3063 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[21] ),
    .X(net6381));
 sg13g2_dlygate4sd3_1 hold3064 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[27] ),
    .X(net6382));
 sg13g2_dlygate4sd3_1 hold3065 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[17] ),
    .X(net6383));
 sg13g2_dlygate4sd3_1 hold3066 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[9] ),
    .X(net6384));
 sg13g2_dlygate4sd3_1 hold3067 (.A(\fpga_top.qspi_if.rdwrch[4] ),
    .X(net6385));
 sg13g2_dlygate4sd3_1 hold3068 (.A(\fpga_top.cpu_top.csr_wadr_mon[3] ),
    .X(net6386));
 sg13g2_dlygate4sd3_1 hold3069 (.A(_04267_),
    .X(net6387));
 sg13g2_dlygate4sd3_1 hold3070 (.A(\fpga_top.io_uart_out.rout_en ),
    .X(net6388));
 sg13g2_dlygate4sd3_1 hold3071 (.A(\fpga_top.cpu_top.execution.alu_sra[31] ),
    .X(net6389));
 sg13g2_dlygate4sd3_1 hold3072 (.A(\fpga_top.cpu_top.alui_shamt[2] ),
    .X(net6390));
 sg13g2_dlygate4sd3_1 hold3073 (.A(\fpga_top.qspi_if.word_data[5] ),
    .X(net6391));
 sg13g2_dlygate4sd3_1 hold3074 (.A(_10165_),
    .X(net6392));
 sg13g2_dlygate4sd3_1 hold3075 (.A(\fpga_top.bus_gather.d_write_data[24] ),
    .X(net6393));
 sg13g2_dlygate4sd3_1 hold3076 (.A(\fpga_top.qspi_if.sck_cntr[3] ),
    .X(net6394));
 sg13g2_dlygate4sd3_1 hold3077 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[5] ),
    .X(net6395));
 sg13g2_dlygate4sd3_1 hold3078 (.A(\fpga_top.bus_gather.u_read_adr[2] ),
    .X(net6396));
 sg13g2_dlygate4sd3_1 hold3079 (.A(\fpga_top.qspi_if.adr_rw[20] ),
    .X(net6397));
 sg13g2_dlygate4sd3_1 hold3080 (.A(_01009_),
    .X(net6398));
 sg13g2_dlygate4sd3_1 hold3081 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[6] ),
    .X(net6399));
 sg13g2_dlygate4sd3_1 hold3082 (.A(\fpga_top.cpu_top.inst_mem_read.imr_stat_dly ),
    .X(net6400));
 sg13g2_dlygate4sd3_1 hold3083 (.A(_09446_),
    .X(net6401));
 sg13g2_dlygate4sd3_1 hold3084 (.A(\fpga_top.cpu_top.csr_wadr_mon[1] ),
    .X(net6402));
 sg13g2_dlygate4sd3_1 hold3085 (.A(_01205_),
    .X(net6403));
 sg13g2_dlygate4sd3_1 hold3086 (.A(\fpga_top.uart_top.uart_if.byte_data[1] ),
    .X(net6404));
 sg13g2_dlygate4sd3_1 hold3087 (.A(_01433_),
    .X(net6405));
 sg13g2_dlygate4sd3_1 hold3088 (.A(\fpga_top.cpu_top.br_ofs[10] ),
    .X(net6406));
 sg13g2_dlygate4sd3_1 hold3089 (.A(\fpga_top.cpu_top.csr_meie ),
    .X(net6407));
 sg13g2_dlygate4sd3_1 hold3090 (.A(\fpga_top.uart_top.uart_if.byte_data[3] ),
    .X(net6408));
 sg13g2_dlygate4sd3_1 hold3091 (.A(_01435_),
    .X(net6409));
 sg13g2_dlygate4sd3_1 hold3092 (.A(\fpga_top.bus_gather.i_read_adr[2] ),
    .X(net6410));
 sg13g2_dlygate4sd3_1 hold3093 (.A(uio_out[7]),
    .X(net6411));
 sg13g2_dlygate4sd3_1 hold3094 (.A(\fpga_top.qspi_if.adr_rw[8] ),
    .X(net6412));
 sg13g2_dlygate4sd3_1 hold3095 (.A(\fpga_top.bus_gather.i_read_adr[25] ),
    .X(net6413));
 sg13g2_dlygate4sd3_1 hold3096 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wen ),
    .X(net6414));
 sg13g2_dlygate4sd3_1 hold3097 (.A(_10576_),
    .X(net6415));
 sg13g2_dlygate4sd3_1 hold3098 (.A(_00211_),
    .X(net6416));
 sg13g2_dlygate4sd3_1 hold3099 (.A(_00085_),
    .X(net6417));
 sg13g2_dlygate4sd3_1 hold3100 (.A(uio_oe[7]),
    .X(net6418));
 sg13g2_dlygate4sd3_1 hold3101 (.A(\fpga_top.uart_top.uart_if.byte_data[0] ),
    .X(net6419));
 sg13g2_dlygate4sd3_1 hold3102 (.A(\fpga_top.qspi_if.cmd_ofs[1] ),
    .X(net6420));
 sg13g2_dlygate4sd3_1 hold3103 (.A(_03177_),
    .X(net6421));
 sg13g2_dlygate4sd3_1 hold3104 (.A(\fpga_top.bus_gather.d_write_data[27] ),
    .X(net6422));
 sg13g2_dlygate4sd3_1 hold3105 (.A(\fpga_top.bus_gather.d_write_data[14] ),
    .X(net6423));
 sg13g2_dlygate4sd3_1 hold3106 (.A(\fpga_top.uart_top.uart_logics.cmd_wadr_cntr[31] ),
    .X(net6424));
 sg13g2_dlygate4sd3_1 hold3107 (.A(\fpga_top.cpu_top.br_ofs[7] ),
    .X(net6425));
 sg13g2_dlygate4sd3_1 hold3108 (.A(_01638_),
    .X(net6426));
 sg13g2_dlygate4sd3_1 hold3109 (.A(\fpga_top.cpu_top.data_rw_mem.data_state[0] ),
    .X(net6427));
 sg13g2_dlygate4sd3_1 hold3110 (.A(_08840_),
    .X(net6428));
 sg13g2_dlygate4sd3_1 hold3111 (.A(_08843_),
    .X(net6429));
 sg13g2_dlygate4sd3_1 hold3112 (.A(\fpga_top.io_spi_lite.sel_mosi[7] ),
    .X(net6430));
 sg13g2_dlygate4sd3_1 hold3113 (.A(\fpga_top.bus_gather.d_write_data[21] ),
    .X(net6431));
 sg13g2_dlygate4sd3_1 hold3114 (.A(\fpga_top.cpu_start_adr[9] ),
    .X(net6432));
 sg13g2_dlygate4sd3_1 hold3115 (.A(\fpga_top.cpu_top.csr_wadr_mon[8] ),
    .X(net6433));
 sg13g2_dlygate4sd3_1 hold3116 (.A(\fpga_top.cpu_top.csr_wadr_mon[2] ),
    .X(net6434));
 sg13g2_dlygate4sd3_1 hold3117 (.A(_01206_),
    .X(net6435));
 sg13g2_dlygate4sd3_1 hold3118 (.A(\fpga_top.qspi_if.adr_rw[18] ),
    .X(net6436));
 sg13g2_dlygate4sd3_1 hold3119 (.A(_03445_),
    .X(net6437));
 sg13g2_dlygate4sd3_1 hold3120 (.A(\fpga_top.cpu_top.br_ofs[12] ),
    .X(net6438));
 sg13g2_dlygate4sd3_1 hold3121 (.A(\fpga_top.cpu_top.decoder.illegal_ops_inst[4] ),
    .X(net6439));
 sg13g2_dlygate4sd3_1 hold3122 (.A(\fpga_top.cpu_top.csr_wadr_mon[6] ),
    .X(net6440));
 sg13g2_dlygate4sd3_1 hold3123 (.A(\fpga_top.uart_top.uart_logics.data_0[5] ),
    .X(net6441));
 sg13g2_dlygate4sd3_1 hold3124 (.A(\fpga_top.io_spi_lite.miso_fifo.radr[1] ),
    .X(net6442));
 sg13g2_dlygate4sd3_1 hold3125 (.A(\fpga_top.qspi_if.adr_rw[6] ),
    .X(net6443));
 sg13g2_dlygate4sd3_1 hold3126 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[13] ),
    .X(net6444));
 sg13g2_dlygate4sd3_1 hold3127 (.A(\fpga_top.cpu_top.br_ofs[5] ),
    .X(net6445));
 sg13g2_dlygate4sd3_1 hold3128 (.A(_01636_),
    .X(net6446));
 sg13g2_dlygate4sd3_1 hold3129 (.A(\fpga_top.uart_top.uart_if.tx_out_cntr[1] ),
    .X(net6447));
 sg13g2_dlygate4sd3_1 hold3130 (.A(\fpga_top.qspi_if.adr_rw[19] ),
    .X(net6448));
 sg13g2_dlygate4sd3_1 hold3131 (.A(\fpga_top.bus_gather.u_read_adr[4] ),
    .X(net6449));
 sg13g2_dlygate4sd3_1 hold3132 (.A(_01403_),
    .X(net6450));
 sg13g2_dlygate4sd3_1 hold3133 (.A(\fpga_top.qspi_if.adr_rw[11] ),
    .X(net6451));
 sg13g2_dlygate4sd3_1 hold3134 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[26] ),
    .X(net6452));
 sg13g2_dlygate4sd3_1 hold3135 (.A(\fpga_top.qspi_if.adr_rw[5] ),
    .X(net6453));
 sg13g2_dlygate4sd3_1 hold3136 (.A(_00994_),
    .X(net6454));
 sg13g2_dlygate4sd3_1 hold3137 (.A(\fpga_top.cpu_top.csr_uimm[3] ),
    .X(net6455));
 sg13g2_dlygate4sd3_1 hold3138 (.A(\fpga_top.cpu_top.alu_code[2] ),
    .X(net6456));
 sg13g2_dlygate4sd3_1 hold3139 (.A(\fpga_top.bus_gather.d_write_data[30] ),
    .X(net6457));
 sg13g2_dlygate4sd3_1 hold3140 (.A(\fpga_top.uart_top.uart_logics.status_dump[0] ),
    .X(net6458));
 sg13g2_dlygate4sd3_1 hold3141 (.A(_06998_),
    .X(net6459));
 sg13g2_dlygate4sd3_1 hold3142 (.A(\fpga_top.uart_top.uart_logics.next_status_dump[0] ),
    .X(net6460));
 sg13g2_dlygate4sd3_1 hold3143 (.A(\fpga_top.qspi_if.adr_rw[10] ),
    .X(net6461));
 sg13g2_dlygate4sd3_1 hold3144 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[12] ),
    .X(net6462));
 sg13g2_dlygate4sd3_1 hold3145 (.A(\fpga_top.cpu_top.alu_code[1] ),
    .X(net6463));
 sg13g2_dlygate4sd3_1 hold3146 (.A(\fpga_top.qspi_if.adr_ofs[0] ),
    .X(net6464));
 sg13g2_dlygate4sd3_1 hold3147 (.A(_01100_),
    .X(net6465));
 sg13g2_dlygate4sd3_1 hold3148 (.A(\fpga_top.qspi_if.adr_ofs[2] ),
    .X(net6466));
 sg13g2_dlygate4sd3_1 hold3149 (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[4] ),
    .X(net6467));
 sg13g2_dlygate4sd3_1 hold3150 (.A(_06953_),
    .X(net6468));
 sg13g2_dlygate4sd3_1 hold3151 (.A(\fpga_top.uart_top.uart_rec_char.g_crlf ),
    .X(net6469));
 sg13g2_dlygate4sd3_1 hold3152 (.A(\fpga_top.cpu_top.br_ofs[8] ),
    .X(net6470));
 sg13g2_dlygate4sd3_1 hold3153 (.A(\fpga_top.qspi_if.adr_rw[15] ),
    .X(net6471));
 sg13g2_dlygate4sd3_1 hold3154 (.A(\fpga_top.cpu_start_adr[3] ),
    .X(net6472));
 sg13g2_dlygate4sd3_1 hold3155 (.A(\fpga_top.qspi_if.rwait_cntr[2] ),
    .X(net6473));
 sg13g2_dlygate4sd3_1 hold3156 (.A(_03524_),
    .X(net6474));
 sg13g2_dlygate4sd3_1 hold3157 (.A(\fpga_top.cpu_top.pc_stage.cpu_adr_ld ),
    .X(net6475));
 sg13g2_dlygate4sd3_1 hold3158 (.A(_01501_),
    .X(net6476));
 sg13g2_dlygate4sd3_1 hold3159 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[22] ),
    .X(net6477));
 sg13g2_dlygate4sd3_1 hold3160 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[28] ),
    .X(net6478));
 sg13g2_dlygate4sd3_1 hold3161 (.A(\fpga_top.bus_gather.i_read_adr[30] ),
    .X(net6479));
 sg13g2_dlygate4sd3_1 hold3162 (.A(\fpga_top.cpu_top.csr_wadr_mon[8] ),
    .X(net6480));
 sg13g2_dlygate4sd3_1 hold3163 (.A(\fpga_top.qspi_if.qspi_state[3] ),
    .X(net6481));
 sg13g2_dlygate4sd3_1 hold3164 (.A(\fpga_top.cpu_top.data_rw_mem.req_w_dly ),
    .X(net6482));
 sg13g2_dlygate4sd3_1 hold3165 (.A(\fpga_top.bus_gather.i_read_adr[5] ),
    .X(net6483));
 sg13g2_dlygate4sd3_1 hold3166 (.A(\fpga_top.io_spi_lite.spi_mode[7] ),
    .X(net6484));
 sg13g2_dlygate4sd3_1 hold3167 (.A(\fpga_top.qspi_if.adr_rw[22] ),
    .X(net6485));
 sg13g2_dlygate4sd3_1 hold3168 (.A(\fpga_top.cpu_top.csr_wdata_mon[1] ),
    .X(net6486));
 sg13g2_dlygate4sd3_1 hold3169 (.A(_01236_),
    .X(net6487));
 sg13g2_dlygate4sd3_1 hold3170 (.A(\fpga_top.bus_gather.i_read_adr[12] ),
    .X(net6488));
 sg13g2_dlygate4sd3_1 hold3171 (.A(\fpga_top.cpu_top.register_file.rfr_state[0] ),
    .X(net6489));
 sg13g2_dlygate4sd3_1 hold3172 (.A(\fpga_top.bus_gather.i_read_adr[31] ),
    .X(net6490));
 sg13g2_dlygate4sd3_1 hold3173 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[1] ),
    .X(net6491));
 sg13g2_dlygate4sd3_1 hold3174 (.A(_00212_),
    .X(net6492));
 sg13g2_dlygate4sd3_1 hold3175 (.A(\fpga_top.bus_gather.i_read_adr[7] ),
    .X(net6493));
 sg13g2_dlygate4sd3_1 hold3176 (.A(\fpga_top.bus_gather.u_read_adr[22] ),
    .X(net6494));
 sg13g2_dlygate4sd3_1 hold3177 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[30] ),
    .X(net6495));
 sg13g2_dlygate4sd3_1 hold3178 (.A(\fpga_top.cpu_top.cpu_state_machine.cpu_state[1] ),
    .X(net6496));
 sg13g2_dlygate4sd3_1 hold3179 (.A(_09456_),
    .X(net6497));
 sg13g2_dlygate4sd3_1 hold3180 (.A(\fpga_top.bus_gather.i_read_adr[4] ),
    .X(net6498));
 sg13g2_dlygate4sd3_1 hold3181 (.A(_01482_),
    .X(net6499));
 sg13g2_dlygate4sd3_1 hold3182 (.A(\fpga_top.qspi_if.adr_rw[21] ),
    .X(net6500));
 sg13g2_dlygate4sd3_1 hold3183 (.A(_03467_),
    .X(net6501));
 sg13g2_dlygate4sd3_1 hold3184 (.A(_01010_),
    .X(net6502));
 sg13g2_dlygate4sd3_1 hold3185 (.A(\fpga_top.qspi_if.cmd_ofs[2] ),
    .X(net6503));
 sg13g2_dlygate4sd3_1 hold3186 (.A(\fpga_top.bus_gather.i_read_adr[14] ),
    .X(net6504));
 sg13g2_dlygate4sd3_1 hold3187 (.A(_01492_),
    .X(net6505));
 sg13g2_dlygate4sd3_1 hold3188 (.A(\fpga_top.bus_gather.i_read_adr[9] ),
    .X(net6506));
 sg13g2_dlygate4sd3_1 hold3189 (.A(\fpga_top.uart_top.uart_send_char.send_cntr[1] ),
    .X(net6507));
 sg13g2_dlygate4sd3_1 hold3190 (.A(_06257_),
    .X(net6508));
 sg13g2_dlygate4sd3_1 hold3191 (.A(_02145_),
    .X(net6509));
 sg13g2_dlygate4sd3_1 hold3192 (.A(\fpga_top.bus_gather.i_read_adr[11] ),
    .X(net6510));
 sg13g2_dlygate4sd3_1 hold3193 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[14] ),
    .X(net6511));
 sg13g2_dlygate4sd3_1 hold3194 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[0] ),
    .X(net6512));
 sg13g2_dlygate4sd3_1 hold3195 (.A(\fpga_top.qspi_if.adr_rw[23] ),
    .X(net6513));
 sg13g2_dlygate4sd3_1 hold3196 (.A(\fpga_top.cpu_top.cpu_state_machine.cpu_state[0] ),
    .X(net6514));
 sg13g2_dlygate4sd3_1 hold3197 (.A(_09447_),
    .X(net6515));
 sg13g2_dlygate4sd3_1 hold3198 (.A(\fpga_top.qspi_if.cmd_ofs[0] ),
    .X(net6516));
 sg13g2_dlygate4sd3_1 hold3199 (.A(\fpga_top.cpu_top.alui_shamt[4] ),
    .X(net6517));
 sg13g2_dlygate4sd3_1 hold3200 (.A(_01635_),
    .X(net6518));
 sg13g2_dlygate4sd3_1 hold3201 (.A(\fpga_top.bus_gather.i_read_adr[15] ),
    .X(net6519));
 sg13g2_dlygate4sd3_1 hold3202 (.A(\fpga_top.cpu_top.alui_shamt[1] ),
    .X(net6520));
 sg13g2_dlygate4sd3_1 hold3203 (.A(\fpga_top.uart_top.uart_if.byte_data[2] ),
    .X(net6521));
 sg13g2_dlygate4sd3_1 hold3204 (.A(\fpga_top.cpu_top.alui_shamt[3] ),
    .X(net6522));
 sg13g2_dlygate4sd3_1 hold3205 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[18] ),
    .X(net6523));
 sg13g2_dlygate4sd3_1 hold3206 (.A(\fpga_top.bus_gather.u_read_adr[31] ),
    .X(net6524));
 sg13g2_dlygate4sd3_1 hold3207 (.A(\fpga_top.uart_top.uart_rec_char.word_valid ),
    .X(net6525));
 sg13g2_dlygate4sd3_1 hold3208 (.A(\fpga_top.uart_top.uart_logics.next_status_dump[1] ),
    .X(net6526));
 sg13g2_dlygate4sd3_1 hold3209 (.A(\fpga_top.bus_gather.u_read_adr[21] ),
    .X(net6527));
 sg13g2_dlygate4sd3_1 hold3210 (.A(_01420_),
    .X(net6528));
 sg13g2_dlygate4sd3_1 hold3211 (.A(\fpga_top.qspi_if.word_adr[24] ),
    .X(net6529));
 sg13g2_dlygate4sd3_1 hold3212 (.A(\fpga_top.bus_gather.i_read_adr[26] ),
    .X(net6530));
 sg13g2_dlygate4sd3_1 hold3213 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[10] ),
    .X(net6531));
 sg13g2_dlygate4sd3_1 hold3214 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[20] ),
    .X(net6532));
 sg13g2_dlygate4sd3_1 hold3215 (.A(\fpga_top.cpu_top.cpu_state_machine.cpu_state[2] ),
    .X(net6533));
 sg13g2_dlygate4sd3_1 hold3216 (.A(_09461_),
    .X(net6534));
 sg13g2_dlygate4sd3_1 hold3217 (.A(\fpga_top.bus_gather.i_read_adr[10] ),
    .X(net6535));
 sg13g2_dlygate4sd3_1 hold3218 (.A(\fpga_top.io_spi_lite.miso_fifo.sfifo_1r1w.ram_wadr[2] ),
    .X(net6536));
 sg13g2_dlygate4sd3_1 hold3219 (.A(_10582_),
    .X(net6537));
 sg13g2_dlygate4sd3_1 hold3220 (.A(\fpga_top.bus_gather.i_read_adr[3] ),
    .X(net6538));
 sg13g2_dlygate4sd3_1 hold3221 (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[0] ),
    .X(net6539));
 sg13g2_dlygate4sd3_1 hold3222 (.A(\fpga_top.bus_gather.i_read_adr[6] ),
    .X(net6540));
 sg13g2_dlygate4sd3_1 hold3223 (.A(_01484_),
    .X(net6541));
 sg13g2_dlygate4sd3_1 hold3224 (.A(\fpga_top.cpu_top.data_rw_mem.data_state[1] ),
    .X(net6542));
 sg13g2_dlygate4sd3_1 hold3225 (.A(_08859_),
    .X(net6543));
 sg13g2_dlygate4sd3_1 hold3226 (.A(\fpga_top.cpu_start ),
    .X(net6544));
 sg13g2_dlygate4sd3_1 hold3227 (.A(\fpga_top.qspi_if.wdata_ofs[2] ),
    .X(net6545));
 sg13g2_dlygate4sd3_1 hold3228 (.A(_03571_),
    .X(net6546));
 sg13g2_dlygate4sd3_1 hold3229 (.A(\fpga_top.bus_gather.i_read_adr[18] ),
    .X(net6547));
 sg13g2_dlygate4sd3_1 hold3230 (.A(_05136_),
    .X(net6548));
 sg13g2_dlygate4sd3_1 hold3231 (.A(\fpga_top.bus_gather.i_read_adr[24] ),
    .X(net6549));
 sg13g2_dlygate4sd3_1 hold3232 (.A(_01502_),
    .X(net6550));
 sg13g2_dlygate4sd3_1 hold3233 (.A(\fpga_top.qspi_if.wdata[12] ),
    .X(net6551));
 sg13g2_dlygate4sd3_1 hold3234 (.A(\fpga_top.bus_gather.i_read_adr[16] ),
    .X(net6552));
 sg13g2_dlygate4sd3_1 hold3235 (.A(_01494_),
    .X(net6553));
 sg13g2_dlygate4sd3_1 hold3236 (.A(\fpga_top.bus_gather.u_read_adr[30] ),
    .X(net6554));
 sg13g2_dlygate4sd3_1 hold3237 (.A(\fpga_top.cpu_top.br_ofs[6] ),
    .X(net6555));
 sg13g2_dlygate4sd3_1 hold3238 (.A(_01637_),
    .X(net6556));
 sg13g2_dlygate4sd3_1 hold3239 (.A(\fpga_top.bus_gather.i_read_adr[17] ),
    .X(net6557));
 sg13g2_dlygate4sd3_1 hold3240 (.A(\fpga_top.bus_gather.i_read_adr[20] ),
    .X(net6558));
 sg13g2_dlygate4sd3_1 hold3241 (.A(\fpga_top.bus_gather.i_read_adr[28] ),
    .X(net6559));
 sg13g2_dlygate4sd3_1 hold3242 (.A(\fpga_top.cpu_start_adr[25] ),
    .X(net6560));
 sg13g2_dlygate4sd3_1 hold3243 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[2] ),
    .X(net6561));
 sg13g2_dlygate4sd3_1 hold3244 (.A(\fpga_top.bus_gather.i_read_adr[21] ),
    .X(net6562));
 sg13g2_dlygate4sd3_1 hold3245 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[7] ),
    .X(net6563));
 sg13g2_dlygate4sd3_1 hold3246 (.A(\fpga_top.bus_gather.i_read_adr[13] ),
    .X(net6564));
 sg13g2_dlygate4sd3_1 hold3247 (.A(\fpga_top.bus_gather.i_read_adr[29] ),
    .X(net6565));
 sg13g2_dlygate4sd3_1 hold3248 (.A(\fpga_top.qspi_if.adr_rw[17] ),
    .X(net6566));
 sg13g2_dlygate4sd3_1 hold3249 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[23] ),
    .X(net6567));
 sg13g2_dlygate4sd3_1 hold3250 (.A(\fpga_top.cpu_top.br_ofs[9] ),
    .X(net6568));
 sg13g2_dlygate4sd3_1 hold3251 (.A(\fpga_top.bus_gather.i_read_adr[27] ),
    .X(net6569));
 sg13g2_dlygate4sd3_1 hold3252 (.A(\fpga_top.qspi_if.qspi_state[6] ),
    .X(net6570));
 sg13g2_dlygate4sd3_1 hold3253 (.A(_09092_),
    .X(net6571));
 sg13g2_dlygate4sd3_1 hold3254 (.A(_09620_),
    .X(net6572));
 sg13g2_dlygate4sd3_1 hold3255 (.A(\fpga_top.uart_top.uart_logics.status_dump[2] ),
    .X(net6573));
 sg13g2_dlygate4sd3_1 hold3256 (.A(\fpga_top.uart_top.uart_logics.radr_enable ),
    .X(net6574));
 sg13g2_dlygate4sd3_1 hold3257 (.A(\fpga_top.cpu_top.csr_wadr_mon[0] ),
    .X(net6575));
 sg13g2_dlygate4sd3_1 hold3258 (.A(_01204_),
    .X(net6576));
 sg13g2_dlygate4sd3_1 hold3259 (.A(\fpga_top.cmd_st_ma ),
    .X(net6577));
 sg13g2_dlygate4sd3_1 hold3260 (.A(_00955_),
    .X(net6578));
 sg13g2_dlygate4sd3_1 hold3261 (.A(\fpga_top.bus_gather.i_read_adr[19] ),
    .X(net6579));
 sg13g2_dlygate4sd3_1 hold3262 (.A(_01497_),
    .X(net6580));
 sg13g2_dlygate4sd3_1 hold3263 (.A(\fpga_top.cpu_top.csr_wdata_mon[0] ),
    .X(net6581));
 sg13g2_dlygate4sd3_1 hold3264 (.A(\fpga_top.cpu_start_adr[2] ),
    .X(net6582));
 sg13g2_dlygate4sd3_1 hold3265 (.A(\fpga_top.bus_gather.i_read_adr[22] ),
    .X(net6583));
 sg13g2_dlygate4sd3_1 hold3266 (.A(\fpga_top.uart_top.uart_send_char.send_cntr[0] ),
    .X(net6584));
 sg13g2_dlygate4sd3_1 hold3267 (.A(\fpga_top.cpu_top.execution.csr_array.rs1_sel[24] ),
    .X(net6585));
 sg13g2_dlygate4sd3_1 hold3268 (.A(\fpga_top.uart_top.uart_rec_char.cmd_status[3] ),
    .X(net6586));
 sg13g2_dlygate4sd3_1 hold3269 (.A(\fpga_top.cpu_start_adr[25] ),
    .X(net6587));
 sg13g2_dlygate4sd3_1 hold3270 (.A(\fpga_top.cpu_start_adr[31] ),
    .X(net6588));
 sg13g2_dlygate4sd3_1 hold3271 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[0] ),
    .X(net6589));
 sg13g2_dlygate4sd3_1 hold3272 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[1] ),
    .X(net6590));
 sg13g2_dlygate4sd3_1 hold3273 (.A(_06267_),
    .X(net6591));
 sg13g2_dlygate4sd3_1 hold3274 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[2] ),
    .X(net6592));
 sg13g2_dlygate4sd3_1 hold3275 (.A(_06273_),
    .X(net6593));
 sg13g2_dlygate4sd3_1 hold3276 (.A(\fpga_top.qspi_if.sck_cntr[9] ),
    .X(net6594));
 sg13g2_dlygate4sd3_1 hold3277 (.A(_09253_),
    .X(net6595));
 sg13g2_dlygate4sd3_1 hold3278 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[26] ),
    .X(net6596));
 sg13g2_dlygate4sd3_1 hold3279 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[2] ),
    .X(net6597));
 sg13g2_dlygate4sd3_1 hold3280 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[0] ),
    .X(net6598));
 sg13g2_dlygate4sd3_1 hold3281 (.A(\fpga_top.uart_top.uart_if.sample_cntr[4] ),
    .X(net6599));
 sg13g2_dlygate4sd3_1 hold3282 (.A(_03639_),
    .X(net6600));
 sg13g2_dlygate4sd3_1 hold3283 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[2] ),
    .X(net6601));
 sg13g2_dlygate4sd3_1 hold3284 (.A(\fpga_top.qspi_if.cmd_ofs[0] ),
    .X(net6602));
 sg13g2_dlygate4sd3_1 hold3285 (.A(\fpga_top.qspi_if.sck_cntr[5] ),
    .X(net6603));
 sg13g2_dlygate4sd3_1 hold3286 (.A(\fpga_top.bus_gather.i_read_adr[6] ),
    .X(net6604));
 sg13g2_dlygate4sd3_1 hold3287 (.A(_05617_),
    .X(net6605));
 sg13g2_dlygate4sd3_1 hold3288 (.A(\fpga_top.io_frc.frc_cntr_val[51] ),
    .X(net6606));
 sg13g2_dlygate4sd3_1 hold3289 (.A(_06182_),
    .X(net6607));
 sg13g2_dlygate4sd3_1 hold3290 (.A(\fpga_top.bus_gather.u_read_adr[30] ),
    .X(net6608));
 sg13g2_dlygate4sd3_1 hold3291 (.A(\fpga_top.uart_top.uart_if.tx_fifo.ram_wadr[1] ),
    .X(net6609));
 sg13g2_dlygate4sd3_1 hold3292 (.A(\fpga_top.io_frc.frc_cntr_val[29] ),
    .X(net6610));
 sg13g2_dlygate4sd3_1 hold3293 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[18] ),
    .X(net6611));
 sg13g2_dlygate4sd3_1 hold3294 (.A(\fpga_top.io_frc.frc_cntr_val[1] ),
    .X(net6612));
 sg13g2_dlygate4sd3_1 hold3295 (.A(\fpga_top.cpu_top.execution.csr_array.csr_mtvec[23] ),
    .X(net6613));
 sg13g2_dlygate4sd3_1 hold3296 (.A(\fpga_top.cpu_top.csr_uimm[2] ),
    .X(net6614));
 sg13g2_dlygate4sd3_1 hold3297 (.A(\fpga_top.cpu_top.br_ofs[8] ),
    .X(net6615));
 sg13g2_dlygate4sd3_1 hold3298 (.A(\fpga_top.qspi_if.qspi_state[11] ),
    .X(net6616));
 sg13g2_dlygate4sd3_1 hold3299 (.A(\fpga_top.io_spi_lite.mosi_fifo.sfifo_1r1w.ram_wadr[0] ),
    .X(net6617));
 sg13g2_dlygate4sd3_1 hold3300 (.A(\fpga_top.cpu_start_adr[25] ),
    .X(net6618));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(rst_n));
 sg13g2_antennanp ANTENNA_3 (.A(_04164_));
 sg13g2_antennanp ANTENNA_4 (.A(\fpga_top.cpu_start_adr[28] ));
 sg13g2_antennanp ANTENNA_5 (.A(\fpga_top.cpu_start_adr[28] ));
 sg13g2_antennanp ANTENNA_6 (.A(\fpga_top.cpu_start_adr[28] ));
 sg13g2_antennanp ANTENNA_7 (.A(\fpga_top.cpu_start_adr[28] ));
 sg13g2_antennanp ANTENNA_8 (.A(\fpga_top.cpu_start_adr[28] ));
 sg13g2_antennanp ANTENNA_9 (.A(\fpga_top.cpu_start_adr[28] ));
 sg13g2_antennanp ANTENNA_10 (.A(\fpga_top.cpu_start_adr[28] ));
 sg13g2_antennanp ANTENNA_11 (.A(\fpga_top.cpu_start_adr[28] ));
 sg13g2_antennanp ANTENNA_12 (.A(\fpga_top.cpu_top.csr_wdata_mon[1] ));
 sg13g2_antennanp ANTENNA_13 (.A(\fpga_top.cpu_top.csr_wdata_mon[1] ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_fill_1 FILLER_0_86 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_fill_2 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_125 ();
 sg13g2_decap_8 FILLER_0_132 ();
 sg13g2_decap_8 FILLER_0_139 ();
 sg13g2_decap_8 FILLER_0_146 ();
 sg13g2_decap_4 FILLER_0_153 ();
 sg13g2_fill_1 FILLER_0_184 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_fill_1 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_fill_2 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_fill_2 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_4 FILLER_0_387 ();
 sg13g2_fill_2 FILLER_0_391 ();
 sg13g2_fill_2 FILLER_0_419 ();
 sg13g2_fill_1 FILLER_0_421 ();
 sg13g2_fill_2 FILLER_0_453 ();
 sg13g2_decap_8 FILLER_0_459 ();
 sg13g2_decap_8 FILLER_0_466 ();
 sg13g2_fill_2 FILLER_0_473 ();
 sg13g2_decap_8 FILLER_0_523 ();
 sg13g2_decap_8 FILLER_0_584 ();
 sg13g2_fill_2 FILLER_0_591 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_4 FILLER_0_630 ();
 sg13g2_fill_2 FILLER_0_634 ();
 sg13g2_decap_4 FILLER_0_644 ();
 sg13g2_fill_1 FILLER_0_648 ();
 sg13g2_decap_8 FILLER_0_653 ();
 sg13g2_decap_8 FILLER_0_660 ();
 sg13g2_decap_8 FILLER_0_667 ();
 sg13g2_decap_8 FILLER_0_674 ();
 sg13g2_decap_8 FILLER_0_681 ();
 sg13g2_decap_8 FILLER_0_688 ();
 sg13g2_fill_2 FILLER_0_695 ();
 sg13g2_decap_8 FILLER_0_725 ();
 sg13g2_decap_8 FILLER_0_732 ();
 sg13g2_decap_8 FILLER_0_739 ();
 sg13g2_decap_8 FILLER_0_746 ();
 sg13g2_decap_4 FILLER_0_753 ();
 sg13g2_fill_1 FILLER_0_757 ();
 sg13g2_fill_2 FILLER_0_763 ();
 sg13g2_fill_1 FILLER_0_765 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_879 ();
 sg13g2_decap_8 FILLER_0_886 ();
 sg13g2_decap_8 FILLER_0_893 ();
 sg13g2_decap_4 FILLER_0_900 ();
 sg13g2_fill_2 FILLER_0_904 ();
 sg13g2_fill_2 FILLER_0_933 ();
 sg13g2_fill_2 FILLER_0_946 ();
 sg13g2_fill_1 FILLER_0_948 ();
 sg13g2_fill_1 FILLER_0_954 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_fill_1 FILLER_0_1018 ();
 sg13g2_fill_2 FILLER_0_1046 ();
 sg13g2_fill_1 FILLER_0_1048 ();
 sg13g2_fill_1 FILLER_0_1052 ();
 sg13g2_decap_8 FILLER_0_1059 ();
 sg13g2_decap_8 FILLER_0_1066 ();
 sg13g2_decap_8 FILLER_0_1073 ();
 sg13g2_decap_8 FILLER_0_1080 ();
 sg13g2_decap_8 FILLER_0_1087 ();
 sg13g2_decap_8 FILLER_0_1094 ();
 sg13g2_decap_4 FILLER_0_1101 ();
 sg13g2_fill_1 FILLER_0_1105 ();
 sg13g2_decap_8 FILLER_0_1133 ();
 sg13g2_decap_8 FILLER_0_1140 ();
 sg13g2_decap_8 FILLER_0_1147 ();
 sg13g2_decap_8 FILLER_0_1154 ();
 sg13g2_decap_8 FILLER_0_1161 ();
 sg13g2_decap_8 FILLER_0_1168 ();
 sg13g2_decap_8 FILLER_0_1175 ();
 sg13g2_decap_8 FILLER_0_1182 ();
 sg13g2_decap_8 FILLER_0_1189 ();
 sg13g2_decap_4 FILLER_0_1196 ();
 sg13g2_fill_1 FILLER_0_1200 ();
 sg13g2_fill_1 FILLER_0_1204 ();
 sg13g2_decap_4 FILLER_0_1231 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_4 FILLER_0_1281 ();
 sg13g2_decap_4 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1298 ();
 sg13g2_decap_8 FILLER_0_1305 ();
 sg13g2_decap_8 FILLER_0_1312 ();
 sg13g2_decap_8 FILLER_0_1319 ();
 sg13g2_decap_8 FILLER_0_1326 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_decap_4 FILLER_0_1372 ();
 sg13g2_fill_2 FILLER_0_1376 ();
 sg13g2_decap_8 FILLER_0_1381 ();
 sg13g2_decap_8 FILLER_0_1388 ();
 sg13g2_decap_4 FILLER_0_1395 ();
 sg13g2_fill_1 FILLER_0_1399 ();
 sg13g2_fill_2 FILLER_0_1436 ();
 sg13g2_decap_8 FILLER_0_1451 ();
 sg13g2_decap_8 FILLER_0_1458 ();
 sg13g2_decap_8 FILLER_0_1465 ();
 sg13g2_decap_8 FILLER_0_1472 ();
 sg13g2_decap_8 FILLER_0_1479 ();
 sg13g2_fill_2 FILLER_0_1486 ();
 sg13g2_fill_2 FILLER_0_1501 ();
 sg13g2_decap_8 FILLER_0_1521 ();
 sg13g2_decap_8 FILLER_0_1528 ();
 sg13g2_decap_8 FILLER_0_1535 ();
 sg13g2_decap_8 FILLER_0_1542 ();
 sg13g2_decap_4 FILLER_0_1549 ();
 sg13g2_decap_8 FILLER_0_1580 ();
 sg13g2_decap_8 FILLER_0_1587 ();
 sg13g2_decap_8 FILLER_0_1594 ();
 sg13g2_decap_8 FILLER_0_1601 ();
 sg13g2_decap_8 FILLER_0_1608 ();
 sg13g2_decap_4 FILLER_0_1615 ();
 sg13g2_fill_2 FILLER_0_1619 ();
 sg13g2_fill_2 FILLER_0_1631 ();
 sg13g2_fill_2 FILLER_0_1636 ();
 sg13g2_decap_8 FILLER_0_1643 ();
 sg13g2_decap_8 FILLER_0_1650 ();
 sg13g2_decap_8 FILLER_0_1657 ();
 sg13g2_decap_8 FILLER_0_1664 ();
 sg13g2_decap_8 FILLER_0_1671 ();
 sg13g2_fill_1 FILLER_0_1678 ();
 sg13g2_decap_8 FILLER_0_1692 ();
 sg13g2_decap_8 FILLER_0_1699 ();
 sg13g2_decap_8 FILLER_0_1706 ();
 sg13g2_decap_8 FILLER_0_1713 ();
 sg13g2_decap_8 FILLER_0_1720 ();
 sg13g2_decap_8 FILLER_0_1727 ();
 sg13g2_decap_8 FILLER_0_1734 ();
 sg13g2_decap_8 FILLER_0_1741 ();
 sg13g2_decap_8 FILLER_0_1748 ();
 sg13g2_decap_8 FILLER_0_1755 ();
 sg13g2_decap_8 FILLER_0_1762 ();
 sg13g2_decap_8 FILLER_0_1769 ();
 sg13g2_decap_8 FILLER_0_1776 ();
 sg13g2_decap_8 FILLER_0_1783 ();
 sg13g2_fill_2 FILLER_0_1798 ();
 sg13g2_decap_8 FILLER_0_1809 ();
 sg13g2_decap_8 FILLER_0_1816 ();
 sg13g2_decap_8 FILLER_0_1823 ();
 sg13g2_decap_8 FILLER_0_1830 ();
 sg13g2_fill_1 FILLER_0_1837 ();
 sg13g2_decap_8 FILLER_0_1865 ();
 sg13g2_decap_8 FILLER_0_1872 ();
 sg13g2_decap_8 FILLER_0_1879 ();
 sg13g2_decap_8 FILLER_0_1886 ();
 sg13g2_decap_8 FILLER_0_1893 ();
 sg13g2_decap_8 FILLER_0_1900 ();
 sg13g2_decap_8 FILLER_0_1907 ();
 sg13g2_decap_8 FILLER_0_1914 ();
 sg13g2_decap_8 FILLER_0_1921 ();
 sg13g2_decap_8 FILLER_0_1928 ();
 sg13g2_decap_8 FILLER_0_1935 ();
 sg13g2_decap_4 FILLER_0_1942 ();
 sg13g2_fill_2 FILLER_0_1946 ();
 sg13g2_decap_8 FILLER_0_1961 ();
 sg13g2_decap_8 FILLER_0_1968 ();
 sg13g2_decap_8 FILLER_0_1975 ();
 sg13g2_fill_2 FILLER_0_1982 ();
 sg13g2_fill_1 FILLER_0_1984 ();
 sg13g2_fill_1 FILLER_0_1998 ();
 sg13g2_decap_4 FILLER_0_2006 ();
 sg13g2_decap_8 FILLER_0_2019 ();
 sg13g2_decap_8 FILLER_0_2026 ();
 sg13g2_decap_4 FILLER_0_2033 ();
 sg13g2_decap_8 FILLER_0_2064 ();
 sg13g2_decap_8 FILLER_0_2071 ();
 sg13g2_decap_8 FILLER_0_2078 ();
 sg13g2_decap_8 FILLER_0_2085 ();
 sg13g2_decap_8 FILLER_0_2092 ();
 sg13g2_decap_8 FILLER_0_2099 ();
 sg13g2_decap_8 FILLER_0_2106 ();
 sg13g2_decap_8 FILLER_0_2113 ();
 sg13g2_decap_8 FILLER_0_2120 ();
 sg13g2_decap_8 FILLER_0_2127 ();
 sg13g2_decap_8 FILLER_0_2134 ();
 sg13g2_decap_8 FILLER_0_2141 ();
 sg13g2_decap_8 FILLER_0_2148 ();
 sg13g2_decap_8 FILLER_0_2155 ();
 sg13g2_decap_8 FILLER_0_2162 ();
 sg13g2_decap_8 FILLER_0_2169 ();
 sg13g2_fill_2 FILLER_0_2176 ();
 sg13g2_fill_2 FILLER_0_2187 ();
 sg13g2_decap_4 FILLER_0_2198 ();
 sg13g2_decap_8 FILLER_0_2206 ();
 sg13g2_decap_8 FILLER_0_2213 ();
 sg13g2_decap_8 FILLER_0_2220 ();
 sg13g2_decap_4 FILLER_0_2227 ();
 sg13g2_fill_1 FILLER_0_2231 ();
 sg13g2_decap_8 FILLER_0_2241 ();
 sg13g2_decap_8 FILLER_0_2248 ();
 sg13g2_decap_8 FILLER_0_2255 ();
 sg13g2_decap_4 FILLER_0_2262 ();
 sg13g2_fill_1 FILLER_0_2266 ();
 sg13g2_decap_8 FILLER_0_2294 ();
 sg13g2_decap_8 FILLER_0_2301 ();
 sg13g2_decap_8 FILLER_0_2308 ();
 sg13g2_decap_8 FILLER_0_2315 ();
 sg13g2_decap_8 FILLER_0_2322 ();
 sg13g2_decap_8 FILLER_0_2329 ();
 sg13g2_decap_8 FILLER_0_2336 ();
 sg13g2_decap_8 FILLER_0_2343 ();
 sg13g2_decap_8 FILLER_0_2350 ();
 sg13g2_decap_8 FILLER_0_2357 ();
 sg13g2_decap_8 FILLER_0_2364 ();
 sg13g2_fill_2 FILLER_0_2371 ();
 sg13g2_decap_8 FILLER_0_2392 ();
 sg13g2_decap_8 FILLER_0_2399 ();
 sg13g2_decap_8 FILLER_0_2406 ();
 sg13g2_decap_8 FILLER_0_2413 ();
 sg13g2_decap_8 FILLER_0_2420 ();
 sg13g2_decap_8 FILLER_0_2427 ();
 sg13g2_decap_8 FILLER_0_2434 ();
 sg13g2_decap_8 FILLER_0_2441 ();
 sg13g2_decap_8 FILLER_0_2448 ();
 sg13g2_decap_4 FILLER_0_2455 ();
 sg13g2_decap_8 FILLER_0_2488 ();
 sg13g2_decap_8 FILLER_0_2495 ();
 sg13g2_decap_8 FILLER_0_2502 ();
 sg13g2_decap_8 FILLER_0_2509 ();
 sg13g2_fill_2 FILLER_0_2526 ();
 sg13g2_fill_1 FILLER_0_2528 ();
 sg13g2_decap_8 FILLER_0_2538 ();
 sg13g2_decap_8 FILLER_0_2545 ();
 sg13g2_decap_8 FILLER_0_2552 ();
 sg13g2_decap_8 FILLER_0_2559 ();
 sg13g2_decap_8 FILLER_0_2566 ();
 sg13g2_decap_8 FILLER_0_2573 ();
 sg13g2_decap_8 FILLER_0_2580 ();
 sg13g2_decap_8 FILLER_0_2587 ();
 sg13g2_decap_8 FILLER_0_2594 ();
 sg13g2_decap_8 FILLER_0_2601 ();
 sg13g2_fill_2 FILLER_0_2608 ();
 sg13g2_decap_8 FILLER_0_2614 ();
 sg13g2_fill_2 FILLER_0_2621 ();
 sg13g2_fill_1 FILLER_0_2623 ();
 sg13g2_decap_8 FILLER_0_2633 ();
 sg13g2_decap_8 FILLER_0_2640 ();
 sg13g2_decap_8 FILLER_0_2647 ();
 sg13g2_decap_8 FILLER_0_2654 ();
 sg13g2_decap_8 FILLER_0_2661 ();
 sg13g2_decap_8 FILLER_0_2668 ();
 sg13g2_decap_8 FILLER_0_2675 ();
 sg13g2_decap_8 FILLER_0_2682 ();
 sg13g2_decap_8 FILLER_0_2689 ();
 sg13g2_decap_4 FILLER_0_2696 ();
 sg13g2_fill_2 FILLER_0_2704 ();
 sg13g2_decap_8 FILLER_0_2725 ();
 sg13g2_decap_8 FILLER_0_2732 ();
 sg13g2_decap_8 FILLER_0_2739 ();
 sg13g2_decap_8 FILLER_0_2746 ();
 sg13g2_decap_8 FILLER_0_2753 ();
 sg13g2_decap_8 FILLER_0_2760 ();
 sg13g2_decap_8 FILLER_0_2767 ();
 sg13g2_decap_8 FILLER_0_2774 ();
 sg13g2_decap_8 FILLER_0_2781 ();
 sg13g2_decap_8 FILLER_0_2788 ();
 sg13g2_decap_4 FILLER_0_2795 ();
 sg13g2_decap_8 FILLER_0_2819 ();
 sg13g2_decap_8 FILLER_0_2826 ();
 sg13g2_decap_8 FILLER_0_2833 ();
 sg13g2_decap_8 FILLER_0_2840 ();
 sg13g2_decap_8 FILLER_0_2847 ();
 sg13g2_fill_2 FILLER_0_2854 ();
 sg13g2_fill_1 FILLER_0_2856 ();
 sg13g2_decap_8 FILLER_0_2884 ();
 sg13g2_decap_8 FILLER_0_2891 ();
 sg13g2_decap_8 FILLER_0_2898 ();
 sg13g2_decap_8 FILLER_0_2905 ();
 sg13g2_decap_4 FILLER_0_2912 ();
 sg13g2_fill_2 FILLER_0_2935 ();
 sg13g2_decap_4 FILLER_0_2947 ();
 sg13g2_fill_1 FILLER_0_2951 ();
 sg13g2_decap_8 FILLER_0_2961 ();
 sg13g2_decap_8 FILLER_0_2968 ();
 sg13g2_decap_8 FILLER_0_2975 ();
 sg13g2_fill_2 FILLER_0_2982 ();
 sg13g2_decap_8 FILLER_0_3011 ();
 sg13g2_decap_8 FILLER_0_3018 ();
 sg13g2_decap_8 FILLER_0_3025 ();
 sg13g2_fill_1 FILLER_0_3032 ();
 sg13g2_decap_8 FILLER_0_3056 ();
 sg13g2_decap_8 FILLER_0_3063 ();
 sg13g2_decap_8 FILLER_0_3070 ();
 sg13g2_decap_8 FILLER_0_3077 ();
 sg13g2_decap_8 FILLER_0_3084 ();
 sg13g2_decap_8 FILLER_0_3091 ();
 sg13g2_decap_8 FILLER_0_3098 ();
 sg13g2_decap_8 FILLER_0_3109 ();
 sg13g2_decap_8 FILLER_0_3116 ();
 sg13g2_decap_8 FILLER_0_3123 ();
 sg13g2_decap_8 FILLER_0_3130 ();
 sg13g2_decap_8 FILLER_0_3137 ();
 sg13g2_decap_8 FILLER_0_3144 ();
 sg13g2_fill_1 FILLER_0_3151 ();
 sg13g2_decap_8 FILLER_0_3179 ();
 sg13g2_decap_8 FILLER_0_3186 ();
 sg13g2_decap_8 FILLER_0_3193 ();
 sg13g2_decap_8 FILLER_0_3200 ();
 sg13g2_decap_8 FILLER_0_3207 ();
 sg13g2_decap_8 FILLER_0_3214 ();
 sg13g2_decap_8 FILLER_0_3221 ();
 sg13g2_decap_8 FILLER_0_3228 ();
 sg13g2_decap_8 FILLER_0_3235 ();
 sg13g2_decap_8 FILLER_0_3242 ();
 sg13g2_decap_8 FILLER_0_3249 ();
 sg13g2_decap_8 FILLER_0_3256 ();
 sg13g2_decap_8 FILLER_0_3263 ();
 sg13g2_decap_8 FILLER_0_3270 ();
 sg13g2_decap_8 FILLER_0_3277 ();
 sg13g2_decap_8 FILLER_0_3284 ();
 sg13g2_decap_8 FILLER_0_3291 ();
 sg13g2_decap_8 FILLER_0_3298 ();
 sg13g2_decap_8 FILLER_0_3305 ();
 sg13g2_decap_8 FILLER_0_3312 ();
 sg13g2_decap_8 FILLER_0_3319 ();
 sg13g2_decap_8 FILLER_0_3326 ();
 sg13g2_decap_8 FILLER_0_3333 ();
 sg13g2_decap_8 FILLER_0_3340 ();
 sg13g2_decap_8 FILLER_0_3347 ();
 sg13g2_decap_8 FILLER_0_3354 ();
 sg13g2_decap_8 FILLER_0_3361 ();
 sg13g2_decap_8 FILLER_0_3368 ();
 sg13g2_decap_8 FILLER_0_3375 ();
 sg13g2_decap_8 FILLER_0_3382 ();
 sg13g2_decap_8 FILLER_0_3389 ();
 sg13g2_decap_8 FILLER_0_3396 ();
 sg13g2_decap_8 FILLER_0_3403 ();
 sg13g2_decap_8 FILLER_0_3410 ();
 sg13g2_decap_8 FILLER_0_3417 ();
 sg13g2_decap_8 FILLER_0_3424 ();
 sg13g2_decap_8 FILLER_0_3431 ();
 sg13g2_decap_8 FILLER_0_3438 ();
 sg13g2_decap_8 FILLER_0_3445 ();
 sg13g2_decap_8 FILLER_0_3452 ();
 sg13g2_decap_8 FILLER_0_3459 ();
 sg13g2_decap_8 FILLER_0_3466 ();
 sg13g2_decap_8 FILLER_0_3473 ();
 sg13g2_decap_8 FILLER_0_3480 ();
 sg13g2_decap_8 FILLER_0_3487 ();
 sg13g2_decap_8 FILLER_0_3494 ();
 sg13g2_decap_8 FILLER_0_3501 ();
 sg13g2_decap_8 FILLER_0_3508 ();
 sg13g2_decap_8 FILLER_0_3515 ();
 sg13g2_decap_8 FILLER_0_3522 ();
 sg13g2_decap_8 FILLER_0_3529 ();
 sg13g2_decap_8 FILLER_0_3536 ();
 sg13g2_decap_8 FILLER_0_3543 ();
 sg13g2_decap_8 FILLER_0_3550 ();
 sg13g2_decap_8 FILLER_0_3557 ();
 sg13g2_decap_8 FILLER_0_3564 ();
 sg13g2_decap_8 FILLER_0_3571 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_fill_2 FILLER_1_99 ();
 sg13g2_fill_2 FILLER_1_128 ();
 sg13g2_fill_1 FILLER_1_130 ();
 sg13g2_fill_1 FILLER_1_144 ();
 sg13g2_fill_1 FILLER_1_149 ();
 sg13g2_fill_2 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_4 FILLER_1_252 ();
 sg13g2_fill_2 FILLER_1_256 ();
 sg13g2_fill_2 FILLER_1_262 ();
 sg13g2_fill_2 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_311 ();
 sg13g2_decap_4 FILLER_1_359 ();
 sg13g2_fill_2 FILLER_1_390 ();
 sg13g2_fill_1 FILLER_1_392 ();
 sg13g2_fill_2 FILLER_1_429 ();
 sg13g2_fill_2 FILLER_1_458 ();
 sg13g2_decap_8 FILLER_1_523 ();
 sg13g2_fill_1 FILLER_1_561 ();
 sg13g2_fill_1 FILLER_1_575 ();
 sg13g2_fill_1 FILLER_1_585 ();
 sg13g2_decap_8 FILLER_1_614 ();
 sg13g2_fill_1 FILLER_1_621 ();
 sg13g2_fill_2 FILLER_1_632 ();
 sg13g2_decap_8 FILLER_1_661 ();
 sg13g2_decap_8 FILLER_1_668 ();
 sg13g2_decap_8 FILLER_1_675 ();
 sg13g2_decap_8 FILLER_1_682 ();
 sg13g2_fill_1 FILLER_1_736 ();
 sg13g2_decap_8 FILLER_1_807 ();
 sg13g2_decap_8 FILLER_1_814 ();
 sg13g2_decap_8 FILLER_1_821 ();
 sg13g2_fill_2 FILLER_1_828 ();
 sg13g2_decap_8 FILLER_1_858 ();
 sg13g2_decap_8 FILLER_1_892 ();
 sg13g2_decap_8 FILLER_1_899 ();
 sg13g2_decap_4 FILLER_1_906 ();
 sg13g2_fill_2 FILLER_1_948 ();
 sg13g2_decap_8 FILLER_1_992 ();
 sg13g2_decap_8 FILLER_1_999 ();
 sg13g2_decap_8 FILLER_1_1006 ();
 sg13g2_fill_2 FILLER_1_1013 ();
 sg13g2_fill_2 FILLER_1_1076 ();
 sg13g2_fill_1 FILLER_1_1105 ();
 sg13g2_decap_4 FILLER_1_1166 ();
 sg13g2_fill_1 FILLER_1_1170 ();
 sg13g2_fill_2 FILLER_1_1232 ();
 sg13g2_decap_8 FILLER_1_1261 ();
 sg13g2_decap_4 FILLER_1_1268 ();
 sg13g2_fill_2 FILLER_1_1272 ();
 sg13g2_fill_2 FILLER_1_1304 ();
 sg13g2_fill_1 FILLER_1_1306 ();
 sg13g2_decap_8 FILLER_1_1313 ();
 sg13g2_decap_4 FILLER_1_1320 ();
 sg13g2_fill_1 FILLER_1_1324 ();
 sg13g2_fill_1 FILLER_1_1382 ();
 sg13g2_decap_4 FILLER_1_1446 ();
 sg13g2_fill_1 FILLER_1_1450 ();
 sg13g2_decap_8 FILLER_1_1464 ();
 sg13g2_decap_8 FILLER_1_1471 ();
 sg13g2_fill_1 FILLER_1_1500 ();
 sg13g2_decap_4 FILLER_1_1528 ();
 sg13g2_fill_1 FILLER_1_1532 ();
 sg13g2_decap_8 FILLER_1_1537 ();
 sg13g2_decap_8 FILLER_1_1544 ();
 sg13g2_fill_2 FILLER_1_1551 ();
 sg13g2_fill_1 FILLER_1_1553 ();
 sg13g2_fill_2 FILLER_1_1581 ();
 sg13g2_fill_1 FILLER_1_1583 ();
 sg13g2_decap_8 FILLER_1_1593 ();
 sg13g2_decap_8 FILLER_1_1600 ();
 sg13g2_decap_4 FILLER_1_1607 ();
 sg13g2_fill_1 FILLER_1_1638 ();
 sg13g2_fill_2 FILLER_1_1648 ();
 sg13g2_fill_2 FILLER_1_1653 ();
 sg13g2_fill_1 FILLER_1_1655 ();
 sg13g2_decap_4 FILLER_1_1660 ();
 sg13g2_fill_1 FILLER_1_1664 ();
 sg13g2_decap_8 FILLER_1_1697 ();
 sg13g2_decap_8 FILLER_1_1704 ();
 sg13g2_decap_4 FILLER_1_1711 ();
 sg13g2_fill_1 FILLER_1_1715 ();
 sg13g2_decap_8 FILLER_1_1743 ();
 sg13g2_decap_8 FILLER_1_1750 ();
 sg13g2_decap_8 FILLER_1_1757 ();
 sg13g2_decap_8 FILLER_1_1764 ();
 sg13g2_decap_8 FILLER_1_1771 ();
 sg13g2_decap_4 FILLER_1_1778 ();
 sg13g2_fill_1 FILLER_1_1782 ();
 sg13g2_decap_8 FILLER_1_1819 ();
 sg13g2_fill_1 FILLER_1_1826 ();
 sg13g2_decap_4 FILLER_1_1830 ();
 sg13g2_fill_1 FILLER_1_1834 ();
 sg13g2_decap_8 FILLER_1_1862 ();
 sg13g2_fill_2 FILLER_1_1869 ();
 sg13g2_decap_8 FILLER_1_1898 ();
 sg13g2_decap_4 FILLER_1_1905 ();
 sg13g2_fill_1 FILLER_1_1909 ();
 sg13g2_decap_8 FILLER_1_1964 ();
 sg13g2_decap_8 FILLER_1_1971 ();
 sg13g2_decap_8 FILLER_1_1978 ();
 sg13g2_decap_4 FILLER_1_1985 ();
 sg13g2_decap_8 FILLER_1_2016 ();
 sg13g2_fill_1 FILLER_1_2023 ();
 sg13g2_decap_8 FILLER_1_2060 ();
 sg13g2_decap_8 FILLER_1_2067 ();
 sg13g2_decap_4 FILLER_1_2074 ();
 sg13g2_fill_2 FILLER_1_2078 ();
 sg13g2_fill_2 FILLER_1_2123 ();
 sg13g2_fill_1 FILLER_1_2125 ();
 sg13g2_decap_4 FILLER_1_2153 ();
 sg13g2_fill_1 FILLER_1_2157 ();
 sg13g2_decap_8 FILLER_1_2161 ();
 sg13g2_decap_4 FILLER_1_2168 ();
 sg13g2_fill_2 FILLER_1_2172 ();
 sg13g2_decap_8 FILLER_1_2241 ();
 sg13g2_decap_8 FILLER_1_2248 ();
 sg13g2_decap_4 FILLER_1_2255 ();
 sg13g2_fill_2 FILLER_1_2259 ();
 sg13g2_decap_8 FILLER_1_2328 ();
 sg13g2_decap_8 FILLER_1_2335 ();
 sg13g2_decap_8 FILLER_1_2342 ();
 sg13g2_decap_4 FILLER_1_2349 ();
 sg13g2_fill_1 FILLER_1_2353 ();
 sg13g2_decap_4 FILLER_1_2391 ();
 sg13g2_fill_1 FILLER_1_2395 ();
 sg13g2_decap_8 FILLER_1_2423 ();
 sg13g2_decap_8 FILLER_1_2430 ();
 sg13g2_fill_2 FILLER_1_2437 ();
 sg13g2_fill_1 FILLER_1_2439 ();
 sg13g2_fill_2 FILLER_1_2450 ();
 sg13g2_fill_1 FILLER_1_2452 ();
 sg13g2_decap_8 FILLER_1_2493 ();
 sg13g2_decap_4 FILLER_1_2500 ();
 sg13g2_fill_2 FILLER_1_2504 ();
 sg13g2_fill_2 FILLER_1_2556 ();
 sg13g2_decap_8 FILLER_1_2585 ();
 sg13g2_decap_4 FILLER_1_2592 ();
 sg13g2_fill_1 FILLER_1_2596 ();
 sg13g2_decap_8 FILLER_1_2645 ();
 sg13g2_decap_8 FILLER_1_2652 ();
 sg13g2_decap_8 FILLER_1_2663 ();
 sg13g2_decap_8 FILLER_1_2670 ();
 sg13g2_decap_8 FILLER_1_2677 ();
 sg13g2_decap_8 FILLER_1_2738 ();
 sg13g2_decap_8 FILLER_1_2745 ();
 sg13g2_decap_4 FILLER_1_2752 ();
 sg13g2_fill_2 FILLER_1_2756 ();
 sg13g2_fill_2 FILLER_1_2781 ();
 sg13g2_decap_8 FILLER_1_2792 ();
 sg13g2_decap_8 FILLER_1_2835 ();
 sg13g2_decap_8 FILLER_1_2842 ();
 sg13g2_fill_1 FILLER_1_2849 ();
 sg13g2_decap_8 FILLER_1_2890 ();
 sg13g2_decap_8 FILLER_1_2897 ();
 sg13g2_fill_1 FILLER_1_2904 ();
 sg13g2_decap_4 FILLER_1_2932 ();
 sg13g2_decap_8 FILLER_1_2967 ();
 sg13g2_decap_4 FILLER_1_2974 ();
 sg13g2_fill_2 FILLER_1_2978 ();
 sg13g2_decap_4 FILLER_1_3025 ();
 sg13g2_decap_8 FILLER_1_3060 ();
 sg13g2_decap_8 FILLER_1_3067 ();
 sg13g2_decap_8 FILLER_1_3074 ();
 sg13g2_fill_1 FILLER_1_3081 ();
 sg13g2_decap_4 FILLER_1_3086 ();
 sg13g2_decap_4 FILLER_1_3127 ();
 sg13g2_decap_8 FILLER_1_3135 ();
 sg13g2_decap_8 FILLER_1_3142 ();
 sg13g2_decap_8 FILLER_1_3185 ();
 sg13g2_decap_8 FILLER_1_3192 ();
 sg13g2_decap_8 FILLER_1_3199 ();
 sg13g2_decap_8 FILLER_1_3206 ();
 sg13g2_decap_8 FILLER_1_3213 ();
 sg13g2_decap_8 FILLER_1_3220 ();
 sg13g2_decap_8 FILLER_1_3227 ();
 sg13g2_decap_8 FILLER_1_3234 ();
 sg13g2_decap_8 FILLER_1_3241 ();
 sg13g2_decap_8 FILLER_1_3248 ();
 sg13g2_decap_8 FILLER_1_3255 ();
 sg13g2_decap_8 FILLER_1_3262 ();
 sg13g2_decap_8 FILLER_1_3269 ();
 sg13g2_decap_8 FILLER_1_3276 ();
 sg13g2_decap_8 FILLER_1_3283 ();
 sg13g2_decap_8 FILLER_1_3290 ();
 sg13g2_decap_8 FILLER_1_3297 ();
 sg13g2_decap_8 FILLER_1_3304 ();
 sg13g2_decap_8 FILLER_1_3311 ();
 sg13g2_decap_8 FILLER_1_3318 ();
 sg13g2_decap_8 FILLER_1_3325 ();
 sg13g2_decap_8 FILLER_1_3332 ();
 sg13g2_decap_8 FILLER_1_3339 ();
 sg13g2_decap_8 FILLER_1_3346 ();
 sg13g2_decap_8 FILLER_1_3353 ();
 sg13g2_decap_8 FILLER_1_3360 ();
 sg13g2_decap_8 FILLER_1_3367 ();
 sg13g2_decap_8 FILLER_1_3374 ();
 sg13g2_decap_8 FILLER_1_3381 ();
 sg13g2_decap_8 FILLER_1_3388 ();
 sg13g2_decap_8 FILLER_1_3395 ();
 sg13g2_decap_8 FILLER_1_3402 ();
 sg13g2_decap_8 FILLER_1_3409 ();
 sg13g2_decap_8 FILLER_1_3416 ();
 sg13g2_decap_8 FILLER_1_3423 ();
 sg13g2_decap_8 FILLER_1_3430 ();
 sg13g2_decap_8 FILLER_1_3437 ();
 sg13g2_decap_8 FILLER_1_3444 ();
 sg13g2_decap_8 FILLER_1_3451 ();
 sg13g2_decap_8 FILLER_1_3458 ();
 sg13g2_decap_8 FILLER_1_3465 ();
 sg13g2_decap_8 FILLER_1_3472 ();
 sg13g2_decap_8 FILLER_1_3479 ();
 sg13g2_decap_8 FILLER_1_3486 ();
 sg13g2_decap_8 FILLER_1_3493 ();
 sg13g2_decap_8 FILLER_1_3500 ();
 sg13g2_decap_8 FILLER_1_3507 ();
 sg13g2_decap_8 FILLER_1_3514 ();
 sg13g2_decap_8 FILLER_1_3521 ();
 sg13g2_decap_8 FILLER_1_3528 ();
 sg13g2_decap_8 FILLER_1_3535 ();
 sg13g2_decap_8 FILLER_1_3542 ();
 sg13g2_decap_8 FILLER_1_3549 ();
 sg13g2_decap_8 FILLER_1_3556 ();
 sg13g2_decap_8 FILLER_1_3563 ();
 sg13g2_decap_8 FILLER_1_3570 ();
 sg13g2_fill_1 FILLER_1_3577 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_49 ();
 sg13g2_fill_1 FILLER_2_51 ();
 sg13g2_fill_1 FILLER_2_92 ();
 sg13g2_fill_2 FILLER_2_133 ();
 sg13g2_fill_1 FILLER_2_144 ();
 sg13g2_fill_2 FILLER_2_181 ();
 sg13g2_fill_1 FILLER_2_183 ();
 sg13g2_fill_2 FILLER_2_194 ();
 sg13g2_fill_1 FILLER_2_196 ();
 sg13g2_fill_1 FILLER_2_210 ();
 sg13g2_fill_1 FILLER_2_239 ();
 sg13g2_fill_2 FILLER_2_365 ();
 sg13g2_fill_2 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_455 ();
 sg13g2_fill_2 FILLER_2_466 ();
 sg13g2_fill_2 FILLER_2_517 ();
 sg13g2_decap_4 FILLER_2_528 ();
 sg13g2_fill_1 FILLER_2_572 ();
 sg13g2_fill_2 FILLER_2_617 ();
 sg13g2_fill_2 FILLER_2_628 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_fill_2 FILLER_2_686 ();
 sg13g2_fill_1 FILLER_2_688 ();
 sg13g2_fill_2 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_4 FILLER_2_826 ();
 sg13g2_fill_2 FILLER_2_830 ();
 sg13g2_fill_1 FILLER_2_850 ();
 sg13g2_decap_8 FILLER_2_897 ();
 sg13g2_decap_8 FILLER_2_904 ();
 sg13g2_decap_4 FILLER_2_911 ();
 sg13g2_fill_2 FILLER_2_915 ();
 sg13g2_fill_2 FILLER_2_947 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_fill_2 FILLER_2_994 ();
 sg13g2_fill_1 FILLER_2_1023 ();
 sg13g2_fill_1 FILLER_2_1107 ();
 sg13g2_decap_8 FILLER_2_1118 ();
 sg13g2_decap_4 FILLER_2_1125 ();
 sg13g2_fill_1 FILLER_2_1129 ();
 sg13g2_decap_4 FILLER_2_1240 ();
 sg13g2_fill_1 FILLER_2_1244 ();
 sg13g2_decap_4 FILLER_2_1264 ();
 sg13g2_fill_1 FILLER_2_1296 ();
 sg13g2_fill_2 FILLER_2_1420 ();
 sg13g2_decap_8 FILLER_2_1460 ();
 sg13g2_decap_8 FILLER_2_1467 ();
 sg13g2_fill_2 FILLER_2_1474 ();
 sg13g2_fill_1 FILLER_2_1476 ();
 sg13g2_fill_2 FILLER_2_1504 ();
 sg13g2_decap_4 FILLER_2_1542 ();
 sg13g2_fill_1 FILLER_2_1578 ();
 sg13g2_decap_8 FILLER_2_1596 ();
 sg13g2_decap_4 FILLER_2_1603 ();
 sg13g2_fill_2 FILLER_2_1607 ();
 sg13g2_fill_1 FILLER_2_1643 ();
 sg13g2_fill_1 FILLER_2_1659 ();
 sg13g2_decap_8 FILLER_2_1699 ();
 sg13g2_decap_4 FILLER_2_1706 ();
 sg13g2_fill_2 FILLER_2_1710 ();
 sg13g2_fill_1 FILLER_2_1746 ();
 sg13g2_fill_1 FILLER_2_1774 ();
 sg13g2_fill_1 FILLER_2_1825 ();
 sg13g2_decap_8 FILLER_2_1979 ();
 sg13g2_fill_2 FILLER_2_1986 ();
 sg13g2_fill_1 FILLER_2_1988 ();
 sg13g2_fill_2 FILLER_2_2016 ();
 sg13g2_decap_8 FILLER_2_2060 ();
 sg13g2_decap_8 FILLER_2_2067 ();
 sg13g2_fill_1 FILLER_2_2074 ();
 sg13g2_fill_2 FILLER_2_2120 ();
 sg13g2_decap_4 FILLER_2_2149 ();
 sg13g2_fill_1 FILLER_2_2153 ();
 sg13g2_decap_4 FILLER_2_2167 ();
 sg13g2_fill_2 FILLER_2_2202 ();
 sg13g2_decap_8 FILLER_2_2325 ();
 sg13g2_decap_8 FILLER_2_2332 ();
 sg13g2_decap_4 FILLER_2_2339 ();
 sg13g2_fill_2 FILLER_2_2383 ();
 sg13g2_fill_1 FILLER_2_2385 ();
 sg13g2_decap_8 FILLER_2_2411 ();
 sg13g2_decap_8 FILLER_2_2418 ();
 sg13g2_decap_8 FILLER_2_2425 ();
 sg13g2_fill_2 FILLER_2_2494 ();
 sg13g2_fill_1 FILLER_2_2496 ();
 sg13g2_fill_1 FILLER_2_2538 ();
 sg13g2_decap_8 FILLER_2_2566 ();
 sg13g2_decap_8 FILLER_2_2573 ();
 sg13g2_decap_8 FILLER_2_2580 ();
 sg13g2_fill_1 FILLER_2_2587 ();
 sg13g2_fill_1 FILLER_2_2629 ();
 sg13g2_fill_2 FILLER_2_2697 ();
 sg13g2_decap_8 FILLER_2_2730 ();
 sg13g2_decap_8 FILLER_2_2737 ();
 sg13g2_decap_8 FILLER_2_2744 ();
 sg13g2_decap_8 FILLER_2_2751 ();
 sg13g2_fill_1 FILLER_2_2758 ();
 sg13g2_fill_2 FILLER_2_2790 ();
 sg13g2_fill_1 FILLER_2_2842 ();
 sg13g2_decap_8 FILLER_2_2890 ();
 sg13g2_fill_2 FILLER_2_2897 ();
 sg13g2_fill_1 FILLER_2_2899 ();
 sg13g2_decap_8 FILLER_2_2962 ();
 sg13g2_fill_2 FILLER_2_2969 ();
 sg13g2_decap_4 FILLER_2_3018 ();
 sg13g2_fill_1 FILLER_2_3022 ();
 sg13g2_decap_8 FILLER_2_3069 ();
 sg13g2_fill_1 FILLER_2_3076 ();
 sg13g2_decap_4 FILLER_2_3140 ();
 sg13g2_decap_8 FILLER_2_3177 ();
 sg13g2_decap_8 FILLER_2_3184 ();
 sg13g2_decap_8 FILLER_2_3191 ();
 sg13g2_decap_8 FILLER_2_3198 ();
 sg13g2_decap_8 FILLER_2_3205 ();
 sg13g2_decap_8 FILLER_2_3212 ();
 sg13g2_decap_8 FILLER_2_3219 ();
 sg13g2_decap_8 FILLER_2_3226 ();
 sg13g2_decap_8 FILLER_2_3233 ();
 sg13g2_decap_8 FILLER_2_3240 ();
 sg13g2_decap_8 FILLER_2_3247 ();
 sg13g2_decap_8 FILLER_2_3254 ();
 sg13g2_decap_8 FILLER_2_3261 ();
 sg13g2_decap_8 FILLER_2_3268 ();
 sg13g2_decap_8 FILLER_2_3275 ();
 sg13g2_decap_8 FILLER_2_3282 ();
 sg13g2_decap_8 FILLER_2_3289 ();
 sg13g2_decap_8 FILLER_2_3296 ();
 sg13g2_decap_8 FILLER_2_3303 ();
 sg13g2_decap_8 FILLER_2_3310 ();
 sg13g2_decap_8 FILLER_2_3317 ();
 sg13g2_decap_8 FILLER_2_3324 ();
 sg13g2_decap_8 FILLER_2_3331 ();
 sg13g2_decap_8 FILLER_2_3338 ();
 sg13g2_decap_8 FILLER_2_3345 ();
 sg13g2_decap_8 FILLER_2_3352 ();
 sg13g2_decap_8 FILLER_2_3359 ();
 sg13g2_decap_8 FILLER_2_3366 ();
 sg13g2_decap_8 FILLER_2_3373 ();
 sg13g2_decap_8 FILLER_2_3380 ();
 sg13g2_decap_8 FILLER_2_3387 ();
 sg13g2_decap_8 FILLER_2_3394 ();
 sg13g2_decap_8 FILLER_2_3401 ();
 sg13g2_decap_8 FILLER_2_3408 ();
 sg13g2_decap_8 FILLER_2_3415 ();
 sg13g2_decap_8 FILLER_2_3422 ();
 sg13g2_decap_8 FILLER_2_3429 ();
 sg13g2_decap_8 FILLER_2_3436 ();
 sg13g2_decap_8 FILLER_2_3443 ();
 sg13g2_decap_8 FILLER_2_3450 ();
 sg13g2_decap_8 FILLER_2_3457 ();
 sg13g2_decap_8 FILLER_2_3464 ();
 sg13g2_decap_8 FILLER_2_3471 ();
 sg13g2_decap_8 FILLER_2_3478 ();
 sg13g2_decap_8 FILLER_2_3485 ();
 sg13g2_decap_8 FILLER_2_3492 ();
 sg13g2_decap_8 FILLER_2_3499 ();
 sg13g2_decap_8 FILLER_2_3506 ();
 sg13g2_decap_8 FILLER_2_3513 ();
 sg13g2_decap_8 FILLER_2_3520 ();
 sg13g2_decap_8 FILLER_2_3527 ();
 sg13g2_decap_8 FILLER_2_3534 ();
 sg13g2_decap_8 FILLER_2_3541 ();
 sg13g2_decap_8 FILLER_2_3548 ();
 sg13g2_decap_8 FILLER_2_3555 ();
 sg13g2_decap_8 FILLER_2_3562 ();
 sg13g2_decap_8 FILLER_2_3569 ();
 sg13g2_fill_2 FILLER_2_3576 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_fill_2 FILLER_3_49 ();
 sg13g2_fill_1 FILLER_3_51 ();
 sg13g2_fill_2 FILLER_3_136 ();
 sg13g2_fill_1 FILLER_3_138 ();
 sg13g2_fill_2 FILLER_3_189 ();
 sg13g2_fill_1 FILLER_3_191 ();
 sg13g2_fill_1 FILLER_3_251 ();
 sg13g2_fill_2 FILLER_3_443 ();
 sg13g2_fill_1 FILLER_3_472 ();
 sg13g2_fill_2 FILLER_3_514 ();
 sg13g2_fill_2 FILLER_3_530 ();
 sg13g2_fill_1 FILLER_3_532 ();
 sg13g2_fill_1 FILLER_3_583 ();
 sg13g2_fill_2 FILLER_3_591 ();
 sg13g2_fill_1 FILLER_3_593 ();
 sg13g2_decap_8 FILLER_3_671 ();
 sg13g2_decap_8 FILLER_3_678 ();
 sg13g2_fill_2 FILLER_3_685 ();
 sg13g2_fill_1 FILLER_3_728 ();
 sg13g2_fill_1 FILLER_3_743 ();
 sg13g2_decap_8 FILLER_3_803 ();
 sg13g2_fill_2 FILLER_3_810 ();
 sg13g2_fill_1 FILLER_3_812 ();
 sg13g2_fill_2 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_856 ();
 sg13g2_fill_2 FILLER_3_866 ();
 sg13g2_fill_1 FILLER_3_868 ();
 sg13g2_decap_8 FILLER_3_905 ();
 sg13g2_decap_8 FILLER_3_912 ();
 sg13g2_fill_2 FILLER_3_963 ();
 sg13g2_fill_1 FILLER_3_965 ();
 sg13g2_decap_8 FILLER_3_1007 ();
 sg13g2_fill_2 FILLER_3_1014 ();
 sg13g2_fill_1 FILLER_3_1026 ();
 sg13g2_fill_1 FILLER_3_1052 ();
 sg13g2_decap_8 FILLER_3_1107 ();
 sg13g2_decap_8 FILLER_3_1114 ();
 sg13g2_decap_8 FILLER_3_1121 ();
 sg13g2_decap_4 FILLER_3_1128 ();
 sg13g2_fill_1 FILLER_3_1132 ();
 sg13g2_fill_2 FILLER_3_1137 ();
 sg13g2_fill_1 FILLER_3_1139 ();
 sg13g2_fill_2 FILLER_3_1153 ();
 sg13g2_fill_1 FILLER_3_1155 ();
 sg13g2_decap_4 FILLER_3_1190 ();
 sg13g2_decap_4 FILLER_3_1203 ();
 sg13g2_fill_1 FILLER_3_1207 ();
 sg13g2_fill_1 FILLER_3_1221 ();
 sg13g2_fill_2 FILLER_3_1309 ();
 sg13g2_decap_4 FILLER_3_1315 ();
 sg13g2_decap_4 FILLER_3_1370 ();
 sg13g2_fill_1 FILLER_3_1374 ();
 sg13g2_decap_4 FILLER_3_1417 ();
 sg13g2_fill_1 FILLER_3_1421 ();
 sg13g2_fill_2 FILLER_3_1440 ();
 sg13g2_fill_1 FILLER_3_1442 ();
 sg13g2_decap_8 FILLER_3_1452 ();
 sg13g2_decap_8 FILLER_3_1459 ();
 sg13g2_decap_8 FILLER_3_1466 ();
 sg13g2_fill_2 FILLER_3_1473 ();
 sg13g2_fill_1 FILLER_3_1511 ();
 sg13g2_fill_1 FILLER_3_1530 ();
 sg13g2_decap_8 FILLER_3_1594 ();
 sg13g2_fill_1 FILLER_3_1601 ();
 sg13g2_fill_2 FILLER_3_1656 ();
 sg13g2_fill_2 FILLER_3_1702 ();
 sg13g2_fill_1 FILLER_3_1704 ();
 sg13g2_fill_1 FILLER_3_1745 ();
 sg13g2_fill_2 FILLER_3_1813 ();
 sg13g2_fill_2 FILLER_3_1871 ();
 sg13g2_fill_1 FILLER_3_1873 ();
 sg13g2_decap_4 FILLER_3_1912 ();
 sg13g2_fill_1 FILLER_3_1979 ();
 sg13g2_decap_8 FILLER_3_2062 ();
 sg13g2_decap_8 FILLER_3_2069 ();
 sg13g2_fill_1 FILLER_3_2089 ();
 sg13g2_fill_2 FILLER_3_2117 ();
 sg13g2_fill_1 FILLER_3_2119 ();
 sg13g2_fill_1 FILLER_3_2154 ();
 sg13g2_decap_8 FILLER_3_2244 ();
 sg13g2_fill_1 FILLER_3_2251 ();
 sg13g2_fill_1 FILLER_3_2285 ();
 sg13g2_fill_2 FILLER_3_2295 ();
 sg13g2_decap_8 FILLER_3_2338 ();
 sg13g2_decap_8 FILLER_3_2345 ();
 sg13g2_fill_1 FILLER_3_2356 ();
 sg13g2_decap_4 FILLER_3_2425 ();
 sg13g2_fill_1 FILLER_3_2429 ();
 sg13g2_fill_2 FILLER_3_2443 ();
 sg13g2_fill_2 FILLER_3_2464 ();
 sg13g2_fill_2 FILLER_3_2493 ();
 sg13g2_fill_1 FILLER_3_2495 ();
 sg13g2_fill_2 FILLER_3_2509 ();
 sg13g2_fill_1 FILLER_3_2511 ();
 sg13g2_fill_2 FILLER_3_2552 ();
 sg13g2_fill_1 FILLER_3_2554 ();
 sg13g2_decap_8 FILLER_3_2574 ();
 sg13g2_decap_8 FILLER_3_2581 ();
 sg13g2_decap_8 FILLER_3_2588 ();
 sg13g2_fill_1 FILLER_3_2646 ();
 sg13g2_decap_4 FILLER_3_2666 ();
 sg13g2_fill_2 FILLER_3_2670 ();
 sg13g2_decap_8 FILLER_3_2725 ();
 sg13g2_fill_1 FILLER_3_2766 ();
 sg13g2_decap_4 FILLER_3_2780 ();
 sg13g2_fill_2 FILLER_3_2784 ();
 sg13g2_fill_2 FILLER_3_2803 ();
 sg13g2_decap_4 FILLER_3_2832 ();
 sg13g2_decap_8 FILLER_3_2849 ();
 sg13g2_fill_1 FILLER_3_2856 ();
 sg13g2_decap_4 FILLER_3_2905 ();
 sg13g2_fill_1 FILLER_3_2913 ();
 sg13g2_fill_2 FILLER_3_2955 ();
 sg13g2_fill_1 FILLER_3_2957 ();
 sg13g2_decap_8 FILLER_3_2967 ();
 sg13g2_decap_4 FILLER_3_2974 ();
 sg13g2_fill_1 FILLER_3_2978 ();
 sg13g2_decap_8 FILLER_3_3019 ();
 sg13g2_fill_2 FILLER_3_3026 ();
 sg13g2_fill_1 FILLER_3_3028 ();
 sg13g2_decap_8 FILLER_3_3060 ();
 sg13g2_decap_8 FILLER_3_3067 ();
 sg13g2_decap_8 FILLER_3_3074 ();
 sg13g2_fill_2 FILLER_3_3111 ();
 sg13g2_fill_1 FILLER_3_3113 ();
 sg13g2_decap_8 FILLER_3_3141 ();
 sg13g2_decap_4 FILLER_3_3148 ();
 sg13g2_fill_2 FILLER_3_3152 ();
 sg13g2_fill_2 FILLER_3_3158 ();
 sg13g2_decap_8 FILLER_3_3185 ();
 sg13g2_decap_8 FILLER_3_3192 ();
 sg13g2_decap_8 FILLER_3_3199 ();
 sg13g2_decap_8 FILLER_3_3206 ();
 sg13g2_decap_8 FILLER_3_3213 ();
 sg13g2_decap_8 FILLER_3_3220 ();
 sg13g2_decap_8 FILLER_3_3227 ();
 sg13g2_decap_8 FILLER_3_3234 ();
 sg13g2_decap_8 FILLER_3_3241 ();
 sg13g2_decap_8 FILLER_3_3248 ();
 sg13g2_decap_8 FILLER_3_3255 ();
 sg13g2_decap_8 FILLER_3_3262 ();
 sg13g2_decap_8 FILLER_3_3269 ();
 sg13g2_decap_8 FILLER_3_3276 ();
 sg13g2_decap_8 FILLER_3_3283 ();
 sg13g2_decap_8 FILLER_3_3290 ();
 sg13g2_decap_8 FILLER_3_3297 ();
 sg13g2_decap_8 FILLER_3_3304 ();
 sg13g2_decap_8 FILLER_3_3311 ();
 sg13g2_decap_8 FILLER_3_3318 ();
 sg13g2_decap_8 FILLER_3_3325 ();
 sg13g2_decap_8 FILLER_3_3332 ();
 sg13g2_decap_8 FILLER_3_3339 ();
 sg13g2_decap_8 FILLER_3_3346 ();
 sg13g2_decap_8 FILLER_3_3353 ();
 sg13g2_decap_8 FILLER_3_3360 ();
 sg13g2_decap_8 FILLER_3_3367 ();
 sg13g2_decap_8 FILLER_3_3374 ();
 sg13g2_decap_8 FILLER_3_3381 ();
 sg13g2_decap_8 FILLER_3_3388 ();
 sg13g2_decap_8 FILLER_3_3395 ();
 sg13g2_decap_8 FILLER_3_3402 ();
 sg13g2_decap_8 FILLER_3_3409 ();
 sg13g2_decap_8 FILLER_3_3416 ();
 sg13g2_decap_8 FILLER_3_3423 ();
 sg13g2_decap_8 FILLER_3_3430 ();
 sg13g2_decap_8 FILLER_3_3437 ();
 sg13g2_decap_8 FILLER_3_3444 ();
 sg13g2_decap_8 FILLER_3_3451 ();
 sg13g2_decap_8 FILLER_3_3458 ();
 sg13g2_decap_8 FILLER_3_3465 ();
 sg13g2_decap_8 FILLER_3_3472 ();
 sg13g2_decap_8 FILLER_3_3479 ();
 sg13g2_decap_8 FILLER_3_3486 ();
 sg13g2_decap_8 FILLER_3_3493 ();
 sg13g2_decap_8 FILLER_3_3500 ();
 sg13g2_decap_8 FILLER_3_3507 ();
 sg13g2_decap_8 FILLER_3_3514 ();
 sg13g2_decap_8 FILLER_3_3521 ();
 sg13g2_decap_8 FILLER_3_3528 ();
 sg13g2_decap_8 FILLER_3_3535 ();
 sg13g2_decap_8 FILLER_3_3542 ();
 sg13g2_decap_8 FILLER_3_3549 ();
 sg13g2_decap_8 FILLER_3_3556 ();
 sg13g2_decap_8 FILLER_3_3563 ();
 sg13g2_decap_8 FILLER_3_3570 ();
 sg13g2_fill_1 FILLER_3_3577 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_fill_2 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_99 ();
 sg13g2_fill_1 FILLER_4_142 ();
 sg13g2_decap_8 FILLER_4_188 ();
 sg13g2_decap_4 FILLER_4_244 ();
 sg13g2_fill_2 FILLER_4_261 ();
 sg13g2_fill_1 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_fill_2 FILLER_4_316 ();
 sg13g2_fill_1 FILLER_4_327 ();
 sg13g2_fill_2 FILLER_4_364 ();
 sg13g2_fill_1 FILLER_4_366 ();
 sg13g2_fill_2 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_406 ();
 sg13g2_fill_2 FILLER_4_421 ();
 sg13g2_fill_1 FILLER_4_423 ();
 sg13g2_fill_1 FILLER_4_443 ();
 sg13g2_fill_2 FILLER_4_476 ();
 sg13g2_fill_1 FILLER_4_478 ();
 sg13g2_fill_1 FILLER_4_516 ();
 sg13g2_decap_8 FILLER_4_526 ();
 sg13g2_fill_1 FILLER_4_556 ();
 sg13g2_fill_2 FILLER_4_575 ();
 sg13g2_decap_8 FILLER_4_601 ();
 sg13g2_fill_2 FILLER_4_608 ();
 sg13g2_fill_1 FILLER_4_610 ();
 sg13g2_decap_8 FILLER_4_675 ();
 sg13g2_decap_8 FILLER_4_682 ();
 sg13g2_decap_8 FILLER_4_689 ();
 sg13g2_fill_1 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_803 ();
 sg13g2_decap_8 FILLER_4_911 ();
 sg13g2_decap_8 FILLER_4_918 ();
 sg13g2_fill_2 FILLER_4_925 ();
 sg13g2_fill_1 FILLER_4_932 ();
 sg13g2_decap_8 FILLER_4_937 ();
 sg13g2_fill_2 FILLER_4_944 ();
 sg13g2_fill_1 FILLER_4_946 ();
 sg13g2_decap_8 FILLER_4_999 ();
 sg13g2_decap_8 FILLER_4_1006 ();
 sg13g2_decap_4 FILLER_4_1013 ();
 sg13g2_decap_8 FILLER_4_1035 ();
 sg13g2_decap_4 FILLER_4_1042 ();
 sg13g2_fill_2 FILLER_4_1088 ();
 sg13g2_fill_2 FILLER_4_1125 ();
 sg13g2_fill_1 FILLER_4_1127 ();
 sg13g2_fill_1 FILLER_4_1166 ();
 sg13g2_decap_8 FILLER_4_1176 ();
 sg13g2_decap_4 FILLER_4_1187 ();
 sg13g2_fill_2 FILLER_4_1191 ();
 sg13g2_decap_4 FILLER_4_1198 ();
 sg13g2_fill_2 FILLER_4_1202 ();
 sg13g2_decap_8 FILLER_4_1217 ();
 sg13g2_decap_8 FILLER_4_1224 ();
 sg13g2_decap_4 FILLER_4_1231 ();
 sg13g2_fill_1 FILLER_4_1235 ();
 sg13g2_decap_4 FILLER_4_1255 ();
 sg13g2_decap_4 FILLER_4_1287 ();
 sg13g2_fill_1 FILLER_4_1291 ();
 sg13g2_fill_2 FILLER_4_1351 ();
 sg13g2_decap_8 FILLER_4_1366 ();
 sg13g2_fill_1 FILLER_4_1373 ();
 sg13g2_fill_2 FILLER_4_1383 ();
 sg13g2_fill_2 FILLER_4_1391 ();
 sg13g2_decap_4 FILLER_4_1434 ();
 sg13g2_fill_1 FILLER_4_1451 ();
 sg13g2_fill_2 FILLER_4_1465 ();
 sg13g2_fill_2 FILLER_4_1507 ();
 sg13g2_fill_1 FILLER_4_1509 ();
 sg13g2_decap_8 FILLER_4_1533 ();
 sg13g2_decap_8 FILLER_4_1540 ();
 sg13g2_decap_4 FILLER_4_1547 ();
 sg13g2_decap_4 FILLER_4_1588 ();
 sg13g2_decap_8 FILLER_4_1596 ();
 sg13g2_decap_8 FILLER_4_1603 ();
 sg13g2_fill_1 FILLER_4_1610 ();
 sg13g2_fill_2 FILLER_4_1630 ();
 sg13g2_fill_2 FILLER_4_1640 ();
 sg13g2_fill_2 FILLER_4_1670 ();
 sg13g2_fill_1 FILLER_4_1672 ();
 sg13g2_decap_8 FILLER_4_1705 ();
 sg13g2_fill_1 FILLER_4_1740 ();
 sg13g2_fill_2 FILLER_4_1750 ();
 sg13g2_fill_1 FILLER_4_1764 ();
 sg13g2_decap_8 FILLER_4_1774 ();
 sg13g2_decap_8 FILLER_4_1781 ();
 sg13g2_fill_1 FILLER_4_1803 ();
 sg13g2_fill_2 FILLER_4_1809 ();
 sg13g2_decap_4 FILLER_4_1820 ();
 sg13g2_fill_1 FILLER_4_1824 ();
 sg13g2_decap_4 FILLER_4_1830 ();
 sg13g2_fill_2 FILLER_4_1853 ();
 sg13g2_fill_1 FILLER_4_1855 ();
 sg13g2_decap_8 FILLER_4_1866 ();
 sg13g2_decap_8 FILLER_4_1873 ();
 sg13g2_decap_8 FILLER_4_1880 ();
 sg13g2_decap_4 FILLER_4_1887 ();
 sg13g2_fill_2 FILLER_4_1891 ();
 sg13g2_fill_2 FILLER_4_1976 ();
 sg13g2_decap_4 FILLER_4_1983 ();
 sg13g2_decap_4 FILLER_4_2008 ();
 sg13g2_fill_1 FILLER_4_2012 ();
 sg13g2_decap_4 FILLER_4_2019 ();
 sg13g2_fill_1 FILLER_4_2023 ();
 sg13g2_decap_8 FILLER_4_2062 ();
 sg13g2_decap_8 FILLER_4_2069 ();
 sg13g2_fill_2 FILLER_4_2076 ();
 sg13g2_fill_1 FILLER_4_2078 ();
 sg13g2_decap_4 FILLER_4_2099 ();
 sg13g2_fill_1 FILLER_4_2103 ();
 sg13g2_fill_2 FILLER_4_2122 ();
 sg13g2_fill_2 FILLER_4_2134 ();
 sg13g2_fill_1 FILLER_4_2136 ();
 sg13g2_fill_2 FILLER_4_2161 ();
 sg13g2_fill_2 FILLER_4_2173 ();
 sg13g2_fill_1 FILLER_4_2175 ();
 sg13g2_fill_2 FILLER_4_2190 ();
 sg13g2_fill_2 FILLER_4_2200 ();
 sg13g2_fill_1 FILLER_4_2202 ();
 sg13g2_fill_2 FILLER_4_2208 ();
 sg13g2_fill_1 FILLER_4_2210 ();
 sg13g2_decap_4 FILLER_4_2224 ();
 sg13g2_fill_2 FILLER_4_2228 ();
 sg13g2_decap_4 FILLER_4_2239 ();
 sg13g2_fill_2 FILLER_4_2243 ();
 sg13g2_decap_4 FILLER_4_2271 ();
 sg13g2_decap_4 FILLER_4_2281 ();
 sg13g2_decap_4 FILLER_4_2292 ();
 sg13g2_fill_1 FILLER_4_2296 ();
 sg13g2_fill_2 FILLER_4_2305 ();
 sg13g2_fill_2 FILLER_4_2313 ();
 sg13g2_decap_8 FILLER_4_2342 ();
 sg13g2_decap_8 FILLER_4_2349 ();
 sg13g2_decap_8 FILLER_4_2356 ();
 sg13g2_fill_2 FILLER_4_2363 ();
 sg13g2_fill_1 FILLER_4_2365 ();
 sg13g2_fill_1 FILLER_4_2370 ();
 sg13g2_decap_4 FILLER_4_2408 ();
 sg13g2_decap_8 FILLER_4_2439 ();
 sg13g2_decap_4 FILLER_4_2446 ();
 sg13g2_decap_4 FILLER_4_2454 ();
 sg13g2_fill_2 FILLER_4_2458 ();
 sg13g2_decap_8 FILLER_4_2481 ();
 sg13g2_decap_8 FILLER_4_2488 ();
 sg13g2_decap_8 FILLER_4_2495 ();
 sg13g2_decap_4 FILLER_4_2502 ();
 sg13g2_fill_2 FILLER_4_2506 ();
 sg13g2_fill_2 FILLER_4_2512 ();
 sg13g2_fill_1 FILLER_4_2514 ();
 sg13g2_decap_8 FILLER_4_2550 ();
 sg13g2_decap_8 FILLER_4_2557 ();
 sg13g2_fill_1 FILLER_4_2564 ();
 sg13g2_decap_8 FILLER_4_2569 ();
 sg13g2_decap_8 FILLER_4_2576 ();
 sg13g2_decap_8 FILLER_4_2583 ();
 sg13g2_decap_4 FILLER_4_2590 ();
 sg13g2_fill_2 FILLER_4_2594 ();
 sg13g2_decap_8 FILLER_4_2632 ();
 sg13g2_decap_8 FILLER_4_2639 ();
 sg13g2_decap_8 FILLER_4_2646 ();
 sg13g2_decap_8 FILLER_4_2653 ();
 sg13g2_decap_8 FILLER_4_2660 ();
 sg13g2_fill_2 FILLER_4_2667 ();
 sg13g2_fill_1 FILLER_4_2683 ();
 sg13g2_decap_8 FILLER_4_2730 ();
 sg13g2_fill_1 FILLER_4_2737 ();
 sg13g2_decap_8 FILLER_4_2765 ();
 sg13g2_decap_8 FILLER_4_2772 ();
 sg13g2_decap_8 FILLER_4_2779 ();
 sg13g2_decap_8 FILLER_4_2786 ();
 sg13g2_fill_2 FILLER_4_2793 ();
 sg13g2_decap_8 FILLER_4_2825 ();
 sg13g2_decap_8 FILLER_4_2832 ();
 sg13g2_decap_8 FILLER_4_2839 ();
 sg13g2_fill_1 FILLER_4_2846 ();
 sg13g2_fill_1 FILLER_4_2857 ();
 sg13g2_decap_8 FILLER_4_2885 ();
 sg13g2_decap_8 FILLER_4_2892 ();
 sg13g2_decap_8 FILLER_4_2899 ();
 sg13g2_decap_8 FILLER_4_2906 ();
 sg13g2_decap_8 FILLER_4_2913 ();
 sg13g2_decap_4 FILLER_4_2920 ();
 sg13g2_decap_8 FILLER_4_2950 ();
 sg13g2_decap_8 FILLER_4_2957 ();
 sg13g2_decap_8 FILLER_4_2964 ();
 sg13g2_fill_2 FILLER_4_2971 ();
 sg13g2_decap_8 FILLER_4_3017 ();
 sg13g2_fill_1 FILLER_4_3024 ();
 sg13g2_fill_2 FILLER_4_3038 ();
 sg13g2_fill_1 FILLER_4_3040 ();
 sg13g2_decap_8 FILLER_4_3071 ();
 sg13g2_decap_8 FILLER_4_3078 ();
 sg13g2_decap_4 FILLER_4_3085 ();
 sg13g2_fill_2 FILLER_4_3089 ();
 sg13g2_fill_2 FILLER_4_3104 ();
 sg13g2_fill_1 FILLER_4_3106 ();
 sg13g2_decap_8 FILLER_4_3137 ();
 sg13g2_fill_2 FILLER_4_3144 ();
 sg13g2_fill_1 FILLER_4_3146 ();
 sg13g2_decap_8 FILLER_4_3211 ();
 sg13g2_decap_8 FILLER_4_3218 ();
 sg13g2_decap_8 FILLER_4_3225 ();
 sg13g2_decap_8 FILLER_4_3232 ();
 sg13g2_decap_8 FILLER_4_3239 ();
 sg13g2_decap_8 FILLER_4_3246 ();
 sg13g2_decap_8 FILLER_4_3253 ();
 sg13g2_decap_8 FILLER_4_3260 ();
 sg13g2_decap_8 FILLER_4_3267 ();
 sg13g2_decap_8 FILLER_4_3274 ();
 sg13g2_decap_8 FILLER_4_3281 ();
 sg13g2_decap_8 FILLER_4_3288 ();
 sg13g2_decap_8 FILLER_4_3295 ();
 sg13g2_decap_8 FILLER_4_3302 ();
 sg13g2_fill_2 FILLER_4_3309 ();
 sg13g2_decap_8 FILLER_4_3315 ();
 sg13g2_decap_8 FILLER_4_3322 ();
 sg13g2_decap_8 FILLER_4_3329 ();
 sg13g2_decap_8 FILLER_4_3336 ();
 sg13g2_decap_8 FILLER_4_3343 ();
 sg13g2_decap_8 FILLER_4_3350 ();
 sg13g2_decap_8 FILLER_4_3357 ();
 sg13g2_decap_8 FILLER_4_3364 ();
 sg13g2_decap_8 FILLER_4_3371 ();
 sg13g2_decap_8 FILLER_4_3378 ();
 sg13g2_decap_8 FILLER_4_3385 ();
 sg13g2_decap_8 FILLER_4_3392 ();
 sg13g2_decap_8 FILLER_4_3399 ();
 sg13g2_decap_8 FILLER_4_3406 ();
 sg13g2_decap_8 FILLER_4_3413 ();
 sg13g2_decap_8 FILLER_4_3420 ();
 sg13g2_decap_8 FILLER_4_3427 ();
 sg13g2_decap_8 FILLER_4_3434 ();
 sg13g2_decap_8 FILLER_4_3441 ();
 sg13g2_decap_8 FILLER_4_3448 ();
 sg13g2_decap_8 FILLER_4_3455 ();
 sg13g2_decap_8 FILLER_4_3462 ();
 sg13g2_decap_8 FILLER_4_3469 ();
 sg13g2_decap_8 FILLER_4_3476 ();
 sg13g2_decap_8 FILLER_4_3483 ();
 sg13g2_decap_8 FILLER_4_3490 ();
 sg13g2_decap_8 FILLER_4_3497 ();
 sg13g2_decap_8 FILLER_4_3504 ();
 sg13g2_decap_8 FILLER_4_3511 ();
 sg13g2_decap_8 FILLER_4_3518 ();
 sg13g2_decap_8 FILLER_4_3525 ();
 sg13g2_decap_8 FILLER_4_3532 ();
 sg13g2_decap_8 FILLER_4_3539 ();
 sg13g2_decap_8 FILLER_4_3546 ();
 sg13g2_decap_8 FILLER_4_3553 ();
 sg13g2_decap_8 FILLER_4_3560 ();
 sg13g2_decap_8 FILLER_4_3567 ();
 sg13g2_decap_4 FILLER_4_3574 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_4 FILLER_5_49 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_143 ();
 sg13g2_decap_8 FILLER_5_150 ();
 sg13g2_decap_4 FILLER_5_157 ();
 sg13g2_fill_1 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_1 FILLER_5_230 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_decap_4 FILLER_5_257 ();
 sg13g2_fill_1 FILLER_5_261 ();
 sg13g2_fill_2 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_fill_2 FILLER_5_331 ();
 sg13g2_fill_1 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_fill_1 FILLER_5_367 ();
 sg13g2_fill_2 FILLER_5_435 ();
 sg13g2_fill_1 FILLER_5_437 ();
 sg13g2_fill_1 FILLER_5_443 ();
 sg13g2_decap_8 FILLER_5_523 ();
 sg13g2_fill_1 FILLER_5_530 ();
 sg13g2_fill_2 FILLER_5_580 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_4 FILLER_5_602 ();
 sg13g2_fill_1 FILLER_5_606 ();
 sg13g2_decap_4 FILLER_5_620 ();
 sg13g2_fill_1 FILLER_5_624 ();
 sg13g2_fill_2 FILLER_5_659 ();
 sg13g2_fill_1 FILLER_5_661 ();
 sg13g2_decap_8 FILLER_5_666 ();
 sg13g2_decap_8 FILLER_5_673 ();
 sg13g2_decap_8 FILLER_5_680 ();
 sg13g2_decap_4 FILLER_5_687 ();
 sg13g2_fill_1 FILLER_5_691 ();
 sg13g2_fill_1 FILLER_5_723 ();
 sg13g2_fill_1 FILLER_5_754 ();
 sg13g2_fill_2 FILLER_5_766 ();
 sg13g2_decap_8 FILLER_5_800 ();
 sg13g2_decap_8 FILLER_5_807 ();
 sg13g2_decap_4 FILLER_5_814 ();
 sg13g2_fill_1 FILLER_5_823 ();
 sg13g2_decap_4 FILLER_5_866 ();
 sg13g2_fill_1 FILLER_5_895 ();
 sg13g2_fill_2 FILLER_5_905 ();
 sg13g2_decap_8 FILLER_5_910 ();
 sg13g2_decap_8 FILLER_5_917 ();
 sg13g2_fill_2 FILLER_5_924 ();
 sg13g2_fill_1 FILLER_5_926 ();
 sg13g2_decap_8 FILLER_5_931 ();
 sg13g2_decap_8 FILLER_5_938 ();
 sg13g2_fill_2 FILLER_5_945 ();
 sg13g2_decap_8 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_fill_1 FILLER_5_1055 ();
 sg13g2_decap_8 FILLER_5_1098 ();
 sg13g2_fill_2 FILLER_5_1105 ();
 sg13g2_fill_1 FILLER_5_1107 ();
 sg13g2_decap_4 FILLER_5_1121 ();
 sg13g2_fill_2 FILLER_5_1125 ();
 sg13g2_decap_4 FILLER_5_1131 ();
 sg13g2_fill_2 FILLER_5_1135 ();
 sg13g2_decap_8 FILLER_5_1198 ();
 sg13g2_decap_8 FILLER_5_1205 ();
 sg13g2_decap_8 FILLER_5_1212 ();
 sg13g2_decap_8 FILLER_5_1219 ();
 sg13g2_decap_8 FILLER_5_1226 ();
 sg13g2_decap_8 FILLER_5_1233 ();
 sg13g2_decap_4 FILLER_5_1240 ();
 sg13g2_fill_1 FILLER_5_1244 ();
 sg13g2_decap_8 FILLER_5_1253 ();
 sg13g2_decap_8 FILLER_5_1260 ();
 sg13g2_decap_8 FILLER_5_1267 ();
 sg13g2_decap_8 FILLER_5_1274 ();
 sg13g2_decap_8 FILLER_5_1281 ();
 sg13g2_decap_8 FILLER_5_1288 ();
 sg13g2_decap_4 FILLER_5_1295 ();
 sg13g2_fill_1 FILLER_5_1299 ();
 sg13g2_fill_2 FILLER_5_1309 ();
 sg13g2_decap_8 FILLER_5_1333 ();
 sg13g2_decap_4 FILLER_5_1340 ();
 sg13g2_fill_1 FILLER_5_1344 ();
 sg13g2_decap_8 FILLER_5_1358 ();
 sg13g2_decap_8 FILLER_5_1365 ();
 sg13g2_decap_4 FILLER_5_1372 ();
 sg13g2_fill_2 FILLER_5_1376 ();
 sg13g2_decap_8 FILLER_5_1381 ();
 sg13g2_fill_2 FILLER_5_1388 ();
 sg13g2_fill_2 FILLER_5_1425 ();
 sg13g2_decap_4 FILLER_5_1437 ();
 sg13g2_fill_2 FILLER_5_1441 ();
 sg13g2_decap_8 FILLER_5_1480 ();
 sg13g2_decap_8 FILLER_5_1533 ();
 sg13g2_decap_8 FILLER_5_1540 ();
 sg13g2_fill_2 FILLER_5_1547 ();
 sg13g2_decap_4 FILLER_5_1554 ();
 sg13g2_decap_8 FILLER_5_1603 ();
 sg13g2_fill_1 FILLER_5_1610 ();
 sg13g2_fill_2 FILLER_5_1635 ();
 sg13g2_fill_1 FILLER_5_1637 ();
 sg13g2_fill_2 FILLER_5_1680 ();
 sg13g2_fill_1 FILLER_5_1682 ();
 sg13g2_decap_8 FILLER_5_1693 ();
 sg13g2_decap_8 FILLER_5_1700 ();
 sg13g2_fill_1 FILLER_5_1744 ();
 sg13g2_fill_2 FILLER_5_1752 ();
 sg13g2_fill_2 FILLER_5_1763 ();
 sg13g2_decap_8 FILLER_5_1771 ();
 sg13g2_decap_8 FILLER_5_1778 ();
 sg13g2_decap_8 FILLER_5_1785 ();
 sg13g2_fill_2 FILLER_5_1792 ();
 sg13g2_fill_1 FILLER_5_1794 ();
 sg13g2_fill_1 FILLER_5_1800 ();
 sg13g2_decap_4 FILLER_5_1820 ();
 sg13g2_fill_1 FILLER_5_1837 ();
 sg13g2_fill_2 FILLER_5_1847 ();
 sg13g2_fill_1 FILLER_5_1855 ();
 sg13g2_decap_4 FILLER_5_1870 ();
 sg13g2_decap_8 FILLER_5_1882 ();
 sg13g2_fill_2 FILLER_5_1889 ();
 sg13g2_decap_4 FILLER_5_1895 ();
 sg13g2_fill_1 FILLER_5_1927 ();
 sg13g2_decap_8 FILLER_5_1967 ();
 sg13g2_decap_8 FILLER_5_1974 ();
 sg13g2_fill_2 FILLER_5_1981 ();
 sg13g2_fill_1 FILLER_5_1983 ();
 sg13g2_decap_8 FILLER_5_1988 ();
 sg13g2_decap_4 FILLER_5_1995 ();
 sg13g2_fill_1 FILLER_5_1999 ();
 sg13g2_decap_8 FILLER_5_2008 ();
 sg13g2_fill_2 FILLER_5_2015 ();
 sg13g2_fill_2 FILLER_5_2025 ();
 sg13g2_decap_4 FILLER_5_2062 ();
 sg13g2_fill_2 FILLER_5_2079 ();
 sg13g2_decap_4 FILLER_5_2133 ();
 sg13g2_fill_1 FILLER_5_2137 ();
 sg13g2_fill_2 FILLER_5_2156 ();
 sg13g2_fill_2 FILLER_5_2161 ();
 sg13g2_fill_1 FILLER_5_2163 ();
 sg13g2_fill_2 FILLER_5_2169 ();
 sg13g2_fill_1 FILLER_5_2180 ();
 sg13g2_fill_2 FILLER_5_2191 ();
 sg13g2_fill_1 FILLER_5_2202 ();
 sg13g2_decap_8 FILLER_5_2215 ();
 sg13g2_decap_8 FILLER_5_2228 ();
 sg13g2_decap_8 FILLER_5_2235 ();
 sg13g2_fill_2 FILLER_5_2242 ();
 sg13g2_fill_1 FILLER_5_2244 ();
 sg13g2_decap_8 FILLER_5_2285 ();
 sg13g2_fill_2 FILLER_5_2292 ();
 sg13g2_fill_1 FILLER_5_2294 ();
 sg13g2_decap_8 FILLER_5_2346 ();
 sg13g2_decap_8 FILLER_5_2353 ();
 sg13g2_decap_8 FILLER_5_2360 ();
 sg13g2_decap_4 FILLER_5_2367 ();
 sg13g2_fill_1 FILLER_5_2371 ();
 sg13g2_fill_2 FILLER_5_2407 ();
 sg13g2_fill_1 FILLER_5_2409 ();
 sg13g2_decap_8 FILLER_5_2444 ();
 sg13g2_decap_8 FILLER_5_2451 ();
 sg13g2_decap_8 FILLER_5_2458 ();
 sg13g2_fill_2 FILLER_5_2484 ();
 sg13g2_decap_8 FILLER_5_2507 ();
 sg13g2_decap_4 FILLER_5_2514 ();
 sg13g2_fill_2 FILLER_5_2518 ();
 sg13g2_decap_8 FILLER_5_2529 ();
 sg13g2_fill_2 FILLER_5_2536 ();
 sg13g2_decap_8 FILLER_5_2548 ();
 sg13g2_fill_1 FILLER_5_2555 ();
 sg13g2_decap_8 FILLER_5_2583 ();
 sg13g2_decap_4 FILLER_5_2590 ();
 sg13g2_decap_4 FILLER_5_2604 ();
 sg13g2_fill_1 FILLER_5_2608 ();
 sg13g2_decap_8 FILLER_5_2632 ();
 sg13g2_decap_8 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_4 FILLER_5_2653 ();
 sg13g2_fill_2 FILLER_5_2657 ();
 sg13g2_decap_8 FILLER_5_2721 ();
 sg13g2_decap_4 FILLER_5_2728 ();
 sg13g2_fill_2 FILLER_5_2732 ();
 sg13g2_decap_8 FILLER_5_2766 ();
 sg13g2_decap_8 FILLER_5_2773 ();
 sg13g2_decap_8 FILLER_5_2780 ();
 sg13g2_decap_8 FILLER_5_2787 ();
 sg13g2_decap_8 FILLER_5_2794 ();
 sg13g2_fill_2 FILLER_5_2801 ();
 sg13g2_fill_1 FILLER_5_2803 ();
 sg13g2_decap_8 FILLER_5_2808 ();
 sg13g2_fill_2 FILLER_5_2815 ();
 sg13g2_decap_8 FILLER_5_2840 ();
 sg13g2_decap_4 FILLER_5_2847 ();
 sg13g2_decap_8 FILLER_5_2855 ();
 sg13g2_fill_1 FILLER_5_2866 ();
 sg13g2_decap_8 FILLER_5_2885 ();
 sg13g2_decap_8 FILLER_5_2892 ();
 sg13g2_decap_4 FILLER_5_2899 ();
 sg13g2_fill_1 FILLER_5_2903 ();
 sg13g2_decap_8 FILLER_5_2925 ();
 sg13g2_decap_8 FILLER_5_2932 ();
 sg13g2_decap_4 FILLER_5_2939 ();
 sg13g2_decap_8 FILLER_5_2953 ();
 sg13g2_decap_8 FILLER_5_2969 ();
 sg13g2_decap_8 FILLER_5_2976 ();
 sg13g2_decap_8 FILLER_5_3017 ();
 sg13g2_decap_8 FILLER_5_3024 ();
 sg13g2_fill_2 FILLER_5_3041 ();
 sg13g2_fill_1 FILLER_5_3043 ();
 sg13g2_decap_8 FILLER_5_3075 ();
 sg13g2_decap_8 FILLER_5_3082 ();
 sg13g2_decap_4 FILLER_5_3098 ();
 sg13g2_fill_1 FILLER_5_3121 ();
 sg13g2_decap_8 FILLER_5_3131 ();
 sg13g2_fill_1 FILLER_5_3138 ();
 sg13g2_decap_8 FILLER_5_3143 ();
 sg13g2_fill_2 FILLER_5_3150 ();
 sg13g2_fill_2 FILLER_5_3165 ();
 sg13g2_fill_1 FILLER_5_3190 ();
 sg13g2_decap_8 FILLER_5_3204 ();
 sg13g2_decap_8 FILLER_5_3211 ();
 sg13g2_decap_8 FILLER_5_3218 ();
 sg13g2_decap_8 FILLER_5_3225 ();
 sg13g2_decap_8 FILLER_5_3232 ();
 sg13g2_decap_8 FILLER_5_3239 ();
 sg13g2_decap_8 FILLER_5_3246 ();
 sg13g2_decap_8 FILLER_5_3253 ();
 sg13g2_fill_2 FILLER_5_3260 ();
 sg13g2_decap_8 FILLER_5_3271 ();
 sg13g2_decap_8 FILLER_5_3278 ();
 sg13g2_decap_8 FILLER_5_3285 ();
 sg13g2_decap_8 FILLER_5_3292 ();
 sg13g2_decap_8 FILLER_5_3299 ();
 sg13g2_decap_8 FILLER_5_3332 ();
 sg13g2_decap_8 FILLER_5_3339 ();
 sg13g2_decap_8 FILLER_5_3346 ();
 sg13g2_decap_8 FILLER_5_3353 ();
 sg13g2_decap_8 FILLER_5_3360 ();
 sg13g2_decap_8 FILLER_5_3367 ();
 sg13g2_decap_8 FILLER_5_3374 ();
 sg13g2_decap_8 FILLER_5_3381 ();
 sg13g2_decap_8 FILLER_5_3388 ();
 sg13g2_decap_8 FILLER_5_3395 ();
 sg13g2_decap_8 FILLER_5_3402 ();
 sg13g2_decap_8 FILLER_5_3409 ();
 sg13g2_decap_8 FILLER_5_3416 ();
 sg13g2_decap_8 FILLER_5_3423 ();
 sg13g2_decap_8 FILLER_5_3430 ();
 sg13g2_decap_8 FILLER_5_3437 ();
 sg13g2_decap_8 FILLER_5_3444 ();
 sg13g2_decap_8 FILLER_5_3451 ();
 sg13g2_decap_8 FILLER_5_3458 ();
 sg13g2_decap_8 FILLER_5_3465 ();
 sg13g2_decap_8 FILLER_5_3472 ();
 sg13g2_decap_8 FILLER_5_3479 ();
 sg13g2_decap_8 FILLER_5_3486 ();
 sg13g2_decap_8 FILLER_5_3493 ();
 sg13g2_decap_8 FILLER_5_3500 ();
 sg13g2_decap_8 FILLER_5_3507 ();
 sg13g2_decap_8 FILLER_5_3514 ();
 sg13g2_decap_8 FILLER_5_3521 ();
 sg13g2_decap_8 FILLER_5_3528 ();
 sg13g2_decap_8 FILLER_5_3535 ();
 sg13g2_decap_8 FILLER_5_3542 ();
 sg13g2_decap_8 FILLER_5_3549 ();
 sg13g2_decap_8 FILLER_5_3556 ();
 sg13g2_decap_8 FILLER_5_3563 ();
 sg13g2_decap_8 FILLER_5_3570 ();
 sg13g2_fill_1 FILLER_5_3577 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_49 ();
 sg13g2_fill_1 FILLER_6_51 ();
 sg13g2_fill_2 FILLER_6_145 ();
 sg13g2_fill_1 FILLER_6_147 ();
 sg13g2_decap_4 FILLER_6_161 ();
 sg13g2_fill_1 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_202 ();
 sg13g2_decap_8 FILLER_6_209 ();
 sg13g2_fill_1 FILLER_6_216 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_decap_4 FILLER_6_235 ();
 sg13g2_fill_2 FILLER_6_239 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_251 ();
 sg13g2_decap_4 FILLER_6_258 ();
 sg13g2_decap_8 FILLER_6_309 ();
 sg13g2_decap_8 FILLER_6_316 ();
 sg13g2_decap_8 FILLER_6_323 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_348 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_fill_1 FILLER_6_376 ();
 sg13g2_fill_1 FILLER_6_381 ();
 sg13g2_fill_2 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_443 ();
 sg13g2_fill_1 FILLER_6_450 ();
 sg13g2_fill_2 FILLER_6_477 ();
 sg13g2_fill_1 FILLER_6_479 ();
 sg13g2_fill_1 FILLER_6_522 ();
 sg13g2_fill_1 FILLER_6_554 ();
 sg13g2_fill_1 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_fill_1 FILLER_6_650 ();
 sg13g2_decap_8 FILLER_6_656 ();
 sg13g2_decap_4 FILLER_6_663 ();
 sg13g2_fill_2 FILLER_6_667 ();
 sg13g2_decap_8 FILLER_6_678 ();
 sg13g2_decap_8 FILLER_6_685 ();
 sg13g2_decap_8 FILLER_6_692 ();
 sg13g2_decap_4 FILLER_6_699 ();
 sg13g2_decap_4 FILLER_6_757 ();
 sg13g2_fill_2 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_4 FILLER_6_826 ();
 sg13g2_fill_2 FILLER_6_830 ();
 sg13g2_fill_1 FILLER_6_837 ();
 sg13g2_fill_2 FILLER_6_846 ();
 sg13g2_decap_8 FILLER_6_857 ();
 sg13g2_decap_8 FILLER_6_864 ();
 sg13g2_fill_2 FILLER_6_876 ();
 sg13g2_fill_1 FILLER_6_878 ();
 sg13g2_fill_2 FILLER_6_916 ();
 sg13g2_fill_2 FILLER_6_946 ();
 sg13g2_fill_1 FILLER_6_992 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_8 FILLER_6_1019 ();
 sg13g2_decap_8 FILLER_6_1026 ();
 sg13g2_decap_4 FILLER_6_1033 ();
 sg13g2_fill_1 FILLER_6_1037 ();
 sg13g2_decap_8 FILLER_6_1047 ();
 sg13g2_decap_4 FILLER_6_1054 ();
 sg13g2_fill_2 FILLER_6_1063 ();
 sg13g2_fill_1 FILLER_6_1098 ();
 sg13g2_decap_8 FILLER_6_1136 ();
 sg13g2_fill_1 FILLER_6_1143 ();
 sg13g2_fill_2 FILLER_6_1148 ();
 sg13g2_decap_8 FILLER_6_1160 ();
 sg13g2_decap_4 FILLER_6_1167 ();
 sg13g2_decap_8 FILLER_6_1184 ();
 sg13g2_decap_8 FILLER_6_1191 ();
 sg13g2_fill_1 FILLER_6_1208 ();
 sg13g2_decap_4 FILLER_6_1222 ();
 sg13g2_fill_2 FILLER_6_1226 ();
 sg13g2_fill_2 FILLER_6_1255 ();
 sg13g2_decap_4 FILLER_6_1266 ();
 sg13g2_fill_1 FILLER_6_1270 ();
 sg13g2_fill_1 FILLER_6_1312 ();
 sg13g2_decap_4 FILLER_6_1350 ();
 sg13g2_fill_2 FILLER_6_1354 ();
 sg13g2_decap_8 FILLER_6_1369 ();
 sg13g2_fill_2 FILLER_6_1376 ();
 sg13g2_fill_1 FILLER_6_1378 ();
 sg13g2_decap_8 FILLER_6_1383 ();
 sg13g2_fill_2 FILLER_6_1390 ();
 sg13g2_fill_2 FILLER_6_1418 ();
 sg13g2_fill_2 FILLER_6_1466 ();
 sg13g2_fill_1 FILLER_6_1468 ();
 sg13g2_decap_4 FILLER_6_1482 ();
 sg13g2_fill_2 FILLER_6_1486 ();
 sg13g2_decap_4 FILLER_6_1525 ();
 sg13g2_fill_2 FILLER_6_1529 ();
 sg13g2_fill_2 FILLER_6_1579 ();
 sg13g2_decap_4 FILLER_6_1593 ();
 sg13g2_fill_2 FILLER_6_1597 ();
 sg13g2_decap_8 FILLER_6_1611 ();
 sg13g2_fill_2 FILLER_6_1661 ();
 sg13g2_fill_1 FILLER_6_1663 ();
 sg13g2_fill_1 FILLER_6_1681 ();
 sg13g2_fill_2 FILLER_6_1687 ();
 sg13g2_fill_1 FILLER_6_1689 ();
 sg13g2_fill_2 FILLER_6_1716 ();
 sg13g2_fill_2 FILLER_6_1724 ();
 sg13g2_fill_1 FILLER_6_1747 ();
 sg13g2_fill_1 FILLER_6_1763 ();
 sg13g2_decap_8 FILLER_6_1790 ();
 sg13g2_decap_8 FILLER_6_1797 ();
 sg13g2_fill_1 FILLER_6_1804 ();
 sg13g2_decap_8 FILLER_6_1818 ();
 sg13g2_decap_8 FILLER_6_1825 ();
 sg13g2_decap_8 FILLER_6_1832 ();
 sg13g2_decap_8 FILLER_6_1839 ();
 sg13g2_decap_8 FILLER_6_1882 ();
 sg13g2_decap_8 FILLER_6_1889 ();
 sg13g2_fill_1 FILLER_6_1896 ();
 sg13g2_fill_2 FILLER_6_1901 ();
 sg13g2_decap_8 FILLER_6_1941 ();
 sg13g2_decap_8 FILLER_6_1948 ();
 sg13g2_decap_8 FILLER_6_1955 ();
 sg13g2_decap_8 FILLER_6_1962 ();
 sg13g2_decap_8 FILLER_6_1969 ();
 sg13g2_fill_1 FILLER_6_1976 ();
 sg13g2_fill_1 FILLER_6_2020 ();
 sg13g2_decap_4 FILLER_6_2037 ();
 sg13g2_decap_8 FILLER_6_2056 ();
 sg13g2_decap_8 FILLER_6_2063 ();
 sg13g2_decap_4 FILLER_6_2070 ();
 sg13g2_fill_1 FILLER_6_2074 ();
 sg13g2_decap_8 FILLER_6_2119 ();
 sg13g2_fill_2 FILLER_6_2130 ();
 sg13g2_decap_8 FILLER_6_2168 ();
 sg13g2_decap_8 FILLER_6_2175 ();
 sg13g2_fill_2 FILLER_6_2187 ();
 sg13g2_decap_8 FILLER_6_2230 ();
 sg13g2_decap_8 FILLER_6_2237 ();
 sg13g2_decap_8 FILLER_6_2244 ();
 sg13g2_decap_4 FILLER_6_2251 ();
 sg13g2_fill_1 FILLER_6_2271 ();
 sg13g2_decap_8 FILLER_6_2291 ();
 sg13g2_decap_8 FILLER_6_2298 ();
 sg13g2_fill_2 FILLER_6_2311 ();
 sg13g2_decap_8 FILLER_6_2354 ();
 sg13g2_decap_8 FILLER_6_2361 ();
 sg13g2_decap_4 FILLER_6_2368 ();
 sg13g2_fill_2 FILLER_6_2394 ();
 sg13g2_decap_4 FILLER_6_2406 ();
 sg13g2_fill_1 FILLER_6_2410 ();
 sg13g2_fill_2 FILLER_6_2431 ();
 sg13g2_fill_1 FILLER_6_2446 ();
 sg13g2_decap_4 FILLER_6_2457 ();
 sg13g2_decap_8 FILLER_6_2507 ();
 sg13g2_decap_8 FILLER_6_2514 ();
 sg13g2_decap_8 FILLER_6_2521 ();
 sg13g2_decap_8 FILLER_6_2528 ();
 sg13g2_fill_1 FILLER_6_2589 ();
 sg13g2_decap_8 FILLER_6_2639 ();
 sg13g2_decap_8 FILLER_6_2646 ();
 sg13g2_decap_4 FILLER_6_2653 ();
 sg13g2_decap_4 FILLER_6_2694 ();
 sg13g2_fill_2 FILLER_6_2698 ();
 sg13g2_decap_8 FILLER_6_2709 ();
 sg13g2_decap_8 FILLER_6_2716 ();
 sg13g2_decap_8 FILLER_6_2723 ();
 sg13g2_decap_8 FILLER_6_2730 ();
 sg13g2_decap_4 FILLER_6_2737 ();
 sg13g2_fill_2 FILLER_6_2741 ();
 sg13g2_decap_8 FILLER_6_2747 ();
 sg13g2_fill_2 FILLER_6_2791 ();
 sg13g2_fill_2 FILLER_6_2820 ();
 sg13g2_decap_8 FILLER_6_2874 ();
 sg13g2_decap_8 FILLER_6_2881 ();
 sg13g2_decap_8 FILLER_6_2888 ();
 sg13g2_decap_4 FILLER_6_2895 ();
 sg13g2_fill_1 FILLER_6_2899 ();
 sg13g2_fill_2 FILLER_6_2927 ();
 sg13g2_decap_8 FILLER_6_2938 ();
 sg13g2_decap_8 FILLER_6_2972 ();
 sg13g2_decap_4 FILLER_6_2979 ();
 sg13g2_fill_1 FILLER_6_2993 ();
 sg13g2_decap_8 FILLER_6_3007 ();
 sg13g2_decap_8 FILLER_6_3014 ();
 sg13g2_decap_8 FILLER_6_3021 ();
 sg13g2_fill_2 FILLER_6_3028 ();
 sg13g2_decap_8 FILLER_6_3040 ();
 sg13g2_fill_1 FILLER_6_3047 ();
 sg13g2_decap_4 FILLER_6_3058 ();
 sg13g2_fill_2 FILLER_6_3062 ();
 sg13g2_decap_4 FILLER_6_3073 ();
 sg13g2_fill_1 FILLER_6_3077 ();
 sg13g2_fill_2 FILLER_6_3105 ();
 sg13g2_decap_4 FILLER_6_3148 ();
 sg13g2_decap_4 FILLER_6_3161 ();
 sg13g2_fill_2 FILLER_6_3165 ();
 sg13g2_decap_8 FILLER_6_3176 ();
 sg13g2_decap_8 FILLER_6_3183 ();
 sg13g2_fill_1 FILLER_6_3194 ();
 sg13g2_decap_8 FILLER_6_3222 ();
 sg13g2_decap_8 FILLER_6_3229 ();
 sg13g2_decap_8 FILLER_6_3236 ();
 sg13g2_decap_8 FILLER_6_3243 ();
 sg13g2_decap_8 FILLER_6_3277 ();
 sg13g2_decap_8 FILLER_6_3284 ();
 sg13g2_decap_8 FILLER_6_3291 ();
 sg13g2_decap_8 FILLER_6_3329 ();
 sg13g2_decap_8 FILLER_6_3336 ();
 sg13g2_decap_8 FILLER_6_3343 ();
 sg13g2_decap_8 FILLER_6_3350 ();
 sg13g2_decap_4 FILLER_6_3357 ();
 sg13g2_decap_8 FILLER_6_3388 ();
 sg13g2_decap_8 FILLER_6_3395 ();
 sg13g2_decap_8 FILLER_6_3402 ();
 sg13g2_decap_8 FILLER_6_3409 ();
 sg13g2_fill_2 FILLER_6_3416 ();
 sg13g2_decap_8 FILLER_6_3427 ();
 sg13g2_decap_8 FILLER_6_3434 ();
 sg13g2_decap_8 FILLER_6_3441 ();
 sg13g2_decap_8 FILLER_6_3448 ();
 sg13g2_decap_8 FILLER_6_3455 ();
 sg13g2_decap_8 FILLER_6_3462 ();
 sg13g2_decap_8 FILLER_6_3469 ();
 sg13g2_decap_8 FILLER_6_3476 ();
 sg13g2_decap_8 FILLER_6_3483 ();
 sg13g2_decap_8 FILLER_6_3490 ();
 sg13g2_decap_8 FILLER_6_3497 ();
 sg13g2_decap_8 FILLER_6_3504 ();
 sg13g2_decap_8 FILLER_6_3511 ();
 sg13g2_decap_8 FILLER_6_3518 ();
 sg13g2_decap_8 FILLER_6_3525 ();
 sg13g2_decap_8 FILLER_6_3532 ();
 sg13g2_decap_8 FILLER_6_3539 ();
 sg13g2_decap_8 FILLER_6_3546 ();
 sg13g2_decap_8 FILLER_6_3553 ();
 sg13g2_decap_8 FILLER_6_3560 ();
 sg13g2_decap_8 FILLER_6_3567 ();
 sg13g2_decap_4 FILLER_6_3574 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_35 ();
 sg13g2_fill_2 FILLER_7_64 ();
 sg13g2_fill_1 FILLER_7_66 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_135 ();
 sg13g2_fill_1 FILLER_7_162 ();
 sg13g2_decap_8 FILLER_7_204 ();
 sg13g2_fill_2 FILLER_7_211 ();
 sg13g2_fill_2 FILLER_7_239 ();
 sg13g2_fill_2 FILLER_7_244 ();
 sg13g2_fill_1 FILLER_7_246 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_fill_2 FILLER_7_325 ();
 sg13g2_fill_2 FILLER_7_330 ();
 sg13g2_fill_1 FILLER_7_332 ();
 sg13g2_fill_2 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_4 FILLER_7_375 ();
 sg13g2_fill_1 FILLER_7_379 ();
 sg13g2_fill_2 FILLER_7_437 ();
 sg13g2_fill_2 FILLER_7_451 ();
 sg13g2_fill_1 FILLER_7_453 ();
 sg13g2_decap_4 FILLER_7_522 ();
 sg13g2_fill_2 FILLER_7_526 ();
 sg13g2_fill_1 FILLER_7_555 ();
 sg13g2_fill_1 FILLER_7_592 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_4 FILLER_7_651 ();
 sg13g2_fill_2 FILLER_7_655 ();
 sg13g2_decap_8 FILLER_7_661 ();
 sg13g2_decap_8 FILLER_7_696 ();
 sg13g2_fill_2 FILLER_7_703 ();
 sg13g2_fill_1 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_750 ();
 sg13g2_decap_8 FILLER_7_757 ();
 sg13g2_decap_4 FILLER_7_764 ();
 sg13g2_fill_2 FILLER_7_768 ();
 sg13g2_decap_8 FILLER_7_773 ();
 sg13g2_fill_2 FILLER_7_780 ();
 sg13g2_fill_1 FILLER_7_782 ();
 sg13g2_decap_8 FILLER_7_792 ();
 sg13g2_decap_8 FILLER_7_799 ();
 sg13g2_decap_8 FILLER_7_806 ();
 sg13g2_decap_8 FILLER_7_813 ();
 sg13g2_fill_1 FILLER_7_825 ();
 sg13g2_fill_2 FILLER_7_830 ();
 sg13g2_decap_8 FILLER_7_841 ();
 sg13g2_decap_8 FILLER_7_848 ();
 sg13g2_decap_4 FILLER_7_855 ();
 sg13g2_fill_1 FILLER_7_859 ();
 sg13g2_fill_2 FILLER_7_870 ();
 sg13g2_fill_2 FILLER_7_941 ();
 sg13g2_fill_2 FILLER_7_948 ();
 sg13g2_fill_1 FILLER_7_950 ();
 sg13g2_fill_2 FILLER_7_983 ();
 sg13g2_decap_8 FILLER_7_999 ();
 sg13g2_decap_8 FILLER_7_1006 ();
 sg13g2_fill_1 FILLER_7_1013 ();
 sg13g2_decap_4 FILLER_7_1024 ();
 sg13g2_fill_2 FILLER_7_1028 ();
 sg13g2_decap_4 FILLER_7_1058 ();
 sg13g2_decap_4 FILLER_7_1069 ();
 sg13g2_fill_1 FILLER_7_1073 ();
 sg13g2_fill_2 FILLER_7_1078 ();
 sg13g2_decap_4 FILLER_7_1102 ();
 sg13g2_fill_2 FILLER_7_1106 ();
 sg13g2_decap_8 FILLER_7_1141 ();
 sg13g2_decap_8 FILLER_7_1148 ();
 sg13g2_decap_8 FILLER_7_1155 ();
 sg13g2_decap_8 FILLER_7_1162 ();
 sg13g2_fill_2 FILLER_7_1169 ();
 sg13g2_fill_1 FILLER_7_1171 ();
 sg13g2_decap_8 FILLER_7_1176 ();
 sg13g2_decap_4 FILLER_7_1183 ();
 sg13g2_fill_1 FILLER_7_1187 ();
 sg13g2_fill_1 FILLER_7_1197 ();
 sg13g2_decap_8 FILLER_7_1211 ();
 sg13g2_decap_4 FILLER_7_1218 ();
 sg13g2_fill_1 FILLER_7_1222 ();
 sg13g2_fill_1 FILLER_7_1263 ();
 sg13g2_fill_2 FILLER_7_1304 ();
 sg13g2_fill_1 FILLER_7_1306 ();
 sg13g2_fill_1 FILLER_7_1325 ();
 sg13g2_decap_4 FILLER_7_1354 ();
 sg13g2_fill_1 FILLER_7_1358 ();
 sg13g2_decap_8 FILLER_7_1369 ();
 sg13g2_fill_1 FILLER_7_1376 ();
 sg13g2_decap_8 FILLER_7_1392 ();
 sg13g2_fill_2 FILLER_7_1409 ();
 sg13g2_fill_1 FILLER_7_1411 ();
 sg13g2_fill_2 FILLER_7_1422 ();
 sg13g2_fill_2 FILLER_7_1452 ();
 sg13g2_fill_1 FILLER_7_1454 ();
 sg13g2_decap_8 FILLER_7_1477 ();
 sg13g2_decap_8 FILLER_7_1484 ();
 sg13g2_decap_4 FILLER_7_1491 ();
 sg13g2_fill_1 FILLER_7_1495 ();
 sg13g2_decap_8 FILLER_7_1519 ();
 sg13g2_decap_4 FILLER_7_1526 ();
 sg13g2_fill_1 FILLER_7_1530 ();
 sg13g2_decap_8 FILLER_7_1614 ();
 sg13g2_decap_8 FILLER_7_1652 ();
 sg13g2_decap_4 FILLER_7_1659 ();
 sg13g2_decap_8 FILLER_7_1786 ();
 sg13g2_fill_1 FILLER_7_1793 ();
 sg13g2_decap_4 FILLER_7_1826 ();
 sg13g2_fill_2 FILLER_7_1875 ();
 sg13g2_fill_2 FILLER_7_1891 ();
 sg13g2_fill_2 FILLER_7_1920 ();
 sg13g2_fill_1 FILLER_7_1922 ();
 sg13g2_decap_8 FILLER_7_1949 ();
 sg13g2_decap_8 FILLER_7_1956 ();
 sg13g2_decap_8 FILLER_7_1963 ();
 sg13g2_fill_1 FILLER_7_1970 ();
 sg13g2_fill_1 FILLER_7_1998 ();
 sg13g2_fill_2 FILLER_7_2065 ();
 sg13g2_fill_1 FILLER_7_2067 ();
 sg13g2_fill_2 FILLER_7_2109 ();
 sg13g2_fill_2 FILLER_7_2152 ();
 sg13g2_decap_8 FILLER_7_2167 ();
 sg13g2_decap_8 FILLER_7_2231 ();
 sg13g2_decap_8 FILLER_7_2238 ();
 sg13g2_fill_2 FILLER_7_2245 ();
 sg13g2_fill_2 FILLER_7_2266 ();
 sg13g2_fill_1 FILLER_7_2268 ();
 sg13g2_decap_8 FILLER_7_2282 ();
 sg13g2_decap_8 FILLER_7_2289 ();
 sg13g2_decap_4 FILLER_7_2301 ();
 sg13g2_fill_1 FILLER_7_2305 ();
 sg13g2_decap_8 FILLER_7_2341 ();
 sg13g2_decap_8 FILLER_7_2348 ();
 sg13g2_decap_8 FILLER_7_2355 ();
 sg13g2_fill_2 FILLER_7_2362 ();
 sg13g2_decap_4 FILLER_7_2391 ();
 sg13g2_fill_1 FILLER_7_2395 ();
 sg13g2_fill_2 FILLER_7_2415 ();
 sg13g2_decap_8 FILLER_7_2515 ();
 sg13g2_decap_4 FILLER_7_2522 ();
 sg13g2_fill_1 FILLER_7_2526 ();
 sg13g2_fill_2 FILLER_7_2586 ();
 sg13g2_decap_8 FILLER_7_2651 ();
 sg13g2_decap_4 FILLER_7_2658 ();
 sg13g2_decap_8 FILLER_7_2666 ();
 sg13g2_fill_1 FILLER_7_2673 ();
 sg13g2_fill_2 FILLER_7_2683 ();
 sg13g2_decap_8 FILLER_7_2694 ();
 sg13g2_decap_4 FILLER_7_2701 ();
 sg13g2_fill_2 FILLER_7_2705 ();
 sg13g2_decap_8 FILLER_7_2736 ();
 sg13g2_decap_4 FILLER_7_2743 ();
 sg13g2_decap_8 FILLER_7_2887 ();
 sg13g2_fill_1 FILLER_7_2894 ();
 sg13g2_fill_2 FILLER_7_2936 ();
 sg13g2_fill_1 FILLER_7_2938 ();
 sg13g2_decap_8 FILLER_7_2970 ();
 sg13g2_decap_8 FILLER_7_2977 ();
 sg13g2_decap_4 FILLER_7_2984 ();
 sg13g2_decap_8 FILLER_7_3015 ();
 sg13g2_decap_4 FILLER_7_3022 ();
 sg13g2_fill_2 FILLER_7_3026 ();
 sg13g2_decap_8 FILLER_7_3059 ();
 sg13g2_decap_8 FILLER_7_3066 ();
 sg13g2_fill_1 FILLER_7_3073 ();
 sg13g2_fill_1 FILLER_7_3110 ();
 sg13g2_decap_8 FILLER_7_3161 ();
 sg13g2_decap_8 FILLER_7_3168 ();
 sg13g2_decap_8 FILLER_7_3175 ();
 sg13g2_fill_2 FILLER_7_3182 ();
 sg13g2_fill_1 FILLER_7_3184 ();
 sg13g2_decap_8 FILLER_7_3223 ();
 sg13g2_decap_8 FILLER_7_3230 ();
 sg13g2_fill_2 FILLER_7_3237 ();
 sg13g2_decap_8 FILLER_7_3280 ();
 sg13g2_decap_8 FILLER_7_3287 ();
 sg13g2_fill_2 FILLER_7_3348 ();
 sg13g2_fill_1 FILLER_7_3350 ();
 sg13g2_decap_8 FILLER_7_3391 ();
 sg13g2_decap_4 FILLER_7_3398 ();
 sg13g2_decap_8 FILLER_7_3429 ();
 sg13g2_decap_8 FILLER_7_3436 ();
 sg13g2_decap_8 FILLER_7_3443 ();
 sg13g2_decap_8 FILLER_7_3450 ();
 sg13g2_decap_8 FILLER_7_3457 ();
 sg13g2_decap_8 FILLER_7_3464 ();
 sg13g2_decap_8 FILLER_7_3471 ();
 sg13g2_decap_8 FILLER_7_3478 ();
 sg13g2_decap_4 FILLER_7_3485 ();
 sg13g2_fill_1 FILLER_7_3489 ();
 sg13g2_decap_4 FILLER_7_3499 ();
 sg13g2_fill_1 FILLER_7_3503 ();
 sg13g2_decap_8 FILLER_7_3523 ();
 sg13g2_decap_8 FILLER_7_3530 ();
 sg13g2_decap_8 FILLER_7_3537 ();
 sg13g2_decap_8 FILLER_7_3544 ();
 sg13g2_decap_8 FILLER_7_3551 ();
 sg13g2_decap_8 FILLER_7_3558 ();
 sg13g2_decap_8 FILLER_7_3565 ();
 sg13g2_decap_4 FILLER_7_3572 ();
 sg13g2_fill_2 FILLER_7_3576 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_4 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_fill_2 FILLER_8_130 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_154 ();
 sg13g2_fill_2 FILLER_8_187 ();
 sg13g2_fill_1 FILLER_8_189 ();
 sg13g2_decap_4 FILLER_8_207 ();
 sg13g2_fill_1 FILLER_8_211 ();
 sg13g2_fill_2 FILLER_8_217 ();
 sg13g2_decap_4 FILLER_8_223 ();
 sg13g2_fill_1 FILLER_8_232 ();
 sg13g2_fill_1 FILLER_8_247 ();
 sg13g2_fill_1 FILLER_8_258 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_fill_1 FILLER_8_346 ();
 sg13g2_decap_4 FILLER_8_374 ();
 sg13g2_fill_1 FILLER_8_378 ();
 sg13g2_fill_1 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_4 FILLER_8_518 ();
 sg13g2_fill_1 FILLER_8_578 ();
 sg13g2_fill_2 FILLER_8_601 ();
 sg13g2_fill_1 FILLER_8_603 ();
 sg13g2_decap_8 FILLER_8_626 ();
 sg13g2_decap_8 FILLER_8_633 ();
 sg13g2_fill_1 FILLER_8_640 ();
 sg13g2_decap_4 FILLER_8_645 ();
 sg13g2_fill_2 FILLER_8_649 ();
 sg13g2_fill_1 FILLER_8_707 ();
 sg13g2_fill_2 FILLER_8_713 ();
 sg13g2_fill_1 FILLER_8_733 ();
 sg13g2_decap_8 FILLER_8_745 ();
 sg13g2_decap_8 FILLER_8_752 ();
 sg13g2_decap_4 FILLER_8_786 ();
 sg13g2_fill_1 FILLER_8_790 ();
 sg13g2_decap_8 FILLER_8_800 ();
 sg13g2_fill_1 FILLER_8_807 ();
 sg13g2_decap_8 FILLER_8_849 ();
 sg13g2_fill_1 FILLER_8_873 ();
 sg13g2_fill_2 FILLER_8_914 ();
 sg13g2_fill_2 FILLER_8_923 ();
 sg13g2_decap_8 FILLER_8_929 ();
 sg13g2_decap_8 FILLER_8_936 ();
 sg13g2_decap_8 FILLER_8_943 ();
 sg13g2_fill_2 FILLER_8_950 ();
 sg13g2_fill_2 FILLER_8_956 ();
 sg13g2_fill_1 FILLER_8_958 ();
 sg13g2_fill_2 FILLER_8_1021 ();
 sg13g2_fill_1 FILLER_8_1023 ();
 sg13g2_decap_8 FILLER_8_1075 ();
 sg13g2_decap_4 FILLER_8_1082 ();
 sg13g2_decap_8 FILLER_8_1095 ();
 sg13g2_fill_1 FILLER_8_1102 ();
 sg13g2_decap_8 FILLER_8_1107 ();
 sg13g2_decap_8 FILLER_8_1114 ();
 sg13g2_decap_4 FILLER_8_1121 ();
 sg13g2_fill_2 FILLER_8_1125 ();
 sg13g2_decap_8 FILLER_8_1140 ();
 sg13g2_decap_8 FILLER_8_1147 ();
 sg13g2_decap_8 FILLER_8_1154 ();
 sg13g2_fill_2 FILLER_8_1165 ();
 sg13g2_fill_1 FILLER_8_1167 ();
 sg13g2_decap_8 FILLER_8_1205 ();
 sg13g2_fill_2 FILLER_8_1212 ();
 sg13g2_fill_1 FILLER_8_1269 ();
 sg13g2_fill_1 FILLER_8_1297 ();
 sg13g2_decap_8 FILLER_8_1346 ();
 sg13g2_decap_8 FILLER_8_1353 ();
 sg13g2_fill_1 FILLER_8_1360 ();
 sg13g2_fill_1 FILLER_8_1399 ();
 sg13g2_decap_4 FILLER_8_1450 ();
 sg13g2_fill_1 FILLER_8_1454 ();
 sg13g2_decap_8 FILLER_8_1468 ();
 sg13g2_fill_1 FILLER_8_1475 ();
 sg13g2_fill_2 FILLER_8_1485 ();
 sg13g2_decap_8 FILLER_8_1518 ();
 sg13g2_fill_2 FILLER_8_1525 ();
 sg13g2_fill_1 FILLER_8_1527 ();
 sg13g2_decap_8 FILLER_8_1533 ();
 sg13g2_fill_2 FILLER_8_1540 ();
 sg13g2_fill_1 FILLER_8_1568 ();
 sg13g2_fill_2 FILLER_8_1592 ();
 sg13g2_fill_1 FILLER_8_1594 ();
 sg13g2_fill_1 FILLER_8_1603 ();
 sg13g2_decap_8 FILLER_8_1609 ();
 sg13g2_decap_8 FILLER_8_1616 ();
 sg13g2_fill_2 FILLER_8_1623 ();
 sg13g2_fill_1 FILLER_8_1625 ();
 sg13g2_fill_1 FILLER_8_1631 ();
 sg13g2_fill_2 FILLER_8_1641 ();
 sg13g2_fill_1 FILLER_8_1643 ();
 sg13g2_decap_8 FILLER_8_1653 ();
 sg13g2_decap_8 FILLER_8_1660 ();
 sg13g2_decap_4 FILLER_8_1667 ();
 sg13g2_decap_4 FILLER_8_1675 ();
 sg13g2_fill_1 FILLER_8_1679 ();
 sg13g2_decap_8 FILLER_8_1696 ();
 sg13g2_fill_2 FILLER_8_1703 ();
 sg13g2_fill_2 FILLER_8_1710 ();
 sg13g2_fill_2 FILLER_8_1720 ();
 sg13g2_fill_1 FILLER_8_1722 ();
 sg13g2_decap_8 FILLER_8_1727 ();
 sg13g2_decap_8 FILLER_8_1734 ();
 sg13g2_fill_1 FILLER_8_1741 ();
 sg13g2_decap_8 FILLER_8_1836 ();
 sg13g2_fill_2 FILLER_8_1843 ();
 sg13g2_fill_2 FILLER_8_1886 ();
 sg13g2_fill_2 FILLER_8_1932 ();
 sg13g2_fill_1 FILLER_8_1934 ();
 sg13g2_fill_2 FILLER_8_1962 ();
 sg13g2_fill_1 FILLER_8_1964 ();
 sg13g2_decap_8 FILLER_8_2022 ();
 sg13g2_decap_8 FILLER_8_2029 ();
 sg13g2_fill_2 FILLER_8_2036 ();
 sg13g2_fill_1 FILLER_8_2038 ();
 sg13g2_decap_4 FILLER_8_2054 ();
 sg13g2_decap_8 FILLER_8_2067 ();
 sg13g2_decap_8 FILLER_8_2074 ();
 sg13g2_decap_8 FILLER_8_2081 ();
 sg13g2_decap_4 FILLER_8_2088 ();
 sg13g2_fill_1 FILLER_8_2097 ();
 sg13g2_fill_2 FILLER_8_2116 ();
 sg13g2_decap_8 FILLER_8_2161 ();
 sg13g2_decap_4 FILLER_8_2168 ();
 sg13g2_fill_1 FILLER_8_2172 ();
 sg13g2_fill_1 FILLER_8_2293 ();
 sg13g2_decap_8 FILLER_8_2299 ();
 sg13g2_decap_8 FILLER_8_2306 ();
 sg13g2_decap_4 FILLER_8_2313 ();
 sg13g2_fill_2 FILLER_8_2317 ();
 sg13g2_decap_8 FILLER_8_2346 ();
 sg13g2_decap_4 FILLER_8_2353 ();
 sg13g2_fill_1 FILLER_8_2357 ();
 sg13g2_decap_8 FILLER_8_2418 ();
 sg13g2_fill_2 FILLER_8_2425 ();
 sg13g2_decap_8 FILLER_8_2432 ();
 sg13g2_fill_2 FILLER_8_2439 ();
 sg13g2_fill_1 FILLER_8_2441 ();
 sg13g2_decap_4 FILLER_8_2459 ();
 sg13g2_decap_8 FILLER_8_2509 ();
 sg13g2_decap_8 FILLER_8_2516 ();
 sg13g2_decap_4 FILLER_8_2523 ();
 sg13g2_fill_2 FILLER_8_2527 ();
 sg13g2_fill_2 FILLER_8_2542 ();
 sg13g2_fill_1 FILLER_8_2548 ();
 sg13g2_decap_8 FILLER_8_2574 ();
 sg13g2_decap_4 FILLER_8_2581 ();
 sg13g2_fill_1 FILLER_8_2612 ();
 sg13g2_decap_8 FILLER_8_2640 ();
 sg13g2_decap_8 FILLER_8_2647 ();
 sg13g2_decap_4 FILLER_8_2654 ();
 sg13g2_fill_2 FILLER_8_2658 ();
 sg13g2_fill_2 FILLER_8_2670 ();
 sg13g2_fill_1 FILLER_8_2672 ();
 sg13g2_decap_4 FILLER_8_2682 ();
 sg13g2_fill_2 FILLER_8_2686 ();
 sg13g2_fill_1 FILLER_8_2698 ();
 sg13g2_decap_4 FILLER_8_2739 ();
 sg13g2_fill_2 FILLER_8_2743 ();
 sg13g2_decap_4 FILLER_8_2768 ();
 sg13g2_fill_1 FILLER_8_2772 ();
 sg13g2_decap_8 FILLER_8_2808 ();
 sg13g2_decap_8 FILLER_8_2815 ();
 sg13g2_fill_1 FILLER_8_2863 ();
 sg13g2_decap_8 FILLER_8_2894 ();
 sg13g2_fill_2 FILLER_8_2901 ();
 sg13g2_fill_1 FILLER_8_2903 ();
 sg13g2_fill_2 FILLER_8_2908 ();
 sg13g2_fill_1 FILLER_8_2910 ();
 sg13g2_fill_1 FILLER_8_2942 ();
 sg13g2_fill_2 FILLER_8_2957 ();
 sg13g2_decap_8 FILLER_8_2968 ();
 sg13g2_decap_4 FILLER_8_2975 ();
 sg13g2_fill_2 FILLER_8_3010 ();
 sg13g2_fill_1 FILLER_8_3012 ();
 sg13g2_fill_2 FILLER_8_3076 ();
 sg13g2_fill_1 FILLER_8_3078 ();
 sg13g2_fill_2 FILLER_8_3119 ();
 sg13g2_decap_8 FILLER_8_3161 ();
 sg13g2_decap_4 FILLER_8_3178 ();
 sg13g2_fill_2 FILLER_8_3182 ();
 sg13g2_decap_8 FILLER_8_3221 ();
 sg13g2_decap_8 FILLER_8_3228 ();
 sg13g2_fill_2 FILLER_8_3245 ();
 sg13g2_decap_8 FILLER_8_3278 ();
 sg13g2_decap_8 FILLER_8_3285 ();
 sg13g2_decap_4 FILLER_8_3292 ();
 sg13g2_decap_4 FILLER_8_3352 ();
 sg13g2_fill_2 FILLER_8_3356 ();
 sg13g2_decap_8 FILLER_8_3387 ();
 sg13g2_decap_8 FILLER_8_3394 ();
 sg13g2_fill_2 FILLER_8_3401 ();
 sg13g2_decap_8 FILLER_8_3451 ();
 sg13g2_decap_8 FILLER_8_3458 ();
 sg13g2_decap_8 FILLER_8_3465 ();
 sg13g2_fill_1 FILLER_8_3472 ();
 sg13g2_decap_4 FILLER_8_3504 ();
 sg13g2_fill_1 FILLER_8_3508 ();
 sg13g2_decap_8 FILLER_8_3536 ();
 sg13g2_decap_8 FILLER_8_3543 ();
 sg13g2_decap_8 FILLER_8_3550 ();
 sg13g2_decap_8 FILLER_8_3557 ();
 sg13g2_decap_8 FILLER_8_3564 ();
 sg13g2_decap_8 FILLER_8_3571 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_4 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_39 ();
 sg13g2_fill_1 FILLER_9_48 ();
 sg13g2_fill_2 FILLER_9_103 ();
 sg13g2_fill_1 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_decap_4 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_138 ();
 sg13g2_fill_2 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_145 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_fill_2 FILLER_9_182 ();
 sg13g2_fill_2 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_205 ();
 sg13g2_fill_1 FILLER_9_216 ();
 sg13g2_fill_1 FILLER_9_241 ();
 sg13g2_fill_2 FILLER_9_256 ();
 sg13g2_decap_4 FILLER_9_297 ();
 sg13g2_fill_1 FILLER_9_309 ();
 sg13g2_fill_2 FILLER_9_318 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_358 ();
 sg13g2_fill_2 FILLER_9_374 ();
 sg13g2_fill_1 FILLER_9_385 ();
 sg13g2_fill_2 FILLER_9_394 ();
 sg13g2_fill_1 FILLER_9_400 ();
 sg13g2_fill_1 FILLER_9_415 ();
 sg13g2_fill_1 FILLER_9_439 ();
 sg13g2_fill_2 FILLER_9_449 ();
 sg13g2_fill_1 FILLER_9_451 ();
 sg13g2_decap_8 FILLER_9_470 ();
 sg13g2_fill_2 FILLER_9_503 ();
 sg13g2_fill_1 FILLER_9_505 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_decap_4 FILLER_9_522 ();
 sg13g2_fill_1 FILLER_9_526 ();
 sg13g2_decap_4 FILLER_9_581 ();
 sg13g2_fill_2 FILLER_9_602 ();
 sg13g2_decap_4 FILLER_9_613 ();
 sg13g2_fill_2 FILLER_9_617 ();
 sg13g2_fill_2 FILLER_9_673 ();
 sg13g2_decap_4 FILLER_9_685 ();
 sg13g2_fill_2 FILLER_9_702 ();
 sg13g2_decap_8 FILLER_9_738 ();
 sg13g2_decap_8 FILLER_9_799 ();
 sg13g2_fill_2 FILLER_9_806 ();
 sg13g2_fill_1 FILLER_9_808 ();
 sg13g2_decap_8 FILLER_9_837 ();
 sg13g2_fill_2 FILLER_9_844 ();
 sg13g2_decap_8 FILLER_9_891 ();
 sg13g2_decap_8 FILLER_9_898 ();
 sg13g2_decap_8 FILLER_9_905 ();
 sg13g2_fill_1 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_923 ();
 sg13g2_decap_8 FILLER_9_930 ();
 sg13g2_fill_2 FILLER_9_937 ();
 sg13g2_fill_1 FILLER_9_939 ();
 sg13g2_decap_8 FILLER_9_943 ();
 sg13g2_decap_8 FILLER_9_950 ();
 sg13g2_decap_8 FILLER_9_957 ();
 sg13g2_fill_1 FILLER_9_964 ();
 sg13g2_fill_2 FILLER_9_983 ();
 sg13g2_fill_1 FILLER_9_985 ();
 sg13g2_decap_8 FILLER_9_1014 ();
 sg13g2_decap_8 FILLER_9_1021 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_2 FILLER_9_1055 ();
 sg13g2_fill_1 FILLER_9_1070 ();
 sg13g2_fill_1 FILLER_9_1103 ();
 sg13g2_fill_1 FILLER_9_1118 ();
 sg13g2_decap_4 FILLER_9_1141 ();
 sg13g2_decap_8 FILLER_9_1149 ();
 sg13g2_decap_8 FILLER_9_1198 ();
 sg13g2_decap_4 FILLER_9_1205 ();
 sg13g2_fill_1 FILLER_9_1209 ();
 sg13g2_fill_2 FILLER_9_1238 ();
 sg13g2_fill_1 FILLER_9_1240 ();
 sg13g2_fill_2 FILLER_9_1268 ();
 sg13g2_fill_2 FILLER_9_1301 ();
 sg13g2_decap_8 FILLER_9_1330 ();
 sg13g2_decap_4 FILLER_9_1337 ();
 sg13g2_fill_2 FILLER_9_1341 ();
 sg13g2_decap_8 FILLER_9_1353 ();
 sg13g2_decap_8 FILLER_9_1360 ();
 sg13g2_decap_8 FILLER_9_1367 ();
 sg13g2_decap_4 FILLER_9_1407 ();
 sg13g2_fill_1 FILLER_9_1411 ();
 sg13g2_decap_8 FILLER_9_1453 ();
 sg13g2_decap_8 FILLER_9_1519 ();
 sg13g2_decap_8 FILLER_9_1531 ();
 sg13g2_decap_8 FILLER_9_1538 ();
 sg13g2_decap_8 FILLER_9_1545 ();
 sg13g2_decap_8 FILLER_9_1552 ();
 sg13g2_fill_1 FILLER_9_1559 ();
 sg13g2_decap_8 FILLER_9_1600 ();
 sg13g2_fill_2 FILLER_9_1607 ();
 sg13g2_decap_8 FILLER_9_1615 ();
 sg13g2_decap_4 FILLER_9_1622 ();
 sg13g2_fill_2 FILLER_9_1653 ();
 sg13g2_fill_1 FILLER_9_1655 ();
 sg13g2_decap_8 FILLER_9_1672 ();
 sg13g2_decap_8 FILLER_9_1679 ();
 sg13g2_fill_2 FILLER_9_1686 ();
 sg13g2_decap_8 FILLER_9_1693 ();
 sg13g2_fill_2 FILLER_9_1700 ();
 sg13g2_decap_8 FILLER_9_1739 ();
 sg13g2_fill_2 FILLER_9_1746 ();
 sg13g2_fill_1 FILLER_9_1748 ();
 sg13g2_decap_4 FILLER_9_1759 ();
 sg13g2_fill_1 FILLER_9_1763 ();
 sg13g2_fill_1 FILLER_9_1770 ();
 sg13g2_decap_4 FILLER_9_1780 ();
 sg13g2_decap_4 FILLER_9_1834 ();
 sg13g2_fill_2 FILLER_9_1838 ();
 sg13g2_fill_1 FILLER_9_1885 ();
 sg13g2_decap_4 FILLER_9_1924 ();
 sg13g2_fill_2 FILLER_9_1928 ();
 sg13g2_fill_1 FILLER_9_1935 ();
 sg13g2_decap_4 FILLER_9_1948 ();
 sg13g2_fill_1 FILLER_9_1952 ();
 sg13g2_decap_8 FILLER_9_2012 ();
 sg13g2_decap_8 FILLER_9_2019 ();
 sg13g2_decap_4 FILLER_9_2026 ();
 sg13g2_fill_1 FILLER_9_2030 ();
 sg13g2_decap_8 FILLER_9_2057 ();
 sg13g2_decap_8 FILLER_9_2064 ();
 sg13g2_decap_8 FILLER_9_2071 ();
 sg13g2_decap_8 FILLER_9_2078 ();
 sg13g2_fill_2 FILLER_9_2085 ();
 sg13g2_fill_2 FILLER_9_2122 ();
 sg13g2_fill_1 FILLER_9_2124 ();
 sg13g2_fill_2 FILLER_9_2135 ();
 sg13g2_fill_2 FILLER_9_2141 ();
 sg13g2_fill_1 FILLER_9_2151 ();
 sg13g2_decap_8 FILLER_9_2161 ();
 sg13g2_decap_8 FILLER_9_2173 ();
 sg13g2_decap_8 FILLER_9_2180 ();
 sg13g2_fill_1 FILLER_9_2197 ();
 sg13g2_fill_1 FILLER_9_2205 ();
 sg13g2_decap_8 FILLER_9_2238 ();
 sg13g2_fill_2 FILLER_9_2245 ();
 sg13g2_fill_1 FILLER_9_2247 ();
 sg13g2_decap_4 FILLER_9_2293 ();
 sg13g2_decap_8 FILLER_9_2346 ();
 sg13g2_decap_8 FILLER_9_2353 ();
 sg13g2_decap_8 FILLER_9_2360 ();
 sg13g2_decap_8 FILLER_9_2424 ();
 sg13g2_decap_8 FILLER_9_2431 ();
 sg13g2_decap_8 FILLER_9_2438 ();
 sg13g2_decap_8 FILLER_9_2445 ();
 sg13g2_decap_8 FILLER_9_2452 ();
 sg13g2_decap_8 FILLER_9_2459 ();
 sg13g2_fill_2 FILLER_9_2466 ();
 sg13g2_decap_8 FILLER_9_2498 ();
 sg13g2_decap_8 FILLER_9_2505 ();
 sg13g2_decap_8 FILLER_9_2512 ();
 sg13g2_decap_4 FILLER_9_2519 ();
 sg13g2_fill_1 FILLER_9_2523 ();
 sg13g2_decap_8 FILLER_9_2555 ();
 sg13g2_decap_8 FILLER_9_2562 ();
 sg13g2_decap_8 FILLER_9_2569 ();
 sg13g2_decap_8 FILLER_9_2576 ();
 sg13g2_decap_8 FILLER_9_2583 ();
 sg13g2_fill_2 FILLER_9_2590 ();
 sg13g2_fill_1 FILLER_9_2592 ();
 sg13g2_decap_4 FILLER_9_2596 ();
 sg13g2_fill_2 FILLER_9_2621 ();
 sg13g2_fill_1 FILLER_9_2623 ();
 sg13g2_decap_8 FILLER_9_2633 ();
 sg13g2_fill_1 FILLER_9_2649 ();
 sg13g2_decap_4 FILLER_9_2681 ();
 sg13g2_fill_1 FILLER_9_2685 ();
 sg13g2_fill_1 FILLER_9_2749 ();
 sg13g2_fill_2 FILLER_9_2754 ();
 sg13g2_fill_1 FILLER_9_2756 ();
 sg13g2_fill_2 FILLER_9_2793 ();
 sg13g2_decap_8 FILLER_9_2804 ();
 sg13g2_decap_8 FILLER_9_2811 ();
 sg13g2_decap_8 FILLER_9_2818 ();
 sg13g2_fill_1 FILLER_9_2825 ();
 sg13g2_decap_8 FILLER_9_2854 ();
 sg13g2_decap_8 FILLER_9_2861 ();
 sg13g2_fill_2 FILLER_9_2868 ();
 sg13g2_fill_1 FILLER_9_2879 ();
 sg13g2_decap_8 FILLER_9_2884 ();
 sg13g2_decap_8 FILLER_9_2891 ();
 sg13g2_decap_8 FILLER_9_2898 ();
 sg13g2_decap_8 FILLER_9_2905 ();
 sg13g2_decap_8 FILLER_9_2912 ();
 sg13g2_fill_2 FILLER_9_2919 ();
 sg13g2_decap_8 FILLER_9_2951 ();
 sg13g2_decap_4 FILLER_9_2971 ();
 sg13g2_fill_1 FILLER_9_3013 ();
 sg13g2_decap_8 FILLER_9_3048 ();
 sg13g2_decap_8 FILLER_9_3055 ();
 sg13g2_decap_8 FILLER_9_3062 ();
 sg13g2_fill_1 FILLER_9_3079 ();
 sg13g2_decap_4 FILLER_9_3124 ();
 sg13g2_fill_1 FILLER_9_3162 ();
 sg13g2_decap_8 FILLER_9_3220 ();
 sg13g2_decap_4 FILLER_9_3227 ();
 sg13g2_decap_8 FILLER_9_3287 ();
 sg13g2_fill_1 FILLER_9_3294 ();
 sg13g2_fill_2 FILLER_9_3314 ();
 sg13g2_fill_1 FILLER_9_3316 ();
 sg13g2_decap_8 FILLER_9_3351 ();
 sg13g2_decap_8 FILLER_9_3358 ();
 sg13g2_decap_8 FILLER_9_3390 ();
 sg13g2_decap_8 FILLER_9_3397 ();
 sg13g2_fill_2 FILLER_9_3404 ();
 sg13g2_fill_1 FILLER_9_3406 ();
 sg13g2_decap_4 FILLER_9_3411 ();
 sg13g2_fill_2 FILLER_9_3469 ();
 sg13g2_fill_1 FILLER_9_3508 ();
 sg13g2_decap_8 FILLER_9_3536 ();
 sg13g2_decap_8 FILLER_9_3543 ();
 sg13g2_decap_8 FILLER_9_3550 ();
 sg13g2_decap_8 FILLER_9_3557 ();
 sg13g2_decap_8 FILLER_9_3564 ();
 sg13g2_decap_8 FILLER_9_3571 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_4 FILLER_10_49 ();
 sg13g2_fill_1 FILLER_10_62 ();
 sg13g2_fill_1 FILLER_10_77 ();
 sg13g2_fill_1 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_fill_1 FILLER_10_165 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_1 FILLER_10_274 ();
 sg13g2_decap_4 FILLER_10_279 ();
 sg13g2_fill_2 FILLER_10_283 ();
 sg13g2_fill_2 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_fill_2 FILLER_10_405 ();
 sg13g2_decap_4 FILLER_10_481 ();
 sg13g2_decap_4 FILLER_10_489 ();
 sg13g2_fill_1 FILLER_10_493 ();
 sg13g2_decap_8 FILLER_10_508 ();
 sg13g2_fill_2 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_555 ();
 sg13g2_decap_8 FILLER_10_562 ();
 sg13g2_decap_8 FILLER_10_577 ();
 sg13g2_fill_2 FILLER_10_584 ();
 sg13g2_fill_1 FILLER_10_586 ();
 sg13g2_fill_2 FILLER_10_615 ();
 sg13g2_fill_1 FILLER_10_677 ();
 sg13g2_fill_1 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_692 ();
 sg13g2_fill_1 FILLER_10_699 ();
 sg13g2_fill_2 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_729 ();
 sg13g2_decap_8 FILLER_10_736 ();
 sg13g2_decap_4 FILLER_10_743 ();
 sg13g2_fill_1 FILLER_10_747 ();
 sg13g2_decap_8 FILLER_10_758 ();
 sg13g2_decap_8 FILLER_10_810 ();
 sg13g2_fill_2 FILLER_10_817 ();
 sg13g2_fill_1 FILLER_10_819 ();
 sg13g2_fill_1 FILLER_10_825 ();
 sg13g2_fill_2 FILLER_10_843 ();
 sg13g2_fill_1 FILLER_10_845 ();
 sg13g2_decap_8 FILLER_10_878 ();
 sg13g2_decap_8 FILLER_10_885 ();
 sg13g2_decap_8 FILLER_10_892 ();
 sg13g2_decap_8 FILLER_10_899 ();
 sg13g2_fill_2 FILLER_10_906 ();
 sg13g2_fill_1 FILLER_10_908 ();
 sg13g2_fill_2 FILLER_10_937 ();
 sg13g2_decap_8 FILLER_10_944 ();
 sg13g2_decap_8 FILLER_10_951 ();
 sg13g2_decap_4 FILLER_10_958 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_decap_8 FILLER_10_1026 ();
 sg13g2_decap_8 FILLER_10_1033 ();
 sg13g2_fill_1 FILLER_10_1040 ();
 sg13g2_fill_1 FILLER_10_1144 ();
 sg13g2_decap_8 FILLER_10_1192 ();
 sg13g2_decap_8 FILLER_10_1199 ();
 sg13g2_decap_8 FILLER_10_1206 ();
 sg13g2_fill_1 FILLER_10_1213 ();
 sg13g2_decap_8 FILLER_10_1265 ();
 sg13g2_decap_8 FILLER_10_1272 ();
 sg13g2_fill_1 FILLER_10_1279 ();
 sg13g2_decap_8 FILLER_10_1334 ();
 sg13g2_decap_8 FILLER_10_1341 ();
 sg13g2_decap_8 FILLER_10_1348 ();
 sg13g2_fill_1 FILLER_10_1355 ();
 sg13g2_decap_4 FILLER_10_1383 ();
 sg13g2_fill_1 FILLER_10_1387 ();
 sg13g2_decap_8 FILLER_10_1410 ();
 sg13g2_decap_8 FILLER_10_1417 ();
 sg13g2_decap_8 FILLER_10_1424 ();
 sg13g2_decap_8 FILLER_10_1431 ();
 sg13g2_decap_8 FILLER_10_1438 ();
 sg13g2_decap_4 FILLER_10_1445 ();
 sg13g2_fill_2 FILLER_10_1458 ();
 sg13g2_fill_1 FILLER_10_1460 ();
 sg13g2_fill_1 FILLER_10_1488 ();
 sg13g2_fill_1 FILLER_10_1501 ();
 sg13g2_fill_2 FILLER_10_1510 ();
 sg13g2_fill_1 FILLER_10_1512 ();
 sg13g2_decap_8 FILLER_10_1522 ();
 sg13g2_decap_4 FILLER_10_1529 ();
 sg13g2_fill_2 FILLER_10_1533 ();
 sg13g2_fill_2 FILLER_10_1540 ();
 sg13g2_fill_1 FILLER_10_1542 ();
 sg13g2_decap_4 FILLER_10_1549 ();
 sg13g2_fill_2 FILLER_10_1558 ();
 sg13g2_fill_2 FILLER_10_1582 ();
 sg13g2_fill_2 FILLER_10_1593 ();
 sg13g2_fill_1 FILLER_10_1595 ();
 sg13g2_decap_8 FILLER_10_1665 ();
 sg13g2_fill_1 FILLER_10_1672 ();
 sg13g2_fill_2 FILLER_10_1691 ();
 sg13g2_decap_8 FILLER_10_1719 ();
 sg13g2_decap_8 FILLER_10_1726 ();
 sg13g2_decap_8 FILLER_10_1733 ();
 sg13g2_decap_8 FILLER_10_1740 ();
 sg13g2_decap_8 FILLER_10_1747 ();
 sg13g2_decap_8 FILLER_10_1754 ();
 sg13g2_decap_8 FILLER_10_1766 ();
 sg13g2_decap_8 FILLER_10_1773 ();
 sg13g2_decap_8 FILLER_10_1780 ();
 sg13g2_fill_2 FILLER_10_1787 ();
 sg13g2_fill_2 FILLER_10_1854 ();
 sg13g2_fill_1 FILLER_10_1880 ();
 sg13g2_fill_1 FILLER_10_1890 ();
 sg13g2_fill_2 FILLER_10_1913 ();
 sg13g2_decap_8 FILLER_10_1923 ();
 sg13g2_decap_8 FILLER_10_1930 ();
 sg13g2_decap_8 FILLER_10_1937 ();
 sg13g2_decap_4 FILLER_10_1944 ();
 sg13g2_fill_2 FILLER_10_1948 ();
 sg13g2_decap_8 FILLER_10_1963 ();
 sg13g2_decap_8 FILLER_10_1970 ();
 sg13g2_decap_8 FILLER_10_2012 ();
 sg13g2_fill_2 FILLER_10_2019 ();
 sg13g2_decap_8 FILLER_10_2060 ();
 sg13g2_decap_4 FILLER_10_2067 ();
 sg13g2_fill_2 FILLER_10_2071 ();
 sg13g2_decap_8 FILLER_10_2100 ();
 sg13g2_fill_2 FILLER_10_2107 ();
 sg13g2_fill_1 FILLER_10_2109 ();
 sg13g2_fill_2 FILLER_10_2115 ();
 sg13g2_decap_8 FILLER_10_2126 ();
 sg13g2_decap_8 FILLER_10_2133 ();
 sg13g2_decap_8 FILLER_10_2140 ();
 sg13g2_decap_8 FILLER_10_2152 ();
 sg13g2_decap_8 FILLER_10_2159 ();
 sg13g2_decap_8 FILLER_10_2166 ();
 sg13g2_decap_8 FILLER_10_2173 ();
 sg13g2_fill_2 FILLER_10_2180 ();
 sg13g2_decap_8 FILLER_10_2192 ();
 sg13g2_fill_2 FILLER_10_2199 ();
 sg13g2_fill_2 FILLER_10_2237 ();
 sg13g2_fill_2 FILLER_10_2245 ();
 sg13g2_fill_1 FILLER_10_2247 ();
 sg13g2_fill_2 FILLER_10_2276 ();
 sg13g2_fill_1 FILLER_10_2278 ();
 sg13g2_decap_4 FILLER_10_2288 ();
 sg13g2_decap_8 FILLER_10_2355 ();
 sg13g2_decap_8 FILLER_10_2362 ();
 sg13g2_fill_1 FILLER_10_2369 ();
 sg13g2_decap_8 FILLER_10_2411 ();
 sg13g2_decap_8 FILLER_10_2418 ();
 sg13g2_decap_8 FILLER_10_2425 ();
 sg13g2_decap_8 FILLER_10_2432 ();
 sg13g2_decap_8 FILLER_10_2439 ();
 sg13g2_decap_8 FILLER_10_2446 ();
 sg13g2_decap_8 FILLER_10_2453 ();
 sg13g2_decap_8 FILLER_10_2460 ();
 sg13g2_decap_4 FILLER_10_2467 ();
 sg13g2_fill_2 FILLER_10_2471 ();
 sg13g2_fill_2 FILLER_10_2477 ();
 sg13g2_fill_1 FILLER_10_2479 ();
 sg13g2_decap_8 FILLER_10_2484 ();
 sg13g2_decap_8 FILLER_10_2491 ();
 sg13g2_decap_8 FILLER_10_2498 ();
 sg13g2_decap_8 FILLER_10_2505 ();
 sg13g2_decap_8 FILLER_10_2512 ();
 sg13g2_decap_8 FILLER_10_2519 ();
 sg13g2_fill_2 FILLER_10_2526 ();
 sg13g2_fill_1 FILLER_10_2528 ();
 sg13g2_decap_8 FILLER_10_2569 ();
 sg13g2_fill_2 FILLER_10_2576 ();
 sg13g2_decap_8 FILLER_10_2583 ();
 sg13g2_decap_8 FILLER_10_2590 ();
 sg13g2_decap_4 FILLER_10_2597 ();
 sg13g2_fill_2 FILLER_10_2601 ();
 sg13g2_decap_4 FILLER_10_2613 ();
 sg13g2_fill_2 FILLER_10_2617 ();
 sg13g2_fill_1 FILLER_10_2629 ();
 sg13g2_decap_8 FILLER_10_2684 ();
 sg13g2_fill_2 FILLER_10_2695 ();
 sg13g2_decap_8 FILLER_10_2743 ();
 sg13g2_decap_8 FILLER_10_2750 ();
 sg13g2_decap_8 FILLER_10_2757 ();
 sg13g2_decap_8 FILLER_10_2764 ();
 sg13g2_fill_1 FILLER_10_2775 ();
 sg13g2_fill_1 FILLER_10_2786 ();
 sg13g2_decap_8 FILLER_10_2791 ();
 sg13g2_decap_8 FILLER_10_2798 ();
 sg13g2_decap_8 FILLER_10_2805 ();
 sg13g2_decap_8 FILLER_10_2812 ();
 sg13g2_decap_8 FILLER_10_2819 ();
 sg13g2_decap_8 FILLER_10_2826 ();
 sg13g2_decap_8 FILLER_10_2833 ();
 sg13g2_decap_8 FILLER_10_2840 ();
 sg13g2_decap_8 FILLER_10_2847 ();
 sg13g2_fill_1 FILLER_10_2854 ();
 sg13g2_decap_8 FILLER_10_2909 ();
 sg13g2_decap_4 FILLER_10_2916 ();
 sg13g2_decap_8 FILLER_10_2966 ();
 sg13g2_decap_8 FILLER_10_2973 ();
 sg13g2_decap_8 FILLER_10_2984 ();
 sg13g2_fill_2 FILLER_10_3001 ();
 sg13g2_decap_8 FILLER_10_3013 ();
 sg13g2_decap_4 FILLER_10_3020 ();
 sg13g2_fill_2 FILLER_10_3024 ();
 sg13g2_decap_8 FILLER_10_3047 ();
 sg13g2_decap_8 FILLER_10_3054 ();
 sg13g2_decap_8 FILLER_10_3061 ();
 sg13g2_decap_8 FILLER_10_3068 ();
 sg13g2_fill_1 FILLER_10_3075 ();
 sg13g2_fill_2 FILLER_10_3080 ();
 sg13g2_fill_1 FILLER_10_3082 ();
 sg13g2_decap_8 FILLER_10_3093 ();
 sg13g2_fill_1 FILLER_10_3100 ();
 sg13g2_decap_8 FILLER_10_3120 ();
 sg13g2_decap_4 FILLER_10_3127 ();
 sg13g2_fill_2 FILLER_10_3131 ();
 sg13g2_decap_4 FILLER_10_3164 ();
 sg13g2_fill_1 FILLER_10_3168 ();
 sg13g2_decap_8 FILLER_10_3213 ();
 sg13g2_decap_8 FILLER_10_3220 ();
 sg13g2_decap_4 FILLER_10_3227 ();
 sg13g2_fill_2 FILLER_10_3253 ();
 sg13g2_decap_8 FILLER_10_3285 ();
 sg13g2_decap_8 FILLER_10_3292 ();
 sg13g2_decap_8 FILLER_10_3299 ();
 sg13g2_fill_2 FILLER_10_3306 ();
 sg13g2_fill_1 FILLER_10_3321 ();
 sg13g2_decap_8 FILLER_10_3332 ();
 sg13g2_decap_8 FILLER_10_3339 ();
 sg13g2_decap_8 FILLER_10_3346 ();
 sg13g2_fill_2 FILLER_10_3399 ();
 sg13g2_fill_1 FILLER_10_3401 ();
 sg13g2_decap_8 FILLER_10_3449 ();
 sg13g2_decap_4 FILLER_10_3465 ();
 sg13g2_fill_2 FILLER_10_3469 ();
 sg13g2_decap_4 FILLER_10_3491 ();
 sg13g2_decap_8 FILLER_10_3524 ();
 sg13g2_decap_8 FILLER_10_3531 ();
 sg13g2_decap_8 FILLER_10_3538 ();
 sg13g2_decap_8 FILLER_10_3545 ();
 sg13g2_decap_8 FILLER_10_3552 ();
 sg13g2_decap_8 FILLER_10_3559 ();
 sg13g2_decap_8 FILLER_10_3566 ();
 sg13g2_decap_4 FILLER_10_3573 ();
 sg13g2_fill_1 FILLER_10_3577 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_43 ();
 sg13g2_fill_1 FILLER_11_45 ();
 sg13g2_decap_8 FILLER_11_55 ();
 sg13g2_fill_1 FILLER_11_62 ();
 sg13g2_decap_4 FILLER_11_156 ();
 sg13g2_fill_2 FILLER_11_160 ();
 sg13g2_fill_1 FILLER_11_198 ();
 sg13g2_decap_4 FILLER_11_235 ();
 sg13g2_fill_2 FILLER_11_239 ();
 sg13g2_decap_8 FILLER_11_254 ();
 sg13g2_fill_1 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_4 FILLER_11_280 ();
 sg13g2_fill_1 FILLER_11_335 ();
 sg13g2_fill_2 FILLER_11_349 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_4 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_431 ();
 sg13g2_fill_1 FILLER_11_433 ();
 sg13g2_fill_1 FILLER_11_474 ();
 sg13g2_fill_1 FILLER_11_491 ();
 sg13g2_fill_2 FILLER_11_496 ();
 sg13g2_fill_1 FILLER_11_498 ();
 sg13g2_decap_8 FILLER_11_503 ();
 sg13g2_fill_2 FILLER_11_510 ();
 sg13g2_fill_1 FILLER_11_512 ();
 sg13g2_decap_8 FILLER_11_554 ();
 sg13g2_decap_8 FILLER_11_561 ();
 sg13g2_decap_8 FILLER_11_568 ();
 sg13g2_fill_1 FILLER_11_575 ();
 sg13g2_decap_4 FILLER_11_622 ();
 sg13g2_fill_2 FILLER_11_626 ();
 sg13g2_decap_4 FILLER_11_637 ();
 sg13g2_fill_2 FILLER_11_641 ();
 sg13g2_fill_2 FILLER_11_667 ();
 sg13g2_decap_8 FILLER_11_710 ();
 sg13g2_decap_4 FILLER_11_717 ();
 sg13g2_fill_1 FILLER_11_721 ();
 sg13g2_fill_2 FILLER_11_727 ();
 sg13g2_fill_2 FILLER_11_765 ();
 sg13g2_fill_2 FILLER_11_772 ();
 sg13g2_fill_2 FILLER_11_805 ();
 sg13g2_fill_1 FILLER_11_807 ();
 sg13g2_decap_8 FILLER_11_813 ();
 sg13g2_decap_8 FILLER_11_820 ();
 sg13g2_decap_4 FILLER_11_827 ();
 sg13g2_fill_1 FILLER_11_831 ();
 sg13g2_decap_4 FILLER_11_841 ();
 sg13g2_fill_2 FILLER_11_845 ();
 sg13g2_decap_8 FILLER_11_876 ();
 sg13g2_decap_8 FILLER_11_883 ();
 sg13g2_decap_8 FILLER_11_890 ();
 sg13g2_decap_8 FILLER_11_897 ();
 sg13g2_decap_4 FILLER_11_904 ();
 sg13g2_fill_1 FILLER_11_908 ();
 sg13g2_fill_1 FILLER_11_922 ();
 sg13g2_fill_2 FILLER_11_928 ();
 sg13g2_fill_1 FILLER_11_930 ();
 sg13g2_fill_1 FILLER_11_959 ();
 sg13g2_fill_2 FILLER_11_986 ();
 sg13g2_decap_8 FILLER_11_1002 ();
 sg13g2_decap_8 FILLER_11_1009 ();
 sg13g2_decap_8 FILLER_11_1016 ();
 sg13g2_decap_8 FILLER_11_1023 ();
 sg13g2_fill_2 FILLER_11_1030 ();
 sg13g2_fill_1 FILLER_11_1032 ();
 sg13g2_decap_4 FILLER_11_1051 ();
 sg13g2_fill_1 FILLER_11_1055 ();
 sg13g2_decap_8 FILLER_11_1074 ();
 sg13g2_fill_2 FILLER_11_1081 ();
 sg13g2_fill_1 FILLER_11_1108 ();
 sg13g2_fill_1 FILLER_11_1117 ();
 sg13g2_decap_4 FILLER_11_1132 ();
 sg13g2_fill_1 FILLER_11_1141 ();
 sg13g2_fill_2 FILLER_11_1147 ();
 sg13g2_fill_1 FILLER_11_1149 ();
 sg13g2_fill_1 FILLER_11_1173 ();
 sg13g2_decap_8 FILLER_11_1195 ();
 sg13g2_fill_2 FILLER_11_1202 ();
 sg13g2_fill_1 FILLER_11_1204 ();
 sg13g2_fill_1 FILLER_11_1226 ();
 sg13g2_fill_2 FILLER_11_1268 ();
 sg13g2_fill_1 FILLER_11_1270 ();
 sg13g2_decap_4 FILLER_11_1276 ();
 sg13g2_decap_8 FILLER_11_1303 ();
 sg13g2_fill_1 FILLER_11_1310 ();
 sg13g2_decap_4 FILLER_11_1338 ();
 sg13g2_fill_2 FILLER_11_1342 ();
 sg13g2_decap_8 FILLER_11_1381 ();
 sg13g2_fill_2 FILLER_11_1388 ();
 sg13g2_fill_1 FILLER_11_1390 ();
 sg13g2_decap_8 FILLER_11_1400 ();
 sg13g2_fill_2 FILLER_11_1407 ();
 sg13g2_decap_4 FILLER_11_1444 ();
 sg13g2_fill_2 FILLER_11_1448 ();
 sg13g2_fill_1 FILLER_11_1489 ();
 sg13g2_decap_8 FILLER_11_1517 ();
 sg13g2_decap_4 FILLER_11_1524 ();
 sg13g2_fill_2 FILLER_11_1556 ();
 sg13g2_fill_1 FILLER_11_1558 ();
 sg13g2_decap_4 FILLER_11_1597 ();
 sg13g2_fill_2 FILLER_11_1601 ();
 sg13g2_fill_2 FILLER_11_1607 ();
 sg13g2_fill_1 FILLER_11_1631 ();
 sg13g2_fill_2 FILLER_11_1689 ();
 sg13g2_decap_8 FILLER_11_1704 ();
 sg13g2_decap_8 FILLER_11_1711 ();
 sg13g2_fill_2 FILLER_11_1718 ();
 sg13g2_fill_2 FILLER_11_1726 ();
 sg13g2_fill_1 FILLER_11_1728 ();
 sg13g2_decap_8 FILLER_11_1765 ();
 sg13g2_decap_8 FILLER_11_1772 ();
 sg13g2_decap_8 FILLER_11_1779 ();
 sg13g2_decap_4 FILLER_11_1786 ();
 sg13g2_fill_1 FILLER_11_1790 ();
 sg13g2_fill_1 FILLER_11_1803 ();
 sg13g2_decap_8 FILLER_11_1817 ();
 sg13g2_decap_8 FILLER_11_1824 ();
 sg13g2_decap_8 FILLER_11_1831 ();
 sg13g2_fill_2 FILLER_11_1838 ();
 sg13g2_decap_8 FILLER_11_1877 ();
 sg13g2_fill_2 FILLER_11_1884 ();
 sg13g2_fill_1 FILLER_11_1886 ();
 sg13g2_fill_2 FILLER_11_1924 ();
 sg13g2_decap_8 FILLER_11_1939 ();
 sg13g2_decap_4 FILLER_11_1946 ();
 sg13g2_fill_1 FILLER_11_1950 ();
 sg13g2_decap_8 FILLER_11_1964 ();
 sg13g2_decap_8 FILLER_11_1971 ();
 sg13g2_fill_2 FILLER_11_1978 ();
 sg13g2_decap_8 FILLER_11_2020 ();
 sg13g2_fill_1 FILLER_11_2027 ();
 sg13g2_fill_2 FILLER_11_2046 ();
 sg13g2_fill_1 FILLER_11_2048 ();
 sg13g2_decap_4 FILLER_11_2062 ();
 sg13g2_fill_1 FILLER_11_2066 ();
 sg13g2_decap_8 FILLER_11_2071 ();
 sg13g2_decap_4 FILLER_11_2095 ();
 sg13g2_fill_1 FILLER_11_2099 ();
 sg13g2_fill_2 FILLER_11_2135 ();
 sg13g2_fill_1 FILLER_11_2137 ();
 sg13g2_decap_4 FILLER_11_2156 ();
 sg13g2_fill_2 FILLER_11_2160 ();
 sg13g2_fill_1 FILLER_11_2171 ();
 sg13g2_decap_8 FILLER_11_2177 ();
 sg13g2_fill_2 FILLER_11_2184 ();
 sg13g2_decap_4 FILLER_11_2207 ();
 sg13g2_decap_4 FILLER_11_2242 ();
 sg13g2_fill_2 FILLER_11_2246 ();
 sg13g2_fill_2 FILLER_11_2263 ();
 sg13g2_fill_1 FILLER_11_2279 ();
 sg13g2_fill_1 FILLER_11_2296 ();
 sg13g2_fill_2 FILLER_11_2311 ();
 sg13g2_fill_1 FILLER_11_2327 ();
 sg13g2_decap_8 FILLER_11_2346 ();
 sg13g2_decap_8 FILLER_11_2353 ();
 sg13g2_decap_8 FILLER_11_2360 ();
 sg13g2_fill_2 FILLER_11_2367 ();
 sg13g2_fill_1 FILLER_11_2369 ();
 sg13g2_decap_8 FILLER_11_2411 ();
 sg13g2_decap_8 FILLER_11_2501 ();
 sg13g2_decap_8 FILLER_11_2508 ();
 sg13g2_decap_8 FILLER_11_2515 ();
 sg13g2_fill_2 FILLER_11_2532 ();
 sg13g2_fill_1 FILLER_11_2534 ();
 sg13g2_fill_1 FILLER_11_2545 ();
 sg13g2_fill_2 FILLER_11_2573 ();
 sg13g2_fill_1 FILLER_11_2575 ();
 sg13g2_fill_2 FILLER_11_2586 ();
 sg13g2_fill_1 FILLER_11_2588 ();
 sg13g2_decap_8 FILLER_11_2643 ();
 sg13g2_decap_4 FILLER_11_2650 ();
 sg13g2_fill_1 FILLER_11_2654 ();
 sg13g2_decap_4 FILLER_11_2669 ();
 sg13g2_fill_1 FILLER_11_2673 ();
 sg13g2_decap_8 FILLER_11_2683 ();
 sg13g2_decap_8 FILLER_11_2690 ();
 sg13g2_decap_4 FILLER_11_2697 ();
 sg13g2_fill_1 FILLER_11_2701 ();
 sg13g2_fill_2 FILLER_11_2706 ();
 sg13g2_decap_8 FILLER_11_2733 ();
 sg13g2_decap_8 FILLER_11_2740 ();
 sg13g2_decap_8 FILLER_11_2747 ();
 sg13g2_decap_4 FILLER_11_2754 ();
 sg13g2_fill_2 FILLER_11_2758 ();
 sg13g2_fill_2 FILLER_11_2787 ();
 sg13g2_fill_1 FILLER_11_2789 ();
 sg13g2_decap_8 FILLER_11_2799 ();
 sg13g2_decap_4 FILLER_11_2806 ();
 sg13g2_fill_2 FILLER_11_2837 ();
 sg13g2_fill_1 FILLER_11_2839 ();
 sg13g2_fill_2 FILLER_11_2867 ();
 sg13g2_decap_8 FILLER_11_2896 ();
 sg13g2_decap_8 FILLER_11_2903 ();
 sg13g2_decap_8 FILLER_11_2910 ();
 sg13g2_fill_1 FILLER_11_2917 ();
 sg13g2_decap_8 FILLER_11_2972 ();
 sg13g2_fill_2 FILLER_11_2979 ();
 sg13g2_decap_8 FILLER_11_3030 ();
 sg13g2_decap_8 FILLER_11_3037 ();
 sg13g2_decap_8 FILLER_11_3044 ();
 sg13g2_decap_8 FILLER_11_3051 ();
 sg13g2_fill_2 FILLER_11_3058 ();
 sg13g2_fill_1 FILLER_11_3060 ();
 sg13g2_decap_4 FILLER_11_3088 ();
 sg13g2_fill_2 FILLER_11_3092 ();
 sg13g2_decap_4 FILLER_11_3131 ();
 sg13g2_fill_2 FILLER_11_3145 ();
 sg13g2_fill_2 FILLER_11_3169 ();
 sg13g2_fill_1 FILLER_11_3171 ();
 sg13g2_fill_2 FILLER_11_3202 ();
 sg13g2_decap_8 FILLER_11_3208 ();
 sg13g2_decap_8 FILLER_11_3215 ();
 sg13g2_decap_8 FILLER_11_3222 ();
 sg13g2_decap_8 FILLER_11_3229 ();
 sg13g2_decap_4 FILLER_11_3236 ();
 sg13g2_fill_2 FILLER_11_3240 ();
 sg13g2_fill_2 FILLER_11_3255 ();
 sg13g2_fill_1 FILLER_11_3257 ();
 sg13g2_fill_1 FILLER_11_3262 ();
 sg13g2_decap_8 FILLER_11_3282 ();
 sg13g2_decap_8 FILLER_11_3289 ();
 sg13g2_decap_8 FILLER_11_3296 ();
 sg13g2_decap_8 FILLER_11_3303 ();
 sg13g2_decap_8 FILLER_11_3310 ();
 sg13g2_fill_1 FILLER_11_3317 ();
 sg13g2_decap_8 FILLER_11_3345 ();
 sg13g2_decap_4 FILLER_11_3352 ();
 sg13g2_fill_1 FILLER_11_3356 ();
 sg13g2_decap_8 FILLER_11_3394 ();
 sg13g2_decap_8 FILLER_11_3401 ();
 sg13g2_decap_4 FILLER_11_3408 ();
 sg13g2_fill_1 FILLER_11_3412 ();
 sg13g2_decap_8 FILLER_11_3445 ();
 sg13g2_decap_8 FILLER_11_3452 ();
 sg13g2_decap_8 FILLER_11_3459 ();
 sg13g2_fill_1 FILLER_11_3466 ();
 sg13g2_fill_1 FILLER_11_3476 ();
 sg13g2_fill_2 FILLER_11_3487 ();
 sg13g2_fill_1 FILLER_11_3489 ();
 sg13g2_fill_1 FILLER_11_3499 ();
 sg13g2_decap_8 FILLER_11_3513 ();
 sg13g2_fill_1 FILLER_11_3520 ();
 sg13g2_decap_8 FILLER_11_3530 ();
 sg13g2_fill_1 FILLER_11_3537 ();
 sg13g2_decap_8 FILLER_11_3547 ();
 sg13g2_decap_8 FILLER_11_3554 ();
 sg13g2_decap_8 FILLER_11_3561 ();
 sg13g2_decap_8 FILLER_11_3568 ();
 sg13g2_fill_2 FILLER_11_3575 ();
 sg13g2_fill_1 FILLER_11_3577 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_59 ();
 sg13g2_decap_8 FILLER_12_66 ();
 sg13g2_decap_4 FILLER_12_73 ();
 sg13g2_fill_2 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_106 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_4 FILLER_12_158 ();
 sg13g2_fill_2 FILLER_12_162 ();
 sg13g2_decap_8 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_195 ();
 sg13g2_fill_2 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_decap_8 FILLER_12_230 ();
 sg13g2_decap_8 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_244 ();
 sg13g2_decap_8 FILLER_12_261 ();
 sg13g2_fill_2 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_decap_4 FILLER_12_276 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_fill_2 FILLER_12_389 ();
 sg13g2_decap_4 FILLER_12_424 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_fill_2 FILLER_12_443 ();
 sg13g2_fill_2 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_fill_1 FILLER_12_574 ();
 sg13g2_fill_1 FILLER_12_593 ();
 sg13g2_fill_1 FILLER_12_599 ();
 sg13g2_fill_2 FILLER_12_605 ();
 sg13g2_fill_1 FILLER_12_607 ();
 sg13g2_decap_8 FILLER_12_618 ();
 sg13g2_decap_8 FILLER_12_625 ();
 sg13g2_decap_4 FILLER_12_632 ();
 sg13g2_fill_2 FILLER_12_647 ();
 sg13g2_fill_1 FILLER_12_649 ();
 sg13g2_fill_2 FILLER_12_656 ();
 sg13g2_fill_1 FILLER_12_658 ();
 sg13g2_fill_1 FILLER_12_687 ();
 sg13g2_decap_4 FILLER_12_692 ();
 sg13g2_fill_2 FILLER_12_696 ();
 sg13g2_fill_2 FILLER_12_743 ();
 sg13g2_fill_1 FILLER_12_745 ();
 sg13g2_decap_4 FILLER_12_762 ();
 sg13g2_decap_4 FILLER_12_771 ();
 sg13g2_fill_2 FILLER_12_775 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_decap_8 FILLER_12_821 ();
 sg13g2_decap_8 FILLER_12_828 ();
 sg13g2_decap_8 FILLER_12_835 ();
 sg13g2_fill_1 FILLER_12_842 ();
 sg13g2_decap_8 FILLER_12_885 ();
 sg13g2_decap_8 FILLER_12_892 ();
 sg13g2_decap_4 FILLER_12_899 ();
 sg13g2_fill_2 FILLER_12_903 ();
 sg13g2_fill_1 FILLER_12_933 ();
 sg13g2_decap_4 FILLER_12_962 ();
 sg13g2_decap_4 FILLER_12_970 ();
 sg13g2_fill_2 FILLER_12_993 ();
 sg13g2_fill_1 FILLER_12_995 ();
 sg13g2_fill_1 FILLER_12_1009 ();
 sg13g2_fill_2 FILLER_12_1015 ();
 sg13g2_fill_1 FILLER_12_1017 ();
 sg13g2_fill_2 FILLER_12_1031 ();
 sg13g2_fill_1 FILLER_12_1033 ();
 sg13g2_decap_8 FILLER_12_1079 ();
 sg13g2_fill_2 FILLER_12_1152 ();
 sg13g2_fill_1 FILLER_12_1154 ();
 sg13g2_decap_8 FILLER_12_1192 ();
 sg13g2_decap_8 FILLER_12_1199 ();
 sg13g2_decap_8 FILLER_12_1206 ();
 sg13g2_fill_1 FILLER_12_1213 ();
 sg13g2_fill_1 FILLER_12_1257 ();
 sg13g2_decap_4 FILLER_12_1263 ();
 sg13g2_fill_1 FILLER_12_1267 ();
 sg13g2_fill_2 FILLER_12_1308 ();
 sg13g2_fill_2 FILLER_12_1326 ();
 sg13g2_fill_1 FILLER_12_1328 ();
 sg13g2_decap_4 FILLER_12_1357 ();
 sg13g2_decap_8 FILLER_12_1370 ();
 sg13g2_decap_8 FILLER_12_1377 ();
 sg13g2_fill_2 FILLER_12_1384 ();
 sg13g2_decap_4 FILLER_12_1436 ();
 sg13g2_decap_8 FILLER_12_1450 ();
 sg13g2_decap_4 FILLER_12_1457 ();
 sg13g2_fill_1 FILLER_12_1466 ();
 sg13g2_decap_4 FILLER_12_1509 ();
 sg13g2_decap_8 FILLER_12_1516 ();
 sg13g2_decap_8 FILLER_12_1523 ();
 sg13g2_fill_2 FILLER_12_1530 ();
 sg13g2_fill_1 FILLER_12_1544 ();
 sg13g2_decap_8 FILLER_12_1560 ();
 sg13g2_decap_8 FILLER_12_1567 ();
 sg13g2_fill_1 FILLER_12_1574 ();
 sg13g2_decap_4 FILLER_12_1579 ();
 sg13g2_fill_1 FILLER_12_1583 ();
 sg13g2_fill_2 FILLER_12_1596 ();
 sg13g2_decap_8 FILLER_12_1603 ();
 sg13g2_decap_4 FILLER_12_1610 ();
 sg13g2_fill_1 FILLER_12_1614 ();
 sg13g2_fill_1 FILLER_12_1627 ();
 sg13g2_fill_2 FILLER_12_1639 ();
 sg13g2_fill_1 FILLER_12_1641 ();
 sg13g2_fill_1 FILLER_12_1708 ();
 sg13g2_fill_1 FILLER_12_1736 ();
 sg13g2_decap_4 FILLER_12_1775 ();
 sg13g2_fill_1 FILLER_12_1779 ();
 sg13g2_decap_8 FILLER_12_1820 ();
 sg13g2_decap_4 FILLER_12_1827 ();
 sg13g2_fill_2 FILLER_12_1831 ();
 sg13g2_decap_8 FILLER_12_1870 ();
 sg13g2_fill_2 FILLER_12_1877 ();
 sg13g2_fill_1 FILLER_12_1879 ();
 sg13g2_decap_4 FILLER_12_1977 ();
 sg13g2_fill_2 FILLER_12_2015 ();
 sg13g2_fill_1 FILLER_12_2017 ();
 sg13g2_fill_1 FILLER_12_2031 ();
 sg13g2_decap_4 FILLER_12_2045 ();
 sg13g2_fill_2 FILLER_12_2049 ();
 sg13g2_fill_2 FILLER_12_2112 ();
 sg13g2_fill_2 FILLER_12_2180 ();
 sg13g2_fill_1 FILLER_12_2182 ();
 sg13g2_fill_2 FILLER_12_2229 ();
 sg13g2_fill_1 FILLER_12_2231 ();
 sg13g2_decap_8 FILLER_12_2241 ();
 sg13g2_decap_4 FILLER_12_2248 ();
 sg13g2_decap_8 FILLER_12_2293 ();
 sg13g2_decap_8 FILLER_12_2300 ();
 sg13g2_fill_2 FILLER_12_2307 ();
 sg13g2_decap_8 FILLER_12_2343 ();
 sg13g2_decap_8 FILLER_12_2350 ();
 sg13g2_decap_8 FILLER_12_2357 ();
 sg13g2_decap_8 FILLER_12_2364 ();
 sg13g2_decap_4 FILLER_12_2371 ();
 sg13g2_fill_2 FILLER_12_2375 ();
 sg13g2_decap_4 FILLER_12_2381 ();
 sg13g2_decap_4 FILLER_12_2412 ();
 sg13g2_fill_1 FILLER_12_2416 ();
 sg13g2_decap_8 FILLER_12_2494 ();
 sg13g2_decap_8 FILLER_12_2501 ();
 sg13g2_fill_1 FILLER_12_2508 ();
 sg13g2_decap_4 FILLER_12_2568 ();
 sg13g2_fill_1 FILLER_12_2572 ();
 sg13g2_fill_1 FILLER_12_2604 ();
 sg13g2_decap_4 FILLER_12_2630 ();
 sg13g2_fill_1 FILLER_12_2634 ();
 sg13g2_decap_8 FILLER_12_2639 ();
 sg13g2_decap_8 FILLER_12_2646 ();
 sg13g2_fill_1 FILLER_12_2653 ();
 sg13g2_decap_8 FILLER_12_2675 ();
 sg13g2_decap_8 FILLER_12_2682 ();
 sg13g2_decap_8 FILLER_12_2689 ();
 sg13g2_decap_8 FILLER_12_2696 ();
 sg13g2_decap_8 FILLER_12_2703 ();
 sg13g2_decap_8 FILLER_12_2710 ();
 sg13g2_decap_4 FILLER_12_2717 ();
 sg13g2_fill_1 FILLER_12_2721 ();
 sg13g2_decap_8 FILLER_12_2726 ();
 sg13g2_decap_8 FILLER_12_2733 ();
 sg13g2_decap_8 FILLER_12_2740 ();
 sg13g2_decap_8 FILLER_12_2747 ();
 sg13g2_fill_2 FILLER_12_2754 ();
 sg13g2_fill_1 FILLER_12_2814 ();
 sg13g2_decap_8 FILLER_12_2819 ();
 sg13g2_decap_8 FILLER_12_2826 ();
 sg13g2_decap_8 FILLER_12_2833 ();
 sg13g2_fill_2 FILLER_12_2840 ();
 sg13g2_decap_4 FILLER_12_2904 ();
 sg13g2_fill_2 FILLER_12_2908 ();
 sg13g2_decap_8 FILLER_12_2969 ();
 sg13g2_fill_1 FILLER_12_2976 ();
 sg13g2_decap_4 FILLER_12_3004 ();
 sg13g2_fill_1 FILLER_12_3008 ();
 sg13g2_decap_8 FILLER_12_3036 ();
 sg13g2_decap_8 FILLER_12_3043 ();
 sg13g2_fill_2 FILLER_12_3050 ();
 sg13g2_decap_8 FILLER_12_3137 ();
 sg13g2_decap_8 FILLER_12_3144 ();
 sg13g2_decap_8 FILLER_12_3151 ();
 sg13g2_fill_1 FILLER_12_3158 ();
 sg13g2_decap_8 FILLER_12_3188 ();
 sg13g2_decap_8 FILLER_12_3195 ();
 sg13g2_decap_8 FILLER_12_3202 ();
 sg13g2_decap_8 FILLER_12_3209 ();
 sg13g2_decap_8 FILLER_12_3216 ();
 sg13g2_decap_4 FILLER_12_3223 ();
 sg13g2_fill_1 FILLER_12_3227 ();
 sg13g2_fill_1 FILLER_12_3242 ();
 sg13g2_decap_8 FILLER_12_3297 ();
 sg13g2_fill_2 FILLER_12_3304 ();
 sg13g2_fill_2 FILLER_12_3343 ();
 sg13g2_fill_1 FILLER_12_3345 ();
 sg13g2_decap_8 FILLER_12_3350 ();
 sg13g2_fill_2 FILLER_12_3357 ();
 sg13g2_fill_1 FILLER_12_3359 ();
 sg13g2_decap_8 FILLER_12_3400 ();
 sg13g2_decap_8 FILLER_12_3407 ();
 sg13g2_decap_8 FILLER_12_3414 ();
 sg13g2_decap_4 FILLER_12_3421 ();
 sg13g2_fill_2 FILLER_12_3425 ();
 sg13g2_decap_4 FILLER_12_3431 ();
 sg13g2_fill_2 FILLER_12_3435 ();
 sg13g2_fill_2 FILLER_12_3452 ();
 sg13g2_decap_8 FILLER_12_3481 ();
 sg13g2_decap_8 FILLER_12_3488 ();
 sg13g2_decap_8 FILLER_12_3495 ();
 sg13g2_decap_8 FILLER_12_3502 ();
 sg13g2_decap_8 FILLER_12_3509 ();
 sg13g2_fill_2 FILLER_12_3516 ();
 sg13g2_decap_4 FILLER_12_3528 ();
 sg13g2_fill_1 FILLER_12_3532 ();
 sg13g2_fill_1 FILLER_12_3537 ();
 sg13g2_decap_8 FILLER_12_3547 ();
 sg13g2_decap_8 FILLER_12_3554 ();
 sg13g2_decap_8 FILLER_12_3561 ();
 sg13g2_decap_8 FILLER_12_3568 ();
 sg13g2_fill_2 FILLER_12_3575 ();
 sg13g2_fill_1 FILLER_12_3577 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_67 ();
 sg13g2_decap_4 FILLER_13_72 ();
 sg13g2_decap_8 FILLER_13_107 ();
 sg13g2_decap_8 FILLER_13_114 ();
 sg13g2_fill_1 FILLER_13_121 ();
 sg13g2_fill_2 FILLER_13_135 ();
 sg13g2_decap_8 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_decap_4 FILLER_13_165 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_decap_8 FILLER_13_177 ();
 sg13g2_decap_8 FILLER_13_184 ();
 sg13g2_decap_8 FILLER_13_191 ();
 sg13g2_decap_8 FILLER_13_215 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_4 FILLER_13_277 ();
 sg13g2_fill_1 FILLER_13_281 ();
 sg13g2_fill_2 FILLER_13_310 ();
 sg13g2_fill_2 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_fill_2 FILLER_13_385 ();
 sg13g2_decap_4 FILLER_13_432 ();
 sg13g2_fill_1 FILLER_13_436 ();
 sg13g2_fill_1 FILLER_13_474 ();
 sg13g2_fill_2 FILLER_13_493 ();
 sg13g2_decap_8 FILLER_13_544 ();
 sg13g2_fill_1 FILLER_13_551 ();
 sg13g2_decap_4 FILLER_13_558 ();
 sg13g2_fill_1 FILLER_13_562 ();
 sg13g2_fill_2 FILLER_13_603 ();
 sg13g2_fill_1 FILLER_13_627 ();
 sg13g2_decap_8 FILLER_13_633 ();
 sg13g2_decap_4 FILLER_13_640 ();
 sg13g2_fill_2 FILLER_13_644 ();
 sg13g2_fill_2 FILLER_13_701 ();
 sg13g2_fill_1 FILLER_13_703 ();
 sg13g2_fill_2 FILLER_13_713 ();
 sg13g2_fill_1 FILLER_13_715 ();
 sg13g2_decap_4 FILLER_13_742 ();
 sg13g2_fill_1 FILLER_13_746 ();
 sg13g2_decap_4 FILLER_13_752 ();
 sg13g2_fill_1 FILLER_13_756 ();
 sg13g2_fill_2 FILLER_13_802 ();
 sg13g2_fill_1 FILLER_13_804 ();
 sg13g2_decap_8 FILLER_13_810 ();
 sg13g2_decap_8 FILLER_13_817 ();
 sg13g2_decap_8 FILLER_13_824 ();
 sg13g2_decap_8 FILLER_13_831 ();
 sg13g2_decap_4 FILLER_13_838 ();
 sg13g2_fill_2 FILLER_13_842 ();
 sg13g2_decap_8 FILLER_13_885 ();
 sg13g2_fill_1 FILLER_13_892 ();
 sg13g2_fill_2 FILLER_13_907 ();
 sg13g2_fill_1 FILLER_13_909 ();
 sg13g2_fill_1 FILLER_13_922 ();
 sg13g2_fill_1 FILLER_13_939 ();
 sg13g2_fill_2 FILLER_13_951 ();
 sg13g2_fill_1 FILLER_13_953 ();
 sg13g2_fill_1 FILLER_13_975 ();
 sg13g2_fill_2 FILLER_13_1004 ();
 sg13g2_fill_1 FILLER_13_1006 ();
 sg13g2_decap_4 FILLER_13_1048 ();
 sg13g2_fill_1 FILLER_13_1090 ();
 sg13g2_fill_1 FILLER_13_1117 ();
 sg13g2_fill_2 FILLER_13_1127 ();
 sg13g2_fill_2 FILLER_13_1180 ();
 sg13g2_decap_8 FILLER_13_1191 ();
 sg13g2_decap_8 FILLER_13_1198 ();
 sg13g2_decap_8 FILLER_13_1205 ();
 sg13g2_decap_4 FILLER_13_1212 ();
 sg13g2_decap_4 FILLER_13_1232 ();
 sg13g2_decap_8 FILLER_13_1259 ();
 sg13g2_decap_8 FILLER_13_1266 ();
 sg13g2_decap_8 FILLER_13_1273 ();
 sg13g2_fill_1 FILLER_13_1280 ();
 sg13g2_decap_8 FILLER_13_1320 ();
 sg13g2_fill_1 FILLER_13_1327 ();
 sg13g2_decap_8 FILLER_13_1337 ();
 sg13g2_decap_4 FILLER_13_1344 ();
 sg13g2_decap_8 FILLER_13_1370 ();
 sg13g2_fill_2 FILLER_13_1377 ();
 sg13g2_fill_1 FILLER_13_1379 ();
 sg13g2_decap_4 FILLER_13_1438 ();
 sg13g2_decap_8 FILLER_13_1479 ();
 sg13g2_decap_4 FILLER_13_1486 ();
 sg13g2_fill_2 FILLER_13_1490 ();
 sg13g2_fill_1 FILLER_13_1506 ();
 sg13g2_decap_8 FILLER_13_1522 ();
 sg13g2_decap_8 FILLER_13_1529 ();
 sg13g2_decap_4 FILLER_13_1540 ();
 sg13g2_decap_4 FILLER_13_1548 ();
 sg13g2_fill_2 FILLER_13_1567 ();
 sg13g2_fill_2 FILLER_13_1580 ();
 sg13g2_fill_1 FILLER_13_1587 ();
 sg13g2_decap_8 FILLER_13_1593 ();
 sg13g2_fill_2 FILLER_13_1600 ();
 sg13g2_decap_8 FILLER_13_1637 ();
 sg13g2_decap_4 FILLER_13_1644 ();
 sg13g2_fill_1 FILLER_13_1648 ();
 sg13g2_fill_1 FILLER_13_1667 ();
 sg13g2_decap_4 FILLER_13_1694 ();
 sg13g2_fill_1 FILLER_13_1698 ();
 sg13g2_fill_2 FILLER_13_1735 ();
 sg13g2_fill_2 FILLER_13_1768 ();
 sg13g2_fill_2 FILLER_13_1775 ();
 sg13g2_fill_1 FILLER_13_1777 ();
 sg13g2_fill_2 FILLER_13_1812 ();
 sg13g2_fill_1 FILLER_13_1814 ();
 sg13g2_fill_1 FILLER_13_1859 ();
 sg13g2_decap_8 FILLER_13_1873 ();
 sg13g2_decap_4 FILLER_13_1880 ();
 sg13g2_fill_1 FILLER_13_1884 ();
 sg13g2_decap_8 FILLER_13_1926 ();
 sg13g2_fill_2 FILLER_13_1933 ();
 sg13g2_decap_8 FILLER_13_1966 ();
 sg13g2_decap_4 FILLER_13_1973 ();
 sg13g2_fill_2 FILLER_13_1977 ();
 sg13g2_decap_8 FILLER_13_2007 ();
 sg13g2_decap_4 FILLER_13_2042 ();
 sg13g2_fill_2 FILLER_13_2046 ();
 sg13g2_decap_8 FILLER_13_2061 ();
 sg13g2_decap_4 FILLER_13_2068 ();
 sg13g2_fill_1 FILLER_13_2072 ();
 sg13g2_fill_2 FILLER_13_2082 ();
 sg13g2_fill_1 FILLER_13_2098 ();
 sg13g2_decap_4 FILLER_13_2125 ();
 sg13g2_fill_1 FILLER_13_2129 ();
 sg13g2_fill_2 FILLER_13_2139 ();
 sg13g2_fill_2 FILLER_13_2186 ();
 sg13g2_fill_1 FILLER_13_2188 ();
 sg13g2_decap_4 FILLER_13_2245 ();
 sg13g2_decap_4 FILLER_13_2296 ();
 sg13g2_fill_1 FILLER_13_2312 ();
 sg13g2_fill_1 FILLER_13_2320 ();
 sg13g2_decap_8 FILLER_13_2348 ();
 sg13g2_decap_8 FILLER_13_2355 ();
 sg13g2_decap_4 FILLER_13_2362 ();
 sg13g2_fill_1 FILLER_13_2366 ();
 sg13g2_decap_8 FILLER_13_2415 ();
 sg13g2_decap_8 FILLER_13_2422 ();
 sg13g2_decap_4 FILLER_13_2469 ();
 sg13g2_fill_1 FILLER_13_2495 ();
 sg13g2_fill_1 FILLER_13_2514 ();
 sg13g2_decap_4 FILLER_13_2519 ();
 sg13g2_fill_2 FILLER_13_2523 ();
 sg13g2_fill_1 FILLER_13_2560 ();
 sg13g2_decap_4 FILLER_13_2574 ();
 sg13g2_fill_2 FILLER_13_2582 ();
 sg13g2_fill_1 FILLER_13_2584 ();
 sg13g2_decap_4 FILLER_13_2604 ();
 sg13g2_fill_2 FILLER_13_2608 ();
 sg13g2_decap_8 FILLER_13_2629 ();
 sg13g2_decap_8 FILLER_13_2640 ();
 sg13g2_decap_8 FILLER_13_2684 ();
 sg13g2_decap_8 FILLER_13_2691 ();
 sg13g2_decap_8 FILLER_13_2698 ();
 sg13g2_decap_8 FILLER_13_2705 ();
 sg13g2_decap_4 FILLER_13_2712 ();
 sg13g2_fill_2 FILLER_13_2716 ();
 sg13g2_decap_8 FILLER_13_2745 ();
 sg13g2_decap_4 FILLER_13_2752 ();
 sg13g2_fill_2 FILLER_13_2756 ();
 sg13g2_fill_2 FILLER_13_2799 ();
 sg13g2_fill_1 FILLER_13_2801 ();
 sg13g2_decap_4 FILLER_13_2816 ();
 sg13g2_decap_8 FILLER_13_2838 ();
 sg13g2_decap_4 FILLER_13_2845 ();
 sg13g2_fill_2 FILLER_13_2883 ();
 sg13g2_fill_1 FILLER_13_2885 ();
 sg13g2_decap_8 FILLER_13_2903 ();
 sg13g2_decap_8 FILLER_13_2910 ();
 sg13g2_decap_8 FILLER_13_2917 ();
 sg13g2_decap_4 FILLER_13_2924 ();
 sg13g2_decap_8 FILLER_13_2959 ();
 sg13g2_decap_8 FILLER_13_2966 ();
 sg13g2_decap_4 FILLER_13_2973 ();
 sg13g2_decap_4 FILLER_13_3027 ();
 sg13g2_fill_1 FILLER_13_3031 ();
 sg13g2_fill_1 FILLER_13_3059 ();
 sg13g2_decap_8 FILLER_13_3133 ();
 sg13g2_fill_2 FILLER_13_3140 ();
 sg13g2_fill_2 FILLER_13_3169 ();
 sg13g2_decap_8 FILLER_13_3207 ();
 sg13g2_decap_8 FILLER_13_3214 ();
 sg13g2_fill_2 FILLER_13_3221 ();
 sg13g2_fill_1 FILLER_13_3223 ();
 sg13g2_decap_8 FILLER_13_3286 ();
 sg13g2_decap_8 FILLER_13_3293 ();
 sg13g2_fill_1 FILLER_13_3300 ();
 sg13g2_decap_8 FILLER_13_3355 ();
 sg13g2_fill_2 FILLER_13_3362 ();
 sg13g2_fill_1 FILLER_13_3364 ();
 sg13g2_fill_1 FILLER_13_3379 ();
 sg13g2_fill_2 FILLER_13_3393 ();
 sg13g2_fill_1 FILLER_13_3395 ();
 sg13g2_decap_8 FILLER_13_3423 ();
 sg13g2_fill_1 FILLER_13_3430 ();
 sg13g2_fill_2 FILLER_13_3471 ();
 sg13g2_fill_1 FILLER_13_3473 ();
 sg13g2_decap_8 FILLER_13_3511 ();
 sg13g2_decap_8 FILLER_13_3555 ();
 sg13g2_decap_8 FILLER_13_3562 ();
 sg13g2_decap_8 FILLER_13_3569 ();
 sg13g2_fill_2 FILLER_13_3576 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_52 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_decap_4 FILLER_14_131 ();
 sg13g2_decap_8 FILLER_14_183 ();
 sg13g2_decap_8 FILLER_14_190 ();
 sg13g2_decap_8 FILLER_14_197 ();
 sg13g2_decap_8 FILLER_14_204 ();
 sg13g2_decap_8 FILLER_14_211 ();
 sg13g2_decap_4 FILLER_14_277 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_decap_8 FILLER_14_295 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_fill_1 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_378 ();
 sg13g2_fill_2 FILLER_14_416 ();
 sg13g2_fill_1 FILLER_14_418 ();
 sg13g2_decap_4 FILLER_14_438 ();
 sg13g2_fill_1 FILLER_14_442 ();
 sg13g2_fill_1 FILLER_14_475 ();
 sg13g2_decap_8 FILLER_14_549 ();
 sg13g2_fill_2 FILLER_14_556 ();
 sg13g2_fill_1 FILLER_14_558 ();
 sg13g2_decap_4 FILLER_14_576 ();
 sg13g2_fill_2 FILLER_14_604 ();
 sg13g2_fill_2 FILLER_14_634 ();
 sg13g2_fill_1 FILLER_14_636 ();
 sg13g2_fill_2 FILLER_14_647 ();
 sg13g2_fill_1 FILLER_14_649 ();
 sg13g2_decap_4 FILLER_14_661 ();
 sg13g2_decap_8 FILLER_14_680 ();
 sg13g2_decap_8 FILLER_14_687 ();
 sg13g2_decap_8 FILLER_14_694 ();
 sg13g2_decap_8 FILLER_14_709 ();
 sg13g2_fill_1 FILLER_14_716 ();
 sg13g2_fill_1 FILLER_14_720 ();
 sg13g2_decap_8 FILLER_14_726 ();
 sg13g2_decap_4 FILLER_14_754 ();
 sg13g2_fill_2 FILLER_14_758 ();
 sg13g2_fill_1 FILLER_14_788 ();
 sg13g2_fill_2 FILLER_14_798 ();
 sg13g2_fill_1 FILLER_14_800 ();
 sg13g2_fill_2 FILLER_14_809 ();
 sg13g2_fill_1 FILLER_14_811 ();
 sg13g2_fill_2 FILLER_14_818 ();
 sg13g2_fill_2 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_836 ();
 sg13g2_decap_8 FILLER_14_843 ();
 sg13g2_fill_2 FILLER_14_850 ();
 sg13g2_fill_1 FILLER_14_852 ();
 sg13g2_fill_1 FILLER_14_879 ();
 sg13g2_decap_4 FILLER_14_884 ();
 sg13g2_fill_2 FILLER_14_891 ();
 sg13g2_fill_2 FILLER_14_922 ();
 sg13g2_fill_1 FILLER_14_924 ();
 sg13g2_decap_4 FILLER_14_957 ();
 sg13g2_fill_1 FILLER_14_961 ();
 sg13g2_fill_2 FILLER_14_970 ();
 sg13g2_fill_2 FILLER_14_1000 ();
 sg13g2_decap_8 FILLER_14_1019 ();
 sg13g2_decap_8 FILLER_14_1026 ();
 sg13g2_decap_8 FILLER_14_1033 ();
 sg13g2_decap_8 FILLER_14_1040 ();
 sg13g2_decap_4 FILLER_14_1047 ();
 sg13g2_fill_2 FILLER_14_1051 ();
 sg13g2_decap_4 FILLER_14_1090 ();
 sg13g2_decap_8 FILLER_14_1126 ();
 sg13g2_decap_4 FILLER_14_1133 ();
 sg13g2_fill_2 FILLER_14_1137 ();
 sg13g2_fill_1 FILLER_14_1142 ();
 sg13g2_fill_2 FILLER_14_1152 ();
 sg13g2_fill_1 FILLER_14_1154 ();
 sg13g2_fill_2 FILLER_14_1173 ();
 sg13g2_decap_8 FILLER_14_1180 ();
 sg13g2_decap_8 FILLER_14_1215 ();
 sg13g2_decap_8 FILLER_14_1267 ();
 sg13g2_fill_2 FILLER_14_1274 ();
 sg13g2_fill_1 FILLER_14_1276 ();
 sg13g2_fill_1 FILLER_14_1306 ();
 sg13g2_decap_8 FILLER_14_1324 ();
 sg13g2_decap_8 FILLER_14_1331 ();
 sg13g2_decap_4 FILLER_14_1338 ();
 sg13g2_fill_2 FILLER_14_1342 ();
 sg13g2_fill_2 FILLER_14_1376 ();
 sg13g2_fill_1 FILLER_14_1405 ();
 sg13g2_decap_8 FILLER_14_1419 ();
 sg13g2_decap_8 FILLER_14_1426 ();
 sg13g2_decap_8 FILLER_14_1433 ();
 sg13g2_fill_2 FILLER_14_1440 ();
 sg13g2_decap_4 FILLER_14_1487 ();
 sg13g2_fill_2 FILLER_14_1491 ();
 sg13g2_fill_2 FILLER_14_1506 ();
 sg13g2_fill_1 FILLER_14_1519 ();
 sg13g2_fill_2 FILLER_14_1536 ();
 sg13g2_fill_1 FILLER_14_1538 ();
 sg13g2_fill_2 FILLER_14_1550 ();
 sg13g2_fill_1 FILLER_14_1552 ();
 sg13g2_fill_2 FILLER_14_1584 ();
 sg13g2_fill_1 FILLER_14_1586 ();
 sg13g2_decap_4 FILLER_14_1594 ();
 sg13g2_fill_1 FILLER_14_1604 ();
 sg13g2_fill_2 FILLER_14_1618 ();
 sg13g2_decap_8 FILLER_14_1642 ();
 sg13g2_decap_4 FILLER_14_1649 ();
 sg13g2_fill_2 FILLER_14_1653 ();
 sg13g2_decap_8 FILLER_14_1686 ();
 sg13g2_decap_4 FILLER_14_1693 ();
 sg13g2_fill_1 FILLER_14_1697 ();
 sg13g2_fill_2 FILLER_14_1707 ();
 sg13g2_fill_1 FILLER_14_1709 ();
 sg13g2_fill_2 FILLER_14_1726 ();
 sg13g2_fill_1 FILLER_14_1742 ();
 sg13g2_fill_2 FILLER_14_1774 ();
 sg13g2_fill_1 FILLER_14_1776 ();
 sg13g2_fill_1 FILLER_14_1781 ();
 sg13g2_decap_4 FILLER_14_1828 ();
 sg13g2_fill_2 FILLER_14_1832 ();
 sg13g2_fill_2 FILLER_14_1839 ();
 sg13g2_fill_1 FILLER_14_1841 ();
 sg13g2_decap_8 FILLER_14_1855 ();
 sg13g2_decap_8 FILLER_14_1862 ();
 sg13g2_decap_8 FILLER_14_1869 ();
 sg13g2_decap_8 FILLER_14_1876 ();
 sg13g2_decap_8 FILLER_14_1928 ();
 sg13g2_fill_2 FILLER_14_1935 ();
 sg13g2_fill_1 FILLER_14_1937 ();
 sg13g2_decap_4 FILLER_14_1972 ();
 sg13g2_fill_1 FILLER_14_1976 ();
 sg13g2_fill_2 FILLER_14_1991 ();
 sg13g2_decap_8 FILLER_14_2005 ();
 sg13g2_decap_8 FILLER_14_2012 ();
 sg13g2_fill_1 FILLER_14_2019 ();
 sg13g2_decap_8 FILLER_14_2070 ();
 sg13g2_decap_4 FILLER_14_2077 ();
 sg13g2_fill_1 FILLER_14_2081 ();
 sg13g2_decap_8 FILLER_14_2109 ();
 sg13g2_decap_8 FILLER_14_2116 ();
 sg13g2_decap_8 FILLER_14_2131 ();
 sg13g2_decap_4 FILLER_14_2138 ();
 sg13g2_fill_1 FILLER_14_2142 ();
 sg13g2_fill_1 FILLER_14_2148 ();
 sg13g2_fill_2 FILLER_14_2158 ();
 sg13g2_fill_1 FILLER_14_2160 ();
 sg13g2_decap_8 FILLER_14_2166 ();
 sg13g2_fill_1 FILLER_14_2173 ();
 sg13g2_fill_2 FILLER_14_2178 ();
 sg13g2_fill_1 FILLER_14_2180 ();
 sg13g2_decap_8 FILLER_14_2226 ();
 sg13g2_decap_8 FILLER_14_2233 ();
 sg13g2_fill_2 FILLER_14_2240 ();
 sg13g2_fill_2 FILLER_14_2247 ();
 sg13g2_decap_8 FILLER_14_2295 ();
 sg13g2_decap_8 FILLER_14_2348 ();
 sg13g2_decap_4 FILLER_14_2355 ();
 sg13g2_fill_1 FILLER_14_2359 ();
 sg13g2_fill_2 FILLER_14_2391 ();
 sg13g2_fill_1 FILLER_14_2393 ();
 sg13g2_decap_8 FILLER_14_2421 ();
 sg13g2_decap_4 FILLER_14_2428 ();
 sg13g2_fill_2 FILLER_14_2432 ();
 sg13g2_decap_4 FILLER_14_2438 ();
 sg13g2_decap_8 FILLER_14_2452 ();
 sg13g2_decap_8 FILLER_14_2459 ();
 sg13g2_decap_8 FILLER_14_2476 ();
 sg13g2_decap_8 FILLER_14_2483 ();
 sg13g2_fill_1 FILLER_14_2490 ();
 sg13g2_decap_8 FILLER_14_2496 ();
 sg13g2_decap_8 FILLER_14_2508 ();
 sg13g2_decap_8 FILLER_14_2519 ();
 sg13g2_fill_2 FILLER_14_2526 ();
 sg13g2_decap_4 FILLER_14_2538 ();
 sg13g2_fill_1 FILLER_14_2542 ();
 sg13g2_fill_2 FILLER_14_2557 ();
 sg13g2_fill_1 FILLER_14_2559 ();
 sg13g2_decap_8 FILLER_14_2569 ();
 sg13g2_decap_8 FILLER_14_2576 ();
 sg13g2_fill_2 FILLER_14_2583 ();
 sg13g2_decap_8 FILLER_14_2598 ();
 sg13g2_fill_2 FILLER_14_2605 ();
 sg13g2_fill_2 FILLER_14_2616 ();
 sg13g2_decap_8 FILLER_14_2637 ();
 sg13g2_decap_8 FILLER_14_2686 ();
 sg13g2_decap_8 FILLER_14_2693 ();
 sg13g2_fill_2 FILLER_14_2700 ();
 sg13g2_fill_1 FILLER_14_2702 ();
 sg13g2_decap_4 FILLER_14_2740 ();
 sg13g2_fill_1 FILLER_14_2744 ();
 sg13g2_decap_8 FILLER_14_2749 ();
 sg13g2_decap_4 FILLER_14_2756 ();
 sg13g2_fill_2 FILLER_14_2760 ();
 sg13g2_fill_1 FILLER_14_2807 ();
 sg13g2_decap_8 FILLER_14_2835 ();
 sg13g2_decap_4 FILLER_14_2842 ();
 sg13g2_fill_2 FILLER_14_2846 ();
 sg13g2_decap_8 FILLER_14_2893 ();
 sg13g2_decap_4 FILLER_14_2900 ();
 sg13g2_fill_2 FILLER_14_2904 ();
 sg13g2_decap_8 FILLER_14_2911 ();
 sg13g2_decap_8 FILLER_14_2918 ();
 sg13g2_fill_1 FILLER_14_2925 ();
 sg13g2_fill_2 FILLER_14_2949 ();
 sg13g2_decap_8 FILLER_14_2960 ();
 sg13g2_decap_8 FILLER_14_2967 ();
 sg13g2_fill_2 FILLER_14_2974 ();
 sg13g2_fill_1 FILLER_14_2976 ();
 sg13g2_fill_2 FILLER_14_3000 ();
 sg13g2_decap_8 FILLER_14_3023 ();
 sg13g2_fill_2 FILLER_14_3030 ();
 sg13g2_fill_1 FILLER_14_3032 ();
 sg13g2_fill_2 FILLER_14_3047 ();
 sg13g2_fill_1 FILLER_14_3049 ();
 sg13g2_fill_2 FILLER_14_3063 ();
 sg13g2_fill_1 FILLER_14_3065 ();
 sg13g2_decap_4 FILLER_14_3070 ();
 sg13g2_fill_1 FILLER_14_3096 ();
 sg13g2_decap_4 FILLER_14_3106 ();
 sg13g2_fill_2 FILLER_14_3110 ();
 sg13g2_decap_8 FILLER_14_3120 ();
 sg13g2_decap_8 FILLER_14_3127 ();
 sg13g2_fill_2 FILLER_14_3134 ();
 sg13g2_decap_4 FILLER_14_3140 ();
 sg13g2_fill_2 FILLER_14_3158 ();
 sg13g2_fill_1 FILLER_14_3214 ();
 sg13g2_fill_2 FILLER_14_3246 ();
 sg13g2_fill_2 FILLER_14_3252 ();
 sg13g2_decap_8 FILLER_14_3273 ();
 sg13g2_fill_1 FILLER_14_3280 ();
 sg13g2_decap_8 FILLER_14_3285 ();
 sg13g2_decap_8 FILLER_14_3292 ();
 sg13g2_decap_8 FILLER_14_3299 ();
 sg13g2_fill_2 FILLER_14_3306 ();
 sg13g2_fill_1 FILLER_14_3308 ();
 sg13g2_decap_8 FILLER_14_3361 ();
 sg13g2_decap_8 FILLER_14_3368 ();
 sg13g2_fill_2 FILLER_14_3375 ();
 sg13g2_decap_8 FILLER_14_3424 ();
 sg13g2_fill_2 FILLER_14_3431 ();
 sg13g2_fill_2 FILLER_14_3517 ();
 sg13g2_decap_8 FILLER_14_3571 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_58 ();
 sg13g2_fill_1 FILLER_15_60 ();
 sg13g2_fill_1 FILLER_15_109 ();
 sg13g2_fill_2 FILLER_15_132 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_4 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_436 ();
 sg13g2_decap_4 FILLER_15_443 ();
 sg13g2_fill_2 FILLER_15_447 ();
 sg13g2_fill_1 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_538 ();
 sg13g2_decap_8 FILLER_15_545 ();
 sg13g2_decap_8 FILLER_15_552 ();
 sg13g2_decap_8 FILLER_15_559 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_fill_1 FILLER_15_578 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_decap_8 FILLER_15_690 ();
 sg13g2_decap_4 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_739 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_fill_1 FILLER_15_753 ();
 sg13g2_fill_2 FILLER_15_771 ();
 sg13g2_fill_2 FILLER_15_778 ();
 sg13g2_fill_2 FILLER_15_802 ();
 sg13g2_decap_4 FILLER_15_836 ();
 sg13g2_fill_1 FILLER_15_840 ();
 sg13g2_fill_1 FILLER_15_855 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_878 ();
 sg13g2_decap_8 FILLER_15_891 ();
 sg13g2_fill_2 FILLER_15_898 ();
 sg13g2_fill_1 FILLER_15_925 ();
 sg13g2_decap_8 FILLER_15_954 ();
 sg13g2_fill_1 FILLER_15_961 ();
 sg13g2_decap_8 FILLER_15_975 ();
 sg13g2_fill_1 FILLER_15_991 ();
 sg13g2_fill_2 FILLER_15_1005 ();
 sg13g2_fill_1 FILLER_15_1007 ();
 sg13g2_decap_8 FILLER_15_1012 ();
 sg13g2_fill_1 FILLER_15_1019 ();
 sg13g2_decap_8 FILLER_15_1046 ();
 sg13g2_decap_8 FILLER_15_1053 ();
 sg13g2_fill_2 FILLER_15_1060 ();
 sg13g2_decap_8 FILLER_15_1065 ();
 sg13g2_decap_4 FILLER_15_1072 ();
 sg13g2_fill_1 FILLER_15_1108 ();
 sg13g2_decap_8 FILLER_15_1122 ();
 sg13g2_decap_8 FILLER_15_1129 ();
 sg13g2_fill_2 FILLER_15_1136 ();
 sg13g2_fill_1 FILLER_15_1138 ();
 sg13g2_fill_1 FILLER_15_1167 ();
 sg13g2_decap_4 FILLER_15_1177 ();
 sg13g2_decap_8 FILLER_15_1215 ();
 sg13g2_decap_8 FILLER_15_1222 ();
 sg13g2_fill_2 FILLER_15_1229 ();
 sg13g2_fill_1 FILLER_15_1231 ();
 sg13g2_fill_1 FILLER_15_1274 ();
 sg13g2_fill_2 FILLER_15_1346 ();
 sg13g2_fill_1 FILLER_15_1348 ();
 sg13g2_decap_8 FILLER_15_1371 ();
 sg13g2_fill_2 FILLER_15_1378 ();
 sg13g2_fill_1 FILLER_15_1380 ();
 sg13g2_fill_2 FILLER_15_1417 ();
 sg13g2_fill_2 FILLER_15_1481 ();
 sg13g2_fill_2 FILLER_15_1492 ();
 sg13g2_fill_2 FILLER_15_1500 ();
 sg13g2_decap_8 FILLER_15_1522 ();
 sg13g2_decap_4 FILLER_15_1548 ();
 sg13g2_decap_4 FILLER_15_1571 ();
 sg13g2_fill_2 FILLER_15_1584 ();
 sg13g2_decap_8 FILLER_15_1593 ();
 sg13g2_decap_8 FILLER_15_1600 ();
 sg13g2_decap_4 FILLER_15_1607 ();
 sg13g2_decap_4 FILLER_15_1647 ();
 sg13g2_fill_2 FILLER_15_1651 ();
 sg13g2_fill_1 FILLER_15_1677 ();
 sg13g2_decap_8 FILLER_15_1693 ();
 sg13g2_decap_4 FILLER_15_1700 ();
 sg13g2_fill_2 FILLER_15_1710 ();
 sg13g2_fill_1 FILLER_15_1712 ();
 sg13g2_fill_2 FILLER_15_1718 ();
 sg13g2_fill_1 FILLER_15_1720 ();
 sg13g2_fill_2 FILLER_15_1727 ();
 sg13g2_fill_1 FILLER_15_1729 ();
 sg13g2_decap_4 FILLER_15_1752 ();
 sg13g2_fill_1 FILLER_15_1782 ();
 sg13g2_decap_8 FILLER_15_1792 ();
 sg13g2_decap_8 FILLER_15_1799 ();
 sg13g2_decap_4 FILLER_15_1806 ();
 sg13g2_fill_1 FILLER_15_1810 ();
 sg13g2_decap_8 FILLER_15_1820 ();
 sg13g2_fill_2 FILLER_15_1827 ();
 sg13g2_fill_1 FILLER_15_1829 ();
 sg13g2_decap_8 FILLER_15_1867 ();
 sg13g2_decap_8 FILLER_15_1874 ();
 sg13g2_decap_4 FILLER_15_1881 ();
 sg13g2_fill_1 FILLER_15_1885 ();
 sg13g2_fill_1 FILLER_15_1892 ();
 sg13g2_decap_8 FILLER_15_1919 ();
 sg13g2_fill_2 FILLER_15_1926 ();
 sg13g2_fill_1 FILLER_15_1928 ();
 sg13g2_decap_4 FILLER_15_1933 ();
 sg13g2_fill_2 FILLER_15_1937 ();
 sg13g2_decap_8 FILLER_15_1970 ();
 sg13g2_decap_4 FILLER_15_1977 ();
 sg13g2_fill_2 FILLER_15_1981 ();
 sg13g2_fill_2 FILLER_15_1993 ();
 sg13g2_fill_1 FILLER_15_1995 ();
 sg13g2_fill_2 FILLER_15_2014 ();
 sg13g2_fill_1 FILLER_15_2016 ();
 sg13g2_decap_4 FILLER_15_2021 ();
 sg13g2_fill_1 FILLER_15_2025 ();
 sg13g2_fill_2 FILLER_15_2049 ();
 sg13g2_fill_1 FILLER_15_2072 ();
 sg13g2_decap_8 FILLER_15_2077 ();
 sg13g2_decap_8 FILLER_15_2084 ();
 sg13g2_decap_4 FILLER_15_2091 ();
 sg13g2_decap_8 FILLER_15_2099 ();
 sg13g2_decap_4 FILLER_15_2106 ();
 sg13g2_fill_1 FILLER_15_2110 ();
 sg13g2_decap_8 FILLER_15_2143 ();
 sg13g2_fill_2 FILLER_15_2150 ();
 sg13g2_fill_1 FILLER_15_2152 ();
 sg13g2_decap_8 FILLER_15_2170 ();
 sg13g2_decap_8 FILLER_15_2177 ();
 sg13g2_decap_8 FILLER_15_2184 ();
 sg13g2_fill_1 FILLER_15_2191 ();
 sg13g2_decap_4 FILLER_15_2197 ();
 sg13g2_fill_1 FILLER_15_2201 ();
 sg13g2_decap_8 FILLER_15_2226 ();
 sg13g2_decap_8 FILLER_15_2233 ();
 sg13g2_fill_1 FILLER_15_2253 ();
 sg13g2_fill_2 FILLER_15_2268 ();
 sg13g2_fill_1 FILLER_15_2270 ();
 sg13g2_decap_4 FILLER_15_2293 ();
 sg13g2_fill_1 FILLER_15_2297 ();
 sg13g2_fill_1 FILLER_15_2303 ();
 sg13g2_fill_1 FILLER_15_2344 ();
 sg13g2_decap_8 FILLER_15_2358 ();
 sg13g2_fill_2 FILLER_15_2365 ();
 sg13g2_decap_8 FILLER_15_2427 ();
 sg13g2_decap_8 FILLER_15_2434 ();
 sg13g2_fill_2 FILLER_15_2441 ();
 sg13g2_decap_4 FILLER_15_2452 ();
 sg13g2_fill_2 FILLER_15_2456 ();
 sg13g2_decap_8 FILLER_15_2477 ();
 sg13g2_decap_8 FILLER_15_2484 ();
 sg13g2_decap_4 FILLER_15_2491 ();
 sg13g2_decap_8 FILLER_15_2500 ();
 sg13g2_fill_2 FILLER_15_2507 ();
 sg13g2_decap_8 FILLER_15_2536 ();
 sg13g2_decap_8 FILLER_15_2552 ();
 sg13g2_decap_8 FILLER_15_2559 ();
 sg13g2_decap_8 FILLER_15_2566 ();
 sg13g2_fill_2 FILLER_15_2573 ();
 sg13g2_fill_1 FILLER_15_2602 ();
 sg13g2_fill_2 FILLER_15_2624 ();
 sg13g2_fill_1 FILLER_15_2626 ();
 sg13g2_fill_2 FILLER_15_2654 ();
 sg13g2_decap_8 FILLER_15_2678 ();
 sg13g2_decap_4 FILLER_15_2685 ();
 sg13g2_fill_2 FILLER_15_2689 ();
 sg13g2_decap_8 FILLER_15_2754 ();
 sg13g2_fill_2 FILLER_15_2761 ();
 sg13g2_decap_8 FILLER_15_2839 ();
 sg13g2_fill_2 FILLER_15_2886 ();
 sg13g2_fill_2 FILLER_15_2898 ();
 sg13g2_decap_8 FILLER_15_2927 ();
 sg13g2_fill_2 FILLER_15_2934 ();
 sg13g2_fill_1 FILLER_15_2936 ();
 sg13g2_decap_8 FILLER_15_2941 ();
 sg13g2_decap_4 FILLER_15_2948 ();
 sg13g2_decap_8 FILLER_15_2961 ();
 sg13g2_decap_8 FILLER_15_2968 ();
 sg13g2_decap_8 FILLER_15_2975 ();
 sg13g2_fill_2 FILLER_15_2982 ();
 sg13g2_decap_8 FILLER_15_3001 ();
 sg13g2_decap_8 FILLER_15_3008 ();
 sg13g2_fill_1 FILLER_15_3015 ();
 sg13g2_fill_1 FILLER_15_3029 ();
 sg13g2_decap_8 FILLER_15_3075 ();
 sg13g2_decap_8 FILLER_15_3082 ();
 sg13g2_decap_8 FILLER_15_3089 ();
 sg13g2_decap_8 FILLER_15_3096 ();
 sg13g2_decap_8 FILLER_15_3103 ();
 sg13g2_decap_4 FILLER_15_3110 ();
 sg13g2_decap_8 FILLER_15_3145 ();
 sg13g2_decap_4 FILLER_15_3152 ();
 sg13g2_fill_1 FILLER_15_3156 ();
 sg13g2_fill_1 FILLER_15_3188 ();
 sg13g2_decap_8 FILLER_15_3193 ();
 sg13g2_decap_8 FILLER_15_3200 ();
 sg13g2_decap_8 FILLER_15_3207 ();
 sg13g2_decap_8 FILLER_15_3214 ();
 sg13g2_fill_2 FILLER_15_3221 ();
 sg13g2_fill_1 FILLER_15_3223 ();
 sg13g2_decap_8 FILLER_15_3256 ();
 sg13g2_decap_4 FILLER_15_3263 ();
 sg13g2_fill_2 FILLER_15_3283 ();
 sg13g2_decap_8 FILLER_15_3295 ();
 sg13g2_decap_8 FILLER_15_3302 ();
 sg13g2_fill_2 FILLER_15_3309 ();
 sg13g2_fill_1 FILLER_15_3311 ();
 sg13g2_fill_1 FILLER_15_3331 ();
 sg13g2_decap_8 FILLER_15_3361 ();
 sg13g2_decap_8 FILLER_15_3368 ();
 sg13g2_decap_8 FILLER_15_3375 ();
 sg13g2_decap_4 FILLER_15_3382 ();
 sg13g2_decap_4 FILLER_15_3390 ();
 sg13g2_fill_1 FILLER_15_3394 ();
 sg13g2_fill_1 FILLER_15_3405 ();
 sg13g2_decap_8 FILLER_15_3431 ();
 sg13g2_decap_4 FILLER_15_3438 ();
 sg13g2_fill_2 FILLER_15_3442 ();
 sg13g2_decap_4 FILLER_15_3471 ();
 sg13g2_fill_1 FILLER_15_3485 ();
 sg13g2_fill_2 FILLER_15_3490 ();
 sg13g2_fill_1 FILLER_15_3492 ();
 sg13g2_decap_4 FILLER_15_3502 ();
 sg13g2_fill_1 FILLER_15_3565 ();
 sg13g2_fill_2 FILLER_15_3575 ();
 sg13g2_fill_1 FILLER_15_3577 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_fill_2 FILLER_16_45 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_fill_2 FILLER_16_67 ();
 sg13g2_fill_1 FILLER_16_69 ();
 sg13g2_decap_8 FILLER_16_124 ();
 sg13g2_decap_4 FILLER_16_131 ();
 sg13g2_fill_1 FILLER_16_199 ();
 sg13g2_fill_2 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_288 ();
 sg13g2_fill_1 FILLER_16_290 ();
 sg13g2_fill_1 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_16_435 ();
 sg13g2_decap_8 FILLER_16_442 ();
 sg13g2_decap_8 FILLER_16_449 ();
 sg13g2_fill_2 FILLER_16_456 ();
 sg13g2_fill_1 FILLER_16_458 ();
 sg13g2_fill_2 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_4 FILLER_16_539 ();
 sg13g2_fill_1 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_580 ();
 sg13g2_decap_8 FILLER_16_587 ();
 sg13g2_decap_8 FILLER_16_594 ();
 sg13g2_decap_8 FILLER_16_601 ();
 sg13g2_decap_8 FILLER_16_608 ();
 sg13g2_decap_8 FILLER_16_615 ();
 sg13g2_decap_8 FILLER_16_622 ();
 sg13g2_decap_4 FILLER_16_685 ();
 sg13g2_fill_1 FILLER_16_717 ();
 sg13g2_fill_2 FILLER_16_764 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_fill_1 FILLER_16_777 ();
 sg13g2_fill_2 FILLER_16_782 ();
 sg13g2_fill_1 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_789 ();
 sg13g2_decap_8 FILLER_16_796 ();
 sg13g2_fill_2 FILLER_16_803 ();
 sg13g2_fill_1 FILLER_16_805 ();
 sg13g2_decap_4 FILLER_16_825 ();
 sg13g2_decap_8 FILLER_16_834 ();
 sg13g2_decap_8 FILLER_16_841 ();
 sg13g2_decap_8 FILLER_16_848 ();
 sg13g2_decap_4 FILLER_16_855 ();
 sg13g2_fill_1 FILLER_16_864 ();
 sg13g2_decap_8 FILLER_16_869 ();
 sg13g2_decap_8 FILLER_16_876 ();
 sg13g2_decap_4 FILLER_16_883 ();
 sg13g2_decap_8 FILLER_16_890 ();
 sg13g2_decap_8 FILLER_16_897 ();
 sg13g2_fill_2 FILLER_16_917 ();
 sg13g2_decap_8 FILLER_16_932 ();
 sg13g2_decap_8 FILLER_16_943 ();
 sg13g2_decap_8 FILLER_16_950 ();
 sg13g2_decap_8 FILLER_16_957 ();
 sg13g2_fill_1 FILLER_16_964 ();
 sg13g2_fill_2 FILLER_16_974 ();
 sg13g2_fill_1 FILLER_16_976 ();
 sg13g2_decap_8 FILLER_16_990 ();
 sg13g2_fill_2 FILLER_16_997 ();
 sg13g2_fill_1 FILLER_16_999 ();
 sg13g2_decap_4 FILLER_16_1042 ();
 sg13g2_fill_1 FILLER_16_1046 ();
 sg13g2_fill_1 FILLER_16_1075 ();
 sg13g2_fill_2 FILLER_16_1085 ();
 sg13g2_decap_8 FILLER_16_1092 ();
 sg13g2_decap_8 FILLER_16_1099 ();
 sg13g2_decap_8 FILLER_16_1106 ();
 sg13g2_decap_8 FILLER_16_1113 ();
 sg13g2_decap_8 FILLER_16_1120 ();
 sg13g2_decap_8 FILLER_16_1127 ();
 sg13g2_decap_8 FILLER_16_1134 ();
 sg13g2_fill_1 FILLER_16_1141 ();
 sg13g2_fill_2 FILLER_16_1165 ();
 sg13g2_fill_1 FILLER_16_1167 ();
 sg13g2_fill_2 FILLER_16_1181 ();
 sg13g2_fill_1 FILLER_16_1183 ();
 sg13g2_decap_8 FILLER_16_1220 ();
 sg13g2_fill_2 FILLER_16_1227 ();
 sg13g2_fill_1 FILLER_16_1229 ();
 sg13g2_decap_8 FILLER_16_1261 ();
 sg13g2_decap_8 FILLER_16_1268 ();
 sg13g2_decap_8 FILLER_16_1275 ();
 sg13g2_fill_1 FILLER_16_1282 ();
 sg13g2_decap_8 FILLER_16_1335 ();
 sg13g2_decap_8 FILLER_16_1377 ();
 sg13g2_decap_8 FILLER_16_1384 ();
 sg13g2_fill_1 FILLER_16_1397 ();
 sg13g2_decap_4 FILLER_16_1404 ();
 sg13g2_fill_1 FILLER_16_1408 ();
 sg13g2_decap_4 FILLER_16_1413 ();
 sg13g2_decap_8 FILLER_16_1436 ();
 sg13g2_decap_8 FILLER_16_1443 ();
 sg13g2_decap_8 FILLER_16_1454 ();
 sg13g2_decap_4 FILLER_16_1488 ();
 sg13g2_decap_8 FILLER_16_1501 ();
 sg13g2_fill_2 FILLER_16_1508 ();
 sg13g2_decap_8 FILLER_16_1514 ();
 sg13g2_decap_8 FILLER_16_1521 ();
 sg13g2_decap_8 FILLER_16_1528 ();
 sg13g2_fill_1 FILLER_16_1535 ();
 sg13g2_decap_8 FILLER_16_1548 ();
 sg13g2_decap_8 FILLER_16_1555 ();
 sg13g2_decap_8 FILLER_16_1590 ();
 sg13g2_decap_4 FILLER_16_1597 ();
 sg13g2_decap_8 FILLER_16_1608 ();
 sg13g2_decap_8 FILLER_16_1615 ();
 sg13g2_fill_2 FILLER_16_1622 ();
 sg13g2_fill_1 FILLER_16_1624 ();
 sg13g2_decap_4 FILLER_16_1656 ();
 sg13g2_fill_2 FILLER_16_1666 ();
 sg13g2_fill_1 FILLER_16_1709 ();
 sg13g2_fill_1 FILLER_16_1717 ();
 sg13g2_fill_2 FILLER_16_1726 ();
 sg13g2_fill_1 FILLER_16_1741 ();
 sg13g2_decap_4 FILLER_16_1761 ();
 sg13g2_fill_2 FILLER_16_1770 ();
 sg13g2_fill_1 FILLER_16_1783 ();
 sg13g2_decap_8 FILLER_16_1816 ();
 sg13g2_decap_8 FILLER_16_1823 ();
 sg13g2_decap_8 FILLER_16_1830 ();
 sg13g2_decap_4 FILLER_16_1874 ();
 sg13g2_fill_1 FILLER_16_1878 ();
 sg13g2_fill_1 FILLER_16_1913 ();
 sg13g2_fill_2 FILLER_16_1968 ();
 sg13g2_fill_1 FILLER_16_1970 ();
 sg13g2_fill_1 FILLER_16_2058 ();
 sg13g2_decap_8 FILLER_16_2095 ();
 sg13g2_decap_4 FILLER_16_2102 ();
 sg13g2_fill_1 FILLER_16_2106 ();
 sg13g2_decap_4 FILLER_16_2142 ();
 sg13g2_fill_2 FILLER_16_2164 ();
 sg13g2_decap_8 FILLER_16_2174 ();
 sg13g2_decap_8 FILLER_16_2181 ();
 sg13g2_decap_8 FILLER_16_2233 ();
 sg13g2_decap_8 FILLER_16_2245 ();
 sg13g2_decap_8 FILLER_16_2279 ();
 sg13g2_decap_8 FILLER_16_2286 ();
 sg13g2_fill_2 FILLER_16_2293 ();
 sg13g2_fill_1 FILLER_16_2309 ();
 sg13g2_fill_1 FILLER_16_2317 ();
 sg13g2_decap_8 FILLER_16_2346 ();
 sg13g2_decap_8 FILLER_16_2353 ();
 sg13g2_decap_8 FILLER_16_2360 ();
 sg13g2_decap_8 FILLER_16_2367 ();
 sg13g2_fill_2 FILLER_16_2374 ();
 sg13g2_decap_8 FILLER_16_2380 ();
 sg13g2_decap_4 FILLER_16_2397 ();
 sg13g2_fill_1 FILLER_16_2401 ();
 sg13g2_decap_8 FILLER_16_2424 ();
 sg13g2_decap_8 FILLER_16_2431 ();
 sg13g2_fill_2 FILLER_16_2438 ();
 sg13g2_fill_2 FILLER_16_2467 ();
 sg13g2_fill_1 FILLER_16_2469 ();
 sg13g2_decap_4 FILLER_16_2491 ();
 sg13g2_decap_4 FILLER_16_2522 ();
 sg13g2_decap_8 FILLER_16_2553 ();
 sg13g2_decap_8 FILLER_16_2560 ();
 sg13g2_fill_1 FILLER_16_2608 ();
 sg13g2_fill_1 FILLER_16_2640 ();
 sg13g2_fill_2 FILLER_16_2645 ();
 sg13g2_decap_4 FILLER_16_2657 ();
 sg13g2_fill_2 FILLER_16_2661 ();
 sg13g2_decap_8 FILLER_16_2672 ();
 sg13g2_decap_8 FILLER_16_2679 ();
 sg13g2_decap_4 FILLER_16_2686 ();
 sg13g2_fill_2 FILLER_16_2690 ();
 sg13g2_fill_2 FILLER_16_2716 ();
 sg13g2_decap_4 FILLER_16_2752 ();
 sg13g2_fill_1 FILLER_16_2756 ();
 sg13g2_decap_8 FILLER_16_2843 ();
 sg13g2_fill_2 FILLER_16_2850 ();
 sg13g2_fill_1 FILLER_16_2852 ();
 sg13g2_fill_1 FILLER_16_2871 ();
 sg13g2_fill_2 FILLER_16_2906 ();
 sg13g2_fill_1 FILLER_16_2908 ();
 sg13g2_decap_8 FILLER_16_2918 ();
 sg13g2_decap_8 FILLER_16_2925 ();
 sg13g2_fill_2 FILLER_16_2932 ();
 sg13g2_decap_8 FILLER_16_2961 ();
 sg13g2_fill_1 FILLER_16_2968 ();
 sg13g2_decap_8 FILLER_16_2996 ();
 sg13g2_decap_8 FILLER_16_3003 ();
 sg13g2_decap_8 FILLER_16_3010 ();
 sg13g2_fill_2 FILLER_16_3017 ();
 sg13g2_decap_8 FILLER_16_3073 ();
 sg13g2_decap_8 FILLER_16_3080 ();
 sg13g2_fill_1 FILLER_16_3100 ();
 sg13g2_fill_1 FILLER_16_3111 ();
 sg13g2_decap_8 FILLER_16_3148 ();
 sg13g2_decap_4 FILLER_16_3155 ();
 sg13g2_fill_2 FILLER_16_3159 ();
 sg13g2_decap_8 FILLER_16_3200 ();
 sg13g2_decap_8 FILLER_16_3220 ();
 sg13g2_fill_2 FILLER_16_3227 ();
 sg13g2_fill_1 FILLER_16_3229 ();
 sg13g2_decap_4 FILLER_16_3243 ();
 sg13g2_fill_2 FILLER_16_3247 ();
 sg13g2_fill_1 FILLER_16_3276 ();
 sg13g2_decap_8 FILLER_16_3304 ();
 sg13g2_decap_8 FILLER_16_3311 ();
 sg13g2_decap_4 FILLER_16_3318 ();
 sg13g2_fill_2 FILLER_16_3322 ();
 sg13g2_decap_8 FILLER_16_3370 ();
 sg13g2_decap_4 FILLER_16_3377 ();
 sg13g2_fill_2 FILLER_16_3381 ();
 sg13g2_decap_8 FILLER_16_3438 ();
 sg13g2_decap_8 FILLER_16_3445 ();
 sg13g2_fill_2 FILLER_16_3452 ();
 sg13g2_fill_1 FILLER_16_3454 ();
 sg13g2_decap_8 FILLER_16_3464 ();
 sg13g2_fill_2 FILLER_16_3471 ();
 sg13g2_decap_8 FILLER_16_3483 ();
 sg13g2_decap_8 FILLER_16_3494 ();
 sg13g2_decap_8 FILLER_16_3501 ();
 sg13g2_decap_4 FILLER_16_3508 ();
 sg13g2_fill_1 FILLER_16_3512 ();
 sg13g2_fill_2 FILLER_16_3526 ();
 sg13g2_fill_2 FILLER_16_3542 ();
 sg13g2_fill_1 FILLER_16_3544 ();
 sg13g2_decap_4 FILLER_16_3572 ();
 sg13g2_fill_2 FILLER_16_3576 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_76 ();
 sg13g2_fill_2 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_114 ();
 sg13g2_decap_4 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_fill_1 FILLER_17_351 ();
 sg13g2_fill_2 FILLER_17_389 ();
 sg13g2_fill_1 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_435 ();
 sg13g2_decap_8 FILLER_17_442 ();
 sg13g2_decap_8 FILLER_17_449 ();
 sg13g2_decap_8 FILLER_17_456 ();
 sg13g2_decap_8 FILLER_17_463 ();
 sg13g2_decap_4 FILLER_17_470 ();
 sg13g2_fill_1 FILLER_17_474 ();
 sg13g2_decap_4 FILLER_17_492 ();
 sg13g2_fill_2 FILLER_17_500 ();
 sg13g2_fill_1 FILLER_17_502 ();
 sg13g2_decap_8 FILLER_17_533 ();
 sg13g2_decap_8 FILLER_17_540 ();
 sg13g2_decap_8 FILLER_17_547 ();
 sg13g2_decap_4 FILLER_17_599 ();
 sg13g2_fill_2 FILLER_17_608 ();
 sg13g2_fill_2 FILLER_17_638 ();
 sg13g2_decap_4 FILLER_17_697 ();
 sg13g2_fill_1 FILLER_17_701 ();
 sg13g2_decap_8 FILLER_17_730 ();
 sg13g2_decap_8 FILLER_17_737 ();
 sg13g2_decap_8 FILLER_17_744 ();
 sg13g2_fill_2 FILLER_17_751 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_fill_2 FILLER_17_774 ();
 sg13g2_fill_1 FILLER_17_776 ();
 sg13g2_decap_8 FILLER_17_782 ();
 sg13g2_decap_4 FILLER_17_789 ();
 sg13g2_fill_1 FILLER_17_793 ();
 sg13g2_decap_8 FILLER_17_834 ();
 sg13g2_fill_1 FILLER_17_841 ();
 sg13g2_decap_4 FILLER_17_846 ();
 sg13g2_decap_4 FILLER_17_865 ();
 sg13g2_fill_1 FILLER_17_869 ();
 sg13g2_decap_8 FILLER_17_876 ();
 sg13g2_decap_8 FILLER_17_883 ();
 sg13g2_decap_4 FILLER_17_890 ();
 sg13g2_fill_2 FILLER_17_894 ();
 sg13g2_decap_8 FILLER_17_936 ();
 sg13g2_decap_8 FILLER_17_943 ();
 sg13g2_decap_8 FILLER_17_950 ();
 sg13g2_fill_2 FILLER_17_957 ();
 sg13g2_fill_1 FILLER_17_987 ();
 sg13g2_decap_4 FILLER_17_992 ();
 sg13g2_fill_2 FILLER_17_996 ();
 sg13g2_decap_8 FILLER_17_1034 ();
 sg13g2_decap_8 FILLER_17_1041 ();
 sg13g2_decap_8 FILLER_17_1048 ();
 sg13g2_decap_8 FILLER_17_1055 ();
 sg13g2_decap_4 FILLER_17_1062 ();
 sg13g2_fill_2 FILLER_17_1093 ();
 sg13g2_fill_1 FILLER_17_1095 ();
 sg13g2_fill_2 FILLER_17_1123 ();
 sg13g2_decap_8 FILLER_17_1153 ();
 sg13g2_decap_8 FILLER_17_1160 ();
 sg13g2_decap_4 FILLER_17_1167 ();
 sg13g2_fill_1 FILLER_17_1203 ();
 sg13g2_fill_2 FILLER_17_1230 ();
 sg13g2_fill_1 FILLER_17_1263 ();
 sg13g2_decap_8 FILLER_17_1269 ();
 sg13g2_decap_8 FILLER_17_1276 ();
 sg13g2_fill_2 FILLER_17_1283 ();
 sg13g2_fill_1 FILLER_17_1285 ();
 sg13g2_fill_2 FILLER_17_1338 ();
 sg13g2_decap_8 FILLER_17_1353 ();
 sg13g2_decap_4 FILLER_17_1360 ();
 sg13g2_decap_8 FILLER_17_1373 ();
 sg13g2_decap_8 FILLER_17_1380 ();
 sg13g2_decap_8 FILLER_17_1387 ();
 sg13g2_fill_2 FILLER_17_1394 ();
 sg13g2_decap_8 FILLER_17_1432 ();
 sg13g2_decap_8 FILLER_17_1439 ();
 sg13g2_decap_4 FILLER_17_1446 ();
 sg13g2_fill_2 FILLER_17_1450 ();
 sg13g2_fill_1 FILLER_17_1492 ();
 sg13g2_fill_2 FILLER_17_1502 ();
 sg13g2_fill_2 FILLER_17_1518 ();
 sg13g2_fill_1 FILLER_17_1520 ();
 sg13g2_decap_8 FILLER_17_1531 ();
 sg13g2_decap_8 FILLER_17_1538 ();
 sg13g2_fill_2 FILLER_17_1545 ();
 sg13g2_decap_8 FILLER_17_1550 ();
 sg13g2_decap_8 FILLER_17_1557 ();
 sg13g2_fill_2 FILLER_17_1564 ();
 sg13g2_fill_1 FILLER_17_1571 ();
 sg13g2_fill_2 FILLER_17_1612 ();
 sg13g2_decap_8 FILLER_17_1619 ();
 sg13g2_decap_4 FILLER_17_1626 ();
 sg13g2_fill_2 FILLER_17_1664 ();
 sg13g2_decap_8 FILLER_17_1698 ();
 sg13g2_decap_4 FILLER_17_1705 ();
 sg13g2_fill_2 FILLER_17_1709 ();
 sg13g2_decap_8 FILLER_17_1716 ();
 sg13g2_decap_4 FILLER_17_1723 ();
 sg13g2_fill_1 FILLER_17_1727 ();
 sg13g2_fill_1 FILLER_17_1769 ();
 sg13g2_fill_1 FILLER_17_1792 ();
 sg13g2_decap_4 FILLER_17_1802 ();
 sg13g2_fill_2 FILLER_17_1806 ();
 sg13g2_fill_2 FILLER_17_1821 ();
 sg13g2_fill_1 FILLER_17_1823 ();
 sg13g2_decap_4 FILLER_17_1837 ();
 sg13g2_decap_8 FILLER_17_1872 ();
 sg13g2_decap_4 FILLER_17_1879 ();
 sg13g2_fill_1 FILLER_17_1883 ();
 sg13g2_fill_1 FILLER_17_1916 ();
 sg13g2_fill_2 FILLER_17_1931 ();
 sg13g2_fill_1 FILLER_17_1933 ();
 sg13g2_fill_2 FILLER_17_1952 ();
 sg13g2_decap_8 FILLER_17_1976 ();
 sg13g2_decap_8 FILLER_17_1983 ();
 sg13g2_decap_8 FILLER_17_1990 ();
 sg13g2_fill_2 FILLER_17_1997 ();
 sg13g2_fill_1 FILLER_17_1999 ();
 sg13g2_decap_8 FILLER_17_2072 ();
 sg13g2_fill_2 FILLER_17_2079 ();
 sg13g2_decap_4 FILLER_17_2094 ();
 sg13g2_fill_1 FILLER_17_2098 ();
 sg13g2_fill_1 FILLER_17_2134 ();
 sg13g2_decap_8 FILLER_17_2148 ();
 sg13g2_fill_2 FILLER_17_2209 ();
 sg13g2_fill_1 FILLER_17_2211 ();
 sg13g2_decap_8 FILLER_17_2226 ();
 sg13g2_decap_8 FILLER_17_2233 ();
 sg13g2_decap_8 FILLER_17_2240 ();
 sg13g2_fill_2 FILLER_17_2247 ();
 sg13g2_fill_1 FILLER_17_2249 ();
 sg13g2_decap_8 FILLER_17_2296 ();
 sg13g2_decap_8 FILLER_17_2303 ();
 sg13g2_decap_8 FILLER_17_2310 ();
 sg13g2_decap_8 FILLER_17_2317 ();
 sg13g2_decap_4 FILLER_17_2324 ();
 sg13g2_decap_8 FILLER_17_2337 ();
 sg13g2_decap_8 FILLER_17_2344 ();
 sg13g2_decap_8 FILLER_17_2351 ();
 sg13g2_decap_8 FILLER_17_2358 ();
 sg13g2_decap_8 FILLER_17_2365 ();
 sg13g2_decap_8 FILLER_17_2372 ();
 sg13g2_decap_8 FILLER_17_2379 ();
 sg13g2_fill_2 FILLER_17_2386 ();
 sg13g2_fill_1 FILLER_17_2388 ();
 sg13g2_decap_8 FILLER_17_2425 ();
 sg13g2_fill_1 FILLER_17_2432 ();
 sg13g2_fill_1 FILLER_17_2468 ();
 sg13g2_decap_4 FILLER_17_2496 ();
 sg13g2_fill_2 FILLER_17_2504 ();
 sg13g2_fill_1 FILLER_17_2506 ();
 sg13g2_decap_8 FILLER_17_2565 ();
 sg13g2_decap_4 FILLER_17_2572 ();
 sg13g2_fill_1 FILLER_17_2576 ();
 sg13g2_fill_1 FILLER_17_2581 ();
 sg13g2_decap_8 FILLER_17_2650 ();
 sg13g2_decap_8 FILLER_17_2657 ();
 sg13g2_decap_4 FILLER_17_2664 ();
 sg13g2_fill_2 FILLER_17_2668 ();
 sg13g2_decap_8 FILLER_17_2683 ();
 sg13g2_decap_8 FILLER_17_2690 ();
 sg13g2_decap_8 FILLER_17_2697 ();
 sg13g2_fill_1 FILLER_17_2740 ();
 sg13g2_decap_8 FILLER_17_2746 ();
 sg13g2_decap_8 FILLER_17_2753 ();
 sg13g2_fill_2 FILLER_17_2760 ();
 sg13g2_fill_1 FILLER_17_2762 ();
 sg13g2_fill_1 FILLER_17_2767 ();
 sg13g2_decap_4 FILLER_17_2797 ();
 sg13g2_fill_1 FILLER_17_2811 ();
 sg13g2_fill_2 FILLER_17_2816 ();
 sg13g2_fill_1 FILLER_17_2818 ();
 sg13g2_decap_8 FILLER_17_2828 ();
 sg13g2_decap_8 FILLER_17_2835 ();
 sg13g2_decap_8 FILLER_17_2842 ();
 sg13g2_decap_8 FILLER_17_2849 ();
 sg13g2_decap_8 FILLER_17_2856 ();
 sg13g2_fill_2 FILLER_17_2873 ();
 sg13g2_fill_1 FILLER_17_2875 ();
 sg13g2_decap_4 FILLER_17_2894 ();
 sg13g2_fill_2 FILLER_17_2903 ();
 sg13g2_fill_1 FILLER_17_2905 ();
 sg13g2_decap_8 FILLER_17_2910 ();
 sg13g2_decap_8 FILLER_17_2917 ();
 sg13g2_decap_8 FILLER_17_2924 ();
 sg13g2_fill_2 FILLER_17_2931 ();
 sg13g2_fill_1 FILLER_17_2933 ();
 sg13g2_decap_8 FILLER_17_2989 ();
 sg13g2_decap_8 FILLER_17_2996 ();
 sg13g2_decap_8 FILLER_17_3003 ();
 sg13g2_decap_4 FILLER_17_3010 ();
 sg13g2_fill_1 FILLER_17_3014 ();
 sg13g2_decap_4 FILLER_17_3056 ();
 sg13g2_decap_8 FILLER_17_3149 ();
 sg13g2_decap_8 FILLER_17_3156 ();
 sg13g2_decap_4 FILLER_17_3163 ();
 sg13g2_fill_2 FILLER_17_3167 ();
 sg13g2_decap_8 FILLER_17_3192 ();
 sg13g2_decap_8 FILLER_17_3212 ();
 sg13g2_decap_8 FILLER_17_3219 ();
 sg13g2_decap_8 FILLER_17_3226 ();
 sg13g2_decap_8 FILLER_17_3233 ();
 sg13g2_fill_2 FILLER_17_3318 ();
 sg13g2_decap_8 FILLER_17_3379 ();
 sg13g2_fill_2 FILLER_17_3386 ();
 sg13g2_fill_1 FILLER_17_3388 ();
 sg13g2_decap_4 FILLER_17_3433 ();
 sg13g2_fill_2 FILLER_17_3437 ();
 sg13g2_decap_4 FILLER_17_3449 ();
 sg13g2_fill_1 FILLER_17_3453 ();
 sg13g2_decap_8 FILLER_17_3481 ();
 sg13g2_fill_2 FILLER_17_3488 ();
 sg13g2_fill_1 FILLER_17_3490 ();
 sg13g2_decap_8 FILLER_17_3500 ();
 sg13g2_fill_2 FILLER_17_3507 ();
 sg13g2_decap_4 FILLER_17_3522 ();
 sg13g2_decap_8 FILLER_17_3556 ();
 sg13g2_decap_8 FILLER_17_3563 ();
 sg13g2_decap_8 FILLER_17_3570 ();
 sg13g2_fill_1 FILLER_17_3577 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_65 ();
 sg13g2_decap_8 FILLER_18_72 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_125 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_4 FILLER_18_189 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_272 ();
 sg13g2_decap_4 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_300 ();
 sg13g2_fill_1 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_4 FILLER_18_353 ();
 sg13g2_decap_4 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_429 ();
 sg13g2_decap_4 FILLER_18_436 ();
 sg13g2_fill_1 FILLER_18_440 ();
 sg13g2_decap_4 FILLER_18_454 ();
 sg13g2_fill_1 FILLER_18_458 ();
 sg13g2_decap_4 FILLER_18_472 ();
 sg13g2_fill_2 FILLER_18_476 ();
 sg13g2_fill_2 FILLER_18_506 ();
 sg13g2_decap_4 FILLER_18_514 ();
 sg13g2_fill_2 FILLER_18_551 ();
 sg13g2_fill_2 FILLER_18_615 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_fill_2 FILLER_18_675 ();
 sg13g2_fill_1 FILLER_18_677 ();
 sg13g2_decap_8 FILLER_18_682 ();
 sg13g2_fill_1 FILLER_18_699 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_fill_2 FILLER_18_783 ();
 sg13g2_fill_2 FILLER_18_821 ();
 sg13g2_fill_1 FILLER_18_823 ();
 sg13g2_fill_2 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_873 ();
 sg13g2_fill_1 FILLER_18_880 ();
 sg13g2_decap_4 FILLER_18_885 ();
 sg13g2_fill_1 FILLER_18_889 ();
 sg13g2_fill_1 FILLER_18_899 ();
 sg13g2_fill_1 FILLER_18_913 ();
 sg13g2_fill_2 FILLER_18_921 ();
 sg13g2_fill_2 FILLER_18_929 ();
 sg13g2_decap_8 FILLER_18_944 ();
 sg13g2_fill_1 FILLER_18_951 ();
 sg13g2_decap_4 FILLER_18_999 ();
 sg13g2_fill_2 FILLER_18_1003 ();
 sg13g2_fill_1 FILLER_18_1009 ();
 sg13g2_decap_8 FILLER_18_1032 ();
 sg13g2_decap_8 FILLER_18_1039 ();
 sg13g2_decap_4 FILLER_18_1046 ();
 sg13g2_fill_1 FILLER_18_1050 ();
 sg13g2_decap_4 FILLER_18_1087 ();
 sg13g2_fill_1 FILLER_18_1109 ();
 sg13g2_decap_8 FILLER_18_1161 ();
 sg13g2_decap_4 FILLER_18_1168 ();
 sg13g2_fill_1 FILLER_18_1172 ();
 sg13g2_fill_1 FILLER_18_1212 ();
 sg13g2_fill_1 FILLER_18_1231 ();
 sg13g2_fill_2 FILLER_18_1242 ();
 sg13g2_fill_1 FILLER_18_1244 ();
 sg13g2_decap_8 FILLER_18_1258 ();
 sg13g2_decap_8 FILLER_18_1265 ();
 sg13g2_decap_8 FILLER_18_1272 ();
 sg13g2_decap_4 FILLER_18_1279 ();
 sg13g2_fill_1 FILLER_18_1283 ();
 sg13g2_fill_1 FILLER_18_1289 ();
 sg13g2_fill_2 FILLER_18_1304 ();
 sg13g2_decap_4 FILLER_18_1319 ();
 sg13g2_fill_2 FILLER_18_1323 ();
 sg13g2_fill_2 FILLER_18_1334 ();
 sg13g2_fill_1 FILLER_18_1336 ();
 sg13g2_decap_8 FILLER_18_1365 ();
 sg13g2_decap_8 FILLER_18_1372 ();
 sg13g2_decap_8 FILLER_18_1379 ();
 sg13g2_decap_4 FILLER_18_1386 ();
 sg13g2_fill_2 FILLER_18_1390 ();
 sg13g2_decap_8 FILLER_18_1437 ();
 sg13g2_decap_8 FILLER_18_1444 ();
 sg13g2_decap_4 FILLER_18_1451 ();
 sg13g2_fill_2 FILLER_18_1455 ();
 sg13g2_decap_8 FILLER_18_1485 ();
 sg13g2_fill_1 FILLER_18_1492 ();
 sg13g2_fill_2 FILLER_18_1498 ();
 sg13g2_fill_1 FILLER_18_1500 ();
 sg13g2_fill_2 FILLER_18_1506 ();
 sg13g2_decap_8 FILLER_18_1540 ();
 sg13g2_decap_8 FILLER_18_1547 ();
 sg13g2_decap_8 FILLER_18_1554 ();
 sg13g2_decap_8 FILLER_18_1561 ();
 sg13g2_decap_8 FILLER_18_1568 ();
 sg13g2_decap_8 FILLER_18_1575 ();
 sg13g2_decap_4 FILLER_18_1582 ();
 sg13g2_fill_2 FILLER_18_1609 ();
 sg13g2_decap_8 FILLER_18_1628 ();
 sg13g2_decap_8 FILLER_18_1635 ();
 sg13g2_decap_8 FILLER_18_1642 ();
 sg13g2_decap_4 FILLER_18_1649 ();
 sg13g2_fill_2 FILLER_18_1653 ();
 sg13g2_fill_2 FILLER_18_1663 ();
 sg13g2_fill_1 FILLER_18_1673 ();
 sg13g2_fill_1 FILLER_18_1683 ();
 sg13g2_decap_8 FILLER_18_1689 ();
 sg13g2_decap_8 FILLER_18_1696 ();
 sg13g2_decap_4 FILLER_18_1703 ();
 sg13g2_decap_8 FILLER_18_1720 ();
 sg13g2_decap_4 FILLER_18_1727 ();
 sg13g2_fill_1 FILLER_18_1731 ();
 sg13g2_fill_1 FILLER_18_1741 ();
 sg13g2_decap_4 FILLER_18_1754 ();
 sg13g2_fill_2 FILLER_18_1758 ();
 sg13g2_decap_4 FILLER_18_1765 ();
 sg13g2_decap_8 FILLER_18_1782 ();
 sg13g2_decap_4 FILLER_18_1789 ();
 sg13g2_fill_1 FILLER_18_1804 ();
 sg13g2_fill_2 FILLER_18_1813 ();
 sg13g2_fill_1 FILLER_18_1815 ();
 sg13g2_decap_8 FILLER_18_1822 ();
 sg13g2_fill_2 FILLER_18_1829 ();
 sg13g2_fill_1 FILLER_18_1846 ();
 sg13g2_fill_2 FILLER_18_1856 ();
 sg13g2_fill_1 FILLER_18_1858 ();
 sg13g2_fill_2 FILLER_18_1868 ();
 sg13g2_fill_1 FILLER_18_1870 ();
 sg13g2_decap_4 FILLER_18_1876 ();
 sg13g2_decap_8 FILLER_18_1908 ();
 sg13g2_decap_8 FILLER_18_1915 ();
 sg13g2_fill_1 FILLER_18_1922 ();
 sg13g2_fill_2 FILLER_18_1936 ();
 sg13g2_fill_1 FILLER_18_1938 ();
 sg13g2_fill_1 FILLER_18_1964 ();
 sg13g2_decap_8 FILLER_18_1991 ();
 sg13g2_decap_4 FILLER_18_1998 ();
 sg13g2_fill_2 FILLER_18_2002 ();
 sg13g2_fill_2 FILLER_18_2013 ();
 sg13g2_fill_1 FILLER_18_2015 ();
 sg13g2_fill_1 FILLER_18_2022 ();
 sg13g2_decap_8 FILLER_18_2069 ();
 sg13g2_decap_8 FILLER_18_2076 ();
 sg13g2_decap_8 FILLER_18_2083 ();
 sg13g2_decap_8 FILLER_18_2090 ();
 sg13g2_fill_2 FILLER_18_2097 ();
 sg13g2_fill_2 FILLER_18_2109 ();
 sg13g2_fill_1 FILLER_18_2111 ();
 sg13g2_decap_8 FILLER_18_2141 ();
 sg13g2_decap_4 FILLER_18_2148 ();
 sg13g2_decap_8 FILLER_18_2163 ();
 sg13g2_fill_1 FILLER_18_2196 ();
 sg13g2_fill_1 FILLER_18_2209 ();
 sg13g2_fill_2 FILLER_18_2246 ();
 sg13g2_fill_2 FILLER_18_2279 ();
 sg13g2_decap_8 FILLER_18_2308 ();
 sg13g2_decap_8 FILLER_18_2315 ();
 sg13g2_decap_8 FILLER_18_2322 ();
 sg13g2_decap_8 FILLER_18_2329 ();
 sg13g2_decap_4 FILLER_18_2336 ();
 sg13g2_fill_2 FILLER_18_2340 ();
 sg13g2_fill_2 FILLER_18_2355 ();
 sg13g2_fill_1 FILLER_18_2357 ();
 sg13g2_fill_2 FILLER_18_2362 ();
 sg13g2_fill_2 FILLER_18_2391 ();
 sg13g2_fill_1 FILLER_18_2393 ();
 sg13g2_fill_1 FILLER_18_2398 ();
 sg13g2_decap_8 FILLER_18_2426 ();
 sg13g2_decap_8 FILLER_18_2433 ();
 sg13g2_fill_2 FILLER_18_2440 ();
 sg13g2_fill_1 FILLER_18_2446 ();
 sg13g2_fill_2 FILLER_18_2474 ();
 sg13g2_fill_2 FILLER_18_2486 ();
 sg13g2_decap_8 FILLER_18_2497 ();
 sg13g2_decap_4 FILLER_18_2504 ();
 sg13g2_fill_1 FILLER_18_2508 ();
 sg13g2_fill_2 FILLER_18_2550 ();
 sg13g2_fill_1 FILLER_18_2552 ();
 sg13g2_decap_8 FILLER_18_2562 ();
 sg13g2_decap_8 FILLER_18_2569 ();
 sg13g2_decap_4 FILLER_18_2576 ();
 sg13g2_decap_4 FILLER_18_2607 ();
 sg13g2_fill_2 FILLER_18_2611 ();
 sg13g2_decap_4 FILLER_18_2649 ();
 sg13g2_decap_8 FILLER_18_2666 ();
 sg13g2_fill_2 FILLER_18_2673 ();
 sg13g2_fill_2 FILLER_18_2727 ();
 sg13g2_decap_8 FILLER_18_2750 ();
 sg13g2_decap_8 FILLER_18_2757 ();
 sg13g2_decap_8 FILLER_18_2764 ();
 sg13g2_decap_8 FILLER_18_2771 ();
 sg13g2_fill_2 FILLER_18_2778 ();
 sg13g2_fill_2 FILLER_18_2808 ();
 sg13g2_decap_8 FILLER_18_2823 ();
 sg13g2_decap_8 FILLER_18_2830 ();
 sg13g2_fill_2 FILLER_18_2837 ();
 sg13g2_fill_1 FILLER_18_2839 ();
 sg13g2_decap_4 FILLER_18_2872 ();
 sg13g2_decap_8 FILLER_18_2881 ();
 sg13g2_decap_8 FILLER_18_2888 ();
 sg13g2_decap_8 FILLER_18_2895 ();
 sg13g2_decap_4 FILLER_18_2902 ();
 sg13g2_fill_1 FILLER_18_2906 ();
 sg13g2_decap_8 FILLER_18_2934 ();
 sg13g2_decap_8 FILLER_18_2941 ();
 sg13g2_fill_2 FILLER_18_2948 ();
 sg13g2_decap_8 FILLER_18_3007 ();
 sg13g2_decap_8 FILLER_18_3014 ();
 sg13g2_fill_2 FILLER_18_3021 ();
 sg13g2_fill_1 FILLER_18_3023 ();
 sg13g2_fill_2 FILLER_18_3028 ();
 sg13g2_decap_8 FILLER_18_3049 ();
 sg13g2_decap_8 FILLER_18_3056 ();
 sg13g2_decap_8 FILLER_18_3063 ();
 sg13g2_decap_4 FILLER_18_3070 ();
 sg13g2_fill_2 FILLER_18_3078 ();
 sg13g2_decap_8 FILLER_18_3140 ();
 sg13g2_decap_8 FILLER_18_3147 ();
 sg13g2_decap_4 FILLER_18_3154 ();
 sg13g2_fill_2 FILLER_18_3158 ();
 sg13g2_fill_2 FILLER_18_3170 ();
 sg13g2_fill_1 FILLER_18_3172 ();
 sg13g2_decap_8 FILLER_18_3220 ();
 sg13g2_decap_8 FILLER_18_3227 ();
 sg13g2_decap_4 FILLER_18_3234 ();
 sg13g2_decap_8 FILLER_18_3255 ();
 sg13g2_fill_1 FILLER_18_3262 ();
 sg13g2_decap_4 FILLER_18_3311 ();
 sg13g2_decap_8 FILLER_18_3383 ();
 sg13g2_decap_8 FILLER_18_3390 ();
 sg13g2_decap_8 FILLER_18_3428 ();
 sg13g2_decap_4 FILLER_18_3435 ();
 sg13g2_fill_1 FILLER_18_3439 ();
 sg13g2_decap_8 FILLER_18_3467 ();
 sg13g2_fill_1 FILLER_18_3474 ();
 sg13g2_decap_8 FILLER_18_3502 ();
 sg13g2_decap_8 FILLER_18_3509 ();
 sg13g2_decap_8 FILLER_18_3516 ();
 sg13g2_fill_2 FILLER_18_3523 ();
 sg13g2_fill_1 FILLER_18_3525 ();
 sg13g2_decap_8 FILLER_18_3562 ();
 sg13g2_decap_8 FILLER_18_3569 ();
 sg13g2_fill_2 FILLER_18_3576 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_57 ();
 sg13g2_decap_8 FILLER_19_64 ();
 sg13g2_fill_2 FILLER_19_71 ();
 sg13g2_decap_8 FILLER_19_78 ();
 sg13g2_decap_4 FILLER_19_85 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_fill_2 FILLER_19_114 ();
 sg13g2_decap_8 FILLER_19_121 ();
 sg13g2_decap_8 FILLER_19_128 ();
 sg13g2_decap_8 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_142 ();
 sg13g2_decap_8 FILLER_19_149 ();
 sg13g2_decap_4 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_decap_4 FILLER_19_299 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_4 FILLER_19_363 ();
 sg13g2_decap_4 FILLER_19_375 ();
 sg13g2_decap_4 FILLER_19_413 ();
 sg13g2_fill_1 FILLER_19_417 ();
 sg13g2_fill_2 FILLER_19_431 ();
 sg13g2_fill_1 FILLER_19_433 ();
 sg13g2_decap_8 FILLER_19_443 ();
 sg13g2_decap_8 FILLER_19_450 ();
 sg13g2_decap_4 FILLER_19_457 ();
 sg13g2_fill_2 FILLER_19_474 ();
 sg13g2_fill_1 FILLER_19_476 ();
 sg13g2_decap_4 FILLER_19_486 ();
 sg13g2_fill_1 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_500 ();
 sg13g2_decap_8 FILLER_19_507 ();
 sg13g2_decap_8 FILLER_19_514 ();
 sg13g2_decap_4 FILLER_19_521 ();
 sg13g2_fill_1 FILLER_19_534 ();
 sg13g2_fill_2 FILLER_19_548 ();
 sg13g2_fill_2 FILLER_19_570 ();
 sg13g2_decap_4 FILLER_19_581 ();
 sg13g2_fill_1 FILLER_19_585 ();
 sg13g2_decap_8 FILLER_19_664 ();
 sg13g2_fill_1 FILLER_19_676 ();
 sg13g2_fill_2 FILLER_19_686 ();
 sg13g2_fill_1 FILLER_19_688 ();
 sg13g2_fill_2 FILLER_19_699 ();
 sg13g2_fill_1 FILLER_19_701 ();
 sg13g2_fill_2 FILLER_19_710 ();
 sg13g2_fill_1 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_fill_1 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_754 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_fill_2 FILLER_19_823 ();
 sg13g2_fill_1 FILLER_19_825 ();
 sg13g2_decap_8 FILLER_19_863 ();
 sg13g2_decap_8 FILLER_19_870 ();
 sg13g2_fill_2 FILLER_19_888 ();
 sg13g2_decap_4 FILLER_19_932 ();
 sg13g2_decap_8 FILLER_19_949 ();
 sg13g2_fill_1 FILLER_19_956 ();
 sg13g2_decap_4 FILLER_19_987 ();
 sg13g2_fill_1 FILLER_19_991 ();
 sg13g2_decap_8 FILLER_19_1036 ();
 sg13g2_decap_8 FILLER_19_1043 ();
 sg13g2_fill_2 FILLER_19_1050 ();
 sg13g2_fill_2 FILLER_19_1092 ();
 sg13g2_fill_2 FILLER_19_1112 ();
 sg13g2_fill_1 FILLER_19_1120 ();
 sg13g2_fill_2 FILLER_19_1137 ();
 sg13g2_fill_1 FILLER_19_1172 ();
 sg13g2_fill_2 FILLER_19_1178 ();
 sg13g2_fill_1 FILLER_19_1180 ();
 sg13g2_fill_2 FILLER_19_1194 ();
 sg13g2_fill_2 FILLER_19_1215 ();
 sg13g2_fill_1 FILLER_19_1230 ();
 sg13g2_decap_8 FILLER_19_1268 ();
 sg13g2_fill_2 FILLER_19_1275 ();
 sg13g2_fill_1 FILLER_19_1277 ();
 sg13g2_decap_4 FILLER_19_1335 ();
 sg13g2_decap_8 FILLER_19_1367 ();
 sg13g2_decap_8 FILLER_19_1374 ();
 sg13g2_decap_8 FILLER_19_1381 ();
 sg13g2_decap_8 FILLER_19_1388 ();
 sg13g2_decap_4 FILLER_19_1395 ();
 sg13g2_fill_2 FILLER_19_1425 ();
 sg13g2_fill_1 FILLER_19_1427 ();
 sg13g2_decap_8 FILLER_19_1446 ();
 sg13g2_decap_8 FILLER_19_1453 ();
 sg13g2_decap_4 FILLER_19_1460 ();
 sg13g2_fill_1 FILLER_19_1464 ();
 sg13g2_decap_8 FILLER_19_1468 ();
 sg13g2_fill_1 FILLER_19_1475 ();
 sg13g2_fill_1 FILLER_19_1494 ();
 sg13g2_fill_2 FILLER_19_1514 ();
 sg13g2_fill_1 FILLER_19_1516 ();
 sg13g2_fill_1 FILLER_19_1536 ();
 sg13g2_decap_8 FILLER_19_1550 ();
 sg13g2_decap_8 FILLER_19_1557 ();
 sg13g2_decap_4 FILLER_19_1564 ();
 sg13g2_decap_4 FILLER_19_1583 ();
 sg13g2_fill_2 FILLER_19_1587 ();
 sg13g2_fill_1 FILLER_19_1629 ();
 sg13g2_decap_4 FILLER_19_1639 ();
 sg13g2_fill_2 FILLER_19_1643 ();
 sg13g2_decap_8 FILLER_19_1658 ();
 sg13g2_fill_2 FILLER_19_1673 ();
 sg13g2_decap_8 FILLER_19_1680 ();
 sg13g2_fill_2 FILLER_19_1687 ();
 sg13g2_decap_8 FILLER_19_1702 ();
 sg13g2_fill_2 FILLER_19_1709 ();
 sg13g2_decap_8 FILLER_19_1715 ();
 sg13g2_fill_1 FILLER_19_1722 ();
 sg13g2_decap_4 FILLER_19_1732 ();
 sg13g2_fill_1 FILLER_19_1736 ();
 sg13g2_decap_8 FILLER_19_1742 ();
 sg13g2_decap_4 FILLER_19_1749 ();
 sg13g2_fill_1 FILLER_19_1753 ();
 sg13g2_decap_8 FILLER_19_1793 ();
 sg13g2_decap_8 FILLER_19_1800 ();
 sg13g2_fill_2 FILLER_19_1816 ();
 sg13g2_decap_4 FILLER_19_1841 ();
 sg13g2_fill_1 FILLER_19_1845 ();
 sg13g2_fill_2 FILLER_19_1856 ();
 sg13g2_fill_2 FILLER_19_1880 ();
 sg13g2_fill_1 FILLER_19_1882 ();
 sg13g2_fill_2 FILLER_19_1892 ();
 sg13g2_fill_1 FILLER_19_1894 ();
 sg13g2_decap_4 FILLER_19_1918 ();
 sg13g2_fill_1 FILLER_19_1922 ();
 sg13g2_decap_8 FILLER_19_1940 ();
 sg13g2_fill_1 FILLER_19_1947 ();
 sg13g2_decap_8 FILLER_19_1989 ();
 sg13g2_fill_1 FILLER_19_1996 ();
 sg13g2_fill_1 FILLER_19_2010 ();
 sg13g2_fill_1 FILLER_19_2017 ();
 sg13g2_fill_1 FILLER_19_2031 ();
 sg13g2_decap_8 FILLER_19_2060 ();
 sg13g2_decap_8 FILLER_19_2067 ();
 sg13g2_decap_4 FILLER_19_2074 ();
 sg13g2_fill_1 FILLER_19_2078 ();
 sg13g2_fill_2 FILLER_19_2107 ();
 sg13g2_fill_2 FILLER_19_2157 ();
 sg13g2_fill_1 FILLER_19_2159 ();
 sg13g2_decap_4 FILLER_19_2172 ();
 sg13g2_fill_2 FILLER_19_2176 ();
 sg13g2_decap_8 FILLER_19_2183 ();
 sg13g2_decap_8 FILLER_19_2190 ();
 sg13g2_decap_8 FILLER_19_2197 ();
 sg13g2_fill_1 FILLER_19_2204 ();
 sg13g2_fill_1 FILLER_19_2210 ();
 sg13g2_fill_1 FILLER_19_2224 ();
 sg13g2_decap_8 FILLER_19_2235 ();
 sg13g2_decap_4 FILLER_19_2242 ();
 sg13g2_fill_2 FILLER_19_2251 ();
 sg13g2_fill_1 FILLER_19_2253 ();
 sg13g2_fill_1 FILLER_19_2305 ();
 sg13g2_decap_4 FILLER_19_2333 ();
 sg13g2_fill_2 FILLER_19_2337 ();
 sg13g2_fill_2 FILLER_19_2408 ();
 sg13g2_decap_8 FILLER_19_2431 ();
 sg13g2_decap_8 FILLER_19_2438 ();
 sg13g2_fill_1 FILLER_19_2445 ();
 sg13g2_decap_8 FILLER_19_2488 ();
 sg13g2_decap_8 FILLER_19_2495 ();
 sg13g2_decap_8 FILLER_19_2502 ();
 sg13g2_decap_8 FILLER_19_2509 ();
 sg13g2_fill_1 FILLER_19_2516 ();
 sg13g2_fill_1 FILLER_19_2530 ();
 sg13g2_decap_4 FILLER_19_2540 ();
 sg13g2_fill_2 FILLER_19_2544 ();
 sg13g2_decap_8 FILLER_19_2550 ();
 sg13g2_decap_8 FILLER_19_2557 ();
 sg13g2_decap_4 FILLER_19_2564 ();
 sg13g2_fill_2 FILLER_19_2568 ();
 sg13g2_fill_2 FILLER_19_2622 ();
 sg13g2_decap_8 FILLER_19_2678 ();
 sg13g2_fill_2 FILLER_19_2685 ();
 sg13g2_decap_8 FILLER_19_2750 ();
 sg13g2_decap_8 FILLER_19_2757 ();
 sg13g2_decap_8 FILLER_19_2764 ();
 sg13g2_decap_4 FILLER_19_2771 ();
 sg13g2_fill_2 FILLER_19_2785 ();
 sg13g2_fill_1 FILLER_19_2787 ();
 sg13g2_decap_4 FILLER_19_2798 ();
 sg13g2_fill_1 FILLER_19_2802 ();
 sg13g2_decap_8 FILLER_19_2830 ();
 sg13g2_fill_2 FILLER_19_2837 ();
 sg13g2_fill_1 FILLER_19_2839 ();
 sg13g2_fill_1 FILLER_19_2880 ();
 sg13g2_decap_8 FILLER_19_2944 ();
 sg13g2_fill_1 FILLER_19_2951 ();
 sg13g2_decap_8 FILLER_19_2994 ();
 sg13g2_decap_8 FILLER_19_3001 ();
 sg13g2_decap_8 FILLER_19_3008 ();
 sg13g2_decap_8 FILLER_19_3015 ();
 sg13g2_decap_8 FILLER_19_3022 ();
 sg13g2_fill_2 FILLER_19_3029 ();
 sg13g2_fill_1 FILLER_19_3031 ();
 sg13g2_decap_8 FILLER_19_3064 ();
 sg13g2_decap_8 FILLER_19_3071 ();
 sg13g2_fill_2 FILLER_19_3078 ();
 sg13g2_decap_8 FILLER_19_3093 ();
 sg13g2_fill_1 FILLER_19_3100 ();
 sg13g2_fill_1 FILLER_19_3113 ();
 sg13g2_decap_4 FILLER_19_3124 ();
 sg13g2_fill_1 FILLER_19_3128 ();
 sg13g2_decap_8 FILLER_19_3138 ();
 sg13g2_decap_8 FILLER_19_3145 ();
 sg13g2_decap_4 FILLER_19_3152 ();
 sg13g2_fill_2 FILLER_19_3156 ();
 sg13g2_decap_8 FILLER_19_3225 ();
 sg13g2_decap_8 FILLER_19_3232 ();
 sg13g2_decap_8 FILLER_19_3239 ();
 sg13g2_decap_4 FILLER_19_3246 ();
 sg13g2_fill_1 FILLER_19_3250 ();
 sg13g2_fill_2 FILLER_19_3278 ();
 sg13g2_fill_1 FILLER_19_3280 ();
 sg13g2_decap_8 FILLER_19_3291 ();
 sg13g2_decap_8 FILLER_19_3298 ();
 sg13g2_decap_8 FILLER_19_3305 ();
 sg13g2_decap_8 FILLER_19_3312 ();
 sg13g2_fill_2 FILLER_19_3319 ();
 sg13g2_decap_8 FILLER_19_3329 ();
 sg13g2_fill_2 FILLER_19_3336 ();
 sg13g2_decap_8 FILLER_19_3381 ();
 sg13g2_decap_8 FILLER_19_3388 ();
 sg13g2_decap_8 FILLER_19_3395 ();
 sg13g2_decap_8 FILLER_19_3402 ();
 sg13g2_decap_8 FILLER_19_3409 ();
 sg13g2_decap_8 FILLER_19_3416 ();
 sg13g2_decap_8 FILLER_19_3423 ();
 sg13g2_decap_8 FILLER_19_3430 ();
 sg13g2_decap_8 FILLER_19_3437 ();
 sg13g2_decap_8 FILLER_19_3506 ();
 sg13g2_decap_8 FILLER_19_3513 ();
 sg13g2_fill_1 FILLER_19_3520 ();
 sg13g2_decap_8 FILLER_19_3571 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_18 ();
 sg13g2_fill_2 FILLER_20_34 ();
 sg13g2_decap_8 FILLER_20_45 ();
 sg13g2_fill_2 FILLER_20_52 ();
 sg13g2_fill_1 FILLER_20_54 ();
 sg13g2_fill_2 FILLER_20_95 ();
 sg13g2_fill_1 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_decap_8 FILLER_20_122 ();
 sg13g2_decap_4 FILLER_20_129 ();
 sg13g2_decap_8 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_decap_8 FILLER_20_187 ();
 sg13g2_fill_2 FILLER_20_194 ();
 sg13g2_fill_1 FILLER_20_196 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_286 ();
 sg13g2_decap_4 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_297 ();
 sg13g2_decap_4 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_decap_4 FILLER_20_340 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_4 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_379 ();
 sg13g2_fill_2 FILLER_20_386 ();
 sg13g2_fill_1 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_decap_8 FILLER_20_407 ();
 sg13g2_fill_2 FILLER_20_414 ();
 sg13g2_fill_1 FILLER_20_416 ();
 sg13g2_decap_4 FILLER_20_445 ();
 sg13g2_decap_8 FILLER_20_477 ();
 sg13g2_decap_8 FILLER_20_484 ();
 sg13g2_decap_8 FILLER_20_491 ();
 sg13g2_fill_2 FILLER_20_498 ();
 sg13g2_fill_1 FILLER_20_500 ();
 sg13g2_fill_1 FILLER_20_542 ();
 sg13g2_decap_4 FILLER_20_552 ();
 sg13g2_fill_1 FILLER_20_556 ();
 sg13g2_decap_4 FILLER_20_609 ();
 sg13g2_fill_2 FILLER_20_613 ();
 sg13g2_decap_4 FILLER_20_620 ();
 sg13g2_fill_1 FILLER_20_624 ();
 sg13g2_fill_2 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_695 ();
 sg13g2_decap_8 FILLER_20_702 ();
 sg13g2_decap_8 FILLER_20_709 ();
 sg13g2_fill_2 FILLER_20_716 ();
 sg13g2_fill_1 FILLER_20_718 ();
 sg13g2_decap_8 FILLER_20_730 ();
 sg13g2_fill_1 FILLER_20_737 ();
 sg13g2_decap_4 FILLER_20_743 ();
 sg13g2_fill_1 FILLER_20_760 ();
 sg13g2_decap_4 FILLER_20_775 ();
 sg13g2_fill_1 FILLER_20_779 ();
 sg13g2_decap_8 FILLER_20_799 ();
 sg13g2_decap_8 FILLER_20_806 ();
 sg13g2_decap_8 FILLER_20_813 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_8 FILLER_20_841 ();
 sg13g2_fill_2 FILLER_20_848 ();
 sg13g2_fill_2 FILLER_20_856 ();
 sg13g2_fill_2 FILLER_20_863 ();
 sg13g2_fill_1 FILLER_20_865 ();
 sg13g2_fill_1 FILLER_20_891 ();
 sg13g2_fill_1 FILLER_20_901 ();
 sg13g2_decap_4 FILLER_20_923 ();
 sg13g2_decap_4 FILLER_20_945 ();
 sg13g2_decap_8 FILLER_20_953 ();
 sg13g2_decap_4 FILLER_20_960 ();
 sg13g2_fill_1 FILLER_20_964 ();
 sg13g2_decap_8 FILLER_20_981 ();
 sg13g2_decap_8 FILLER_20_988 ();
 sg13g2_decap_8 FILLER_20_995 ();
 sg13g2_decap_8 FILLER_20_1002 ();
 sg13g2_decap_4 FILLER_20_1009 ();
 sg13g2_decap_8 FILLER_20_1041 ();
 sg13g2_decap_4 FILLER_20_1048 ();
 sg13g2_fill_1 FILLER_20_1052 ();
 sg13g2_fill_2 FILLER_20_1078 ();
 sg13g2_fill_1 FILLER_20_1086 ();
 sg13g2_decap_4 FILLER_20_1101 ();
 sg13g2_decap_8 FILLER_20_1110 ();
 sg13g2_fill_1 FILLER_20_1117 ();
 sg13g2_fill_2 FILLER_20_1180 ();
 sg13g2_fill_1 FILLER_20_1182 ();
 sg13g2_decap_8 FILLER_20_1192 ();
 sg13g2_fill_2 FILLER_20_1214 ();
 sg13g2_fill_2 FILLER_20_1312 ();
 sg13g2_decap_8 FILLER_20_1342 ();
 sg13g2_decap_8 FILLER_20_1349 ();
 sg13g2_decap_8 FILLER_20_1356 ();
 sg13g2_decap_8 FILLER_20_1363 ();
 sg13g2_fill_1 FILLER_20_1436 ();
 sg13g2_decap_8 FILLER_20_1446 ();
 sg13g2_decap_8 FILLER_20_1453 ();
 sg13g2_decap_8 FILLER_20_1460 ();
 sg13g2_decap_8 FILLER_20_1467 ();
 sg13g2_fill_2 FILLER_20_1474 ();
 sg13g2_fill_2 FILLER_20_1493 ();
 sg13g2_fill_2 FILLER_20_1504 ();
 sg13g2_fill_1 FILLER_20_1506 ();
 sg13g2_fill_2 FILLER_20_1544 ();
 sg13g2_fill_1 FILLER_20_1546 ();
 sg13g2_fill_2 FILLER_20_1555 ();
 sg13g2_fill_1 FILLER_20_1557 ();
 sg13g2_fill_2 FILLER_20_1586 ();
 sg13g2_fill_2 FILLER_20_1592 ();
 sg13g2_fill_2 FILLER_20_1607 ();
 sg13g2_fill_1 FILLER_20_1627 ();
 sg13g2_decap_8 FILLER_20_1634 ();
 sg13g2_decap_8 FILLER_20_1641 ();
 sg13g2_decap_8 FILLER_20_1648 ();
 sg13g2_decap_8 FILLER_20_1655 ();
 sg13g2_fill_2 FILLER_20_1662 ();
 sg13g2_fill_1 FILLER_20_1664 ();
 sg13g2_fill_2 FILLER_20_1675 ();
 sg13g2_fill_1 FILLER_20_1677 ();
 sg13g2_decap_4 FILLER_20_1683 ();
 sg13g2_fill_2 FILLER_20_1687 ();
 sg13g2_decap_8 FILLER_20_1702 ();
 sg13g2_decap_4 FILLER_20_1709 ();
 sg13g2_fill_2 FILLER_20_1718 ();
 sg13g2_fill_1 FILLER_20_1720 ();
 sg13g2_decap_8 FILLER_20_1726 ();
 sg13g2_decap_8 FILLER_20_1737 ();
 sg13g2_decap_4 FILLER_20_1744 ();
 sg13g2_decap_8 FILLER_20_1774 ();
 sg13g2_fill_2 FILLER_20_1794 ();
 sg13g2_fill_1 FILLER_20_1796 ();
 sg13g2_decap_8 FILLER_20_1810 ();
 sg13g2_decap_8 FILLER_20_1817 ();
 sg13g2_decap_8 FILLER_20_1824 ();
 sg13g2_fill_2 FILLER_20_1831 ();
 sg13g2_fill_1 FILLER_20_1833 ();
 sg13g2_fill_2 FILLER_20_1857 ();
 sg13g2_fill_1 FILLER_20_1859 ();
 sg13g2_decap_4 FILLER_20_1864 ();
 sg13g2_fill_2 FILLER_20_1881 ();
 sg13g2_fill_1 FILLER_20_1883 ();
 sg13g2_fill_1 FILLER_20_1889 ();
 sg13g2_fill_2 FILLER_20_1895 ();
 sg13g2_fill_1 FILLER_20_1897 ();
 sg13g2_decap_8 FILLER_20_1907 ();
 sg13g2_decap_8 FILLER_20_1914 ();
 sg13g2_decap_8 FILLER_20_1921 ();
 sg13g2_decap_8 FILLER_20_1928 ();
 sg13g2_decap_4 FILLER_20_1935 ();
 sg13g2_fill_2 FILLER_20_1939 ();
 sg13g2_fill_2 FILLER_20_1946 ();
 sg13g2_fill_1 FILLER_20_1948 ();
 sg13g2_fill_2 FILLER_20_1961 ();
 sg13g2_fill_1 FILLER_20_1963 ();
 sg13g2_decap_4 FILLER_20_1973 ();
 sg13g2_fill_1 FILLER_20_1977 ();
 sg13g2_decap_8 FILLER_20_1988 ();
 sg13g2_decap_4 FILLER_20_1995 ();
 sg13g2_fill_2 FILLER_20_1999 ();
 sg13g2_fill_2 FILLER_20_2006 ();
 sg13g2_fill_1 FILLER_20_2008 ();
 sg13g2_fill_2 FILLER_20_2019 ();
 sg13g2_fill_1 FILLER_20_2021 ();
 sg13g2_fill_1 FILLER_20_2040 ();
 sg13g2_decap_8 FILLER_20_2067 ();
 sg13g2_fill_2 FILLER_20_2074 ();
 sg13g2_fill_1 FILLER_20_2076 ();
 sg13g2_fill_2 FILLER_20_2090 ();
 sg13g2_fill_1 FILLER_20_2092 ();
 sg13g2_decap_4 FILLER_20_2103 ();
 sg13g2_decap_8 FILLER_20_2115 ();
 sg13g2_fill_2 FILLER_20_2122 ();
 sg13g2_fill_2 FILLER_20_2187 ();
 sg13g2_fill_1 FILLER_20_2189 ();
 sg13g2_decap_8 FILLER_20_2195 ();
 sg13g2_fill_2 FILLER_20_2202 ();
 sg13g2_fill_2 FILLER_20_2246 ();
 sg13g2_fill_2 FILLER_20_2271 ();
 sg13g2_fill_1 FILLER_20_2273 ();
 sg13g2_fill_2 FILLER_20_2287 ();
 sg13g2_decap_4 FILLER_20_2316 ();
 sg13g2_decap_8 FILLER_20_2325 ();
 sg13g2_decap_8 FILLER_20_2332 ();
 sg13g2_decap_8 FILLER_20_2339 ();
 sg13g2_decap_8 FILLER_20_2346 ();
 sg13g2_decap_4 FILLER_20_2353 ();
 sg13g2_fill_2 FILLER_20_2357 ();
 sg13g2_decap_4 FILLER_20_2363 ();
 sg13g2_fill_2 FILLER_20_2367 ();
 sg13g2_fill_2 FILLER_20_2373 ();
 sg13g2_decap_4 FILLER_20_2394 ();
 sg13g2_fill_2 FILLER_20_2412 ();
 sg13g2_decap_8 FILLER_20_2423 ();
 sg13g2_decap_8 FILLER_20_2493 ();
 sg13g2_decap_8 FILLER_20_2500 ();
 sg13g2_fill_2 FILLER_20_2507 ();
 sg13g2_fill_1 FILLER_20_2509 ();
 sg13g2_fill_2 FILLER_20_2520 ();
 sg13g2_fill_1 FILLER_20_2522 ();
 sg13g2_decap_8 FILLER_20_2559 ();
 sg13g2_decap_8 FILLER_20_2566 ();
 sg13g2_fill_1 FILLER_20_2573 ();
 sg13g2_decap_8 FILLER_20_2616 ();
 sg13g2_fill_2 FILLER_20_2623 ();
 sg13g2_fill_2 FILLER_20_2643 ();
 sg13g2_decap_4 FILLER_20_2659 ();
 sg13g2_decap_8 FILLER_20_2672 ();
 sg13g2_decap_8 FILLER_20_2679 ();
 sg13g2_decap_4 FILLER_20_2686 ();
 sg13g2_fill_1 FILLER_20_2690 ();
 sg13g2_fill_2 FILLER_20_2720 ();
 sg13g2_decap_8 FILLER_20_2759 ();
 sg13g2_fill_2 FILLER_20_2766 ();
 sg13g2_fill_2 FILLER_20_2772 ();
 sg13g2_decap_8 FILLER_20_2828 ();
 sg13g2_fill_2 FILLER_20_2861 ();
 sg13g2_fill_1 FILLER_20_2863 ();
 sg13g2_fill_2 FILLER_20_2922 ();
 sg13g2_decap_8 FILLER_20_2937 ();
 sg13g2_decap_8 FILLER_20_2944 ();
 sg13g2_fill_2 FILLER_20_2951 ();
 sg13g2_decap_8 FILLER_20_2989 ();
 sg13g2_decap_8 FILLER_20_2996 ();
 sg13g2_decap_4 FILLER_20_3003 ();
 sg13g2_fill_2 FILLER_20_3007 ();
 sg13g2_decap_8 FILLER_20_3067 ();
 sg13g2_decap_8 FILLER_20_3074 ();
 sg13g2_decap_8 FILLER_20_3081 ();
 sg13g2_decap_8 FILLER_20_3088 ();
 sg13g2_decap_8 FILLER_20_3095 ();
 sg13g2_fill_2 FILLER_20_3102 ();
 sg13g2_fill_1 FILLER_20_3104 ();
 sg13g2_fill_2 FILLER_20_3115 ();
 sg13g2_decap_8 FILLER_20_3143 ();
 sg13g2_decap_8 FILLER_20_3150 ();
 sg13g2_decap_4 FILLER_20_3157 ();
 sg13g2_fill_2 FILLER_20_3161 ();
 sg13g2_decap_4 FILLER_20_3167 ();
 sg13g2_fill_2 FILLER_20_3171 ();
 sg13g2_decap_8 FILLER_20_3221 ();
 sg13g2_decap_8 FILLER_20_3228 ();
 sg13g2_decap_8 FILLER_20_3235 ();
 sg13g2_fill_2 FILLER_20_3242 ();
 sg13g2_fill_1 FILLER_20_3244 ();
 sg13g2_fill_1 FILLER_20_3262 ();
 sg13g2_decap_4 FILLER_20_3273 ();
 sg13g2_decap_8 FILLER_20_3286 ();
 sg13g2_decap_8 FILLER_20_3293 ();
 sg13g2_fill_1 FILLER_20_3300 ();
 sg13g2_decap_8 FILLER_20_3311 ();
 sg13g2_decap_8 FILLER_20_3318 ();
 sg13g2_fill_2 FILLER_20_3325 ();
 sg13g2_fill_1 FILLER_20_3327 ();
 sg13g2_decap_4 FILLER_20_3341 ();
 sg13g2_fill_1 FILLER_20_3345 ();
 sg13g2_decap_8 FILLER_20_3377 ();
 sg13g2_decap_8 FILLER_20_3384 ();
 sg13g2_decap_4 FILLER_20_3391 ();
 sg13g2_fill_2 FILLER_20_3395 ();
 sg13g2_decap_8 FILLER_20_3410 ();
 sg13g2_fill_1 FILLER_20_3417 ();
 sg13g2_decap_4 FILLER_20_3441 ();
 sg13g2_fill_1 FILLER_20_3445 ();
 sg13g2_decap_8 FILLER_20_3495 ();
 sg13g2_decap_8 FILLER_20_3502 ();
 sg13g2_fill_1 FILLER_20_3509 ();
 sg13g2_decap_4 FILLER_20_3574 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_39 ();
 sg13g2_decap_4 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_fill_2 FILLER_21_88 ();
 sg13g2_fill_1 FILLER_21_90 ();
 sg13g2_decap_8 FILLER_21_118 ();
 sg13g2_fill_2 FILLER_21_125 ();
 sg13g2_fill_1 FILLER_21_127 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_4 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_2 FILLER_21_240 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_282 ();
 sg13g2_decap_8 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_296 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_fill_2 FILLER_21_326 ();
 sg13g2_fill_2 FILLER_21_341 ();
 sg13g2_fill_1 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_fill_1 FILLER_21_396 ();
 sg13g2_fill_1 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_440 ();
 sg13g2_decap_4 FILLER_21_447 ();
 sg13g2_fill_1 FILLER_21_451 ();
 sg13g2_fill_2 FILLER_21_461 ();
 sg13g2_decap_4 FILLER_21_477 ();
 sg13g2_decap_8 FILLER_21_494 ();
 sg13g2_decap_8 FILLER_21_501 ();
 sg13g2_fill_2 FILLER_21_541 ();
 sg13g2_fill_1 FILLER_21_546 ();
 sg13g2_fill_2 FILLER_21_578 ();
 sg13g2_fill_2 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_fill_2 FILLER_21_630 ();
 sg13g2_fill_2 FILLER_21_635 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_fill_2 FILLER_21_686 ();
 sg13g2_fill_1 FILLER_21_688 ();
 sg13g2_fill_1 FILLER_21_710 ();
 sg13g2_fill_1 FILLER_21_752 ();
 sg13g2_fill_2 FILLER_21_766 ();
 sg13g2_fill_1 FILLER_21_768 ();
 sg13g2_decap_4 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_810 ();
 sg13g2_fill_2 FILLER_21_817 ();
 sg13g2_fill_2 FILLER_21_829 ();
 sg13g2_fill_1 FILLER_21_831 ();
 sg13g2_fill_1 FILLER_21_840 ();
 sg13g2_decap_4 FILLER_21_856 ();
 sg13g2_fill_1 FILLER_21_860 ();
 sg13g2_fill_2 FILLER_21_866 ();
 sg13g2_decap_8 FILLER_21_889 ();
 sg13g2_decap_8 FILLER_21_896 ();
 sg13g2_decap_8 FILLER_21_903 ();
 sg13g2_decap_8 FILLER_21_910 ();
 sg13g2_fill_2 FILLER_21_917 ();
 sg13g2_fill_1 FILLER_21_919 ();
 sg13g2_fill_2 FILLER_21_925 ();
 sg13g2_fill_1 FILLER_21_927 ();
 sg13g2_decap_4 FILLER_21_942 ();
 sg13g2_fill_1 FILLER_21_946 ();
 sg13g2_decap_8 FILLER_21_952 ();
 sg13g2_fill_2 FILLER_21_959 ();
 sg13g2_decap_8 FILLER_21_981 ();
 sg13g2_decap_8 FILLER_21_988 ();
 sg13g2_decap_8 FILLER_21_995 ();
 sg13g2_decap_8 FILLER_21_1002 ();
 sg13g2_decap_8 FILLER_21_1009 ();
 sg13g2_decap_4 FILLER_21_1016 ();
 sg13g2_fill_1 FILLER_21_1020 ();
 sg13g2_decap_8 FILLER_21_1045 ();
 sg13g2_fill_2 FILLER_21_1052 ();
 sg13g2_decap_4 FILLER_21_1074 ();
 sg13g2_fill_2 FILLER_21_1104 ();
 sg13g2_fill_1 FILLER_21_1106 ();
 sg13g2_decap_4 FILLER_21_1120 ();
 sg13g2_fill_2 FILLER_21_1124 ();
 sg13g2_fill_2 FILLER_21_1139 ();
 sg13g2_fill_2 FILLER_21_1169 ();
 sg13g2_decap_8 FILLER_21_1199 ();
 sg13g2_fill_2 FILLER_21_1260 ();
 sg13g2_fill_2 FILLER_21_1268 ();
 sg13g2_fill_1 FILLER_21_1284 ();
 sg13g2_decap_4 FILLER_21_1335 ();
 sg13g2_fill_1 FILLER_21_1339 ();
 sg13g2_decap_8 FILLER_21_1349 ();
 sg13g2_decap_8 FILLER_21_1356 ();
 sg13g2_decap_4 FILLER_21_1363 ();
 sg13g2_fill_2 FILLER_21_1386 ();
 sg13g2_fill_1 FILLER_21_1388 ();
 sg13g2_fill_1 FILLER_21_1403 ();
 sg13g2_decap_8 FILLER_21_1446 ();
 sg13g2_decap_8 FILLER_21_1453 ();
 sg13g2_fill_2 FILLER_21_1460 ();
 sg13g2_decap_8 FILLER_21_1506 ();
 sg13g2_decap_4 FILLER_21_1527 ();
 sg13g2_decap_8 FILLER_21_1545 ();
 sg13g2_fill_2 FILLER_21_1552 ();
 sg13g2_decap_4 FILLER_21_1595 ();
 sg13g2_fill_1 FILLER_21_1612 ();
 sg13g2_fill_2 FILLER_21_1649 ();
 sg13g2_decap_4 FILLER_21_1706 ();
 sg13g2_fill_1 FILLER_21_1710 ();
 sg13g2_decap_4 FILLER_21_1776 ();
 sg13g2_fill_1 FILLER_21_1780 ();
 sg13g2_decap_8 FILLER_21_1798 ();
 sg13g2_decap_8 FILLER_21_1805 ();
 sg13g2_decap_8 FILLER_21_1812 ();
 sg13g2_decap_8 FILLER_21_1819 ();
 sg13g2_fill_1 FILLER_21_1826 ();
 sg13g2_decap_8 FILLER_21_1863 ();
 sg13g2_decap_8 FILLER_21_1870 ();
 sg13g2_decap_8 FILLER_21_1924 ();
 sg13g2_fill_2 FILLER_21_1931 ();
 sg13g2_decap_8 FILLER_21_1982 ();
 sg13g2_decap_8 FILLER_21_1989 ();
 sg13g2_fill_1 FILLER_21_1996 ();
 sg13g2_fill_1 FILLER_21_2016 ();
 sg13g2_fill_1 FILLER_21_2030 ();
 sg13g2_fill_2 FILLER_21_2050 ();
 sg13g2_fill_1 FILLER_21_2052 ();
 sg13g2_decap_8 FILLER_21_2071 ();
 sg13g2_fill_2 FILLER_21_2112 ();
 sg13g2_fill_1 FILLER_21_2114 ();
 sg13g2_decap_8 FILLER_21_2126 ();
 sg13g2_fill_2 FILLER_21_2133 ();
 sg13g2_fill_2 FILLER_21_2157 ();
 sg13g2_fill_1 FILLER_21_2159 ();
 sg13g2_decap_8 FILLER_21_2165 ();
 sg13g2_decap_8 FILLER_21_2172 ();
 sg13g2_decap_4 FILLER_21_2179 ();
 sg13g2_fill_1 FILLER_21_2183 ();
 sg13g2_fill_1 FILLER_21_2245 ();
 sg13g2_decap_8 FILLER_21_2259 ();
 sg13g2_fill_2 FILLER_21_2266 ();
 sg13g2_fill_1 FILLER_21_2287 ();
 sg13g2_decap_8 FILLER_21_2339 ();
 sg13g2_decap_8 FILLER_21_2346 ();
 sg13g2_fill_1 FILLER_21_2353 ();
 sg13g2_decap_8 FILLER_21_2404 ();
 sg13g2_fill_2 FILLER_21_2411 ();
 sg13g2_fill_1 FILLER_21_2413 ();
 sg13g2_decap_8 FILLER_21_2423 ();
 sg13g2_fill_2 FILLER_21_2430 ();
 sg13g2_fill_1 FILLER_21_2459 ();
 sg13g2_decap_4 FILLER_21_2500 ();
 sg13g2_decap_8 FILLER_21_2562 ();
 sg13g2_decap_8 FILLER_21_2569 ();
 sg13g2_decap_8 FILLER_21_2576 ();
 sg13g2_decap_8 FILLER_21_2583 ();
 sg13g2_decap_8 FILLER_21_2590 ();
 sg13g2_fill_1 FILLER_21_2597 ();
 sg13g2_fill_2 FILLER_21_2607 ();
 sg13g2_fill_1 FILLER_21_2609 ();
 sg13g2_decap_8 FILLER_21_2637 ();
 sg13g2_decap_8 FILLER_21_2644 ();
 sg13g2_decap_8 FILLER_21_2651 ();
 sg13g2_decap_8 FILLER_21_2658 ();
 sg13g2_fill_2 FILLER_21_2665 ();
 sg13g2_decap_8 FILLER_21_2694 ();
 sg13g2_decap_8 FILLER_21_2701 ();
 sg13g2_decap_4 FILLER_21_2708 ();
 sg13g2_fill_2 FILLER_21_2712 ();
 sg13g2_fill_2 FILLER_21_2718 ();
 sg13g2_fill_1 FILLER_21_2720 ();
 sg13g2_fill_2 FILLER_21_2731 ();
 sg13g2_fill_1 FILLER_21_2733 ();
 sg13g2_decap_8 FILLER_21_2756 ();
 sg13g2_decap_8 FILLER_21_2828 ();
 sg13g2_decap_8 FILLER_21_2835 ();
 sg13g2_fill_2 FILLER_21_2842 ();
 sg13g2_fill_1 FILLER_21_2844 ();
 sg13g2_fill_2 FILLER_21_2849 ();
 sg13g2_fill_1 FILLER_21_2851 ();
 sg13g2_fill_2 FILLER_21_2893 ();
 sg13g2_fill_1 FILLER_21_2895 ();
 sg13g2_fill_2 FILLER_21_2915 ();
 sg13g2_decap_8 FILLER_21_2994 ();
 sg13g2_decap_4 FILLER_21_3001 ();
 sg13g2_fill_2 FILLER_21_3005 ();
 sg13g2_fill_1 FILLER_21_3044 ();
 sg13g2_decap_8 FILLER_21_3072 ();
 sg13g2_decap_4 FILLER_21_3079 ();
 sg13g2_decap_8 FILLER_21_3147 ();
 sg13g2_decap_8 FILLER_21_3154 ();
 sg13g2_decap_4 FILLER_21_3161 ();
 sg13g2_fill_1 FILLER_21_3174 ();
 sg13g2_decap_8 FILLER_21_3188 ();
 sg13g2_decap_8 FILLER_21_3208 ();
 sg13g2_decap_8 FILLER_21_3215 ();
 sg13g2_decap_8 FILLER_21_3222 ();
 sg13g2_decap_8 FILLER_21_3229 ();
 sg13g2_fill_1 FILLER_21_3236 ();
 sg13g2_decap_8 FILLER_21_3287 ();
 sg13g2_decap_8 FILLER_21_3330 ();
 sg13g2_decap_8 FILLER_21_3337 ();
 sg13g2_fill_2 FILLER_21_3344 ();
 sg13g2_fill_2 FILLER_21_3356 ();
 sg13g2_fill_1 FILLER_21_3358 ();
 sg13g2_fill_1 FILLER_21_3378 ();
 sg13g2_decap_8 FILLER_21_3388 ();
 sg13g2_decap_4 FILLER_21_3395 ();
 sg13g2_decap_4 FILLER_21_3409 ();
 sg13g2_fill_2 FILLER_21_3413 ();
 sg13g2_fill_1 FILLER_21_3451 ();
 sg13g2_fill_1 FILLER_21_3465 ();
 sg13g2_fill_2 FILLER_21_3475 ();
 sg13g2_fill_1 FILLER_21_3477 ();
 sg13g2_decap_8 FILLER_21_3490 ();
 sg13g2_decap_8 FILLER_21_3497 ();
 sg13g2_decap_8 FILLER_21_3504 ();
 sg13g2_decap_8 FILLER_21_3511 ();
 sg13g2_decap_4 FILLER_21_3518 ();
 sg13g2_fill_2 FILLER_21_3522 ();
 sg13g2_decap_4 FILLER_21_3572 ();
 sg13g2_fill_2 FILLER_21_3576 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_11 ();
 sg13g2_fill_2 FILLER_22_40 ();
 sg13g2_fill_2 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_183 ();
 sg13g2_fill_2 FILLER_22_190 ();
 sg13g2_decap_4 FILLER_22_232 ();
 sg13g2_decap_8 FILLER_22_240 ();
 sg13g2_decap_4 FILLER_22_247 ();
 sg13g2_decap_4 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_304 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_4 FILLER_22_396 ();
 sg13g2_fill_2 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_461 ();
 sg13g2_fill_1 FILLER_22_463 ();
 sg13g2_fill_2 FILLER_22_492 ();
 sg13g2_fill_2 FILLER_22_511 ();
 sg13g2_decap_4 FILLER_22_543 ();
 sg13g2_decap_4 FILLER_22_569 ();
 sg13g2_decap_8 FILLER_22_603 ();
 sg13g2_decap_8 FILLER_22_610 ();
 sg13g2_fill_2 FILLER_22_617 ();
 sg13g2_fill_1 FILLER_22_619 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_fill_2 FILLER_22_694 ();
 sg13g2_fill_1 FILLER_22_705 ();
 sg13g2_decap_4 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_fill_2 FILLER_22_847 ();
 sg13g2_fill_1 FILLER_22_849 ();
 sg13g2_fill_2 FILLER_22_861 ();
 sg13g2_decap_4 FILLER_22_881 ();
 sg13g2_decap_8 FILLER_22_889 ();
 sg13g2_decap_8 FILLER_22_896 ();
 sg13g2_decap_8 FILLER_22_903 ();
 sg13g2_fill_1 FILLER_22_910 ();
 sg13g2_fill_1 FILLER_22_923 ();
 sg13g2_decap_8 FILLER_22_962 ();
 sg13g2_fill_2 FILLER_22_969 ();
 sg13g2_fill_1 FILLER_22_971 ();
 sg13g2_decap_8 FILLER_22_1017 ();
 sg13g2_decap_8 FILLER_22_1024 ();
 sg13g2_decap_8 FILLER_22_1031 ();
 sg13g2_fill_2 FILLER_22_1038 ();
 sg13g2_fill_1 FILLER_22_1040 ();
 sg13g2_decap_8 FILLER_22_1045 ();
 sg13g2_decap_4 FILLER_22_1052 ();
 sg13g2_fill_1 FILLER_22_1056 ();
 sg13g2_decap_4 FILLER_22_1108 ();
 sg13g2_fill_1 FILLER_22_1112 ();
 sg13g2_fill_2 FILLER_22_1160 ();
 sg13g2_fill_2 FILLER_22_1208 ();
 sg13g2_fill_1 FILLER_22_1210 ();
 sg13g2_decap_4 FILLER_22_1216 ();
 sg13g2_fill_1 FILLER_22_1236 ();
 sg13g2_fill_1 FILLER_22_1251 ();
 sg13g2_decap_4 FILLER_22_1263 ();
 sg13g2_decap_8 FILLER_22_1272 ();
 sg13g2_fill_2 FILLER_22_1279 ();
 sg13g2_fill_1 FILLER_22_1281 ();
 sg13g2_decap_4 FILLER_22_1345 ();
 sg13g2_decap_8 FILLER_22_1362 ();
 sg13g2_decap_4 FILLER_22_1369 ();
 sg13g2_fill_2 FILLER_22_1410 ();
 sg13g2_decap_8 FILLER_22_1445 ();
 sg13g2_decap_8 FILLER_22_1452 ();
 sg13g2_decap_8 FILLER_22_1459 ();
 sg13g2_fill_2 FILLER_22_1466 ();
 sg13g2_decap_8 FILLER_22_1495 ();
 sg13g2_decap_8 FILLER_22_1502 ();
 sg13g2_decap_4 FILLER_22_1509 ();
 sg13g2_fill_1 FILLER_22_1513 ();
 sg13g2_decap_8 FILLER_22_1550 ();
 sg13g2_decap_8 FILLER_22_1557 ();
 sg13g2_decap_4 FILLER_22_1591 ();
 sg13g2_fill_1 FILLER_22_1595 ();
 sg13g2_decap_4 FILLER_22_1609 ();
 sg13g2_decap_8 FILLER_22_1633 ();
 sg13g2_decap_4 FILLER_22_1649 ();
 sg13g2_fill_2 FILLER_22_1653 ();
 sg13g2_fill_1 FILLER_22_1692 ();
 sg13g2_decap_4 FILLER_22_1702 ();
 sg13g2_fill_1 FILLER_22_1719 ();
 sg13g2_fill_1 FILLER_22_1724 ();
 sg13g2_decap_8 FILLER_22_1730 ();
 sg13g2_decap_8 FILLER_22_1737 ();
 sg13g2_decap_8 FILLER_22_1744 ();
 sg13g2_decap_4 FILLER_22_1755 ();
 sg13g2_fill_2 FILLER_22_1768 ();
 sg13g2_fill_1 FILLER_22_1770 ();
 sg13g2_decap_8 FILLER_22_1812 ();
 sg13g2_decap_8 FILLER_22_1819 ();
 sg13g2_fill_2 FILLER_22_1826 ();
 sg13g2_decap_8 FILLER_22_1857 ();
 sg13g2_decap_8 FILLER_22_1864 ();
 sg13g2_decap_8 FILLER_22_1871 ();
 sg13g2_fill_2 FILLER_22_1878 ();
 sg13g2_fill_1 FILLER_22_1880 ();
 sg13g2_fill_2 FILLER_22_1919 ();
 sg13g2_fill_1 FILLER_22_1921 ();
 sg13g2_fill_2 FILLER_22_1932 ();
 sg13g2_decap_8 FILLER_22_1983 ();
 sg13g2_decap_4 FILLER_22_1990 ();
 sg13g2_decap_4 FILLER_22_2026 ();
 sg13g2_fill_2 FILLER_22_2030 ();
 sg13g2_fill_2 FILLER_22_2042 ();
 sg13g2_fill_1 FILLER_22_2082 ();
 sg13g2_fill_2 FILLER_22_2119 ();
 sg13g2_decap_4 FILLER_22_2135 ();
 sg13g2_decap_8 FILLER_22_2169 ();
 sg13g2_fill_2 FILLER_22_2176 ();
 sg13g2_fill_1 FILLER_22_2178 ();
 sg13g2_decap_8 FILLER_22_2183 ();
 sg13g2_decap_4 FILLER_22_2190 ();
 sg13g2_fill_2 FILLER_22_2194 ();
 sg13g2_decap_8 FILLER_22_2234 ();
 sg13g2_decap_8 FILLER_22_2241 ();
 sg13g2_decap_8 FILLER_22_2248 ();
 sg13g2_decap_8 FILLER_22_2255 ();
 sg13g2_fill_1 FILLER_22_2262 ();
 sg13g2_decap_8 FILLER_22_2267 ();
 sg13g2_fill_2 FILLER_22_2283 ();
 sg13g2_fill_1 FILLER_22_2285 ();
 sg13g2_decap_4 FILLER_22_2289 ();
 sg13g2_fill_1 FILLER_22_2293 ();
 sg13g2_fill_1 FILLER_22_2301 ();
 sg13g2_decap_8 FILLER_22_2347 ();
 sg13g2_decap_8 FILLER_22_2354 ();
 sg13g2_decap_8 FILLER_22_2361 ();
 sg13g2_fill_2 FILLER_22_2368 ();
 sg13g2_fill_1 FILLER_22_2370 ();
 sg13g2_decap_8 FILLER_22_2408 ();
 sg13g2_fill_2 FILLER_22_2424 ();
 sg13g2_fill_1 FILLER_22_2439 ();
 sg13g2_fill_2 FILLER_22_2505 ();
 sg13g2_fill_1 FILLER_22_2507 ();
 sg13g2_decap_8 FILLER_22_2575 ();
 sg13g2_decap_4 FILLER_22_2582 ();
 sg13g2_fill_1 FILLER_22_2586 ();
 sg13g2_decap_4 FILLER_22_2624 ();
 sg13g2_fill_1 FILLER_22_2628 ();
 sg13g2_decap_8 FILLER_22_2642 ();
 sg13g2_decap_8 FILLER_22_2649 ();
 sg13g2_decap_4 FILLER_22_2656 ();
 sg13g2_decap_8 FILLER_22_2700 ();
 sg13g2_fill_2 FILLER_22_2707 ();
 sg13g2_decap_8 FILLER_22_2736 ();
 sg13g2_decap_8 FILLER_22_2743 ();
 sg13g2_decap_8 FILLER_22_2750 ();
 sg13g2_fill_2 FILLER_22_2757 ();
 sg13g2_fill_2 FILLER_22_2779 ();
 sg13g2_fill_1 FILLER_22_2781 ();
 sg13g2_decap_8 FILLER_22_2791 ();
 sg13g2_fill_1 FILLER_22_2798 ();
 sg13g2_decap_4 FILLER_22_2812 ();
 sg13g2_fill_1 FILLER_22_2816 ();
 sg13g2_decap_8 FILLER_22_2830 ();
 sg13g2_decap_8 FILLER_22_2837 ();
 sg13g2_decap_4 FILLER_22_2844 ();
 sg13g2_decap_8 FILLER_22_2861 ();
 sg13g2_decap_4 FILLER_22_2868 ();
 sg13g2_fill_1 FILLER_22_2872 ();
 sg13g2_fill_2 FILLER_22_2896 ();
 sg13g2_fill_2 FILLER_22_2907 ();
 sg13g2_decap_8 FILLER_22_2917 ();
 sg13g2_decap_8 FILLER_22_2924 ();
 sg13g2_fill_2 FILLER_22_2935 ();
 sg13g2_fill_1 FILLER_22_2985 ();
 sg13g2_decap_8 FILLER_22_2999 ();
 sg13g2_decap_4 FILLER_22_3006 ();
 sg13g2_fill_2 FILLER_22_3010 ();
 sg13g2_fill_1 FILLER_22_3020 ();
 sg13g2_decap_8 FILLER_22_3065 ();
 sg13g2_fill_1 FILLER_22_3072 ();
 sg13g2_fill_1 FILLER_22_3119 ();
 sg13g2_decap_4 FILLER_22_3124 ();
 sg13g2_decap_8 FILLER_22_3137 ();
 sg13g2_decap_8 FILLER_22_3144 ();
 sg13g2_decap_8 FILLER_22_3151 ();
 sg13g2_decap_4 FILLER_22_3158 ();
 sg13g2_decap_8 FILLER_22_3189 ();
 sg13g2_decap_8 FILLER_22_3196 ();
 sg13g2_decap_8 FILLER_22_3203 ();
 sg13g2_decap_4 FILLER_22_3210 ();
 sg13g2_fill_2 FILLER_22_3214 ();
 sg13g2_fill_2 FILLER_22_3220 ();
 sg13g2_decap_8 FILLER_22_3270 ();
 sg13g2_decap_4 FILLER_22_3277 ();
 sg13g2_decap_8 FILLER_22_3329 ();
 sg13g2_fill_2 FILLER_22_3336 ();
 sg13g2_fill_1 FILLER_22_3396 ();
 sg13g2_decap_4 FILLER_22_3469 ();
 sg13g2_decap_8 FILLER_22_3513 ();
 sg13g2_decap_8 FILLER_22_3520 ();
 sg13g2_fill_2 FILLER_22_3547 ();
 sg13g2_fill_2 FILLER_22_3576 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_11 ();
 sg13g2_fill_1 FILLER_23_13 ();
 sg13g2_fill_2 FILLER_23_59 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_118 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_decap_8 FILLER_23_178 ();
 sg13g2_decap_8 FILLER_23_185 ();
 sg13g2_decap_8 FILLER_23_192 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_4 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_decap_8 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_307 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_2 FILLER_23_354 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_fill_2 FILLER_23_390 ();
 sg13g2_fill_2 FILLER_23_411 ();
 sg13g2_fill_1 FILLER_23_413 ();
 sg13g2_fill_2 FILLER_23_446 ();
 sg13g2_fill_1 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_458 ();
 sg13g2_fill_1 FILLER_23_465 ();
 sg13g2_decap_4 FILLER_23_503 ();
 sg13g2_fill_2 FILLER_23_507 ();
 sg13g2_decap_8 FILLER_23_514 ();
 sg13g2_decap_8 FILLER_23_521 ();
 sg13g2_fill_1 FILLER_23_528 ();
 sg13g2_fill_1 FILLER_23_547 ();
 sg13g2_decap_4 FILLER_23_608 ();
 sg13g2_fill_2 FILLER_23_653 ();
 sg13g2_fill_1 FILLER_23_655 ();
 sg13g2_fill_2 FILLER_23_669 ();
 sg13g2_decap_8 FILLER_23_680 ();
 sg13g2_decap_4 FILLER_23_687 ();
 sg13g2_fill_2 FILLER_23_691 ();
 sg13g2_decap_4 FILLER_23_701 ();
 sg13g2_fill_2 FILLER_23_705 ();
 sg13g2_fill_2 FILLER_23_743 ();
 sg13g2_decap_8 FILLER_23_803 ();
 sg13g2_decap_8 FILLER_23_857 ();
 sg13g2_decap_8 FILLER_23_872 ();
 sg13g2_fill_2 FILLER_23_879 ();
 sg13g2_fill_1 FILLER_23_881 ();
 sg13g2_decap_8 FILLER_23_891 ();
 sg13g2_fill_1 FILLER_23_911 ();
 sg13g2_fill_2 FILLER_23_923 ();
 sg13g2_decap_8 FILLER_23_1049 ();
 sg13g2_decap_8 FILLER_23_1056 ();
 sg13g2_decap_8 FILLER_23_1063 ();
 sg13g2_fill_2 FILLER_23_1070 ();
 sg13g2_decap_8 FILLER_23_1109 ();
 sg13g2_fill_2 FILLER_23_1170 ();
 sg13g2_fill_1 FILLER_23_1172 ();
 sg13g2_decap_8 FILLER_23_1256 ();
 sg13g2_decap_8 FILLER_23_1263 ();
 sg13g2_decap_8 FILLER_23_1270 ();
 sg13g2_fill_2 FILLER_23_1277 ();
 sg13g2_fill_1 FILLER_23_1279 ();
 sg13g2_decap_8 FILLER_23_1304 ();
 sg13g2_decap_4 FILLER_23_1328 ();
 sg13g2_fill_2 FILLER_23_1377 ();
 sg13g2_fill_1 FILLER_23_1379 ();
 sg13g2_fill_1 FILLER_23_1384 ();
 sg13g2_decap_4 FILLER_23_1393 ();
 sg13g2_fill_2 FILLER_23_1402 ();
 sg13g2_fill_2 FILLER_23_1438 ();
 sg13g2_decap_8 FILLER_23_1449 ();
 sg13g2_decap_8 FILLER_23_1456 ();
 sg13g2_fill_2 FILLER_23_1463 ();
 sg13g2_fill_1 FILLER_23_1465 ();
 sg13g2_fill_2 FILLER_23_1501 ();
 sg13g2_decap_8 FILLER_23_1506 ();
 sg13g2_fill_2 FILLER_23_1513 ();
 sg13g2_decap_8 FILLER_23_1543 ();
 sg13g2_decap_8 FILLER_23_1550 ();
 sg13g2_decap_8 FILLER_23_1557 ();
 sg13g2_decap_4 FILLER_23_1564 ();
 sg13g2_fill_2 FILLER_23_1568 ();
 sg13g2_fill_2 FILLER_23_1582 ();
 sg13g2_fill_1 FILLER_23_1588 ();
 sg13g2_decap_8 FILLER_23_1593 ();
 sg13g2_decap_8 FILLER_23_1600 ();
 sg13g2_decap_8 FILLER_23_1607 ();
 sg13g2_decap_8 FILLER_23_1614 ();
 sg13g2_fill_1 FILLER_23_1621 ();
 sg13g2_decap_4 FILLER_23_1631 ();
 sg13g2_fill_2 FILLER_23_1635 ();
 sg13g2_decap_8 FILLER_23_1642 ();
 sg13g2_fill_2 FILLER_23_1649 ();
 sg13g2_fill_1 FILLER_23_1651 ();
 sg13g2_fill_2 FILLER_23_1665 ();
 sg13g2_fill_1 FILLER_23_1667 ();
 sg13g2_decap_8 FILLER_23_1683 ();
 sg13g2_decap_4 FILLER_23_1690 ();
 sg13g2_fill_2 FILLER_23_1694 ();
 sg13g2_decap_4 FILLER_23_1701 ();
 sg13g2_fill_2 FILLER_23_1705 ();
 sg13g2_fill_2 FILLER_23_1725 ();
 sg13g2_fill_1 FILLER_23_1727 ();
 sg13g2_fill_1 FILLER_23_1735 ();
 sg13g2_decap_4 FILLER_23_1759 ();
 sg13g2_fill_1 FILLER_23_1763 ();
 sg13g2_fill_1 FILLER_23_1769 ();
 sg13g2_fill_1 FILLER_23_1793 ();
 sg13g2_decap_8 FILLER_23_1809 ();
 sg13g2_decap_8 FILLER_23_1816 ();
 sg13g2_decap_4 FILLER_23_1823 ();
 sg13g2_fill_1 FILLER_23_1827 ();
 sg13g2_fill_1 FILLER_23_1855 ();
 sg13g2_decap_4 FILLER_23_1864 ();
 sg13g2_fill_2 FILLER_23_1868 ();
 sg13g2_fill_1 FILLER_23_1875 ();
 sg13g2_fill_1 FILLER_23_1885 ();
 sg13g2_fill_2 FILLER_23_1918 ();
 sg13g2_fill_1 FILLER_23_1920 ();
 sg13g2_fill_1 FILLER_23_1964 ();
 sg13g2_fill_2 FILLER_23_1984 ();
 sg13g2_decap_8 FILLER_23_2025 ();
 sg13g2_decap_4 FILLER_23_2032 ();
 sg13g2_fill_1 FILLER_23_2050 ();
 sg13g2_fill_2 FILLER_23_2064 ();
 sg13g2_fill_1 FILLER_23_2066 ();
 sg13g2_fill_1 FILLER_23_2104 ();
 sg13g2_decap_8 FILLER_23_2137 ();
 sg13g2_decap_8 FILLER_23_2144 ();
 sg13g2_decap_4 FILLER_23_2156 ();
 sg13g2_decap_8 FILLER_23_2170 ();
 sg13g2_decap_8 FILLER_23_2177 ();
 sg13g2_decap_8 FILLER_23_2184 ();
 sg13g2_decap_8 FILLER_23_2191 ();
 sg13g2_decap_4 FILLER_23_2198 ();
 sg13g2_fill_1 FILLER_23_2202 ();
 sg13g2_decap_8 FILLER_23_2239 ();
 sg13g2_fill_1 FILLER_23_2251 ();
 sg13g2_fill_1 FILLER_23_2257 ();
 sg13g2_decap_4 FILLER_23_2286 ();
 sg13g2_fill_2 FILLER_23_2290 ();
 sg13g2_decap_8 FILLER_23_2352 ();
 sg13g2_decap_8 FILLER_23_2359 ();
 sg13g2_fill_2 FILLER_23_2366 ();
 sg13g2_fill_1 FILLER_23_2368 ();
 sg13g2_fill_1 FILLER_23_2396 ();
 sg13g2_decap_8 FILLER_23_2428 ();
 sg13g2_decap_4 FILLER_23_2435 ();
 sg13g2_fill_1 FILLER_23_2447 ();
 sg13g2_fill_2 FILLER_23_2452 ();
 sg13g2_fill_1 FILLER_23_2454 ();
 sg13g2_decap_8 FILLER_23_2490 ();
 sg13g2_decap_4 FILLER_23_2497 ();
 sg13g2_decap_4 FILLER_23_2514 ();
 sg13g2_fill_1 FILLER_23_2518 ();
 sg13g2_decap_8 FILLER_23_2569 ();
 sg13g2_fill_2 FILLER_23_2576 ();
 sg13g2_fill_1 FILLER_23_2625 ();
 sg13g2_fill_2 FILLER_23_2686 ();
 sg13g2_decap_8 FILLER_23_2728 ();
 sg13g2_decap_8 FILLER_23_2735 ();
 sg13g2_decap_8 FILLER_23_2742 ();
 sg13g2_decap_4 FILLER_23_2786 ();
 sg13g2_fill_2 FILLER_23_2790 ();
 sg13g2_decap_8 FILLER_23_2805 ();
 sg13g2_decap_8 FILLER_23_2812 ();
 sg13g2_fill_2 FILLER_23_2819 ();
 sg13g2_fill_1 FILLER_23_2821 ();
 sg13g2_fill_1 FILLER_23_2832 ();
 sg13g2_decap_8 FILLER_23_2855 ();
 sg13g2_decap_8 FILLER_23_2862 ();
 sg13g2_decap_4 FILLER_23_2869 ();
 sg13g2_fill_2 FILLER_23_2873 ();
 sg13g2_decap_8 FILLER_23_2911 ();
 sg13g2_decap_8 FILLER_23_2918 ();
 sg13g2_fill_2 FILLER_23_2934 ();
 sg13g2_decap_8 FILLER_23_2946 ();
 sg13g2_fill_1 FILLER_23_2953 ();
 sg13g2_decap_8 FILLER_23_2991 ();
 sg13g2_decap_8 FILLER_23_2998 ();
 sg13g2_decap_8 FILLER_23_3005 ();
 sg13g2_decap_8 FILLER_23_3012 ();
 sg13g2_decap_8 FILLER_23_3019 ();
 sg13g2_decap_4 FILLER_23_3026 ();
 sg13g2_fill_2 FILLER_23_3030 ();
 sg13g2_decap_4 FILLER_23_3041 ();
 sg13g2_decap_4 FILLER_23_3055 ();
 sg13g2_fill_2 FILLER_23_3059 ();
 sg13g2_fill_1 FILLER_23_3097 ();
 sg13g2_decap_4 FILLER_23_3128 ();
 sg13g2_fill_1 FILLER_23_3132 ();
 sg13g2_decap_4 FILLER_23_3143 ();
 sg13g2_decap_8 FILLER_23_3197 ();
 sg13g2_decap_8 FILLER_23_3204 ();
 sg13g2_fill_1 FILLER_23_3242 ();
 sg13g2_decap_8 FILLER_23_3270 ();
 sg13g2_fill_2 FILLER_23_3277 ();
 sg13g2_fill_2 FILLER_23_3293 ();
 sg13g2_fill_1 FILLER_23_3295 ();
 sg13g2_decap_4 FILLER_23_3327 ();
 sg13g2_fill_2 FILLER_23_3331 ();
 sg13g2_decap_8 FILLER_23_3360 ();
 sg13g2_decap_8 FILLER_23_3394 ();
 sg13g2_fill_1 FILLER_23_3401 ();
 sg13g2_decap_8 FILLER_23_3450 ();
 sg13g2_decap_8 FILLER_23_3457 ();
 sg13g2_decap_8 FILLER_23_3464 ();
 sg13g2_decap_8 FILLER_23_3471 ();
 sg13g2_decap_4 FILLER_23_3478 ();
 sg13g2_fill_1 FILLER_23_3482 ();
 sg13g2_decap_8 FILLER_23_3570 ();
 sg13g2_fill_1 FILLER_23_3577 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_52 ();
 sg13g2_fill_1 FILLER_24_54 ();
 sg13g2_fill_2 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_fill_2 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_fill_2 FILLER_24_141 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_decap_8 FILLER_24_185 ();
 sg13g2_decap_8 FILLER_24_192 ();
 sg13g2_decap_8 FILLER_24_199 ();
 sg13g2_fill_2 FILLER_24_206 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_232 ();
 sg13g2_decap_4 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_4 FILLER_24_359 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_fill_2 FILLER_24_369 ();
 sg13g2_fill_1 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_fill_2 FILLER_24_391 ();
 sg13g2_fill_2 FILLER_24_403 ();
 sg13g2_fill_1 FILLER_24_434 ();
 sg13g2_fill_1 FILLER_24_439 ();
 sg13g2_decap_8 FILLER_24_446 ();
 sg13g2_fill_2 FILLER_24_453 ();
 sg13g2_decap_8 FILLER_24_461 ();
 sg13g2_decap_8 FILLER_24_468 ();
 sg13g2_fill_2 FILLER_24_475 ();
 sg13g2_decap_8 FILLER_24_505 ();
 sg13g2_decap_8 FILLER_24_512 ();
 sg13g2_fill_2 FILLER_24_519 ();
 sg13g2_fill_1 FILLER_24_521 ();
 sg13g2_decap_8 FILLER_24_563 ();
 sg13g2_fill_2 FILLER_24_618 ();
 sg13g2_fill_2 FILLER_24_634 ();
 sg13g2_decap_8 FILLER_24_687 ();
 sg13g2_decap_8 FILLER_24_694 ();
 sg13g2_decap_8 FILLER_24_701 ();
 sg13g2_decap_4 FILLER_24_708 ();
 sg13g2_fill_2 FILLER_24_737 ();
 sg13g2_fill_1 FILLER_24_752 ();
 sg13g2_fill_2 FILLER_24_785 ();
 sg13g2_fill_1 FILLER_24_787 ();
 sg13g2_decap_8 FILLER_24_802 ();
 sg13g2_decap_4 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_857 ();
 sg13g2_fill_2 FILLER_24_864 ();
 sg13g2_fill_1 FILLER_24_866 ();
 sg13g2_decap_8 FILLER_24_876 ();
 sg13g2_decap_8 FILLER_24_883 ();
 sg13g2_decap_8 FILLER_24_890 ();
 sg13g2_decap_8 FILLER_24_897 ();
 sg13g2_decap_4 FILLER_24_904 ();
 sg13g2_fill_1 FILLER_24_908 ();
 sg13g2_fill_2 FILLER_24_924 ();
 sg13g2_fill_1 FILLER_24_935 ();
 sg13g2_decap_4 FILLER_24_949 ();
 sg13g2_fill_1 FILLER_24_953 ();
 sg13g2_decap_8 FILLER_24_963 ();
 sg13g2_fill_2 FILLER_24_970 ();
 sg13g2_fill_1 FILLER_24_972 ();
 sg13g2_fill_1 FILLER_24_978 ();
 sg13g2_decap_8 FILLER_24_997 ();
 sg13g2_decap_8 FILLER_24_1004 ();
 sg13g2_decap_8 FILLER_24_1011 ();
 sg13g2_fill_2 FILLER_24_1018 ();
 sg13g2_fill_1 FILLER_24_1020 ();
 sg13g2_fill_2 FILLER_24_1030 ();
 sg13g2_decap_8 FILLER_24_1053 ();
 sg13g2_decap_4 FILLER_24_1073 ();
 sg13g2_fill_2 FILLER_24_1077 ();
 sg13g2_fill_2 FILLER_24_1092 ();
 sg13g2_fill_1 FILLER_24_1094 ();
 sg13g2_decap_8 FILLER_24_1105 ();
 sg13g2_decap_8 FILLER_24_1112 ();
 sg13g2_decap_8 FILLER_24_1119 ();
 sg13g2_fill_2 FILLER_24_1126 ();
 sg13g2_fill_1 FILLER_24_1146 ();
 sg13g2_fill_1 FILLER_24_1154 ();
 sg13g2_fill_2 FILLER_24_1175 ();
 sg13g2_fill_1 FILLER_24_1177 ();
 sg13g2_decap_4 FILLER_24_1196 ();
 sg13g2_fill_1 FILLER_24_1200 ();
 sg13g2_decap_8 FILLER_24_1229 ();
 sg13g2_decap_8 FILLER_24_1236 ();
 sg13g2_decap_8 FILLER_24_1261 ();
 sg13g2_fill_2 FILLER_24_1268 ();
 sg13g2_fill_1 FILLER_24_1270 ();
 sg13g2_decap_8 FILLER_24_1304 ();
 sg13g2_decap_8 FILLER_24_1311 ();
 sg13g2_decap_8 FILLER_24_1318 ();
 sg13g2_decap_8 FILLER_24_1325 ();
 sg13g2_decap_8 FILLER_24_1332 ();
 sg13g2_decap_8 FILLER_24_1339 ();
 sg13g2_decap_4 FILLER_24_1346 ();
 sg13g2_fill_1 FILLER_24_1350 ();
 sg13g2_decap_8 FILLER_24_1453 ();
 sg13g2_decap_8 FILLER_24_1460 ();
 sg13g2_decap_4 FILLER_24_1467 ();
 sg13g2_fill_2 FILLER_24_1471 ();
 sg13g2_fill_2 FILLER_24_1482 ();
 sg13g2_fill_1 FILLER_24_1496 ();
 sg13g2_decap_8 FILLER_24_1542 ();
 sg13g2_decap_8 FILLER_24_1549 ();
 sg13g2_decap_8 FILLER_24_1556 ();
 sg13g2_decap_4 FILLER_24_1563 ();
 sg13g2_fill_2 FILLER_24_1567 ();
 sg13g2_fill_2 FILLER_24_1584 ();
 sg13g2_decap_8 FILLER_24_1600 ();
 sg13g2_fill_2 FILLER_24_1607 ();
 sg13g2_fill_1 FILLER_24_1609 ();
 sg13g2_fill_2 FILLER_24_1639 ();
 sg13g2_fill_1 FILLER_24_1641 ();
 sg13g2_decap_4 FILLER_24_1647 ();
 sg13g2_fill_1 FILLER_24_1651 ();
 sg13g2_decap_8 FILLER_24_1677 ();
 sg13g2_fill_2 FILLER_24_1684 ();
 sg13g2_decap_8 FILLER_24_1691 ();
 sg13g2_decap_4 FILLER_24_1698 ();
 sg13g2_fill_2 FILLER_24_1702 ();
 sg13g2_fill_2 FILLER_24_1722 ();
 sg13g2_fill_2 FILLER_24_1729 ();
 sg13g2_decap_8 FILLER_24_1749 ();
 sg13g2_decap_4 FILLER_24_1756 ();
 sg13g2_decap_8 FILLER_24_1809 ();
 sg13g2_decap_4 FILLER_24_1816 ();
 sg13g2_fill_2 FILLER_24_1869 ();
 sg13g2_decap_4 FILLER_24_1876 ();
 sg13g2_fill_1 FILLER_24_1880 ();
 sg13g2_decap_4 FILLER_24_1929 ();
 sg13g2_fill_2 FILLER_24_1942 ();
 sg13g2_fill_1 FILLER_24_1976 ();
 sg13g2_fill_1 FILLER_24_1990 ();
 sg13g2_decap_8 FILLER_24_2022 ();
 sg13g2_decap_8 FILLER_24_2029 ();
 sg13g2_fill_2 FILLER_24_2036 ();
 sg13g2_fill_1 FILLER_24_2038 ();
 sg13g2_fill_2 FILLER_24_2048 ();
 sg13g2_decap_8 FILLER_24_2077 ();
 sg13g2_decap_8 FILLER_24_2084 ();
 sg13g2_decap_4 FILLER_24_2091 ();
 sg13g2_decap_8 FILLER_24_2113 ();
 sg13g2_decap_8 FILLER_24_2120 ();
 sg13g2_decap_8 FILLER_24_2127 ();
 sg13g2_decap_8 FILLER_24_2134 ();
 sg13g2_decap_8 FILLER_24_2141 ();
 sg13g2_decap_4 FILLER_24_2158 ();
 sg13g2_decap_8 FILLER_24_2167 ();
 sg13g2_decap_4 FILLER_24_2174 ();
 sg13g2_fill_1 FILLER_24_2178 ();
 sg13g2_decap_8 FILLER_24_2192 ();
 sg13g2_decap_4 FILLER_24_2199 ();
 sg13g2_fill_1 FILLER_24_2203 ();
 sg13g2_fill_2 FILLER_24_2223 ();
 sg13g2_fill_1 FILLER_24_2225 ();
 sg13g2_fill_2 FILLER_24_2246 ();
 sg13g2_fill_1 FILLER_24_2285 ();
 sg13g2_fill_2 FILLER_24_2299 ();
 sg13g2_fill_1 FILLER_24_2301 ();
 sg13g2_fill_2 FILLER_24_2324 ();
 sg13g2_fill_1 FILLER_24_2326 ();
 sg13g2_fill_2 FILLER_24_2336 ();
 sg13g2_decap_8 FILLER_24_2360 ();
 sg13g2_fill_2 FILLER_24_2367 ();
 sg13g2_fill_1 FILLER_24_2369 ();
 sg13g2_fill_2 FILLER_24_2378 ();
 sg13g2_decap_8 FILLER_24_2411 ();
 sg13g2_decap_8 FILLER_24_2418 ();
 sg13g2_decap_8 FILLER_24_2425 ();
 sg13g2_decap_8 FILLER_24_2432 ();
 sg13g2_decap_8 FILLER_24_2439 ();
 sg13g2_decap_8 FILLER_24_2446 ();
 sg13g2_fill_2 FILLER_24_2453 ();
 sg13g2_fill_1 FILLER_24_2473 ();
 sg13g2_decap_8 FILLER_24_2487 ();
 sg13g2_decap_8 FILLER_24_2494 ();
 sg13g2_decap_8 FILLER_24_2501 ();
 sg13g2_decap_8 FILLER_24_2508 ();
 sg13g2_decap_8 FILLER_24_2515 ();
 sg13g2_decap_4 FILLER_24_2526 ();
 sg13g2_decap_8 FILLER_24_2568 ();
 sg13g2_fill_1 FILLER_24_2575 ();
 sg13g2_fill_2 FILLER_24_2593 ();
 sg13g2_fill_1 FILLER_24_2595 ();
 sg13g2_decap_8 FILLER_24_2635 ();
 sg13g2_fill_2 FILLER_24_2642 ();
 sg13g2_fill_1 FILLER_24_2658 ();
 sg13g2_fill_2 FILLER_24_2672 ();
 sg13g2_decap_4 FILLER_24_2683 ();
 sg13g2_decap_4 FILLER_24_2714 ();
 sg13g2_fill_1 FILLER_24_2718 ();
 sg13g2_decap_8 FILLER_24_2723 ();
 sg13g2_decap_8 FILLER_24_2730 ();
 sg13g2_fill_2 FILLER_24_2737 ();
 sg13g2_fill_1 FILLER_24_2743 ();
 sg13g2_decap_8 FILLER_24_2793 ();
 sg13g2_decap_8 FILLER_24_2800 ();
 sg13g2_fill_1 FILLER_24_2817 ();
 sg13g2_decap_8 FILLER_24_2855 ();
 sg13g2_decap_4 FILLER_24_2862 ();
 sg13g2_fill_2 FILLER_24_2866 ();
 sg13g2_decap_8 FILLER_24_2997 ();
 sg13g2_decap_8 FILLER_24_3004 ();
 sg13g2_decap_8 FILLER_24_3011 ();
 sg13g2_fill_1 FILLER_24_3045 ();
 sg13g2_decap_8 FILLER_24_3059 ();
 sg13g2_decap_8 FILLER_24_3066 ();
 sg13g2_fill_2 FILLER_24_3073 ();
 sg13g2_fill_2 FILLER_24_3079 ();
 sg13g2_decap_8 FILLER_24_3113 ();
 sg13g2_decap_8 FILLER_24_3120 ();
 sg13g2_decap_4 FILLER_24_3127 ();
 sg13g2_fill_1 FILLER_24_3172 ();
 sg13g2_decap_8 FILLER_24_3200 ();
 sg13g2_decap_8 FILLER_24_3207 ();
 sg13g2_decap_4 FILLER_24_3214 ();
 sg13g2_fill_1 FILLER_24_3218 ();
 sg13g2_decap_8 FILLER_24_3275 ();
 sg13g2_decap_8 FILLER_24_3282 ();
 sg13g2_decap_4 FILLER_24_3289 ();
 sg13g2_fill_1 FILLER_24_3293 ();
 sg13g2_fill_2 FILLER_24_3327 ();
 sg13g2_fill_1 FILLER_24_3329 ();
 sg13g2_fill_1 FILLER_24_3377 ();
 sg13g2_decap_8 FILLER_24_3387 ();
 sg13g2_decap_8 FILLER_24_3394 ();
 sg13g2_decap_8 FILLER_24_3401 ();
 sg13g2_fill_1 FILLER_24_3408 ();
 sg13g2_decap_8 FILLER_24_3458 ();
 sg13g2_decap_8 FILLER_24_3465 ();
 sg13g2_decap_8 FILLER_24_3472 ();
 sg13g2_fill_2 FILLER_24_3479 ();
 sg13g2_fill_1 FILLER_24_3481 ();
 sg13g2_fill_2 FILLER_24_3500 ();
 sg13g2_decap_4 FILLER_24_3524 ();
 sg13g2_decap_8 FILLER_24_3565 ();
 sg13g2_decap_4 FILLER_24_3572 ();
 sg13g2_fill_2 FILLER_24_3576 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_1 FILLER_25_33 ();
 sg13g2_decap_8 FILLER_25_55 ();
 sg13g2_decap_4 FILLER_25_62 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_decap_8 FILLER_25_107 ();
 sg13g2_fill_2 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_decap_8 FILLER_25_183 ();
 sg13g2_decap_8 FILLER_25_190 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_278 ();
 sg13g2_decap_4 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_289 ();
 sg13g2_decap_4 FILLER_25_293 ();
 sg13g2_fill_2 FILLER_25_297 ();
 sg13g2_decap_8 FILLER_25_302 ();
 sg13g2_decap_8 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_decap_4 FILLER_25_345 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_375 ();
 sg13g2_decap_4 FILLER_25_386 ();
 sg13g2_fill_2 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_430 ();
 sg13g2_decap_4 FILLER_25_437 ();
 sg13g2_fill_1 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_447 ();
 sg13g2_decap_8 FILLER_25_454 ();
 sg13g2_decap_8 FILLER_25_461 ();
 sg13g2_fill_1 FILLER_25_473 ();
 sg13g2_decap_8 FILLER_25_506 ();
 sg13g2_decap_8 FILLER_25_513 ();
 sg13g2_decap_8 FILLER_25_520 ();
 sg13g2_decap_8 FILLER_25_527 ();
 sg13g2_decap_8 FILLER_25_561 ();
 sg13g2_decap_8 FILLER_25_568 ();
 sg13g2_fill_2 FILLER_25_575 ();
 sg13g2_fill_1 FILLER_25_577 ();
 sg13g2_fill_1 FILLER_25_583 ();
 sg13g2_decap_8 FILLER_25_592 ();
 sg13g2_decap_8 FILLER_25_608 ();
 sg13g2_decap_4 FILLER_25_615 ();
 sg13g2_fill_1 FILLER_25_619 ();
 sg13g2_fill_2 FILLER_25_625 ();
 sg13g2_fill_1 FILLER_25_681 ();
 sg13g2_decap_8 FILLER_25_691 ();
 sg13g2_decap_8 FILLER_25_698 ();
 sg13g2_decap_8 FILLER_25_705 ();
 sg13g2_decap_8 FILLER_25_712 ();
 sg13g2_decap_8 FILLER_25_761 ();
 sg13g2_fill_1 FILLER_25_768 ();
 sg13g2_fill_2 FILLER_25_780 ();
 sg13g2_decap_8 FILLER_25_790 ();
 sg13g2_decap_8 FILLER_25_797 ();
 sg13g2_decap_8 FILLER_25_804 ();
 sg13g2_fill_1 FILLER_25_811 ();
 sg13g2_fill_1 FILLER_25_843 ();
 sg13g2_fill_2 FILLER_25_870 ();
 sg13g2_fill_2 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_25_884 ();
 sg13g2_decap_8 FILLER_25_891 ();
 sg13g2_decap_8 FILLER_25_898 ();
 sg13g2_fill_2 FILLER_25_905 ();
 sg13g2_fill_1 FILLER_25_925 ();
 sg13g2_decap_8 FILLER_25_947 ();
 sg13g2_decap_8 FILLER_25_954 ();
 sg13g2_decap_8 FILLER_25_961 ();
 sg13g2_decap_8 FILLER_25_968 ();
 sg13g2_fill_1 FILLER_25_987 ();
 sg13g2_decap_4 FILLER_25_996 ();
 sg13g2_fill_2 FILLER_25_1009 ();
 sg13g2_fill_1 FILLER_25_1011 ();
 sg13g2_fill_2 FILLER_25_1044 ();
 sg13g2_decap_8 FILLER_25_1059 ();
 sg13g2_decap_8 FILLER_25_1066 ();
 sg13g2_decap_4 FILLER_25_1073 ();
 sg13g2_fill_1 FILLER_25_1077 ();
 sg13g2_decap_8 FILLER_25_1106 ();
 sg13g2_fill_2 FILLER_25_1113 ();
 sg13g2_fill_1 FILLER_25_1115 ();
 sg13g2_fill_2 FILLER_25_1120 ();
 sg13g2_fill_2 FILLER_25_1158 ();
 sg13g2_fill_1 FILLER_25_1160 ();
 sg13g2_decap_8 FILLER_25_1204 ();
 sg13g2_decap_4 FILLER_25_1211 ();
 sg13g2_fill_1 FILLER_25_1215 ();
 sg13g2_decap_8 FILLER_25_1229 ();
 sg13g2_decap_8 FILLER_25_1236 ();
 sg13g2_fill_2 FILLER_25_1243 ();
 sg13g2_fill_1 FILLER_25_1245 ();
 sg13g2_decap_4 FILLER_25_1250 ();
 sg13g2_fill_1 FILLER_25_1254 ();
 sg13g2_decap_8 FILLER_25_1268 ();
 sg13g2_fill_1 FILLER_25_1290 ();
 sg13g2_fill_1 FILLER_25_1296 ();
 sg13g2_decap_8 FILLER_25_1310 ();
 sg13g2_decap_8 FILLER_25_1317 ();
 sg13g2_decap_8 FILLER_25_1324 ();
 sg13g2_decap_8 FILLER_25_1331 ();
 sg13g2_decap_4 FILLER_25_1338 ();
 sg13g2_fill_2 FILLER_25_1355 ();
 sg13g2_fill_1 FILLER_25_1357 ();
 sg13g2_fill_1 FILLER_25_1373 ();
 sg13g2_fill_1 FILLER_25_1402 ();
 sg13g2_fill_2 FILLER_25_1425 ();
 sg13g2_fill_2 FILLER_25_1446 ();
 sg13g2_fill_1 FILLER_25_1448 ();
 sg13g2_decap_8 FILLER_25_1462 ();
 sg13g2_fill_1 FILLER_25_1477 ();
 sg13g2_decap_8 FILLER_25_1484 ();
 sg13g2_fill_2 FILLER_25_1491 ();
 sg13g2_fill_1 FILLER_25_1493 ();
 sg13g2_decap_8 FILLER_25_1534 ();
 sg13g2_decap_8 FILLER_25_1541 ();
 sg13g2_decap_8 FILLER_25_1548 ();
 sg13g2_decap_4 FILLER_25_1555 ();
 sg13g2_fill_1 FILLER_25_1559 ();
 sg13g2_fill_2 FILLER_25_1606 ();
 sg13g2_fill_1 FILLER_25_1608 ();
 sg13g2_decap_4 FILLER_25_1627 ();
 sg13g2_decap_4 FILLER_25_1651 ();
 sg13g2_fill_2 FILLER_25_1655 ();
 sg13g2_decap_8 FILLER_25_1672 ();
 sg13g2_decap_4 FILLER_25_1684 ();
 sg13g2_fill_2 FILLER_25_1688 ();
 sg13g2_fill_1 FILLER_25_1696 ();
 sg13g2_decap_4 FILLER_25_1708 ();
 sg13g2_fill_2 FILLER_25_1720 ();
 sg13g2_fill_2 FILLER_25_1727 ();
 sg13g2_decap_8 FILLER_25_1752 ();
 sg13g2_decap_8 FILLER_25_1759 ();
 sg13g2_fill_2 FILLER_25_1794 ();
 sg13g2_decap_4 FILLER_25_1822 ();
 sg13g2_decap_4 FILLER_25_1863 ();
 sg13g2_decap_8 FILLER_25_1938 ();
 sg13g2_decap_8 FILLER_25_1945 ();
 sg13g2_fill_1 FILLER_25_1952 ();
 sg13g2_decap_4 FILLER_25_1985 ();
 sg13g2_fill_1 FILLER_25_1989 ();
 sg13g2_fill_2 FILLER_25_2017 ();
 sg13g2_decap_4 FILLER_25_2038 ();
 sg13g2_fill_1 FILLER_25_2061 ();
 sg13g2_decap_8 FILLER_25_2089 ();
 sg13g2_fill_1 FILLER_25_2096 ();
 sg13g2_decap_8 FILLER_25_2123 ();
 sg13g2_decap_8 FILLER_25_2130 ();
 sg13g2_fill_1 FILLER_25_2137 ();
 sg13g2_decap_8 FILLER_25_2142 ();
 sg13g2_decap_8 FILLER_25_2149 ();
 sg13g2_decap_8 FILLER_25_2156 ();
 sg13g2_fill_2 FILLER_25_2163 ();
 sg13g2_fill_1 FILLER_25_2165 ();
 sg13g2_decap_8 FILLER_25_2188 ();
 sg13g2_decap_8 FILLER_25_2195 ();
 sg13g2_decap_8 FILLER_25_2202 ();
 sg13g2_fill_2 FILLER_25_2209 ();
 sg13g2_fill_1 FILLER_25_2211 ();
 sg13g2_fill_2 FILLER_25_2217 ();
 sg13g2_decap_8 FILLER_25_2239 ();
 sg13g2_decap_4 FILLER_25_2246 ();
 sg13g2_fill_1 FILLER_25_2250 ();
 sg13g2_fill_1 FILLER_25_2288 ();
 sg13g2_fill_1 FILLER_25_2311 ();
 sg13g2_fill_2 FILLER_25_2317 ();
 sg13g2_fill_1 FILLER_25_2319 ();
 sg13g2_fill_2 FILLER_25_2325 ();
 sg13g2_decap_8 FILLER_25_2355 ();
 sg13g2_decap_8 FILLER_25_2362 ();
 sg13g2_decap_8 FILLER_25_2369 ();
 sg13g2_decap_8 FILLER_25_2376 ();
 sg13g2_fill_2 FILLER_25_2383 ();
 sg13g2_fill_1 FILLER_25_2385 ();
 sg13g2_fill_2 FILLER_25_2405 ();
 sg13g2_fill_1 FILLER_25_2407 ();
 sg13g2_decap_8 FILLER_25_2444 ();
 sg13g2_fill_2 FILLER_25_2451 ();
 sg13g2_decap_8 FILLER_25_2495 ();
 sg13g2_decap_8 FILLER_25_2502 ();
 sg13g2_decap_8 FILLER_25_2557 ();
 sg13g2_decap_8 FILLER_25_2564 ();
 sg13g2_decap_8 FILLER_25_2571 ();
 sg13g2_decap_4 FILLER_25_2578 ();
 sg13g2_fill_1 FILLER_25_2582 ();
 sg13g2_fill_2 FILLER_25_2593 ();
 sg13g2_fill_1 FILLER_25_2595 ();
 sg13g2_decap_8 FILLER_25_2645 ();
 sg13g2_decap_4 FILLER_25_2652 ();
 sg13g2_fill_2 FILLER_25_2656 ();
 sg13g2_decap_8 FILLER_25_2671 ();
 sg13g2_decap_4 FILLER_25_2678 ();
 sg13g2_fill_1 FILLER_25_2682 ();
 sg13g2_decap_8 FILLER_25_2716 ();
 sg13g2_decap_8 FILLER_25_2723 ();
 sg13g2_decap_4 FILLER_25_2730 ();
 sg13g2_fill_2 FILLER_25_2761 ();
 sg13g2_fill_1 FILLER_25_2834 ();
 sg13g2_decap_8 FILLER_25_2862 ();
 sg13g2_decap_8 FILLER_25_2869 ();
 sg13g2_decap_8 FILLER_25_2907 ();
 sg13g2_decap_8 FILLER_25_2914 ();
 sg13g2_decap_8 FILLER_25_2925 ();
 sg13g2_decap_8 FILLER_25_2932 ();
 sg13g2_decap_4 FILLER_25_2939 ();
 sg13g2_decap_8 FILLER_25_3000 ();
 sg13g2_fill_2 FILLER_25_3007 ();
 sg13g2_fill_1 FILLER_25_3009 ();
 sg13g2_fill_2 FILLER_25_3041 ();
 sg13g2_fill_1 FILLER_25_3043 ();
 sg13g2_decap_8 FILLER_25_3065 ();
 sg13g2_decap_8 FILLER_25_3072 ();
 sg13g2_fill_2 FILLER_25_3079 ();
 sg13g2_fill_1 FILLER_25_3081 ();
 sg13g2_decap_8 FILLER_25_3109 ();
 sg13g2_decap_4 FILLER_25_3116 ();
 sg13g2_fill_2 FILLER_25_3120 ();
 sg13g2_decap_4 FILLER_25_3131 ();
 sg13g2_fill_1 FILLER_25_3135 ();
 sg13g2_fill_1 FILLER_25_3149 ();
 sg13g2_fill_2 FILLER_25_3193 ();
 sg13g2_fill_1 FILLER_25_3195 ();
 sg13g2_decap_8 FILLER_25_3209 ();
 sg13g2_decap_8 FILLER_25_3216 ();
 sg13g2_decap_4 FILLER_25_3223 ();
 sg13g2_fill_2 FILLER_25_3240 ();
 sg13g2_fill_2 FILLER_25_3252 ();
 sg13g2_fill_1 FILLER_25_3254 ();
 sg13g2_decap_8 FILLER_25_3271 ();
 sg13g2_decap_8 FILLER_25_3278 ();
 sg13g2_decap_8 FILLER_25_3285 ();
 sg13g2_decap_8 FILLER_25_3292 ();
 sg13g2_decap_8 FILLER_25_3299 ();
 sg13g2_fill_2 FILLER_25_3310 ();
 sg13g2_fill_1 FILLER_25_3312 ();
 sg13g2_decap_8 FILLER_25_3317 ();
 sg13g2_decap_8 FILLER_25_3324 ();
 sg13g2_decap_4 FILLER_25_3331 ();
 sg13g2_fill_2 FILLER_25_3335 ();
 sg13g2_decap_4 FILLER_25_3347 ();
 sg13g2_fill_2 FILLER_25_3351 ();
 sg13g2_decap_8 FILLER_25_3375 ();
 sg13g2_decap_8 FILLER_25_3382 ();
 sg13g2_decap_8 FILLER_25_3389 ();
 sg13g2_decap_8 FILLER_25_3396 ();
 sg13g2_decap_8 FILLER_25_3403 ();
 sg13g2_decap_8 FILLER_25_3410 ();
 sg13g2_fill_1 FILLER_25_3417 ();
 sg13g2_fill_1 FILLER_25_3428 ();
 sg13g2_decap_4 FILLER_25_3438 ();
 sg13g2_decap_4 FILLER_25_3452 ();
 sg13g2_fill_1 FILLER_25_3456 ();
 sg13g2_decap_8 FILLER_25_3466 ();
 sg13g2_decap_8 FILLER_25_3473 ();
 sg13g2_decap_8 FILLER_25_3480 ();
 sg13g2_decap_4 FILLER_25_3487 ();
 sg13g2_decap_8 FILLER_25_3501 ();
 sg13g2_decap_8 FILLER_25_3526 ();
 sg13g2_fill_1 FILLER_25_3533 ();
 sg13g2_fill_1 FILLER_25_3544 ();
 sg13g2_decap_4 FILLER_25_3572 ();
 sg13g2_fill_2 FILLER_25_3576 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_decap_4 FILLER_26_59 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_fill_2 FILLER_26_69 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_decap_8 FILLER_26_99 ();
 sg13g2_decap_8 FILLER_26_106 ();
 sg13g2_decap_4 FILLER_26_113 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_fill_2 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_405 ();
 sg13g2_fill_2 FILLER_26_412 ();
 sg13g2_fill_1 FILLER_26_428 ();
 sg13g2_fill_2 FILLER_26_437 ();
 sg13g2_fill_2 FILLER_26_467 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_fill_2 FILLER_26_525 ();
 sg13g2_fill_1 FILLER_26_527 ();
 sg13g2_fill_2 FILLER_26_533 ();
 sg13g2_fill_1 FILLER_26_535 ();
 sg13g2_decap_8 FILLER_26_562 ();
 sg13g2_decap_8 FILLER_26_569 ();
 sg13g2_decap_8 FILLER_26_576 ();
 sg13g2_fill_2 FILLER_26_583 ();
 sg13g2_decap_8 FILLER_26_593 ();
 sg13g2_decap_8 FILLER_26_600 ();
 sg13g2_decap_8 FILLER_26_607 ();
 sg13g2_decap_8 FILLER_26_614 ();
 sg13g2_decap_8 FILLER_26_621 ();
 sg13g2_decap_8 FILLER_26_628 ();
 sg13g2_decap_8 FILLER_26_635 ();
 sg13g2_fill_1 FILLER_26_642 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_4 FILLER_26_700 ();
 sg13g2_fill_1 FILLER_26_704 ();
 sg13g2_decap_4 FILLER_26_733 ();
 sg13g2_fill_1 FILLER_26_737 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_4 FILLER_26_803 ();
 sg13g2_fill_2 FILLER_26_807 ();
 sg13g2_decap_4 FILLER_26_837 ();
 sg13g2_fill_2 FILLER_26_841 ();
 sg13g2_fill_1 FILLER_26_856 ();
 sg13g2_decap_8 FILLER_26_883 ();
 sg13g2_decap_4 FILLER_26_890 ();
 sg13g2_fill_1 FILLER_26_894 ();
 sg13g2_fill_1 FILLER_26_979 ();
 sg13g2_fill_1 FILLER_26_991 ();
 sg13g2_fill_2 FILLER_26_1018 ();
 sg13g2_fill_1 FILLER_26_1020 ();
 sg13g2_decap_8 FILLER_26_1058 ();
 sg13g2_decap_8 FILLER_26_1065 ();
 sg13g2_fill_1 FILLER_26_1072 ();
 sg13g2_fill_1 FILLER_26_1149 ();
 sg13g2_fill_1 FILLER_26_1173 ();
 sg13g2_fill_1 FILLER_26_1179 ();
 sg13g2_decap_8 FILLER_26_1184 ();
 sg13g2_decap_8 FILLER_26_1191 ();
 sg13g2_decap_8 FILLER_26_1208 ();
 sg13g2_decap_8 FILLER_26_1215 ();
 sg13g2_decap_8 FILLER_26_1222 ();
 sg13g2_decap_4 FILLER_26_1229 ();
 sg13g2_fill_2 FILLER_26_1233 ();
 sg13g2_fill_2 FILLER_26_1248 ();
 sg13g2_decap_8 FILLER_26_1263 ();
 sg13g2_fill_2 FILLER_26_1270 ();
 sg13g2_fill_1 FILLER_26_1300 ();
 sg13g2_fill_2 FILLER_26_1309 ();
 sg13g2_fill_2 FILLER_26_1333 ();
 sg13g2_fill_1 FILLER_26_1335 ();
 sg13g2_decap_8 FILLER_26_1340 ();
 sg13g2_decap_8 FILLER_26_1347 ();
 sg13g2_decap_4 FILLER_26_1400 ();
 sg13g2_fill_1 FILLER_26_1412 ();
 sg13g2_decap_4 FILLER_26_1453 ();
 sg13g2_fill_2 FILLER_26_1457 ();
 sg13g2_decap_8 FILLER_26_1487 ();
 sg13g2_decap_4 FILLER_26_1494 ();
 sg13g2_fill_1 FILLER_26_1498 ();
 sg13g2_fill_2 FILLER_26_1507 ();
 sg13g2_decap_8 FILLER_26_1544 ();
 sg13g2_decap_8 FILLER_26_1551 ();
 sg13g2_decap_4 FILLER_26_1558 ();
 sg13g2_fill_1 FILLER_26_1562 ();
 sg13g2_fill_1 FILLER_26_1596 ();
 sg13g2_fill_2 FILLER_26_1625 ();
 sg13g2_fill_1 FILLER_26_1627 ();
 sg13g2_decap_8 FILLER_26_1643 ();
 sg13g2_fill_2 FILLER_26_1662 ();
 sg13g2_decap_8 FILLER_26_1669 ();
 sg13g2_fill_2 FILLER_26_1676 ();
 sg13g2_fill_1 FILLER_26_1678 ();
 sg13g2_decap_4 FILLER_26_1695 ();
 sg13g2_fill_2 FILLER_26_1705 ();
 sg13g2_fill_1 FILLER_26_1707 ();
 sg13g2_fill_2 FILLER_26_1733 ();
 sg13g2_decap_8 FILLER_26_1754 ();
 sg13g2_decap_8 FILLER_26_1761 ();
 sg13g2_fill_2 FILLER_26_1768 ();
 sg13g2_fill_2 FILLER_26_1776 ();
 sg13g2_fill_1 FILLER_26_1778 ();
 sg13g2_fill_1 FILLER_26_1793 ();
 sg13g2_fill_1 FILLER_26_1798 ();
 sg13g2_fill_2 FILLER_26_1803 ();
 sg13g2_fill_1 FILLER_26_1805 ();
 sg13g2_decap_8 FILLER_26_1819 ();
 sg13g2_decap_4 FILLER_26_1826 ();
 sg13g2_fill_1 FILLER_26_1842 ();
 sg13g2_decap_8 FILLER_26_1861 ();
 sg13g2_fill_2 FILLER_26_1931 ();
 sg13g2_fill_1 FILLER_26_1933 ();
 sg13g2_decap_4 FILLER_26_1943 ();
 sg13g2_fill_1 FILLER_26_1947 ();
 sg13g2_decap_4 FILLER_26_1953 ();
 sg13g2_fill_1 FILLER_26_1957 ();
 sg13g2_fill_1 FILLER_26_1966 ();
 sg13g2_decap_8 FILLER_26_1975 ();
 sg13g2_decap_8 FILLER_26_1982 ();
 sg13g2_decap_8 FILLER_26_1989 ();
 sg13g2_decap_4 FILLER_26_1996 ();
 sg13g2_decap_8 FILLER_26_2021 ();
 sg13g2_fill_1 FILLER_26_2028 ();
 sg13g2_decap_8 FILLER_26_2034 ();
 sg13g2_decap_4 FILLER_26_2041 ();
 sg13g2_fill_1 FILLER_26_2045 ();
 sg13g2_decap_8 FILLER_26_2077 ();
 sg13g2_decap_8 FILLER_26_2084 ();
 sg13g2_fill_2 FILLER_26_2091 ();
 sg13g2_decap_8 FILLER_26_2130 ();
 sg13g2_fill_2 FILLER_26_2137 ();
 sg13g2_fill_1 FILLER_26_2159 ();
 sg13g2_fill_1 FILLER_26_2165 ();
 sg13g2_decap_8 FILLER_26_2196 ();
 sg13g2_decap_8 FILLER_26_2237 ();
 sg13g2_decap_8 FILLER_26_2244 ();
 sg13g2_decap_4 FILLER_26_2251 ();
 sg13g2_fill_1 FILLER_26_2273 ();
 sg13g2_fill_1 FILLER_26_2297 ();
 sg13g2_fill_2 FILLER_26_2308 ();
 sg13g2_decap_8 FILLER_26_2360 ();
 sg13g2_decap_8 FILLER_26_2367 ();
 sg13g2_decap_8 FILLER_26_2374 ();
 sg13g2_decap_4 FILLER_26_2381 ();
 sg13g2_decap_4 FILLER_26_2403 ();
 sg13g2_fill_2 FILLER_26_2417 ();
 sg13g2_fill_1 FILLER_26_2419 ();
 sg13g2_decap_8 FILLER_26_2443 ();
 sg13g2_decap_4 FILLER_26_2450 ();
 sg13g2_fill_2 FILLER_26_2454 ();
 sg13g2_decap_8 FILLER_26_2498 ();
 sg13g2_fill_1 FILLER_26_2532 ();
 sg13g2_fill_2 FILLER_26_2537 ();
 sg13g2_decap_8 FILLER_26_2566 ();
 sg13g2_decap_4 FILLER_26_2573 ();
 sg13g2_fill_1 FILLER_26_2577 ();
 sg13g2_decap_4 FILLER_26_2604 ();
 sg13g2_fill_1 FILLER_26_2608 ();
 sg13g2_fill_2 FILLER_26_2619 ();
 sg13g2_fill_1 FILLER_26_2621 ();
 sg13g2_fill_2 FILLER_26_2632 ();
 sg13g2_decap_8 FILLER_26_2659 ();
 sg13g2_decap_4 FILLER_26_2666 ();
 sg13g2_fill_2 FILLER_26_2675 ();
 sg13g2_fill_1 FILLER_26_2677 ();
 sg13g2_decap_8 FILLER_26_2711 ();
 sg13g2_decap_8 FILLER_26_2718 ();
 sg13g2_decap_4 FILLER_26_2725 ();
 sg13g2_fill_2 FILLER_26_2729 ();
 sg13g2_fill_2 FILLER_26_2763 ();
 sg13g2_decap_8 FILLER_26_2792 ();
 sg13g2_decap_8 FILLER_26_2799 ();
 sg13g2_fill_2 FILLER_26_2806 ();
 sg13g2_fill_2 FILLER_26_2861 ();
 sg13g2_decap_8 FILLER_26_2866 ();
 sg13g2_decap_8 FILLER_26_2873 ();
 sg13g2_decap_4 FILLER_26_2936 ();
 sg13g2_fill_2 FILLER_26_2940 ();
 sg13g2_decap_8 FILLER_26_2979 ();
 sg13g2_decap_8 FILLER_26_2986 ();
 sg13g2_decap_8 FILLER_26_2993 ();
 sg13g2_decap_4 FILLER_26_3000 ();
 sg13g2_fill_1 FILLER_26_3004 ();
 sg13g2_fill_2 FILLER_26_3019 ();
 sg13g2_fill_2 FILLER_26_3048 ();
 sg13g2_decap_4 FILLER_26_3077 ();
 sg13g2_fill_2 FILLER_26_3081 ();
 sg13g2_decap_8 FILLER_26_3141 ();
 sg13g2_decap_8 FILLER_26_3148 ();
 sg13g2_fill_1 FILLER_26_3159 ();
 sg13g2_fill_1 FILLER_26_3184 ();
 sg13g2_decap_8 FILLER_26_3194 ();
 sg13g2_decap_8 FILLER_26_3201 ();
 sg13g2_decap_4 FILLER_26_3208 ();
 sg13g2_fill_1 FILLER_26_3212 ();
 sg13g2_decap_8 FILLER_26_3226 ();
 sg13g2_fill_2 FILLER_26_3233 ();
 sg13g2_fill_1 FILLER_26_3235 ();
 sg13g2_fill_2 FILLER_26_3249 ();
 sg13g2_fill_1 FILLER_26_3265 ();
 sg13g2_decap_8 FILLER_26_3271 ();
 sg13g2_decap_8 FILLER_26_3278 ();
 sg13g2_fill_2 FILLER_26_3285 ();
 sg13g2_decap_8 FILLER_26_3314 ();
 sg13g2_decap_8 FILLER_26_3321 ();
 sg13g2_decap_8 FILLER_26_3328 ();
 sg13g2_decap_8 FILLER_26_3335 ();
 sg13g2_fill_2 FILLER_26_3342 ();
 sg13g2_fill_1 FILLER_26_3344 ();
 sg13g2_decap_4 FILLER_26_3386 ();
 sg13g2_fill_1 FILLER_26_3390 ();
 sg13g2_decap_8 FILLER_26_3400 ();
 sg13g2_decap_8 FILLER_26_3407 ();
 sg13g2_decap_8 FILLER_26_3414 ();
 sg13g2_decap_4 FILLER_26_3421 ();
 sg13g2_fill_2 FILLER_26_3425 ();
 sg13g2_decap_4 FILLER_26_3437 ();
 sg13g2_decap_8 FILLER_26_3468 ();
 sg13g2_decap_8 FILLER_26_3475 ();
 sg13g2_decap_8 FILLER_26_3482 ();
 sg13g2_decap_8 FILLER_26_3516 ();
 sg13g2_decap_4 FILLER_26_3523 ();
 sg13g2_fill_2 FILLER_26_3527 ();
 sg13g2_decap_8 FILLER_26_3566 ();
 sg13g2_decap_4 FILLER_26_3573 ();
 sg13g2_fill_1 FILLER_26_3577 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_decap_4 FILLER_27_53 ();
 sg13g2_decap_8 FILLER_27_111 ();
 sg13g2_fill_2 FILLER_27_118 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_fill_2 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_337 ();
 sg13g2_decap_4 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_fill_1 FILLER_27_399 ();
 sg13g2_fill_1 FILLER_27_416 ();
 sg13g2_fill_2 FILLER_27_437 ();
 sg13g2_fill_1 FILLER_27_439 ();
 sg13g2_fill_2 FILLER_27_462 ();
 sg13g2_fill_1 FILLER_27_464 ();
 sg13g2_fill_2 FILLER_27_483 ();
 sg13g2_fill_1 FILLER_27_485 ();
 sg13g2_decap_8 FILLER_27_508 ();
 sg13g2_decap_8 FILLER_27_515 ();
 sg13g2_fill_2 FILLER_27_522 ();
 sg13g2_fill_1 FILLER_27_524 ();
 sg13g2_fill_2 FILLER_27_572 ();
 sg13g2_fill_1 FILLER_27_574 ();
 sg13g2_fill_2 FILLER_27_608 ();
 sg13g2_decap_8 FILLER_27_626 ();
 sg13g2_decap_8 FILLER_27_633 ();
 sg13g2_decap_8 FILLER_27_640 ();
 sg13g2_fill_1 FILLER_27_647 ();
 sg13g2_fill_2 FILLER_27_679 ();
 sg13g2_decap_4 FILLER_27_690 ();
 sg13g2_fill_1 FILLER_27_736 ();
 sg13g2_decap_8 FILLER_27_774 ();
 sg13g2_decap_4 FILLER_27_781 ();
 sg13g2_decap_8 FILLER_27_790 ();
 sg13g2_decap_8 FILLER_27_797 ();
 sg13g2_decap_8 FILLER_27_822 ();
 sg13g2_decap_4 FILLER_27_829 ();
 sg13g2_fill_1 FILLER_27_833 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_885 ();
 sg13g2_decap_8 FILLER_27_892 ();
 sg13g2_fill_2 FILLER_27_899 ();
 sg13g2_fill_1 FILLER_27_901 ();
 sg13g2_fill_2 FILLER_27_1004 ();
 sg13g2_fill_1 FILLER_27_1006 ();
 sg13g2_decap_8 FILLER_27_1049 ();
 sg13g2_decap_8 FILLER_27_1056 ();
 sg13g2_fill_1 FILLER_27_1063 ();
 sg13g2_fill_2 FILLER_27_1114 ();
 sg13g2_decap_4 FILLER_27_1157 ();
 sg13g2_decap_4 FILLER_27_1166 ();
 sg13g2_decap_4 FILLER_27_1211 ();
 sg13g2_fill_2 FILLER_27_1215 ();
 sg13g2_fill_2 FILLER_27_1245 ();
 sg13g2_decap_4 FILLER_27_1289 ();
 sg13g2_fill_2 FILLER_27_1293 ();
 sg13g2_fill_1 FILLER_27_1305 ();
 sg13g2_decap_4 FILLER_27_1357 ();
 sg13g2_fill_2 FILLER_27_1361 ();
 sg13g2_fill_1 FILLER_27_1394 ();
 sg13g2_decap_8 FILLER_27_1404 ();
 sg13g2_decap_8 FILLER_27_1411 ();
 sg13g2_fill_2 FILLER_27_1418 ();
 sg13g2_fill_1 FILLER_27_1420 ();
 sg13g2_fill_1 FILLER_27_1439 ();
 sg13g2_decap_4 FILLER_27_1444 ();
 sg13g2_fill_2 FILLER_27_1448 ();
 sg13g2_decap_8 FILLER_27_1492 ();
 sg13g2_decap_8 FILLER_27_1499 ();
 sg13g2_fill_1 FILLER_27_1506 ();
 sg13g2_decap_8 FILLER_27_1534 ();
 sg13g2_decap_4 FILLER_27_1541 ();
 sg13g2_fill_1 FILLER_27_1545 ();
 sg13g2_fill_1 FILLER_27_1573 ();
 sg13g2_decap_8 FILLER_27_1584 ();
 sg13g2_decap_8 FILLER_27_1591 ();
 sg13g2_decap_8 FILLER_27_1598 ();
 sg13g2_decap_4 FILLER_27_1605 ();
 sg13g2_fill_2 FILLER_27_1609 ();
 sg13g2_decap_8 FILLER_27_1620 ();
 sg13g2_decap_8 FILLER_27_1632 ();
 sg13g2_decap_8 FILLER_27_1639 ();
 sg13g2_decap_8 FILLER_27_1646 ();
 sg13g2_decap_4 FILLER_27_1653 ();
 sg13g2_fill_2 FILLER_27_1657 ();
 sg13g2_decap_4 FILLER_27_1683 ();
 sg13g2_fill_2 FILLER_27_1687 ();
 sg13g2_fill_1 FILLER_27_1708 ();
 sg13g2_fill_2 FILLER_27_1718 ();
 sg13g2_fill_1 FILLER_27_1720 ();
 sg13g2_decap_4 FILLER_27_1749 ();
 sg13g2_fill_2 FILLER_27_1771 ();
 sg13g2_fill_1 FILLER_27_1773 ();
 sg13g2_decap_8 FILLER_27_1787 ();
 sg13g2_decap_8 FILLER_27_1794 ();
 sg13g2_decap_8 FILLER_27_1801 ();
 sg13g2_decap_8 FILLER_27_1808 ();
 sg13g2_decap_8 FILLER_27_1815 ();
 sg13g2_decap_8 FILLER_27_1822 ();
 sg13g2_decap_4 FILLER_27_1829 ();
 sg13g2_fill_1 FILLER_27_1833 ();
 sg13g2_fill_2 FILLER_27_1842 ();
 sg13g2_decap_8 FILLER_27_1858 ();
 sg13g2_decap_4 FILLER_27_1865 ();
 sg13g2_fill_2 FILLER_27_1869 ();
 sg13g2_fill_2 FILLER_27_1888 ();
 sg13g2_fill_2 FILLER_27_1899 ();
 sg13g2_fill_1 FILLER_27_1901 ();
 sg13g2_fill_2 FILLER_27_1910 ();
 sg13g2_fill_1 FILLER_27_1921 ();
 sg13g2_fill_2 FILLER_27_1927 ();
 sg13g2_fill_1 FILLER_27_1929 ();
 sg13g2_decap_4 FILLER_27_1935 ();
 sg13g2_fill_1 FILLER_27_1939 ();
 sg13g2_fill_1 FILLER_27_1956 ();
 sg13g2_decap_8 FILLER_27_1965 ();
 sg13g2_decap_8 FILLER_27_1972 ();
 sg13g2_fill_1 FILLER_27_1979 ();
 sg13g2_decap_4 FILLER_27_1988 ();
 sg13g2_fill_2 FILLER_27_2005 ();
 sg13g2_decap_4 FILLER_27_2037 ();
 sg13g2_fill_2 FILLER_27_2041 ();
 sg13g2_fill_1 FILLER_27_2047 ();
 sg13g2_decap_8 FILLER_27_2076 ();
 sg13g2_decap_8 FILLER_27_2083 ();
 sg13g2_fill_2 FILLER_27_2102 ();
 sg13g2_fill_2 FILLER_27_2109 ();
 sg13g2_decap_8 FILLER_27_2137 ();
 sg13g2_fill_2 FILLER_27_2144 ();
 sg13g2_fill_1 FILLER_27_2146 ();
 sg13g2_fill_2 FILLER_27_2173 ();
 sg13g2_decap_4 FILLER_27_2198 ();
 sg13g2_fill_2 FILLER_27_2202 ();
 sg13g2_fill_2 FILLER_27_2222 ();
 sg13g2_decap_8 FILLER_27_2229 ();
 sg13g2_decap_8 FILLER_27_2236 ();
 sg13g2_decap_8 FILLER_27_2243 ();
 sg13g2_decap_8 FILLER_27_2250 ();
 sg13g2_fill_2 FILLER_27_2257 ();
 sg13g2_fill_1 FILLER_27_2259 ();
 sg13g2_fill_1 FILLER_27_2292 ();
 sg13g2_fill_1 FILLER_27_2310 ();
 sg13g2_fill_2 FILLER_27_2320 ();
 sg13g2_fill_1 FILLER_27_2337 ();
 sg13g2_decap_8 FILLER_27_2366 ();
 sg13g2_decap_8 FILLER_27_2373 ();
 sg13g2_fill_2 FILLER_27_2380 ();
 sg13g2_decap_4 FILLER_27_2409 ();
 sg13g2_fill_2 FILLER_27_2413 ();
 sg13g2_decap_8 FILLER_27_2436 ();
 sg13g2_fill_2 FILLER_27_2453 ();
 sg13g2_fill_1 FILLER_27_2455 ();
 sg13g2_decap_8 FILLER_27_2493 ();
 sg13g2_decap_8 FILLER_27_2500 ();
 sg13g2_fill_2 FILLER_27_2507 ();
 sg13g2_fill_1 FILLER_27_2509 ();
 sg13g2_fill_2 FILLER_27_2574 ();
 sg13g2_decap_8 FILLER_27_2656 ();
 sg13g2_decap_8 FILLER_27_2663 ();
 sg13g2_fill_2 FILLER_27_2674 ();
 sg13g2_decap_4 FILLER_27_2703 ();
 sg13g2_fill_1 FILLER_27_2707 ();
 sg13g2_decap_4 FILLER_27_2735 ();
 sg13g2_fill_1 FILLER_27_2739 ();
 sg13g2_decap_8 FILLER_27_2778 ();
 sg13g2_fill_2 FILLER_27_2785 ();
 sg13g2_decap_8 FILLER_27_2796 ();
 sg13g2_decap_8 FILLER_27_2803 ();
 sg13g2_decap_4 FILLER_27_2810 ();
 sg13g2_fill_2 FILLER_27_2814 ();
 sg13g2_decap_4 FILLER_27_2830 ();
 sg13g2_decap_8 FILLER_27_2855 ();
 sg13g2_decap_8 FILLER_27_2862 ();
 sg13g2_decap_8 FILLER_27_2874 ();
 sg13g2_decap_8 FILLER_27_2881 ();
 sg13g2_fill_2 FILLER_27_2888 ();
 sg13g2_fill_1 FILLER_27_2890 ();
 sg13g2_decap_8 FILLER_27_2913 ();
 sg13g2_decap_8 FILLER_27_2920 ();
 sg13g2_decap_4 FILLER_27_2927 ();
 sg13g2_fill_2 FILLER_27_2931 ();
 sg13g2_decap_8 FILLER_27_2983 ();
 sg13g2_decap_8 FILLER_27_2990 ();
 sg13g2_decap_8 FILLER_27_2997 ();
 sg13g2_decap_8 FILLER_27_3004 ();
 sg13g2_fill_1 FILLER_27_3044 ();
 sg13g2_decap_8 FILLER_27_3073 ();
 sg13g2_decap_8 FILLER_27_3080 ();
 sg13g2_fill_1 FILLER_27_3087 ();
 sg13g2_decap_8 FILLER_27_3092 ();
 sg13g2_fill_2 FILLER_27_3099 ();
 sg13g2_fill_1 FILLER_27_3101 ();
 sg13g2_fill_2 FILLER_27_3129 ();
 sg13g2_decap_8 FILLER_27_3141 ();
 sg13g2_fill_2 FILLER_27_3148 ();
 sg13g2_fill_1 FILLER_27_3171 ();
 sg13g2_decap_8 FILLER_27_3208 ();
 sg13g2_fill_1 FILLER_27_3215 ();
 sg13g2_decap_8 FILLER_27_3272 ();
 sg13g2_fill_2 FILLER_27_3279 ();
 sg13g2_fill_1 FILLER_27_3281 ();
 sg13g2_fill_2 FILLER_27_3377 ();
 sg13g2_fill_1 FILLER_27_3379 ();
 sg13g2_fill_2 FILLER_27_3407 ();
 sg13g2_fill_1 FILLER_27_3409 ();
 sg13g2_decap_4 FILLER_27_3480 ();
 sg13g2_fill_2 FILLER_27_3542 ();
 sg13g2_fill_1 FILLER_27_3548 ();
 sg13g2_decap_8 FILLER_27_3567 ();
 sg13g2_decap_4 FILLER_27_3574 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_43 ();
 sg13g2_decap_8 FILLER_28_50 ();
 sg13g2_decap_4 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_fill_2 FILLER_28_106 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_4 FILLER_28_201 ();
 sg13g2_decap_4 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_331 ();
 sg13g2_decap_4 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_342 ();
 sg13g2_fill_2 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_4 FILLER_28_391 ();
 sg13g2_fill_2 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_418 ();
 sg13g2_decap_8 FILLER_28_425 ();
 sg13g2_decap_8 FILLER_28_432 ();
 sg13g2_fill_2 FILLER_28_439 ();
 sg13g2_fill_2 FILLER_28_467 ();
 sg13g2_decap_8 FILLER_28_505 ();
 sg13g2_decap_8 FILLER_28_512 ();
 sg13g2_fill_1 FILLER_28_626 ();
 sg13g2_decap_8 FILLER_28_647 ();
 sg13g2_fill_1 FILLER_28_654 ();
 sg13g2_fill_1 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_670 ();
 sg13g2_decap_4 FILLER_28_677 ();
 sg13g2_fill_2 FILLER_28_706 ();
 sg13g2_decap_4 FILLER_28_718 ();
 sg13g2_fill_2 FILLER_28_740 ();
 sg13g2_fill_1 FILLER_28_742 ();
 sg13g2_fill_1 FILLER_28_788 ();
 sg13g2_decap_8 FILLER_28_817 ();
 sg13g2_decap_8 FILLER_28_824 ();
 sg13g2_decap_8 FILLER_28_831 ();
 sg13g2_decap_8 FILLER_28_838 ();
 sg13g2_decap_8 FILLER_28_874 ();
 sg13g2_decap_8 FILLER_28_881 ();
 sg13g2_decap_8 FILLER_28_888 ();
 sg13g2_decap_8 FILLER_28_895 ();
 sg13g2_fill_2 FILLER_28_931 ();
 sg13g2_fill_1 FILLER_28_933 ();
 sg13g2_decap_8 FILLER_28_951 ();
 sg13g2_fill_2 FILLER_28_958 ();
 sg13g2_fill_1 FILLER_28_960 ();
 sg13g2_fill_2 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1051 ();
 sg13g2_decap_8 FILLER_28_1058 ();
 sg13g2_decap_4 FILLER_28_1065 ();
 sg13g2_decap_8 FILLER_28_1157 ();
 sg13g2_fill_2 FILLER_28_1164 ();
 sg13g2_fill_1 FILLER_28_1193 ();
 sg13g2_decap_8 FILLER_28_1238 ();
 sg13g2_fill_1 FILLER_28_1259 ();
 sg13g2_decap_8 FILLER_28_1269 ();
 sg13g2_decap_8 FILLER_28_1276 ();
 sg13g2_fill_2 FILLER_28_1283 ();
 sg13g2_decap_8 FILLER_28_1356 ();
 sg13g2_decap_8 FILLER_28_1363 ();
 sg13g2_decap_4 FILLER_28_1370 ();
 sg13g2_fill_1 FILLER_28_1374 ();
 sg13g2_decap_8 FILLER_28_1397 ();
 sg13g2_decap_8 FILLER_28_1404 ();
 sg13g2_decap_8 FILLER_28_1411 ();
 sg13g2_fill_2 FILLER_28_1418 ();
 sg13g2_fill_1 FILLER_28_1420 ();
 sg13g2_decap_8 FILLER_28_1431 ();
 sg13g2_decap_8 FILLER_28_1438 ();
 sg13g2_decap_4 FILLER_28_1445 ();
 sg13g2_decap_8 FILLER_28_1495 ();
 sg13g2_decap_8 FILLER_28_1502 ();
 sg13g2_decap_8 FILLER_28_1509 ();
 sg13g2_fill_2 FILLER_28_1516 ();
 sg13g2_fill_1 FILLER_28_1518 ();
 sg13g2_decap_8 FILLER_28_1532 ();
 sg13g2_decap_8 FILLER_28_1579 ();
 sg13g2_decap_8 FILLER_28_1586 ();
 sg13g2_fill_2 FILLER_28_1593 ();
 sg13g2_decap_4 FILLER_28_1625 ();
 sg13g2_fill_2 FILLER_28_1629 ();
 sg13g2_decap_8 FILLER_28_1644 ();
 sg13g2_fill_1 FILLER_28_1651 ();
 sg13g2_fill_1 FILLER_28_1679 ();
 sg13g2_decap_4 FILLER_28_1693 ();
 sg13g2_fill_2 FILLER_28_1697 ();
 sg13g2_decap_8 FILLER_28_1726 ();
 sg13g2_decap_4 FILLER_28_1733 ();
 sg13g2_fill_2 FILLER_28_1737 ();
 sg13g2_decap_8 FILLER_28_1793 ();
 sg13g2_decap_4 FILLER_28_1800 ();
 sg13g2_fill_2 FILLER_28_1804 ();
 sg13g2_decap_4 FILLER_28_1825 ();
 sg13g2_fill_1 FILLER_28_1829 ();
 sg13g2_fill_2 FILLER_28_1834 ();
 sg13g2_fill_1 FILLER_28_1836 ();
 sg13g2_decap_8 FILLER_28_1848 ();
 sg13g2_decap_8 FILLER_28_1855 ();
 sg13g2_decap_8 FILLER_28_1862 ();
 sg13g2_decap_8 FILLER_28_1869 ();
 sg13g2_decap_4 FILLER_28_1876 ();
 sg13g2_fill_2 FILLER_28_1880 ();
 sg13g2_decap_4 FILLER_28_1921 ();
 sg13g2_fill_2 FILLER_28_1925 ();
 sg13g2_decap_4 FILLER_28_1931 ();
 sg13g2_fill_1 FILLER_28_1935 ();
 sg13g2_fill_2 FILLER_28_1983 ();
 sg13g2_decap_8 FILLER_28_1993 ();
 sg13g2_decap_8 FILLER_28_2000 ();
 sg13g2_fill_1 FILLER_28_2019 ();
 sg13g2_decap_4 FILLER_28_2033 ();
 sg13g2_fill_1 FILLER_28_2037 ();
 sg13g2_decap_8 FILLER_28_2065 ();
 sg13g2_decap_8 FILLER_28_2072 ();
 sg13g2_decap_8 FILLER_28_2079 ();
 sg13g2_decap_8 FILLER_28_2086 ();
 sg13g2_decap_4 FILLER_28_2093 ();
 sg13g2_fill_2 FILLER_28_2102 ();
 sg13g2_decap_4 FILLER_28_2109 ();
 sg13g2_decap_8 FILLER_28_2128 ();
 sg13g2_fill_1 FILLER_28_2135 ();
 sg13g2_fill_2 FILLER_28_2154 ();
 sg13g2_fill_2 FILLER_28_2161 ();
 sg13g2_fill_2 FILLER_28_2168 ();
 sg13g2_fill_2 FILLER_28_2180 ();
 sg13g2_fill_1 FILLER_28_2182 ();
 sg13g2_decap_4 FILLER_28_2192 ();
 sg13g2_fill_1 FILLER_28_2196 ();
 sg13g2_decap_8 FILLER_28_2222 ();
 sg13g2_decap_8 FILLER_28_2229 ();
 sg13g2_decap_8 FILLER_28_2236 ();
 sg13g2_decap_8 FILLER_28_2243 ();
 sg13g2_decap_4 FILLER_28_2250 ();
 sg13g2_fill_1 FILLER_28_2254 ();
 sg13g2_fill_2 FILLER_28_2315 ();
 sg13g2_fill_1 FILLER_28_2322 ();
 sg13g2_decap_8 FILLER_28_2369 ();
 sg13g2_fill_2 FILLER_28_2376 ();
 sg13g2_decap_4 FILLER_28_2405 ();
 sg13g2_fill_2 FILLER_28_2473 ();
 sg13g2_fill_1 FILLER_28_2475 ();
 sg13g2_decap_8 FILLER_28_2485 ();
 sg13g2_decap_8 FILLER_28_2492 ();
 sg13g2_decap_8 FILLER_28_2499 ();
 sg13g2_decap_8 FILLER_28_2506 ();
 sg13g2_decap_8 FILLER_28_2513 ();
 sg13g2_decap_8 FILLER_28_2520 ();
 sg13g2_fill_1 FILLER_28_2536 ();
 sg13g2_fill_1 FILLER_28_2554 ();
 sg13g2_decap_8 FILLER_28_2585 ();
 sg13g2_fill_2 FILLER_28_2592 ();
 sg13g2_fill_1 FILLER_28_2594 ();
 sg13g2_fill_2 FILLER_28_2612 ();
 sg13g2_decap_4 FILLER_28_2659 ();
 sg13g2_fill_2 FILLER_28_2663 ();
 sg13g2_fill_1 FILLER_28_2696 ();
 sg13g2_decap_8 FILLER_28_2734 ();
 sg13g2_decap_8 FILLER_28_2767 ();
 sg13g2_decap_4 FILLER_28_2774 ();
 sg13g2_fill_1 FILLER_28_2778 ();
 sg13g2_decap_8 FILLER_28_2789 ();
 sg13g2_fill_1 FILLER_28_2796 ();
 sg13g2_fill_2 FILLER_28_2820 ();
 sg13g2_fill_1 FILLER_28_2822 ();
 sg13g2_decap_8 FILLER_28_2827 ();
 sg13g2_fill_1 FILLER_28_2834 ();
 sg13g2_decap_8 FILLER_28_2844 ();
 sg13g2_decap_4 FILLER_28_2861 ();
 sg13g2_fill_1 FILLER_28_2865 ();
 sg13g2_fill_2 FILLER_28_2875 ();
 sg13g2_decap_8 FILLER_28_2887 ();
 sg13g2_fill_2 FILLER_28_2894 ();
 sg13g2_decap_8 FILLER_28_2909 ();
 sg13g2_decap_8 FILLER_28_2916 ();
 sg13g2_decap_8 FILLER_28_2923 ();
 sg13g2_decap_8 FILLER_28_2930 ();
 sg13g2_fill_2 FILLER_28_2964 ();
 sg13g2_decap_8 FILLER_28_2992 ();
 sg13g2_decap_8 FILLER_28_2999 ();
 sg13g2_fill_1 FILLER_28_3038 ();
 sg13g2_decap_8 FILLER_28_3062 ();
 sg13g2_decap_8 FILLER_28_3069 ();
 sg13g2_decap_8 FILLER_28_3076 ();
 sg13g2_fill_2 FILLER_28_3083 ();
 sg13g2_decap_8 FILLER_28_3094 ();
 sg13g2_fill_2 FILLER_28_3159 ();
 sg13g2_decap_8 FILLER_28_3202 ();
 sg13g2_fill_2 FILLER_28_3209 ();
 sg13g2_fill_1 FILLER_28_3224 ();
 sg13g2_decap_8 FILLER_28_3252 ();
 sg13g2_decap_8 FILLER_28_3259 ();
 sg13g2_decap_8 FILLER_28_3266 ();
 sg13g2_fill_2 FILLER_28_3273 ();
 sg13g2_decap_8 FILLER_28_3327 ();
 sg13g2_fill_2 FILLER_28_3334 ();
 sg13g2_fill_2 FILLER_28_3350 ();
 sg13g2_fill_2 FILLER_28_3356 ();
 sg13g2_decap_4 FILLER_28_3393 ();
 sg13g2_fill_2 FILLER_28_3397 ();
 sg13g2_decap_8 FILLER_28_3480 ();
 sg13g2_decap_4 FILLER_28_3487 ();
 sg13g2_fill_1 FILLER_28_3505 ();
 sg13g2_fill_2 FILLER_28_3519 ();
 sg13g2_decap_8 FILLER_28_3542 ();
 sg13g2_fill_1 FILLER_28_3549 ();
 sg13g2_decap_8 FILLER_28_3554 ();
 sg13g2_decap_8 FILLER_28_3561 ();
 sg13g2_decap_8 FILLER_28_3568 ();
 sg13g2_fill_2 FILLER_28_3575 ();
 sg13g2_fill_1 FILLER_28_3577 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_18 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_decap_8 FILLER_29_45 ();
 sg13g2_decap_8 FILLER_29_52 ();
 sg13g2_decap_8 FILLER_29_59 ();
 sg13g2_fill_2 FILLER_29_66 ();
 sg13g2_fill_2 FILLER_29_85 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_205 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_decap_4 FILLER_29_255 ();
 sg13g2_fill_2 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_321 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_fill_2 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_decap_8 FILLER_29_416 ();
 sg13g2_decap_8 FILLER_29_423 ();
 sg13g2_decap_8 FILLER_29_430 ();
 sg13g2_decap_8 FILLER_29_437 ();
 sg13g2_fill_1 FILLER_29_444 ();
 sg13g2_decap_4 FILLER_29_455 ();
 sg13g2_fill_1 FILLER_29_472 ();
 sg13g2_decap_8 FILLER_29_506 ();
 sg13g2_decap_8 FILLER_29_513 ();
 sg13g2_decap_8 FILLER_29_520 ();
 sg13g2_fill_2 FILLER_29_572 ();
 sg13g2_fill_1 FILLER_29_592 ();
 sg13g2_fill_1 FILLER_29_599 ();
 sg13g2_fill_2 FILLER_29_614 ();
 sg13g2_fill_1 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_648 ();
 sg13g2_decap_4 FILLER_29_655 ();
 sg13g2_fill_2 FILLER_29_659 ();
 sg13g2_fill_2 FILLER_29_664 ();
 sg13g2_fill_2 FILLER_29_694 ();
 sg13g2_decap_8 FILLER_29_701 ();
 sg13g2_fill_2 FILLER_29_708 ();
 sg13g2_fill_1 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_724 ();
 sg13g2_decap_4 FILLER_29_731 ();
 sg13g2_fill_2 FILLER_29_748 ();
 sg13g2_fill_1 FILLER_29_750 ();
 sg13g2_decap_8 FILLER_29_773 ();
 sg13g2_decap_4 FILLER_29_780 ();
 sg13g2_decap_8 FILLER_29_824 ();
 sg13g2_decap_8 FILLER_29_831 ();
 sg13g2_decap_8 FILLER_29_838 ();
 sg13g2_fill_2 FILLER_29_845 ();
 sg13g2_fill_2 FILLER_29_873 ();
 sg13g2_fill_2 FILLER_29_880 ();
 sg13g2_fill_1 FILLER_29_887 ();
 sg13g2_fill_1 FILLER_29_892 ();
 sg13g2_decap_4 FILLER_29_903 ();
 sg13g2_fill_2 FILLER_29_907 ();
 sg13g2_decap_8 FILLER_29_945 ();
 sg13g2_decap_8 FILLER_29_952 ();
 sg13g2_fill_2 FILLER_29_994 ();
 sg13g2_fill_1 FILLER_29_1001 ();
 sg13g2_decap_4 FILLER_29_1038 ();
 sg13g2_fill_1 FILLER_29_1042 ();
 sg13g2_decap_8 FILLER_29_1052 ();
 sg13g2_decap_8 FILLER_29_1059 ();
 sg13g2_fill_2 FILLER_29_1098 ();
 sg13g2_fill_1 FILLER_29_1100 ();
 sg13g2_decap_4 FILLER_29_1123 ();
 sg13g2_fill_2 FILLER_29_1127 ();
 sg13g2_fill_1 FILLER_29_1144 ();
 sg13g2_decap_8 FILLER_29_1148 ();
 sg13g2_decap_4 FILLER_29_1155 ();
 sg13g2_fill_2 FILLER_29_1159 ();
 sg13g2_fill_2 FILLER_29_1188 ();
 sg13g2_fill_1 FILLER_29_1190 ();
 sg13g2_decap_4 FILLER_29_1214 ();
 sg13g2_fill_2 FILLER_29_1218 ();
 sg13g2_decap_8 FILLER_29_1229 ();
 sg13g2_decap_8 FILLER_29_1236 ();
 sg13g2_decap_4 FILLER_29_1243 ();
 sg13g2_decap_8 FILLER_29_1275 ();
 sg13g2_decap_8 FILLER_29_1282 ();
 sg13g2_decap_8 FILLER_29_1289 ();
 sg13g2_fill_1 FILLER_29_1296 ();
 sg13g2_fill_1 FILLER_29_1343 ();
 sg13g2_decap_8 FILLER_29_1359 ();
 sg13g2_decap_8 FILLER_29_1366 ();
 sg13g2_decap_4 FILLER_29_1410 ();
 sg13g2_fill_1 FILLER_29_1414 ();
 sg13g2_fill_2 FILLER_29_1436 ();
 sg13g2_fill_1 FILLER_29_1438 ();
 sg13g2_decap_8 FILLER_29_1444 ();
 sg13g2_decap_8 FILLER_29_1451 ();
 sg13g2_fill_1 FILLER_29_1495 ();
 sg13g2_fill_2 FILLER_29_1504 ();
 sg13g2_decap_8 FILLER_29_1532 ();
 sg13g2_fill_2 FILLER_29_1539 ();
 sg13g2_fill_1 FILLER_29_1541 ();
 sg13g2_fill_2 FILLER_29_1561 ();
 sg13g2_fill_1 FILLER_29_1563 ();
 sg13g2_decap_8 FILLER_29_1586 ();
 sg13g2_decap_4 FILLER_29_1593 ();
 sg13g2_fill_1 FILLER_29_1597 ();
 sg13g2_fill_2 FILLER_29_1634 ();
 sg13g2_fill_1 FILLER_29_1636 ();
 sg13g2_decap_8 FILLER_29_1656 ();
 sg13g2_decap_8 FILLER_29_1676 ();
 sg13g2_fill_2 FILLER_29_1683 ();
 sg13g2_fill_1 FILLER_29_1685 ();
 sg13g2_decap_8 FILLER_29_1695 ();
 sg13g2_fill_2 FILLER_29_1702 ();
 sg13g2_fill_2 FILLER_29_1714 ();
 sg13g2_fill_1 FILLER_29_1716 ();
 sg13g2_decap_8 FILLER_29_1733 ();
 sg13g2_decap_8 FILLER_29_1740 ();
 sg13g2_decap_8 FILLER_29_1747 ();
 sg13g2_decap_4 FILLER_29_1754 ();
 sg13g2_fill_2 FILLER_29_1758 ();
 sg13g2_fill_1 FILLER_29_1764 ();
 sg13g2_decap_8 FILLER_29_1807 ();
 sg13g2_decap_8 FILLER_29_1814 ();
 sg13g2_decap_8 FILLER_29_1821 ();
 sg13g2_fill_2 FILLER_29_1828 ();
 sg13g2_decap_8 FILLER_29_1861 ();
 sg13g2_decap_8 FILLER_29_1868 ();
 sg13g2_decap_8 FILLER_29_1875 ();
 sg13g2_decap_8 FILLER_29_1882 ();
 sg13g2_decap_4 FILLER_29_1889 ();
 sg13g2_decap_8 FILLER_29_1931 ();
 sg13g2_decap_4 FILLER_29_1938 ();
 sg13g2_fill_1 FILLER_29_1942 ();
 sg13g2_decap_8 FILLER_29_1958 ();
 sg13g2_decap_8 FILLER_29_1965 ();
 sg13g2_decap_8 FILLER_29_1972 ();
 sg13g2_fill_1 FILLER_29_1979 ();
 sg13g2_decap_4 FILLER_29_1984 ();
 sg13g2_decap_4 FILLER_29_1992 ();
 sg13g2_fill_2 FILLER_29_1996 ();
 sg13g2_fill_2 FILLER_29_2003 ();
 sg13g2_decap_8 FILLER_29_2013 ();
 sg13g2_decap_8 FILLER_29_2020 ();
 sg13g2_decap_4 FILLER_29_2027 ();
 sg13g2_fill_2 FILLER_29_2031 ();
 sg13g2_fill_1 FILLER_29_2056 ();
 sg13g2_decap_8 FILLER_29_2071 ();
 sg13g2_decap_8 FILLER_29_2078 ();
 sg13g2_decap_8 FILLER_29_2085 ();
 sg13g2_decap_8 FILLER_29_2092 ();
 sg13g2_fill_1 FILLER_29_2099 ();
 sg13g2_fill_1 FILLER_29_2117 ();
 sg13g2_decap_4 FILLER_29_2144 ();
 sg13g2_decap_8 FILLER_29_2163 ();
 sg13g2_fill_2 FILLER_29_2170 ();
 sg13g2_fill_2 FILLER_29_2177 ();
 sg13g2_fill_1 FILLER_29_2179 ();
 sg13g2_decap_8 FILLER_29_2185 ();
 sg13g2_fill_1 FILLER_29_2192 ();
 sg13g2_fill_1 FILLER_29_2198 ();
 sg13g2_decap_4 FILLER_29_2223 ();
 sg13g2_fill_1 FILLER_29_2227 ();
 sg13g2_fill_2 FILLER_29_2232 ();
 sg13g2_fill_1 FILLER_29_2234 ();
 sg13g2_fill_1 FILLER_29_2325 ();
 sg13g2_decap_8 FILLER_29_2353 ();
 sg13g2_fill_1 FILLER_29_2360 ();
 sg13g2_decap_8 FILLER_29_2374 ();
 sg13g2_fill_2 FILLER_29_2381 ();
 sg13g2_fill_1 FILLER_29_2383 ();
 sg13g2_fill_1 FILLER_29_2439 ();
 sg13g2_decap_8 FILLER_29_2453 ();
 sg13g2_decap_4 FILLER_29_2469 ();
 sg13g2_decap_8 FILLER_29_2481 ();
 sg13g2_decap_8 FILLER_29_2488 ();
 sg13g2_decap_8 FILLER_29_2495 ();
 sg13g2_decap_8 FILLER_29_2502 ();
 sg13g2_decap_8 FILLER_29_2509 ();
 sg13g2_fill_1 FILLER_29_2516 ();
 sg13g2_decap_8 FILLER_29_2526 ();
 sg13g2_fill_2 FILLER_29_2533 ();
 sg13g2_fill_2 FILLER_29_2545 ();
 sg13g2_decap_8 FILLER_29_2556 ();
 sg13g2_decap_4 FILLER_29_2563 ();
 sg13g2_fill_2 FILLER_29_2567 ();
 sg13g2_decap_8 FILLER_29_2582 ();
 sg13g2_decap_8 FILLER_29_2589 ();
 sg13g2_decap_8 FILLER_29_2596 ();
 sg13g2_decap_8 FILLER_29_2603 ();
 sg13g2_decap_8 FILLER_29_2610 ();
 sg13g2_decap_4 FILLER_29_2617 ();
 sg13g2_fill_1 FILLER_29_2621 ();
 sg13g2_decap_8 FILLER_29_2649 ();
 sg13g2_decap_8 FILLER_29_2656 ();
 sg13g2_decap_4 FILLER_29_2663 ();
 sg13g2_fill_1 FILLER_29_2667 ();
 sg13g2_fill_2 FILLER_29_2678 ();
 sg13g2_fill_1 FILLER_29_2699 ();
 sg13g2_fill_2 FILLER_29_2710 ();
 sg13g2_fill_1 FILLER_29_2712 ();
 sg13g2_decap_8 FILLER_29_2735 ();
 sg13g2_decap_4 FILLER_29_2742 ();
 sg13g2_decap_4 FILLER_29_2759 ();
 sg13g2_fill_1 FILLER_29_2763 ();
 sg13g2_fill_1 FILLER_29_2791 ();
 sg13g2_decap_8 FILLER_29_2832 ();
 sg13g2_decap_4 FILLER_29_2839 ();
 sg13g2_fill_2 FILLER_29_2843 ();
 sg13g2_fill_2 FILLER_29_2881 ();
 sg13g2_decap_8 FILLER_29_2919 ();
 sg13g2_decap_8 FILLER_29_2926 ();
 sg13g2_decap_8 FILLER_29_2933 ();
 sg13g2_fill_1 FILLER_29_2940 ();
 sg13g2_decap_8 FILLER_29_2972 ();
 sg13g2_decap_8 FILLER_29_2979 ();
 sg13g2_decap_8 FILLER_29_2986 ();
 sg13g2_decap_4 FILLER_29_2993 ();
 sg13g2_fill_2 FILLER_29_3001 ();
 sg13g2_fill_1 FILLER_29_3003 ();
 sg13g2_fill_1 FILLER_29_3041 ();
 sg13g2_decap_4 FILLER_29_3096 ();
 sg13g2_fill_1 FILLER_29_3100 ();
 sg13g2_fill_1 FILLER_29_3141 ();
 sg13g2_decap_4 FILLER_29_3191 ();
 sg13g2_fill_2 FILLER_29_3195 ();
 sg13g2_decap_8 FILLER_29_3206 ();
 sg13g2_fill_2 FILLER_29_3213 ();
 sg13g2_decap_8 FILLER_29_3261 ();
 sg13g2_decap_8 FILLER_29_3268 ();
 sg13g2_decap_8 FILLER_29_3275 ();
 sg13g2_fill_1 FILLER_29_3282 ();
 sg13g2_fill_1 FILLER_29_3322 ();
 sg13g2_decap_8 FILLER_29_3332 ();
 sg13g2_decap_4 FILLER_29_3339 ();
 sg13g2_decap_8 FILLER_29_3393 ();
 sg13g2_decap_4 FILLER_29_3400 ();
 sg13g2_fill_2 FILLER_29_3404 ();
 sg13g2_decap_4 FILLER_29_3416 ();
 sg13g2_decap_4 FILLER_29_3429 ();
 sg13g2_fill_1 FILLER_29_3433 ();
 sg13g2_decap_8 FILLER_29_3485 ();
 sg13g2_fill_2 FILLER_29_3515 ();
 sg13g2_fill_2 FILLER_29_3547 ();
 sg13g2_fill_1 FILLER_29_3549 ();
 sg13g2_decap_8 FILLER_29_3558 ();
 sg13g2_decap_8 FILLER_29_3565 ();
 sg13g2_decap_4 FILLER_29_3572 ();
 sg13g2_fill_2 FILLER_29_3576 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_18 ();
 sg13g2_fill_2 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_31 ();
 sg13g2_decap_8 FILLER_30_53 ();
 sg13g2_decap_8 FILLER_30_60 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_decap_8 FILLER_30_114 ();
 sg13g2_decap_8 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_190 ();
 sg13g2_decap_8 FILLER_30_197 ();
 sg13g2_decap_8 FILLER_30_204 ();
 sg13g2_decap_8 FILLER_30_211 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_decap_8 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_decap_4 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_fill_2 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_fill_2 FILLER_30_333 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_fill_1 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_8 FILLER_30_424 ();
 sg13g2_decap_8 FILLER_30_431 ();
 sg13g2_decap_4 FILLER_30_438 ();
 sg13g2_fill_2 FILLER_30_442 ();
 sg13g2_fill_1 FILLER_30_472 ();
 sg13g2_fill_2 FILLER_30_486 ();
 sg13g2_decap_8 FILLER_30_506 ();
 sg13g2_decap_8 FILLER_30_513 ();
 sg13g2_decap_4 FILLER_30_520 ();
 sg13g2_fill_1 FILLER_30_524 ();
 sg13g2_fill_2 FILLER_30_538 ();
 sg13g2_fill_1 FILLER_30_540 ();
 sg13g2_fill_1 FILLER_30_589 ();
 sg13g2_decap_4 FILLER_30_599 ();
 sg13g2_fill_2 FILLER_30_613 ();
 sg13g2_fill_1 FILLER_30_615 ();
 sg13g2_decap_4 FILLER_30_621 ();
 sg13g2_fill_2 FILLER_30_625 ();
 sg13g2_fill_1 FILLER_30_632 ();
 sg13g2_decap_8 FILLER_30_641 ();
 sg13g2_decap_4 FILLER_30_648 ();
 sg13g2_fill_2 FILLER_30_665 ();
 sg13g2_fill_1 FILLER_30_667 ();
 sg13g2_fill_2 FILLER_30_681 ();
 sg13g2_decap_8 FILLER_30_696 ();
 sg13g2_decap_4 FILLER_30_707 ();
 sg13g2_fill_1 FILLER_30_711 ();
 sg13g2_fill_2 FILLER_30_716 ();
 sg13g2_fill_1 FILLER_30_718 ();
 sg13g2_decap_8 FILLER_30_732 ();
 sg13g2_decap_8 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_fill_2 FILLER_30_781 ();
 sg13g2_fill_1 FILLER_30_783 ();
 sg13g2_fill_2 FILLER_30_819 ();
 sg13g2_fill_1 FILLER_30_821 ();
 sg13g2_decap_4 FILLER_30_836 ();
 sg13g2_fill_2 FILLER_30_840 ();
 sg13g2_decap_4 FILLER_30_875 ();
 sg13g2_fill_1 FILLER_30_879 ();
 sg13g2_fill_2 FILLER_30_896 ();
 sg13g2_fill_1 FILLER_30_898 ();
 sg13g2_decap_4 FILLER_30_904 ();
 sg13g2_fill_2 FILLER_30_913 ();
 sg13g2_fill_1 FILLER_30_930 ();
 sg13g2_decap_8 FILLER_30_935 ();
 sg13g2_decap_8 FILLER_30_942 ();
 sg13g2_decap_4 FILLER_30_949 ();
 sg13g2_fill_1 FILLER_30_953 ();
 sg13g2_decap_8 FILLER_30_958 ();
 sg13g2_fill_2 FILLER_30_965 ();
 sg13g2_fill_2 FILLER_30_989 ();
 sg13g2_fill_1 FILLER_30_995 ();
 sg13g2_fill_2 FILLER_30_1000 ();
 sg13g2_fill_1 FILLER_30_1002 ();
 sg13g2_decap_4 FILLER_30_1012 ();
 sg13g2_decap_8 FILLER_30_1025 ();
 sg13g2_decap_8 FILLER_30_1032 ();
 sg13g2_decap_8 FILLER_30_1039 ();
 sg13g2_decap_8 FILLER_30_1046 ();
 sg13g2_decap_8 FILLER_30_1053 ();
 sg13g2_fill_2 FILLER_30_1060 ();
 sg13g2_fill_1 FILLER_30_1062 ();
 sg13g2_fill_1 FILLER_30_1091 ();
 sg13g2_fill_1 FILLER_30_1113 ();
 sg13g2_decap_8 FILLER_30_1127 ();
 sg13g2_decap_8 FILLER_30_1134 ();
 sg13g2_decap_8 FILLER_30_1141 ();
 sg13g2_fill_2 FILLER_30_1148 ();
 sg13g2_fill_1 FILLER_30_1150 ();
 sg13g2_fill_1 FILLER_30_1179 ();
 sg13g2_fill_2 FILLER_30_1194 ();
 sg13g2_decap_4 FILLER_30_1210 ();
 sg13g2_fill_1 FILLER_30_1214 ();
 sg13g2_decap_8 FILLER_30_1230 ();
 sg13g2_decap_8 FILLER_30_1285 ();
 sg13g2_fill_1 FILLER_30_1292 ();
 sg13g2_decap_4 FILLER_30_1303 ();
 sg13g2_fill_2 FILLER_30_1330 ();
 sg13g2_fill_1 FILLER_30_1332 ();
 sg13g2_fill_1 FILLER_30_1353 ();
 sg13g2_decap_8 FILLER_30_1359 ();
 sg13g2_decap_8 FILLER_30_1366 ();
 sg13g2_decap_8 FILLER_30_1373 ();
 sg13g2_decap_8 FILLER_30_1386 ();
 sg13g2_decap_8 FILLER_30_1393 ();
 sg13g2_fill_2 FILLER_30_1400 ();
 sg13g2_decap_4 FILLER_30_1437 ();
 sg13g2_fill_1 FILLER_30_1441 ();
 sg13g2_decap_8 FILLER_30_1450 ();
 sg13g2_decap_8 FILLER_30_1457 ();
 sg13g2_decap_4 FILLER_30_1464 ();
 sg13g2_fill_1 FILLER_30_1468 ();
 sg13g2_decap_8 FILLER_30_1508 ();
 sg13g2_decap_8 FILLER_30_1515 ();
 sg13g2_decap_8 FILLER_30_1522 ();
 sg13g2_decap_8 FILLER_30_1529 ();
 sg13g2_decap_8 FILLER_30_1536 ();
 sg13g2_fill_2 FILLER_30_1553 ();
 sg13g2_fill_1 FILLER_30_1555 ();
 sg13g2_fill_2 FILLER_30_1571 ();
 sg13g2_fill_1 FILLER_30_1573 ();
 sg13g2_decap_4 FILLER_30_1624 ();
 sg13g2_fill_2 FILLER_30_1628 ();
 sg13g2_fill_2 FILLER_30_1648 ();
 sg13g2_decap_8 FILLER_30_1655 ();
 sg13g2_fill_1 FILLER_30_1676 ();
 sg13g2_decap_8 FILLER_30_1682 ();
 sg13g2_fill_2 FILLER_30_1689 ();
 sg13g2_decap_8 FILLER_30_1706 ();
 sg13g2_fill_1 FILLER_30_1718 ();
 sg13g2_fill_1 FILLER_30_1724 ();
 sg13g2_decap_8 FILLER_30_1731 ();
 sg13g2_decap_8 FILLER_30_1738 ();
 sg13g2_decap_4 FILLER_30_1745 ();
 sg13g2_fill_2 FILLER_30_1749 ();
 sg13g2_fill_1 FILLER_30_1790 ();
 sg13g2_decap_4 FILLER_30_1816 ();
 sg13g2_fill_1 FILLER_30_1820 ();
 sg13g2_decap_8 FILLER_30_1853 ();
 sg13g2_decap_8 FILLER_30_1860 ();
 sg13g2_decap_8 FILLER_30_1867 ();
 sg13g2_decap_8 FILLER_30_1874 ();
 sg13g2_decap_8 FILLER_30_1881 ();
 sg13g2_decap_4 FILLER_30_1888 ();
 sg13g2_fill_1 FILLER_30_1892 ();
 sg13g2_fill_2 FILLER_30_1903 ();
 sg13g2_decap_8 FILLER_30_1916 ();
 sg13g2_decap_8 FILLER_30_1923 ();
 sg13g2_decap_8 FILLER_30_1930 ();
 sg13g2_decap_4 FILLER_30_1937 ();
 sg13g2_fill_2 FILLER_30_1959 ();
 sg13g2_fill_1 FILLER_30_1961 ();
 sg13g2_fill_2 FILLER_30_1989 ();
 sg13g2_fill_1 FILLER_30_1991 ();
 sg13g2_fill_2 FILLER_30_1997 ();
 sg13g2_decap_8 FILLER_30_2020 ();
 sg13g2_decap_4 FILLER_30_2027 ();
 sg13g2_fill_1 FILLER_30_2031 ();
 sg13g2_decap_4 FILLER_30_2061 ();
 sg13g2_decap_4 FILLER_30_2070 ();
 sg13g2_decap_8 FILLER_30_2079 ();
 sg13g2_fill_2 FILLER_30_2086 ();
 sg13g2_fill_1 FILLER_30_2088 ();
 sg13g2_fill_1 FILLER_30_2094 ();
 sg13g2_fill_1 FILLER_30_2108 ();
 sg13g2_decap_8 FILLER_30_2126 ();
 sg13g2_decap_4 FILLER_30_2133 ();
 sg13g2_decap_8 FILLER_30_2142 ();
 sg13g2_decap_4 FILLER_30_2149 ();
 sg13g2_fill_1 FILLER_30_2153 ();
 sg13g2_decap_8 FILLER_30_2159 ();
 sg13g2_fill_2 FILLER_30_2176 ();
 sg13g2_decap_4 FILLER_30_2203 ();
 sg13g2_fill_2 FILLER_30_2233 ();
 sg13g2_fill_1 FILLER_30_2235 ();
 sg13g2_fill_1 FILLER_30_2245 ();
 sg13g2_decap_8 FILLER_30_2255 ();
 sg13g2_decap_4 FILLER_30_2262 ();
 sg13g2_fill_2 FILLER_30_2266 ();
 sg13g2_fill_1 FILLER_30_2272 ();
 sg13g2_fill_1 FILLER_30_2297 ();
 sg13g2_decap_8 FILLER_30_2353 ();
 sg13g2_decap_8 FILLER_30_2360 ();
 sg13g2_decap_8 FILLER_30_2367 ();
 sg13g2_decap_8 FILLER_30_2374 ();
 sg13g2_decap_8 FILLER_30_2381 ();
 sg13g2_fill_2 FILLER_30_2388 ();
 sg13g2_fill_1 FILLER_30_2390 ();
 sg13g2_decap_8 FILLER_30_2404 ();
 sg13g2_fill_1 FILLER_30_2420 ();
 sg13g2_decap_8 FILLER_30_2434 ();
 sg13g2_decap_8 FILLER_30_2441 ();
 sg13g2_decap_8 FILLER_30_2448 ();
 sg13g2_decap_8 FILLER_30_2455 ();
 sg13g2_decap_8 FILLER_30_2462 ();
 sg13g2_decap_8 FILLER_30_2469 ();
 sg13g2_decap_8 FILLER_30_2476 ();
 sg13g2_decap_8 FILLER_30_2483 ();
 sg13g2_decap_8 FILLER_30_2490 ();
 sg13g2_fill_2 FILLER_30_2497 ();
 sg13g2_decap_8 FILLER_30_2536 ();
 sg13g2_fill_1 FILLER_30_2543 ();
 sg13g2_decap_8 FILLER_30_2557 ();
 sg13g2_decap_8 FILLER_30_2564 ();
 sg13g2_decap_4 FILLER_30_2571 ();
 sg13g2_fill_2 FILLER_30_2575 ();
 sg13g2_decap_8 FILLER_30_2604 ();
 sg13g2_decap_8 FILLER_30_2611 ();
 sg13g2_decap_8 FILLER_30_2618 ();
 sg13g2_fill_2 FILLER_30_2625 ();
 sg13g2_fill_1 FILLER_30_2627 ();
 sg13g2_decap_8 FILLER_30_2632 ();
 sg13g2_decap_8 FILLER_30_2639 ();
 sg13g2_decap_8 FILLER_30_2646 ();
 sg13g2_decap_8 FILLER_30_2653 ();
 sg13g2_decap_8 FILLER_30_2660 ();
 sg13g2_fill_2 FILLER_30_2667 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_decap_4 FILLER_30_2680 ();
 sg13g2_fill_1 FILLER_30_2684 ();
 sg13g2_decap_8 FILLER_30_2703 ();
 sg13g2_decap_8 FILLER_30_2710 ();
 sg13g2_decap_8 FILLER_30_2721 ();
 sg13g2_decap_8 FILLER_30_2728 ();
 sg13g2_decap_4 FILLER_30_2745 ();
 sg13g2_fill_2 FILLER_30_2758 ();
 sg13g2_decap_8 FILLER_30_2773 ();
 sg13g2_fill_1 FILLER_30_2780 ();
 sg13g2_decap_8 FILLER_30_2832 ();
 sg13g2_decap_8 FILLER_30_2839 ();
 sg13g2_fill_2 FILLER_30_2907 ();
 sg13g2_decap_8 FILLER_30_2944 ();
 sg13g2_decap_8 FILLER_30_2955 ();
 sg13g2_decap_8 FILLER_30_2975 ();
 sg13g2_decap_8 FILLER_30_2982 ();
 sg13g2_fill_2 FILLER_30_2989 ();
 sg13g2_fill_1 FILLER_30_2991 ();
 sg13g2_decap_8 FILLER_30_3055 ();
 sg13g2_decap_4 FILLER_30_3062 ();
 sg13g2_fill_2 FILLER_30_3080 ();
 sg13g2_fill_1 FILLER_30_3082 ();
 sg13g2_decap_8 FILLER_30_3104 ();
 sg13g2_decap_8 FILLER_30_3111 ();
 sg13g2_decap_8 FILLER_30_3118 ();
 sg13g2_decap_8 FILLER_30_3125 ();
 sg13g2_decap_8 FILLER_30_3132 ();
 sg13g2_decap_8 FILLER_30_3139 ();
 sg13g2_fill_2 FILLER_30_3146 ();
 sg13g2_fill_2 FILLER_30_3175 ();
 sg13g2_decap_8 FILLER_30_3214 ();
 sg13g2_decap_8 FILLER_30_3221 ();
 sg13g2_fill_2 FILLER_30_3228 ();
 sg13g2_fill_2 FILLER_30_3234 ();
 sg13g2_decap_8 FILLER_30_3273 ();
 sg13g2_decap_8 FILLER_30_3280 ();
 sg13g2_fill_2 FILLER_30_3323 ();
 sg13g2_fill_1 FILLER_30_3325 ();
 sg13g2_decap_8 FILLER_30_3334 ();
 sg13g2_decap_8 FILLER_30_3341 ();
 sg13g2_fill_2 FILLER_30_3348 ();
 sg13g2_decap_8 FILLER_30_3385 ();
 sg13g2_decap_8 FILLER_30_3392 ();
 sg13g2_decap_8 FILLER_30_3399 ();
 sg13g2_fill_2 FILLER_30_3406 ();
 sg13g2_decap_4 FILLER_30_3439 ();
 sg13g2_fill_1 FILLER_30_3443 ();
 sg13g2_fill_2 FILLER_30_3461 ();
 sg13g2_fill_1 FILLER_30_3467 ();
 sg13g2_decap_4 FILLER_30_3481 ();
 sg13g2_fill_2 FILLER_30_3485 ();
 sg13g2_fill_1 FILLER_30_3500 ();
 sg13g2_fill_2 FILLER_30_3532 ();
 sg13g2_fill_1 FILLER_30_3534 ();
 sg13g2_decap_4 FILLER_30_3572 ();
 sg13g2_fill_2 FILLER_30_3576 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_decap_4 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_129 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_214 ();
 sg13g2_decap_4 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_333 ();
 sg13g2_decap_8 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_decap_8 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_31_436 ();
 sg13g2_fill_2 FILLER_31_443 ();
 sg13g2_decap_8 FILLER_31_460 ();
 sg13g2_decap_8 FILLER_31_467 ();
 sg13g2_decap_8 FILLER_31_474 ();
 sg13g2_decap_4 FILLER_31_481 ();
 sg13g2_fill_1 FILLER_31_485 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_4 FILLER_31_511 ();
 sg13g2_fill_2 FILLER_31_515 ();
 sg13g2_decap_4 FILLER_31_544 ();
 sg13g2_fill_2 FILLER_31_548 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_fill_2 FILLER_31_560 ();
 sg13g2_fill_1 FILLER_31_562 ();
 sg13g2_fill_1 FILLER_31_568 ();
 sg13g2_fill_2 FILLER_31_597 ();
 sg13g2_fill_2 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_625 ();
 sg13g2_decap_8 FILLER_31_636 ();
 sg13g2_fill_2 FILLER_31_643 ();
 sg13g2_fill_2 FILLER_31_668 ();
 sg13g2_decap_8 FILLER_31_683 ();
 sg13g2_fill_2 FILLER_31_690 ();
 sg13g2_fill_1 FILLER_31_692 ();
 sg13g2_fill_1 FILLER_31_703 ();
 sg13g2_decap_8 FILLER_31_751 ();
 sg13g2_fill_2 FILLER_31_758 ();
 sg13g2_fill_1 FILLER_31_760 ();
 sg13g2_decap_4 FILLER_31_774 ();
 sg13g2_decap_4 FILLER_31_789 ();
 sg13g2_fill_2 FILLER_31_793 ();
 sg13g2_fill_1 FILLER_31_835 ();
 sg13g2_decap_4 FILLER_31_886 ();
 sg13g2_fill_2 FILLER_31_890 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_fill_1 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_991 ();
 sg13g2_decap_8 FILLER_31_998 ();
 sg13g2_decap_8 FILLER_31_1005 ();
 sg13g2_decap_4 FILLER_31_1012 ();
 sg13g2_fill_1 FILLER_31_1016 ();
 sg13g2_decap_8 FILLER_31_1041 ();
 sg13g2_decap_8 FILLER_31_1048 ();
 sg13g2_decap_8 FILLER_31_1055 ();
 sg13g2_decap_4 FILLER_31_1062 ();
 sg13g2_fill_1 FILLER_31_1066 ();
 sg13g2_decap_4 FILLER_31_1076 ();
 sg13g2_fill_2 FILLER_31_1080 ();
 sg13g2_decap_8 FILLER_31_1123 ();
 sg13g2_decap_8 FILLER_31_1130 ();
 sg13g2_decap_8 FILLER_31_1137 ();
 sg13g2_decap_8 FILLER_31_1144 ();
 sg13g2_decap_8 FILLER_31_1151 ();
 sg13g2_fill_1 FILLER_31_1158 ();
 sg13g2_decap_8 FILLER_31_1200 ();
 sg13g2_decap_8 FILLER_31_1207 ();
 sg13g2_decap_4 FILLER_31_1214 ();
 sg13g2_fill_1 FILLER_31_1218 ();
 sg13g2_decap_8 FILLER_31_1229 ();
 sg13g2_decap_8 FILLER_31_1236 ();
 sg13g2_decap_8 FILLER_31_1243 ();
 sg13g2_decap_4 FILLER_31_1250 ();
 sg13g2_fill_1 FILLER_31_1254 ();
 sg13g2_fill_2 FILLER_31_1268 ();
 sg13g2_fill_2 FILLER_31_1278 ();
 sg13g2_decap_8 FILLER_31_1289 ();
 sg13g2_decap_4 FILLER_31_1296 ();
 sg13g2_fill_1 FILLER_31_1312 ();
 sg13g2_fill_1 FILLER_31_1324 ();
 sg13g2_decap_4 FILLER_31_1349 ();
 sg13g2_decap_8 FILLER_31_1358 ();
 sg13g2_decap_8 FILLER_31_1365 ();
 sg13g2_decap_8 FILLER_31_1372 ();
 sg13g2_decap_8 FILLER_31_1379 ();
 sg13g2_decap_8 FILLER_31_1386 ();
 sg13g2_decap_8 FILLER_31_1393 ();
 sg13g2_decap_4 FILLER_31_1404 ();
 sg13g2_fill_2 FILLER_31_1408 ();
 sg13g2_fill_1 FILLER_31_1436 ();
 sg13g2_fill_1 FILLER_31_1455 ();
 sg13g2_fill_2 FILLER_31_1472 ();
 sg13g2_fill_2 FILLER_31_1491 ();
 sg13g2_fill_1 FILLER_31_1493 ();
 sg13g2_fill_2 FILLER_31_1599 ();
 sg13g2_fill_1 FILLER_31_1601 ();
 sg13g2_fill_2 FILLER_31_1647 ();
 sg13g2_fill_1 FILLER_31_1649 ();
 sg13g2_fill_2 FILLER_31_1655 ();
 sg13g2_fill_2 FILLER_31_1662 ();
 sg13g2_fill_1 FILLER_31_1664 ();
 sg13g2_decap_8 FILLER_31_1680 ();
 sg13g2_decap_4 FILLER_31_1687 ();
 sg13g2_fill_1 FILLER_31_1691 ();
 sg13g2_decap_4 FILLER_31_1701 ();
 sg13g2_decap_8 FILLER_31_1735 ();
 sg13g2_decap_8 FILLER_31_1742 ();
 sg13g2_decap_4 FILLER_31_1749 ();
 sg13g2_fill_2 FILLER_31_1753 ();
 sg13g2_fill_2 FILLER_31_1764 ();
 sg13g2_fill_1 FILLER_31_1771 ();
 sg13g2_decap_8 FILLER_31_1849 ();
 sg13g2_decap_8 FILLER_31_1856 ();
 sg13g2_decap_4 FILLER_31_1863 ();
 sg13g2_fill_2 FILLER_31_1867 ();
 sg13g2_fill_1 FILLER_31_1910 ();
 sg13g2_decap_8 FILLER_31_1921 ();
 sg13g2_decap_8 FILLER_31_1928 ();
 sg13g2_decap_8 FILLER_31_1935 ();
 sg13g2_fill_2 FILLER_31_1942 ();
 sg13g2_decap_8 FILLER_31_1949 ();
 sg13g2_fill_2 FILLER_31_1969 ();
 sg13g2_fill_2 FILLER_31_2021 ();
 sg13g2_fill_2 FILLER_31_2027 ();
 sg13g2_decap_4 FILLER_31_2063 ();
 sg13g2_fill_1 FILLER_31_2067 ();
 sg13g2_fill_2 FILLER_31_2074 ();
 sg13g2_fill_1 FILLER_31_2115 ();
 sg13g2_decap_8 FILLER_31_2134 ();
 sg13g2_decap_8 FILLER_31_2141 ();
 sg13g2_fill_1 FILLER_31_2174 ();
 sg13g2_fill_1 FILLER_31_2180 ();
 sg13g2_decap_8 FILLER_31_2194 ();
 sg13g2_decap_8 FILLER_31_2201 ();
 sg13g2_fill_2 FILLER_31_2208 ();
 sg13g2_fill_1 FILLER_31_2210 ();
 sg13g2_decap_4 FILLER_31_2229 ();
 sg13g2_decap_4 FILLER_31_2238 ();
 sg13g2_fill_1 FILLER_31_2242 ();
 sg13g2_decap_8 FILLER_31_2247 ();
 sg13g2_decap_8 FILLER_31_2254 ();
 sg13g2_decap_8 FILLER_31_2261 ();
 sg13g2_decap_8 FILLER_31_2268 ();
 sg13g2_fill_1 FILLER_31_2275 ();
 sg13g2_fill_2 FILLER_31_2281 ();
 sg13g2_fill_1 FILLER_31_2283 ();
 sg13g2_fill_2 FILLER_31_2293 ();
 sg13g2_fill_1 FILLER_31_2331 ();
 sg13g2_decap_8 FILLER_31_2349 ();
 sg13g2_decap_8 FILLER_31_2356 ();
 sg13g2_decap_8 FILLER_31_2363 ();
 sg13g2_decap_8 FILLER_31_2370 ();
 sg13g2_decap_8 FILLER_31_2377 ();
 sg13g2_fill_2 FILLER_31_2384 ();
 sg13g2_fill_2 FILLER_31_2396 ();
 sg13g2_fill_1 FILLER_31_2398 ();
 sg13g2_decap_8 FILLER_31_2409 ();
 sg13g2_decap_8 FILLER_31_2416 ();
 sg13g2_decap_8 FILLER_31_2423 ();
 sg13g2_decap_4 FILLER_31_2430 ();
 sg13g2_fill_2 FILLER_31_2434 ();
 sg13g2_fill_2 FILLER_31_2446 ();
 sg13g2_fill_1 FILLER_31_2448 ();
 sg13g2_decap_8 FILLER_31_2458 ();
 sg13g2_decap_8 FILLER_31_2465 ();
 sg13g2_decap_8 FILLER_31_2472 ();
 sg13g2_decap_8 FILLER_31_2479 ();
 sg13g2_decap_4 FILLER_31_2499 ();
 sg13g2_decap_8 FILLER_31_2549 ();
 sg13g2_decap_4 FILLER_31_2556 ();
 sg13g2_fill_2 FILLER_31_2560 ();
 sg13g2_fill_2 FILLER_31_2593 ();
 sg13g2_decap_8 FILLER_31_2616 ();
 sg13g2_fill_2 FILLER_31_2623 ();
 sg13g2_decap_8 FILLER_31_2647 ();
 sg13g2_decap_4 FILLER_31_2654 ();
 sg13g2_fill_2 FILLER_31_2658 ();
 sg13g2_decap_8 FILLER_31_2708 ();
 sg13g2_decap_8 FILLER_31_2715 ();
 sg13g2_fill_2 FILLER_31_2722 ();
 sg13g2_fill_2 FILLER_31_2728 ();
 sg13g2_fill_1 FILLER_31_2730 ();
 sg13g2_decap_4 FILLER_31_2768 ();
 sg13g2_fill_2 FILLER_31_2772 ();
 sg13g2_fill_2 FILLER_31_2787 ();
 sg13g2_fill_1 FILLER_31_2789 ();
 sg13g2_fill_2 FILLER_31_2838 ();
 sg13g2_decap_4 FILLER_31_2845 ();
 sg13g2_fill_1 FILLER_31_2849 ();
 sg13g2_decap_4 FILLER_31_2894 ();
 sg13g2_decap_8 FILLER_31_2948 ();
 sg13g2_decap_8 FILLER_31_2955 ();
 sg13g2_decap_4 FILLER_31_2962 ();
 sg13g2_fill_1 FILLER_31_2966 ();
 sg13g2_decap_8 FILLER_31_2980 ();
 sg13g2_decap_8 FILLER_31_2987 ();
 sg13g2_decap_8 FILLER_31_2994 ();
 sg13g2_decap_4 FILLER_31_3001 ();
 sg13g2_fill_2 FILLER_31_3005 ();
 sg13g2_fill_1 FILLER_31_3046 ();
 sg13g2_decap_8 FILLER_31_3051 ();
 sg13g2_decap_8 FILLER_31_3058 ();
 sg13g2_decap_4 FILLER_31_3065 ();
 sg13g2_fill_1 FILLER_31_3069 ();
 sg13g2_fill_2 FILLER_31_3101 ();
 sg13g2_fill_1 FILLER_31_3103 ();
 sg13g2_decap_8 FILLER_31_3131 ();
 sg13g2_decap_8 FILLER_31_3138 ();
 sg13g2_decap_8 FILLER_31_3145 ();
 sg13g2_fill_1 FILLER_31_3152 ();
 sg13g2_fill_1 FILLER_31_3157 ();
 sg13g2_decap_4 FILLER_31_3163 ();
 sg13g2_fill_2 FILLER_31_3167 ();
 sg13g2_decap_8 FILLER_31_3182 ();
 sg13g2_fill_2 FILLER_31_3189 ();
 sg13g2_fill_1 FILLER_31_3191 ();
 sg13g2_decap_8 FILLER_31_3196 ();
 sg13g2_decap_8 FILLER_31_3203 ();
 sg13g2_decap_8 FILLER_31_3210 ();
 sg13g2_fill_2 FILLER_31_3217 ();
 sg13g2_fill_1 FILLER_31_3219 ();
 sg13g2_decap_8 FILLER_31_3273 ();
 sg13g2_decap_8 FILLER_31_3280 ();
 sg13g2_decap_8 FILLER_31_3287 ();
 sg13g2_decap_8 FILLER_31_3294 ();
 sg13g2_decap_8 FILLER_31_3301 ();
 sg13g2_fill_2 FILLER_31_3308 ();
 sg13g2_fill_2 FILLER_31_3337 ();
 sg13g2_fill_1 FILLER_31_3365 ();
 sg13g2_decap_8 FILLER_31_3375 ();
 sg13g2_decap_8 FILLER_31_3382 ();
 sg13g2_decap_8 FILLER_31_3389 ();
 sg13g2_fill_2 FILLER_31_3396 ();
 sg13g2_fill_1 FILLER_31_3398 ();
 sg13g2_fill_2 FILLER_31_3439 ();
 sg13g2_decap_8 FILLER_31_3446 ();
 sg13g2_decap_4 FILLER_31_3453 ();
 sg13g2_fill_1 FILLER_31_3457 ();
 sg13g2_decap_8 FILLER_31_3471 ();
 sg13g2_decap_8 FILLER_31_3478 ();
 sg13g2_decap_8 FILLER_31_3485 ();
 sg13g2_decap_8 FILLER_31_3492 ();
 sg13g2_decap_8 FILLER_31_3499 ();
 sg13g2_decap_4 FILLER_31_3529 ();
 sg13g2_fill_2 FILLER_31_3533 ();
 sg13g2_decap_4 FILLER_31_3572 ();
 sg13g2_fill_2 FILLER_31_3576 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_55 ();
 sg13g2_fill_2 FILLER_32_83 ();
 sg13g2_fill_1 FILLER_32_85 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_decap_8 FILLER_32_127 ();
 sg13g2_decap_4 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_decap_4 FILLER_32_281 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_decap_4 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_4 FILLER_32_434 ();
 sg13g2_fill_1 FILLER_32_469 ();
 sg13g2_decap_4 FILLER_32_497 ();
 sg13g2_fill_1 FILLER_32_501 ();
 sg13g2_decap_8 FILLER_32_508 ();
 sg13g2_fill_1 FILLER_32_515 ();
 sg13g2_decap_8 FILLER_32_534 ();
 sg13g2_fill_2 FILLER_32_541 ();
 sg13g2_fill_2 FILLER_32_547 ();
 sg13g2_fill_1 FILLER_32_565 ();
 sg13g2_fill_1 FILLER_32_569 ();
 sg13g2_decap_8 FILLER_32_576 ();
 sg13g2_fill_2 FILLER_32_620 ();
 sg13g2_fill_1 FILLER_32_622 ();
 sg13g2_decap_8 FILLER_32_628 ();
 sg13g2_decap_8 FILLER_32_635 ();
 sg13g2_decap_4 FILLER_32_642 ();
 sg13g2_decap_4 FILLER_32_684 ();
 sg13g2_fill_2 FILLER_32_688 ();
 sg13g2_decap_4 FILLER_32_746 ();
 sg13g2_fill_2 FILLER_32_750 ();
 sg13g2_decap_8 FILLER_32_778 ();
 sg13g2_decap_8 FILLER_32_785 ();
 sg13g2_decap_4 FILLER_32_792 ();
 sg13g2_fill_2 FILLER_32_796 ();
 sg13g2_fill_1 FILLER_32_825 ();
 sg13g2_fill_2 FILLER_32_846 ();
 sg13g2_fill_1 FILLER_32_848 ();
 sg13g2_fill_2 FILLER_32_864 ();
 sg13g2_fill_1 FILLER_32_866 ();
 sg13g2_decap_8 FILLER_32_880 ();
 sg13g2_decap_8 FILLER_32_887 ();
 sg13g2_fill_1 FILLER_32_894 ();
 sg13g2_decap_8 FILLER_32_941 ();
 sg13g2_decap_8 FILLER_32_948 ();
 sg13g2_decap_4 FILLER_32_955 ();
 sg13g2_fill_1 FILLER_32_993 ();
 sg13g2_decap_4 FILLER_32_1007 ();
 sg13g2_fill_1 FILLER_32_1011 ();
 sg13g2_decap_4 FILLER_32_1028 ();
 sg13g2_fill_1 FILLER_32_1032 ();
 sg13g2_decap_4 FILLER_32_1046 ();
 sg13g2_fill_2 FILLER_32_1078 ();
 sg13g2_fill_1 FILLER_32_1080 ();
 sg13g2_decap_4 FILLER_32_1085 ();
 sg13g2_fill_2 FILLER_32_1089 ();
 sg13g2_fill_2 FILLER_32_1134 ();
 sg13g2_fill_1 FILLER_32_1136 ();
 sg13g2_decap_8 FILLER_32_1147 ();
 sg13g2_decap_8 FILLER_32_1154 ();
 sg13g2_fill_2 FILLER_32_1161 ();
 sg13g2_fill_1 FILLER_32_1180 ();
 sg13g2_fill_2 FILLER_32_1196 ();
 sg13g2_fill_1 FILLER_32_1198 ();
 sg13g2_decap_8 FILLER_32_1206 ();
 sg13g2_decap_4 FILLER_32_1213 ();
 sg13g2_fill_1 FILLER_32_1251 ();
 sg13g2_decap_8 FILLER_32_1268 ();
 sg13g2_decap_8 FILLER_32_1275 ();
 sg13g2_decap_8 FILLER_32_1282 ();
 sg13g2_decap_8 FILLER_32_1289 ();
 sg13g2_fill_2 FILLER_32_1296 ();
 sg13g2_decap_8 FILLER_32_1357 ();
 sg13g2_decap_8 FILLER_32_1364 ();
 sg13g2_decap_8 FILLER_32_1379 ();
 sg13g2_decap_8 FILLER_32_1386 ();
 sg13g2_fill_1 FILLER_32_1393 ();
 sg13g2_fill_2 FILLER_32_1405 ();
 sg13g2_fill_2 FILLER_32_1431 ();
 sg13g2_decap_4 FILLER_32_1439 ();
 sg13g2_fill_2 FILLER_32_1443 ();
 sg13g2_decap_4 FILLER_32_1449 ();
 sg13g2_fill_1 FILLER_32_1453 ();
 sg13g2_decap_8 FILLER_32_1472 ();
 sg13g2_fill_2 FILLER_32_1479 ();
 sg13g2_fill_2 FILLER_32_1499 ();
 sg13g2_fill_1 FILLER_32_1501 ();
 sg13g2_fill_2 FILLER_32_1518 ();
 sg13g2_fill_1 FILLER_32_1524 ();
 sg13g2_decap_8 FILLER_32_1544 ();
 sg13g2_decap_4 FILLER_32_1551 ();
 sg13g2_fill_1 FILLER_32_1555 ();
 sg13g2_fill_2 FILLER_32_1561 ();
 sg13g2_fill_1 FILLER_32_1563 ();
 sg13g2_decap_8 FILLER_32_1591 ();
 sg13g2_decap_4 FILLER_32_1598 ();
 sg13g2_decap_8 FILLER_32_1641 ();
 sg13g2_decap_4 FILLER_32_1648 ();
 sg13g2_fill_2 FILLER_32_1673 ();
 sg13g2_decap_8 FILLER_32_1688 ();
 sg13g2_decap_4 FILLER_32_1695 ();
 sg13g2_fill_1 FILLER_32_1699 ();
 sg13g2_fill_2 FILLER_32_1705 ();
 sg13g2_fill_2 FILLER_32_1725 ();
 sg13g2_decap_8 FILLER_32_1733 ();
 sg13g2_decap_4 FILLER_32_1740 ();
 sg13g2_fill_2 FILLER_32_1744 ();
 sg13g2_fill_2 FILLER_32_1751 ();
 sg13g2_fill_1 FILLER_32_1753 ();
 sg13g2_decap_8 FILLER_32_1783 ();
 sg13g2_decap_8 FILLER_32_1790 ();
 sg13g2_decap_8 FILLER_32_1797 ();
 sg13g2_decap_8 FILLER_32_1804 ();
 sg13g2_fill_2 FILLER_32_1811 ();
 sg13g2_decap_8 FILLER_32_1822 ();
 sg13g2_fill_2 FILLER_32_1834 ();
 sg13g2_fill_1 FILLER_32_1836 ();
 sg13g2_fill_1 FILLER_32_1902 ();
 sg13g2_fill_2 FILLER_32_1916 ();
 sg13g2_fill_2 FILLER_32_1931 ();
 sg13g2_fill_1 FILLER_32_1933 ();
 sg13g2_decap_8 FILLER_32_1947 ();
 sg13g2_fill_2 FILLER_32_1967 ();
 sg13g2_fill_2 FILLER_32_1985 ();
 sg13g2_fill_2 FILLER_32_1996 ();
 sg13g2_fill_2 FILLER_32_2024 ();
 sg13g2_fill_2 FILLER_32_2035 ();
 sg13g2_decap_4 FILLER_32_2060 ();
 sg13g2_fill_2 FILLER_32_2074 ();
 sg13g2_fill_1 FILLER_32_2080 ();
 sg13g2_fill_2 FILLER_32_2085 ();
 sg13g2_fill_1 FILLER_32_2100 ();
 sg13g2_fill_2 FILLER_32_2106 ();
 sg13g2_fill_1 FILLER_32_2108 ();
 sg13g2_fill_1 FILLER_32_2135 ();
 sg13g2_fill_1 FILLER_32_2156 ();
 sg13g2_fill_2 FILLER_32_2175 ();
 sg13g2_fill_2 FILLER_32_2186 ();
 sg13g2_fill_1 FILLER_32_2188 ();
 sg13g2_decap_8 FILLER_32_2198 ();
 sg13g2_decap_8 FILLER_32_2205 ();
 sg13g2_decap_8 FILLER_32_2212 ();
 sg13g2_decap_8 FILLER_32_2219 ();
 sg13g2_decap_4 FILLER_32_2226 ();
 sg13g2_decap_8 FILLER_32_2262 ();
 sg13g2_decap_8 FILLER_32_2269 ();
 sg13g2_decap_8 FILLER_32_2276 ();
 sg13g2_fill_2 FILLER_32_2309 ();
 sg13g2_decap_4 FILLER_32_2328 ();
 sg13g2_decap_8 FILLER_32_2354 ();
 sg13g2_decap_8 FILLER_32_2361 ();
 sg13g2_decap_4 FILLER_32_2368 ();
 sg13g2_fill_2 FILLER_32_2412 ();
 sg13g2_fill_2 FILLER_32_2423 ();
 sg13g2_fill_1 FILLER_32_2425 ();
 sg13g2_fill_1 FILLER_32_2430 ();
 sg13g2_decap_4 FILLER_32_2468 ();
 sg13g2_fill_1 FILLER_32_2522 ();
 sg13g2_fill_2 FILLER_32_2567 ();
 sg13g2_fill_1 FILLER_32_2579 ();
 sg13g2_fill_1 FILLER_32_2607 ();
 sg13g2_decap_4 FILLER_32_2645 ();
 sg13g2_fill_2 FILLER_32_2649 ();
 sg13g2_fill_2 FILLER_32_2678 ();
 sg13g2_fill_1 FILLER_32_2680 ();
 sg13g2_decap_8 FILLER_32_2708 ();
 sg13g2_decap_4 FILLER_32_2715 ();
 sg13g2_fill_1 FILLER_32_2756 ();
 sg13g2_decap_8 FILLER_32_2784 ();
 sg13g2_decap_4 FILLER_32_2791 ();
 sg13g2_fill_2 FILLER_32_2795 ();
 sg13g2_fill_1 FILLER_32_2829 ();
 sg13g2_decap_4 FILLER_32_2849 ();
 sg13g2_fill_1 FILLER_32_2853 ();
 sg13g2_decap_8 FILLER_32_2883 ();
 sg13g2_decap_4 FILLER_32_2890 ();
 sg13g2_fill_1 FILLER_32_2913 ();
 sg13g2_decap_8 FILLER_32_2946 ();
 sg13g2_fill_2 FILLER_32_2953 ();
 sg13g2_decap_8 FILLER_32_2992 ();
 sg13g2_decap_8 FILLER_32_2999 ();
 sg13g2_decap_8 FILLER_32_3006 ();
 sg13g2_decap_8 FILLER_32_3013 ();
 sg13g2_fill_1 FILLER_32_3020 ();
 sg13g2_decap_8 FILLER_32_3052 ();
 sg13g2_decap_4 FILLER_32_3059 ();
 sg13g2_fill_1 FILLER_32_3076 ();
 sg13g2_fill_2 FILLER_32_3087 ();
 sg13g2_fill_1 FILLER_32_3089 ();
 sg13g2_decap_4 FILLER_32_3126 ();
 sg13g2_fill_1 FILLER_32_3130 ();
 sg13g2_decap_8 FILLER_32_3161 ();
 sg13g2_decap_8 FILLER_32_3168 ();
 sg13g2_decap_8 FILLER_32_3175 ();
 sg13g2_decap_8 FILLER_32_3182 ();
 sg13g2_decap_8 FILLER_32_3189 ();
 sg13g2_decap_8 FILLER_32_3196 ();
 sg13g2_decap_4 FILLER_32_3203 ();
 sg13g2_fill_2 FILLER_32_3207 ();
 sg13g2_fill_2 FILLER_32_3213 ();
 sg13g2_fill_2 FILLER_32_3259 ();
 sg13g2_decap_8 FILLER_32_3270 ();
 sg13g2_fill_1 FILLER_32_3277 ();
 sg13g2_decap_8 FILLER_32_3291 ();
 sg13g2_decap_8 FILLER_32_3298 ();
 sg13g2_decap_4 FILLER_32_3332 ();
 sg13g2_fill_2 FILLER_32_3336 ();
 sg13g2_decap_8 FILLER_32_3378 ();
 sg13g2_decap_4 FILLER_32_3385 ();
 sg13g2_fill_2 FILLER_32_3389 ();
 sg13g2_decap_4 FILLER_32_3432 ();
 sg13g2_fill_1 FILLER_32_3436 ();
 sg13g2_decap_8 FILLER_32_3450 ();
 sg13g2_decap_8 FILLER_32_3457 ();
 sg13g2_decap_8 FILLER_32_3464 ();
 sg13g2_decap_4 FILLER_32_3481 ();
 sg13g2_fill_2 FILLER_32_3485 ();
 sg13g2_decap_8 FILLER_32_3496 ();
 sg13g2_fill_2 FILLER_32_3503 ();
 sg13g2_fill_1 FILLER_32_3505 ();
 sg13g2_decap_8 FILLER_32_3516 ();
 sg13g2_fill_2 FILLER_32_3523 ();
 sg13g2_fill_1 FILLER_32_3525 ();
 sg13g2_decap_8 FILLER_32_3544 ();
 sg13g2_decap_4 FILLER_32_3551 ();
 sg13g2_decap_8 FILLER_32_3564 ();
 sg13g2_decap_8 FILLER_32_3571 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_143 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_184 ();
 sg13g2_decap_8 FILLER_33_223 ();
 sg13g2_decap_8 FILLER_33_230 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_292 ();
 sg13g2_decap_8 FILLER_33_352 ();
 sg13g2_decap_4 FILLER_33_359 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_decap_4 FILLER_33_402 ();
 sg13g2_decap_4 FILLER_33_412 ();
 sg13g2_decap_4 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_425 ();
 sg13g2_decap_4 FILLER_33_436 ();
 sg13g2_decap_8 FILLER_33_456 ();
 sg13g2_decap_8 FILLER_33_514 ();
 sg13g2_decap_8 FILLER_33_521 ();
 sg13g2_decap_4 FILLER_33_528 ();
 sg13g2_fill_2 FILLER_33_532 ();
 sg13g2_fill_1 FILLER_33_554 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_fill_2 FILLER_33_588 ();
 sg13g2_decap_4 FILLER_33_603 ();
 sg13g2_fill_2 FILLER_33_620 ();
 sg13g2_fill_1 FILLER_33_622 ();
 sg13g2_fill_2 FILLER_33_628 ();
 sg13g2_fill_1 FILLER_33_630 ();
 sg13g2_fill_1 FILLER_33_638 ();
 sg13g2_decap_8 FILLER_33_676 ();
 sg13g2_fill_1 FILLER_33_701 ();
 sg13g2_decap_4 FILLER_33_746 ();
 sg13g2_fill_1 FILLER_33_750 ();
 sg13g2_decap_4 FILLER_33_757 ();
 sg13g2_fill_2 FILLER_33_765 ();
 sg13g2_fill_1 FILLER_33_767 ();
 sg13g2_decap_8 FILLER_33_773 ();
 sg13g2_fill_1 FILLER_33_780 ();
 sg13g2_fill_1 FILLER_33_794 ();
 sg13g2_fill_1 FILLER_33_808 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_decap_8 FILLER_33_846 ();
 sg13g2_decap_4 FILLER_33_853 ();
 sg13g2_fill_2 FILLER_33_879 ();
 sg13g2_fill_1 FILLER_33_894 ();
 sg13g2_decap_4 FILLER_33_909 ();
 sg13g2_fill_1 FILLER_33_926 ();
 sg13g2_decap_8 FILLER_33_935 ();
 sg13g2_decap_8 FILLER_33_942 ();
 sg13g2_decap_8 FILLER_33_949 ();
 sg13g2_fill_2 FILLER_33_956 ();
 sg13g2_fill_1 FILLER_33_958 ();
 sg13g2_fill_1 FILLER_33_992 ();
 sg13g2_fill_2 FILLER_33_998 ();
 sg13g2_fill_2 FILLER_33_1017 ();
 sg13g2_fill_1 FILLER_33_1019 ();
 sg13g2_fill_1 FILLER_33_1036 ();
 sg13g2_fill_1 FILLER_33_1050 ();
 sg13g2_fill_2 FILLER_33_1088 ();
 sg13g2_fill_1 FILLER_33_1107 ();
 sg13g2_decap_8 FILLER_33_1132 ();
 sg13g2_decap_4 FILLER_33_1139 ();
 sg13g2_fill_1 FILLER_33_1143 ();
 sg13g2_decap_8 FILLER_33_1151 ();
 sg13g2_decap_8 FILLER_33_1158 ();
 sg13g2_decap_8 FILLER_33_1165 ();
 sg13g2_fill_2 FILLER_33_1172 ();
 sg13g2_decap_8 FILLER_33_1200 ();
 sg13g2_decap_8 FILLER_33_1207 ();
 sg13g2_fill_2 FILLER_33_1214 ();
 sg13g2_fill_1 FILLER_33_1216 ();
 sg13g2_fill_2 FILLER_33_1245 ();
 sg13g2_fill_1 FILLER_33_1247 ();
 sg13g2_fill_2 FILLER_33_1293 ();
 sg13g2_fill_1 FILLER_33_1295 ();
 sg13g2_fill_1 FILLER_33_1329 ();
 sg13g2_decap_8 FILLER_33_1349 ();
 sg13g2_decap_8 FILLER_33_1356 ();
 sg13g2_decap_4 FILLER_33_1363 ();
 sg13g2_fill_1 FILLER_33_1367 ();
 sg13g2_fill_2 FILLER_33_1396 ();
 sg13g2_decap_8 FILLER_33_1404 ();
 sg13g2_fill_1 FILLER_33_1439 ();
 sg13g2_fill_2 FILLER_33_1448 ();
 sg13g2_fill_1 FILLER_33_1462 ();
 sg13g2_decap_4 FILLER_33_1521 ();
 sg13g2_fill_1 FILLER_33_1525 ();
 sg13g2_decap_4 FILLER_33_1572 ();
 sg13g2_decap_4 FILLER_33_1581 ();
 sg13g2_decap_8 FILLER_33_1598 ();
 sg13g2_fill_1 FILLER_33_1605 ();
 sg13g2_decap_8 FILLER_33_1632 ();
 sg13g2_decap_8 FILLER_33_1639 ();
 sg13g2_decap_4 FILLER_33_1646 ();
 sg13g2_decap_8 FILLER_33_1692 ();
 sg13g2_decap_8 FILLER_33_1699 ();
 sg13g2_decap_4 FILLER_33_1706 ();
 sg13g2_decap_8 FILLER_33_1727 ();
 sg13g2_fill_2 FILLER_33_1734 ();
 sg13g2_fill_1 FILLER_33_1736 ();
 sg13g2_fill_2 FILLER_33_1763 ();
 sg13g2_fill_1 FILLER_33_1765 ();
 sg13g2_decap_8 FILLER_33_1785 ();
 sg13g2_decap_8 FILLER_33_1792 ();
 sg13g2_decap_8 FILLER_33_1799 ();
 sg13g2_decap_4 FILLER_33_1811 ();
 sg13g2_fill_1 FILLER_33_1815 ();
 sg13g2_fill_2 FILLER_33_1857 ();
 sg13g2_fill_1 FILLER_33_1859 ();
 sg13g2_fill_2 FILLER_33_1865 ();
 sg13g2_decap_8 FILLER_33_1873 ();
 sg13g2_decap_8 FILLER_33_1890 ();
 sg13g2_fill_2 FILLER_33_1897 ();
 sg13g2_fill_1 FILLER_33_1913 ();
 sg13g2_decap_4 FILLER_33_1922 ();
 sg13g2_fill_1 FILLER_33_1926 ();
 sg13g2_fill_2 FILLER_33_1953 ();
 sg13g2_fill_2 FILLER_33_1960 ();
 sg13g2_fill_1 FILLER_33_1962 ();
 sg13g2_decap_8 FILLER_33_1976 ();
 sg13g2_decap_8 FILLER_33_1983 ();
 sg13g2_decap_8 FILLER_33_1990 ();
 sg13g2_decap_4 FILLER_33_2038 ();
 sg13g2_fill_1 FILLER_33_2042 ();
 sg13g2_decap_8 FILLER_33_2071 ();
 sg13g2_fill_2 FILLER_33_2078 ();
 sg13g2_decap_8 FILLER_33_2088 ();
 sg13g2_decap_8 FILLER_33_2095 ();
 sg13g2_decap_8 FILLER_33_2102 ();
 sg13g2_decap_4 FILLER_33_2109 ();
 sg13g2_fill_1 FILLER_33_2113 ();
 sg13g2_decap_4 FILLER_33_2127 ();
 sg13g2_fill_2 FILLER_33_2131 ();
 sg13g2_fill_1 FILLER_33_2157 ();
 sg13g2_fill_2 FILLER_33_2167 ();
 sg13g2_decap_8 FILLER_33_2176 ();
 sg13g2_decap_4 FILLER_33_2183 ();
 sg13g2_decap_4 FILLER_33_2215 ();
 sg13g2_fill_1 FILLER_33_2219 ();
 sg13g2_fill_2 FILLER_33_2333 ();
 sg13g2_decap_8 FILLER_33_2344 ();
 sg13g2_decap_8 FILLER_33_2351 ();
 sg13g2_decap_4 FILLER_33_2358 ();
 sg13g2_decap_4 FILLER_33_2498 ();
 sg13g2_fill_2 FILLER_33_2519 ();
 sg13g2_fill_2 FILLER_33_2604 ();
 sg13g2_decap_8 FILLER_33_2644 ();
 sg13g2_decap_8 FILLER_33_2705 ();
 sg13g2_decap_8 FILLER_33_2712 ();
 sg13g2_fill_2 FILLER_33_2719 ();
 sg13g2_fill_1 FILLER_33_2721 ();
 sg13g2_decap_8 FILLER_33_2772 ();
 sg13g2_fill_1 FILLER_33_2779 ();
 sg13g2_decap_8 FILLER_33_2851 ();
 sg13g2_decap_4 FILLER_33_2858 ();
 sg13g2_fill_2 FILLER_33_2862 ();
 sg13g2_decap_8 FILLER_33_2868 ();
 sg13g2_decap_8 FILLER_33_2875 ();
 sg13g2_decap_8 FILLER_33_2882 ();
 sg13g2_decap_4 FILLER_33_2889 ();
 sg13g2_fill_1 FILLER_33_2893 ();
 sg13g2_fill_1 FILLER_33_2908 ();
 sg13g2_fill_2 FILLER_33_2936 ();
 sg13g2_fill_1 FILLER_33_2938 ();
 sg13g2_decap_4 FILLER_33_2952 ();
 sg13g2_decap_4 FILLER_33_3002 ();
 sg13g2_fill_1 FILLER_33_3048 ();
 sg13g2_fill_1 FILLER_33_3053 ();
 sg13g2_fill_2 FILLER_33_3126 ();
 sg13g2_decap_4 FILLER_33_3141 ();
 sg13g2_fill_2 FILLER_33_3145 ();
 sg13g2_fill_2 FILLER_33_3178 ();
 sg13g2_fill_1 FILLER_33_3180 ();
 sg13g2_fill_1 FILLER_33_3185 ();
 sg13g2_decap_8 FILLER_33_3190 ();
 sg13g2_decap_8 FILLER_33_3197 ();
 sg13g2_fill_2 FILLER_33_3257 ();
 sg13g2_fill_1 FILLER_33_3259 ();
 sg13g2_decap_4 FILLER_33_3331 ();
 sg13g2_fill_1 FILLER_33_3335 ();
 sg13g2_decap_4 FILLER_33_3380 ();
 sg13g2_fill_2 FILLER_33_3384 ();
 sg13g2_fill_2 FILLER_33_3399 ();
 sg13g2_decap_8 FILLER_33_3441 ();
 sg13g2_decap_8 FILLER_33_3448 ();
 sg13g2_decap_8 FILLER_33_3455 ();
 sg13g2_decap_8 FILLER_33_3462 ();
 sg13g2_fill_2 FILLER_33_3469 ();
 sg13g2_fill_1 FILLER_33_3471 ();
 sg13g2_fill_2 FILLER_33_3499 ();
 sg13g2_fill_2 FILLER_33_3514 ();
 sg13g2_decap_8 FILLER_33_3543 ();
 sg13g2_decap_4 FILLER_33_3550 ();
 sg13g2_fill_1 FILLER_33_3554 ();
 sg13g2_decap_8 FILLER_33_3564 ();
 sg13g2_decap_8 FILLER_33_3571 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_11 ();
 sg13g2_decap_4 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_53 ();
 sg13g2_fill_1 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_2 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_decap_4 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_fill_2 FILLER_34_159 ();
 sg13g2_decap_4 FILLER_34_183 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_decap_4 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_decap_8 FILLER_34_282 ();
 sg13g2_decap_8 FILLER_34_289 ();
 sg13g2_decap_8 FILLER_34_296 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_decap_4 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_358 ();
 sg13g2_decap_4 FILLER_34_365 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_392 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_fill_2 FILLER_34_426 ();
 sg13g2_decap_4 FILLER_34_436 ();
 sg13g2_fill_1 FILLER_34_440 ();
 sg13g2_decap_8 FILLER_34_463 ();
 sg13g2_decap_4 FILLER_34_496 ();
 sg13g2_fill_1 FILLER_34_510 ();
 sg13g2_fill_2 FILLER_34_538 ();
 sg13g2_fill_1 FILLER_34_540 ();
 sg13g2_decap_8 FILLER_34_576 ();
 sg13g2_decap_8 FILLER_34_583 ();
 sg13g2_decap_8 FILLER_34_590 ();
 sg13g2_fill_1 FILLER_34_597 ();
 sg13g2_decap_8 FILLER_34_608 ();
 sg13g2_decap_8 FILLER_34_615 ();
 sg13g2_decap_8 FILLER_34_622 ();
 sg13g2_decap_4 FILLER_34_629 ();
 sg13g2_fill_2 FILLER_34_633 ();
 sg13g2_fill_1 FILLER_34_670 ();
 sg13g2_decap_8 FILLER_34_680 ();
 sg13g2_decap_8 FILLER_34_687 ();
 sg13g2_decap_4 FILLER_34_694 ();
 sg13g2_fill_2 FILLER_34_706 ();
 sg13g2_fill_1 FILLER_34_721 ();
 sg13g2_fill_1 FILLER_34_726 ();
 sg13g2_fill_1 FILLER_34_745 ();
 sg13g2_decap_8 FILLER_34_752 ();
 sg13g2_fill_2 FILLER_34_759 ();
 sg13g2_fill_1 FILLER_34_761 ();
 sg13g2_fill_1 FILLER_34_795 ();
 sg13g2_fill_1 FILLER_34_832 ();
 sg13g2_decap_4 FILLER_34_838 ();
 sg13g2_fill_1 FILLER_34_848 ();
 sg13g2_decap_8 FILLER_34_867 ();
 sg13g2_decap_8 FILLER_34_874 ();
 sg13g2_fill_1 FILLER_34_923 ();
 sg13g2_decap_8 FILLER_34_937 ();
 sg13g2_decap_8 FILLER_34_944 ();
 sg13g2_fill_2 FILLER_34_951 ();
 sg13g2_fill_1 FILLER_34_953 ();
 sg13g2_fill_1 FILLER_34_988 ();
 sg13g2_fill_1 FILLER_34_1035 ();
 sg13g2_decap_8 FILLER_34_1053 ();
 sg13g2_fill_2 FILLER_34_1060 ();
 sg13g2_decap_4 FILLER_34_1065 ();
 sg13g2_fill_1 FILLER_34_1069 ();
 sg13g2_decap_8 FILLER_34_1138 ();
 sg13g2_fill_2 FILLER_34_1150 ();
 sg13g2_fill_1 FILLER_34_1152 ();
 sg13g2_decap_8 FILLER_34_1161 ();
 sg13g2_decap_8 FILLER_34_1168 ();
 sg13g2_fill_2 FILLER_34_1175 ();
 sg13g2_fill_1 FILLER_34_1177 ();
 sg13g2_fill_2 FILLER_34_1192 ();
 sg13g2_fill_1 FILLER_34_1200 ();
 sg13g2_decap_8 FILLER_34_1210 ();
 sg13g2_fill_2 FILLER_34_1226 ();
 sg13g2_fill_2 FILLER_34_1247 ();
 sg13g2_fill_2 FILLER_34_1255 ();
 sg13g2_fill_2 FILLER_34_1285 ();
 sg13g2_fill_1 FILLER_34_1287 ();
 sg13g2_decap_4 FILLER_34_1331 ();
 sg13g2_decap_8 FILLER_34_1345 ();
 sg13g2_decap_8 FILLER_34_1352 ();
 sg13g2_decap_8 FILLER_34_1359 ();
 sg13g2_decap_8 FILLER_34_1366 ();
 sg13g2_decap_8 FILLER_34_1373 ();
 sg13g2_decap_8 FILLER_34_1380 ();
 sg13g2_decap_8 FILLER_34_1387 ();
 sg13g2_fill_2 FILLER_34_1407 ();
 sg13g2_decap_8 FILLER_34_1436 ();
 sg13g2_decap_4 FILLER_34_1451 ();
 sg13g2_fill_1 FILLER_34_1455 ();
 sg13g2_decap_8 FILLER_34_1461 ();
 sg13g2_decap_8 FILLER_34_1468 ();
 sg13g2_decap_8 FILLER_34_1475 ();
 sg13g2_decap_8 FILLER_34_1482 ();
 sg13g2_decap_8 FILLER_34_1499 ();
 sg13g2_fill_1 FILLER_34_1506 ();
 sg13g2_decap_8 FILLER_34_1516 ();
 sg13g2_decap_8 FILLER_34_1523 ();
 sg13g2_decap_8 FILLER_34_1530 ();
 sg13g2_decap_8 FILLER_34_1537 ();
 sg13g2_decap_4 FILLER_34_1544 ();
 sg13g2_fill_1 FILLER_34_1548 ();
 sg13g2_decap_8 FILLER_34_1556 ();
 sg13g2_decap_8 FILLER_34_1563 ();
 sg13g2_decap_8 FILLER_34_1570 ();
 sg13g2_decap_8 FILLER_34_1577 ();
 sg13g2_decap_8 FILLER_34_1584 ();
 sg13g2_decap_4 FILLER_34_1591 ();
 sg13g2_fill_2 FILLER_34_1595 ();
 sg13g2_fill_2 FILLER_34_1611 ();
 sg13g2_fill_1 FILLER_34_1613 ();
 sg13g2_fill_1 FILLER_34_1623 ();
 sg13g2_fill_2 FILLER_34_1654 ();
 sg13g2_fill_1 FILLER_34_1656 ();
 sg13g2_decap_8 FILLER_34_1692 ();
 sg13g2_decap_8 FILLER_34_1699 ();
 sg13g2_decap_8 FILLER_34_1706 ();
 sg13g2_decap_8 FILLER_34_1713 ();
 sg13g2_decap_8 FILLER_34_1720 ();
 sg13g2_decap_4 FILLER_34_1727 ();
 sg13g2_fill_2 FILLER_34_1731 ();
 sg13g2_decap_4 FILLER_34_1752 ();
 sg13g2_fill_2 FILLER_34_1768 ();
 sg13g2_fill_1 FILLER_34_1770 ();
 sg13g2_fill_2 FILLER_34_1777 ();
 sg13g2_decap_8 FILLER_34_1783 ();
 sg13g2_decap_8 FILLER_34_1790 ();
 sg13g2_decap_8 FILLER_34_1797 ();
 sg13g2_fill_2 FILLER_34_1804 ();
 sg13g2_decap_8 FILLER_34_1854 ();
 sg13g2_decap_8 FILLER_34_1861 ();
 sg13g2_fill_1 FILLER_34_1868 ();
 sg13g2_fill_1 FILLER_34_1890 ();
 sg13g2_decap_4 FILLER_34_1901 ();
 sg13g2_decap_8 FILLER_34_1923 ();
 sg13g2_decap_4 FILLER_34_1930 ();
 sg13g2_fill_1 FILLER_34_1934 ();
 sg13g2_decap_8 FILLER_34_1939 ();
 sg13g2_fill_2 FILLER_34_1946 ();
 sg13g2_fill_1 FILLER_34_1948 ();
 sg13g2_decap_8 FILLER_34_1962 ();
 sg13g2_fill_2 FILLER_34_1969 ();
 sg13g2_fill_1 FILLER_34_1971 ();
 sg13g2_decap_8 FILLER_34_1975 ();
 sg13g2_fill_2 FILLER_34_1982 ();
 sg13g2_fill_1 FILLER_34_1984 ();
 sg13g2_decap_8 FILLER_34_1998 ();
 sg13g2_decap_4 FILLER_34_2005 ();
 sg13g2_decap_8 FILLER_34_2021 ();
 sg13g2_decap_8 FILLER_34_2028 ();
 sg13g2_decap_8 FILLER_34_2035 ();
 sg13g2_fill_1 FILLER_34_2042 ();
 sg13g2_fill_2 FILLER_34_2048 ();
 sg13g2_fill_1 FILLER_34_2050 ();
 sg13g2_decap_8 FILLER_34_2055 ();
 sg13g2_decap_8 FILLER_34_2062 ();
 sg13g2_decap_8 FILLER_34_2069 ();
 sg13g2_decap_8 FILLER_34_2076 ();
 sg13g2_decap_8 FILLER_34_2083 ();
 sg13g2_decap_8 FILLER_34_2090 ();
 sg13g2_decap_8 FILLER_34_2097 ();
 sg13g2_decap_4 FILLER_34_2104 ();
 sg13g2_fill_1 FILLER_34_2108 ();
 sg13g2_fill_1 FILLER_34_2118 ();
 sg13g2_decap_8 FILLER_34_2123 ();
 sg13g2_decap_4 FILLER_34_2130 ();
 sg13g2_fill_1 FILLER_34_2134 ();
 sg13g2_fill_2 FILLER_34_2157 ();
 sg13g2_fill_1 FILLER_34_2159 ();
 sg13g2_fill_2 FILLER_34_2178 ();
 sg13g2_decap_8 FILLER_34_2185 ();
 sg13g2_fill_1 FILLER_34_2192 ();
 sg13g2_decap_8 FILLER_34_2202 ();
 sg13g2_decap_8 FILLER_34_2209 ();
 sg13g2_decap_8 FILLER_34_2216 ();
 sg13g2_decap_8 FILLER_34_2223 ();
 sg13g2_fill_1 FILLER_34_2230 ();
 sg13g2_decap_8 FILLER_34_2267 ();
 sg13g2_fill_2 FILLER_34_2274 ();
 sg13g2_decap_8 FILLER_34_2344 ();
 sg13g2_decap_8 FILLER_34_2351 ();
 sg13g2_decap_4 FILLER_34_2358 ();
 sg13g2_fill_1 FILLER_34_2362 ();
 sg13g2_fill_2 FILLER_34_2394 ();
 sg13g2_decap_4 FILLER_34_2417 ();
 sg13g2_fill_2 FILLER_34_2421 ();
 sg13g2_fill_2 FILLER_34_2433 ();
 sg13g2_decap_4 FILLER_34_2484 ();
 sg13g2_fill_2 FILLER_34_2488 ();
 sg13g2_decap_8 FILLER_34_2494 ();
 sg13g2_decap_8 FILLER_34_2501 ();
 sg13g2_decap_8 FILLER_34_2508 ();
 sg13g2_decap_8 FILLER_34_2515 ();
 sg13g2_decap_8 FILLER_34_2522 ();
 sg13g2_decap_8 FILLER_34_2529 ();
 sg13g2_decap_8 FILLER_34_2549 ();
 sg13g2_fill_2 FILLER_34_2556 ();
 sg13g2_fill_1 FILLER_34_2558 ();
 sg13g2_decap_8 FILLER_34_2569 ();
 sg13g2_fill_2 FILLER_34_2576 ();
 sg13g2_decap_8 FILLER_34_2606 ();
 sg13g2_decap_8 FILLER_34_2613 ();
 sg13g2_decap_8 FILLER_34_2620 ();
 sg13g2_decap_4 FILLER_34_2627 ();
 sg13g2_fill_2 FILLER_34_2631 ();
 sg13g2_decap_4 FILLER_34_2656 ();
 sg13g2_fill_1 FILLER_34_2660 ();
 sg13g2_fill_2 FILLER_34_2675 ();
 sg13g2_decap_8 FILLER_34_2696 ();
 sg13g2_decap_8 FILLER_34_2703 ();
 sg13g2_fill_2 FILLER_34_2710 ();
 sg13g2_fill_1 FILLER_34_2712 ();
 sg13g2_decap_8 FILLER_34_2765 ();
 sg13g2_decap_8 FILLER_34_2772 ();
 sg13g2_decap_8 FILLER_34_2779 ();
 sg13g2_decap_8 FILLER_34_2786 ();
 sg13g2_decap_4 FILLER_34_2793 ();
 sg13g2_fill_1 FILLER_34_2797 ();
 sg13g2_decap_8 FILLER_34_2802 ();
 sg13g2_decap_8 FILLER_34_2809 ();
 sg13g2_fill_2 FILLER_34_2816 ();
 sg13g2_fill_1 FILLER_34_2818 ();
 sg13g2_decap_8 FILLER_34_2865 ();
 sg13g2_decap_4 FILLER_34_2872 ();
 sg13g2_fill_2 FILLER_34_2876 ();
 sg13g2_decap_8 FILLER_34_2886 ();
 sg13g2_decap_4 FILLER_34_2893 ();
 sg13g2_fill_2 FILLER_34_2897 ();
 sg13g2_decap_4 FILLER_34_2939 ();
 sg13g2_fill_2 FILLER_34_2943 ();
 sg13g2_decap_8 FILLER_34_2990 ();
 sg13g2_decap_4 FILLER_34_2997 ();
 sg13g2_fill_1 FILLER_34_3001 ();
 sg13g2_fill_2 FILLER_34_3044 ();
 sg13g2_fill_1 FILLER_34_3046 ();
 sg13g2_decap_4 FILLER_34_3074 ();
 sg13g2_fill_2 FILLER_34_3078 ();
 sg13g2_decap_4 FILLER_34_3106 ();
 sg13g2_decap_8 FILLER_34_3128 ();
 sg13g2_fill_2 FILLER_34_3135 ();
 sg13g2_fill_2 FILLER_34_3183 ();
 sg13g2_fill_1 FILLER_34_3185 ();
 sg13g2_decap_8 FILLER_34_3191 ();
 sg13g2_decap_4 FILLER_34_3198 ();
 sg13g2_fill_1 FILLER_34_3202 ();
 sg13g2_fill_1 FILLER_34_3243 ();
 sg13g2_decap_8 FILLER_34_3254 ();
 sg13g2_decap_4 FILLER_34_3261 ();
 sg13g2_fill_2 FILLER_34_3275 ();
 sg13g2_fill_2 FILLER_34_3303 ();
 sg13g2_fill_1 FILLER_34_3305 ();
 sg13g2_decap_8 FILLER_34_3371 ();
 sg13g2_decap_8 FILLER_34_3378 ();
 sg13g2_fill_1 FILLER_34_3385 ();
 sg13g2_fill_2 FILLER_34_3405 ();
 sg13g2_fill_1 FILLER_34_3407 ();
 sg13g2_decap_8 FILLER_34_3427 ();
 sg13g2_decap_8 FILLER_34_3434 ();
 sg13g2_decap_8 FILLER_34_3441 ();
 sg13g2_fill_2 FILLER_34_3448 ();
 sg13g2_decap_4 FILLER_34_3504 ();
 sg13g2_fill_1 FILLER_34_3508 ();
 sg13g2_decap_8 FILLER_34_3549 ();
 sg13g2_decap_8 FILLER_34_3556 ();
 sg13g2_decap_8 FILLER_34_3563 ();
 sg13g2_decap_8 FILLER_34_3570 ();
 sg13g2_fill_1 FILLER_34_3577 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_decap_8 FILLER_35_55 ();
 sg13g2_fill_1 FILLER_35_62 ();
 sg13g2_fill_2 FILLER_35_143 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_4 FILLER_35_211 ();
 sg13g2_fill_2 FILLER_35_215 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_305 ();
 sg13g2_fill_2 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_4 FILLER_35_396 ();
 sg13g2_fill_2 FILLER_35_400 ();
 sg13g2_decap_4 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_35_411 ();
 sg13g2_fill_1 FILLER_35_425 ();
 sg13g2_decap_8 FILLER_35_465 ();
 sg13g2_decap_4 FILLER_35_472 ();
 sg13g2_fill_2 FILLER_35_476 ();
 sg13g2_fill_2 FILLER_35_482 ();
 sg13g2_fill_1 FILLER_35_489 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_4 FILLER_35_532 ();
 sg13g2_fill_2 FILLER_35_536 ();
 sg13g2_fill_1 FILLER_35_547 ();
 sg13g2_fill_1 FILLER_35_557 ();
 sg13g2_decap_8 FILLER_35_570 ();
 sg13g2_decap_8 FILLER_35_577 ();
 sg13g2_decap_8 FILLER_35_584 ();
 sg13g2_decap_8 FILLER_35_591 ();
 sg13g2_decap_8 FILLER_35_598 ();
 sg13g2_decap_8 FILLER_35_605 ();
 sg13g2_decap_8 FILLER_35_612 ();
 sg13g2_fill_1 FILLER_35_619 ();
 sg13g2_decap_8 FILLER_35_625 ();
 sg13g2_fill_2 FILLER_35_632 ();
 sg13g2_fill_2 FILLER_35_647 ();
 sg13g2_fill_2 FILLER_35_669 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_fill_2 FILLER_35_686 ();
 sg13g2_fill_1 FILLER_35_688 ();
 sg13g2_decap_8 FILLER_35_751 ();
 sg13g2_decap_8 FILLER_35_758 ();
 sg13g2_fill_1 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_783 ();
 sg13g2_decap_8 FILLER_35_790 ();
 sg13g2_decap_8 FILLER_35_797 ();
 sg13g2_decap_8 FILLER_35_804 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_decap_8 FILLER_35_818 ();
 sg13g2_decap_4 FILLER_35_825 ();
 sg13g2_fill_2 FILLER_35_829 ();
 sg13g2_fill_1 FILLER_35_851 ();
 sg13g2_decap_8 FILLER_35_870 ();
 sg13g2_decap_4 FILLER_35_877 ();
 sg13g2_fill_1 FILLER_35_881 ();
 sg13g2_fill_1 FILLER_35_887 ();
 sg13g2_fill_2 FILLER_35_902 ();
 sg13g2_decap_8 FILLER_35_921 ();
 sg13g2_decap_8 FILLER_35_928 ();
 sg13g2_decap_8 FILLER_35_935 ();
 sg13g2_fill_2 FILLER_35_942 ();
 sg13g2_decap_4 FILLER_35_948 ();
 sg13g2_fill_1 FILLER_35_952 ();
 sg13g2_decap_4 FILLER_35_958 ();
 sg13g2_fill_2 FILLER_35_962 ();
 sg13g2_decap_4 FILLER_35_992 ();
 sg13g2_fill_2 FILLER_35_996 ();
 sg13g2_decap_4 FILLER_35_1011 ();
 sg13g2_fill_2 FILLER_35_1015 ();
 sg13g2_fill_2 FILLER_35_1030 ();
 sg13g2_decap_8 FILLER_35_1044 ();
 sg13g2_decap_8 FILLER_35_1051 ();
 sg13g2_decap_8 FILLER_35_1058 ();
 sg13g2_decap_8 FILLER_35_1065 ();
 sg13g2_fill_2 FILLER_35_1072 ();
 sg13g2_fill_1 FILLER_35_1074 ();
 sg13g2_fill_2 FILLER_35_1083 ();
 sg13g2_fill_1 FILLER_35_1085 ();
 sg13g2_fill_1 FILLER_35_1095 ();
 sg13g2_fill_2 FILLER_35_1110 ();
 sg13g2_fill_2 FILLER_35_1122 ();
 sg13g2_fill_2 FILLER_35_1128 ();
 sg13g2_fill_2 FILLER_35_1143 ();
 sg13g2_fill_1 FILLER_35_1145 ();
 sg13g2_fill_1 FILLER_35_1150 ();
 sg13g2_decap_4 FILLER_35_1160 ();
 sg13g2_fill_1 FILLER_35_1164 ();
 sg13g2_decap_4 FILLER_35_1169 ();
 sg13g2_decap_8 FILLER_35_1220 ();
 sg13g2_fill_2 FILLER_35_1227 ();
 sg13g2_decap_8 FILLER_35_1239 ();
 sg13g2_fill_2 FILLER_35_1301 ();
 sg13g2_decap_8 FILLER_35_1346 ();
 sg13g2_decap_8 FILLER_35_1353 ();
 sg13g2_decap_8 FILLER_35_1360 ();
 sg13g2_fill_2 FILLER_35_1367 ();
 sg13g2_fill_2 FILLER_35_1374 ();
 sg13g2_fill_1 FILLER_35_1376 ();
 sg13g2_decap_4 FILLER_35_1381 ();
 sg13g2_fill_1 FILLER_35_1409 ();
 sg13g2_decap_8 FILLER_35_1414 ();
 sg13g2_fill_1 FILLER_35_1421 ();
 sg13g2_decap_8 FILLER_35_1427 ();
 sg13g2_decap_4 FILLER_35_1434 ();
 sg13g2_decap_8 FILLER_35_1444 ();
 sg13g2_decap_8 FILLER_35_1451 ();
 sg13g2_decap_8 FILLER_35_1458 ();
 sg13g2_decap_8 FILLER_35_1465 ();
 sg13g2_decap_8 FILLER_35_1472 ();
 sg13g2_fill_1 FILLER_35_1479 ();
 sg13g2_decap_8 FILLER_35_1512 ();
 sg13g2_fill_2 FILLER_35_1519 ();
 sg13g2_fill_1 FILLER_35_1521 ();
 sg13g2_decap_4 FILLER_35_1530 ();
 sg13g2_fill_1 FILLER_35_1534 ();
 sg13g2_fill_2 FILLER_35_1560 ();
 sg13g2_decap_8 FILLER_35_1566 ();
 sg13g2_decap_8 FILLER_35_1573 ();
 sg13g2_decap_8 FILLER_35_1580 ();
 sg13g2_decap_4 FILLER_35_1587 ();
 sg13g2_fill_2 FILLER_35_1591 ();
 sg13g2_decap_4 FILLER_35_1626 ();
 sg13g2_fill_2 FILLER_35_1630 ();
 sg13g2_fill_2 FILLER_35_1688 ();
 sg13g2_fill_1 FILLER_35_1690 ();
 sg13g2_decap_8 FILLER_35_1703 ();
 sg13g2_fill_2 FILLER_35_1710 ();
 sg13g2_fill_1 FILLER_35_1712 ();
 sg13g2_fill_1 FILLER_35_1722 ();
 sg13g2_fill_1 FILLER_35_1767 ();
 sg13g2_decap_8 FILLER_35_1796 ();
 sg13g2_decap_8 FILLER_35_1803 ();
 sg13g2_decap_8 FILLER_35_1810 ();
 sg13g2_decap_8 FILLER_35_1817 ();
 sg13g2_decap_8 FILLER_35_1824 ();
 sg13g2_decap_4 FILLER_35_1831 ();
 sg13g2_decap_8 FILLER_35_1840 ();
 sg13g2_decap_8 FILLER_35_1847 ();
 sg13g2_decap_8 FILLER_35_1854 ();
 sg13g2_fill_1 FILLER_35_1861 ();
 sg13g2_fill_1 FILLER_35_1884 ();
 sg13g2_decap_8 FILLER_35_1890 ();
 sg13g2_decap_8 FILLER_35_1897 ();
 sg13g2_fill_1 FILLER_35_1904 ();
 sg13g2_fill_2 FILLER_35_1913 ();
 sg13g2_fill_2 FILLER_35_1932 ();
 sg13g2_fill_1 FILLER_35_1934 ();
 sg13g2_fill_2 FILLER_35_1948 ();
 sg13g2_fill_1 FILLER_35_1950 ();
 sg13g2_decap_8 FILLER_35_1993 ();
 sg13g2_fill_1 FILLER_35_2000 ();
 sg13g2_decap_4 FILLER_35_2029 ();
 sg13g2_fill_1 FILLER_35_2033 ();
 sg13g2_fill_1 FILLER_35_2047 ();
 sg13g2_fill_1 FILLER_35_2058 ();
 sg13g2_decap_8 FILLER_35_2063 ();
 sg13g2_decap_8 FILLER_35_2070 ();
 sg13g2_fill_2 FILLER_35_2077 ();
 sg13g2_fill_1 FILLER_35_2079 ();
 sg13g2_fill_2 FILLER_35_2108 ();
 sg13g2_decap_8 FILLER_35_2121 ();
 sg13g2_decap_8 FILLER_35_2128 ();
 sg13g2_decap_4 FILLER_35_2135 ();
 sg13g2_fill_2 FILLER_35_2139 ();
 sg13g2_fill_1 FILLER_35_2163 ();
 sg13g2_fill_1 FILLER_35_2202 ();
 sg13g2_decap_8 FILLER_35_2212 ();
 sg13g2_decap_8 FILLER_35_2219 ();
 sg13g2_decap_4 FILLER_35_2226 ();
 sg13g2_fill_1 FILLER_35_2230 ();
 sg13g2_decap_8 FILLER_35_2264 ();
 sg13g2_decap_8 FILLER_35_2271 ();
 sg13g2_fill_2 FILLER_35_2278 ();
 sg13g2_fill_1 FILLER_35_2289 ();
 sg13g2_fill_1 FILLER_35_2317 ();
 sg13g2_decap_8 FILLER_35_2354 ();
 sg13g2_decap_8 FILLER_35_2361 ();
 sg13g2_decap_8 FILLER_35_2372 ();
 sg13g2_fill_1 FILLER_35_2379 ();
 sg13g2_decap_8 FILLER_35_2409 ();
 sg13g2_decap_8 FILLER_35_2416 ();
 sg13g2_decap_8 FILLER_35_2423 ();
 sg13g2_decap_8 FILLER_35_2430 ();
 sg13g2_fill_2 FILLER_35_2437 ();
 sg13g2_fill_1 FILLER_35_2448 ();
 sg13g2_decap_8 FILLER_35_2474 ();
 sg13g2_decap_4 FILLER_35_2485 ();
 sg13g2_decap_8 FILLER_35_2498 ();
 sg13g2_decap_8 FILLER_35_2505 ();
 sg13g2_decap_8 FILLER_35_2512 ();
 sg13g2_decap_8 FILLER_35_2519 ();
 sg13g2_decap_8 FILLER_35_2526 ();
 sg13g2_fill_2 FILLER_35_2533 ();
 sg13g2_decap_8 FILLER_35_2548 ();
 sg13g2_decap_8 FILLER_35_2591 ();
 sg13g2_decap_8 FILLER_35_2598 ();
 sg13g2_fill_1 FILLER_35_2605 ();
 sg13g2_decap_4 FILLER_35_2619 ();
 sg13g2_decap_4 FILLER_35_2637 ();
 sg13g2_decap_8 FILLER_35_2654 ();
 sg13g2_decap_8 FILLER_35_2661 ();
 sg13g2_fill_2 FILLER_35_2668 ();
 sg13g2_fill_1 FILLER_35_2670 ();
 sg13g2_fill_2 FILLER_35_2684 ();
 sg13g2_fill_1 FILLER_35_2686 ();
 sg13g2_decap_4 FILLER_35_2691 ();
 sg13g2_fill_1 FILLER_35_2695 ();
 sg13g2_fill_2 FILLER_35_2724 ();
 sg13g2_fill_1 FILLER_35_2761 ();
 sg13g2_decap_8 FILLER_35_2767 ();
 sg13g2_decap_8 FILLER_35_2774 ();
 sg13g2_decap_8 FILLER_35_2781 ();
 sg13g2_fill_1 FILLER_35_2788 ();
 sg13g2_fill_2 FILLER_35_2794 ();
 sg13g2_decap_8 FILLER_35_2809 ();
 sg13g2_fill_2 FILLER_35_2816 ();
 sg13g2_decap_8 FILLER_35_2866 ();
 sg13g2_decap_8 FILLER_35_2873 ();
 sg13g2_decap_8 FILLER_35_2880 ();
 sg13g2_decap_4 FILLER_35_2887 ();
 sg13g2_fill_1 FILLER_35_2891 ();
 sg13g2_decap_8 FILLER_35_2931 ();
 sg13g2_decap_8 FILLER_35_2938 ();
 sg13g2_decap_4 FILLER_35_2945 ();
 sg13g2_fill_1 FILLER_35_2949 ();
 sg13g2_decap_8 FILLER_35_2995 ();
 sg13g2_fill_2 FILLER_35_3002 ();
 sg13g2_fill_1 FILLER_35_3004 ();
 sg13g2_fill_1 FILLER_35_3013 ();
 sg13g2_fill_2 FILLER_35_3031 ();
 sg13g2_fill_1 FILLER_35_3033 ();
 sg13g2_decap_8 FILLER_35_3071 ();
 sg13g2_decap_8 FILLER_35_3078 ();
 sg13g2_fill_2 FILLER_35_3085 ();
 sg13g2_fill_1 FILLER_35_3087 ();
 sg13g2_fill_1 FILLER_35_3164 ();
 sg13g2_decap_4 FILLER_35_3186 ();
 sg13g2_fill_2 FILLER_35_3200 ();
 sg13g2_fill_2 FILLER_35_3229 ();
 sg13g2_decap_8 FILLER_35_3250 ();
 sg13g2_fill_1 FILLER_35_3257 ();
 sg13g2_decap_4 FILLER_35_3284 ();
 sg13g2_fill_1 FILLER_35_3288 ();
 sg13g2_decap_8 FILLER_35_3302 ();
 sg13g2_fill_1 FILLER_35_3309 ();
 sg13g2_fill_2 FILLER_35_3320 ();
 sg13g2_fill_1 FILLER_35_3322 ();
 sg13g2_fill_2 FILLER_35_3332 ();
 sg13g2_fill_1 FILLER_35_3334 ();
 sg13g2_decap_8 FILLER_35_3356 ();
 sg13g2_decap_8 FILLER_35_3363 ();
 sg13g2_decap_8 FILLER_35_3370 ();
 sg13g2_decap_4 FILLER_35_3377 ();
 sg13g2_fill_1 FILLER_35_3381 ();
 sg13g2_decap_8 FILLER_35_3418 ();
 sg13g2_decap_8 FILLER_35_3425 ();
 sg13g2_decap_8 FILLER_35_3432 ();
 sg13g2_decap_4 FILLER_35_3439 ();
 sg13g2_decap_8 FILLER_35_3498 ();
 sg13g2_fill_2 FILLER_35_3505 ();
 sg13g2_fill_1 FILLER_35_3507 ();
 sg13g2_decap_4 FILLER_35_3539 ();
 sg13g2_fill_1 FILLER_35_3543 ();
 sg13g2_decap_8 FILLER_35_3571 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_68 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_fill_2 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_decap_4 FILLER_36_355 ();
 sg13g2_fill_2 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_8 FILLER_36_403 ();
 sg13g2_decap_4 FILLER_36_410 ();
 sg13g2_fill_2 FILLER_36_414 ();
 sg13g2_decap_4 FILLER_36_421 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_decap_8 FILLER_36_458 ();
 sg13g2_decap_8 FILLER_36_465 ();
 sg13g2_decap_8 FILLER_36_472 ();
 sg13g2_decap_8 FILLER_36_479 ();
 sg13g2_decap_8 FILLER_36_486 ();
 sg13g2_decap_4 FILLER_36_493 ();
 sg13g2_fill_1 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_decap_8 FILLER_36_511 ();
 sg13g2_fill_2 FILLER_36_518 ();
 sg13g2_decap_8 FILLER_36_533 ();
 sg13g2_decap_4 FILLER_36_540 ();
 sg13g2_fill_2 FILLER_36_566 ();
 sg13g2_decap_8 FILLER_36_579 ();
 sg13g2_decap_8 FILLER_36_586 ();
 sg13g2_decap_4 FILLER_36_593 ();
 sg13g2_fill_2 FILLER_36_597 ();
 sg13g2_decap_8 FILLER_36_635 ();
 sg13g2_fill_2 FILLER_36_642 ();
 sg13g2_fill_1 FILLER_36_644 ();
 sg13g2_decap_8 FILLER_36_667 ();
 sg13g2_decap_8 FILLER_36_674 ();
 sg13g2_decap_4 FILLER_36_681 ();
 sg13g2_fill_1 FILLER_36_709 ();
 sg13g2_decap_8 FILLER_36_747 ();
 sg13g2_fill_1 FILLER_36_754 ();
 sg13g2_decap_8 FILLER_36_773 ();
 sg13g2_decap_8 FILLER_36_780 ();
 sg13g2_decap_8 FILLER_36_787 ();
 sg13g2_decap_8 FILLER_36_794 ();
 sg13g2_fill_2 FILLER_36_801 ();
 sg13g2_fill_1 FILLER_36_803 ();
 sg13g2_fill_2 FILLER_36_814 ();
 sg13g2_fill_2 FILLER_36_829 ();
 sg13g2_fill_1 FILLER_36_831 ();
 sg13g2_fill_1 FILLER_36_837 ();
 sg13g2_fill_1 FILLER_36_846 ();
 sg13g2_fill_2 FILLER_36_855 ();
 sg13g2_fill_2 FILLER_36_885 ();
 sg13g2_fill_1 FILLER_36_887 ();
 sg13g2_decap_4 FILLER_36_932 ();
 sg13g2_fill_1 FILLER_36_936 ();
 sg13g2_decap_4 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1011 ();
 sg13g2_decap_8 FILLER_36_1018 ();
 sg13g2_decap_8 FILLER_36_1025 ();
 sg13g2_fill_2 FILLER_36_1032 ();
 sg13g2_decap_8 FILLER_36_1047 ();
 sg13g2_decap_8 FILLER_36_1054 ();
 sg13g2_decap_8 FILLER_36_1061 ();
 sg13g2_decap_4 FILLER_36_1068 ();
 sg13g2_fill_2 FILLER_36_1072 ();
 sg13g2_decap_4 FILLER_36_1093 ();
 sg13g2_fill_1 FILLER_36_1101 ();
 sg13g2_decap_4 FILLER_36_1127 ();
 sg13g2_fill_1 FILLER_36_1131 ();
 sg13g2_fill_2 FILLER_36_1144 ();
 sg13g2_fill_1 FILLER_36_1169 ();
 sg13g2_fill_1 FILLER_36_1184 ();
 sg13g2_fill_2 FILLER_36_1203 ();
 sg13g2_fill_2 FILLER_36_1217 ();
 sg13g2_fill_1 FILLER_36_1219 ();
 sg13g2_fill_2 FILLER_36_1230 ();
 sg13g2_decap_8 FILLER_36_1236 ();
 sg13g2_decap_4 FILLER_36_1243 ();
 sg13g2_fill_2 FILLER_36_1252 ();
 sg13g2_fill_1 FILLER_36_1254 ();
 sg13g2_decap_8 FILLER_36_1291 ();
 sg13g2_fill_1 FILLER_36_1298 ();
 sg13g2_decap_4 FILLER_36_1320 ();
 sg13g2_decap_8 FILLER_36_1337 ();
 sg13g2_decap_8 FILLER_36_1344 ();
 sg13g2_decap_8 FILLER_36_1351 ();
 sg13g2_fill_2 FILLER_36_1358 ();
 sg13g2_fill_1 FILLER_36_1360 ();
 sg13g2_fill_2 FILLER_36_1398 ();
 sg13g2_decap_4 FILLER_36_1420 ();
 sg13g2_fill_2 FILLER_36_1424 ();
 sg13g2_fill_1 FILLER_36_1431 ();
 sg13g2_decap_4 FILLER_36_1448 ();
 sg13g2_decap_8 FILLER_36_1468 ();
 sg13g2_fill_1 FILLER_36_1475 ();
 sg13g2_decap_4 FILLER_36_1533 ();
 sg13g2_decap_4 FILLER_36_1565 ();
 sg13g2_fill_2 FILLER_36_1569 ();
 sg13g2_fill_2 FILLER_36_1591 ();
 sg13g2_decap_8 FILLER_36_1598 ();
 sg13g2_decap_8 FILLER_36_1605 ();
 sg13g2_decap_4 FILLER_36_1612 ();
 sg13g2_fill_2 FILLER_36_1616 ();
 sg13g2_decap_8 FILLER_36_1630 ();
 sg13g2_decap_8 FILLER_36_1637 ();
 sg13g2_decap_8 FILLER_36_1644 ();
 sg13g2_decap_4 FILLER_36_1651 ();
 sg13g2_fill_2 FILLER_36_1655 ();
 sg13g2_decap_8 FILLER_36_1670 ();
 sg13g2_decap_8 FILLER_36_1677 ();
 sg13g2_decap_4 FILLER_36_1684 ();
 sg13g2_fill_1 FILLER_36_1688 ();
 sg13g2_fill_1 FILLER_36_1702 ();
 sg13g2_decap_4 FILLER_36_1716 ();
 sg13g2_fill_1 FILLER_36_1720 ();
 sg13g2_decap_8 FILLER_36_1797 ();
 sg13g2_fill_1 FILLER_36_1804 ();
 sg13g2_decap_8 FILLER_36_1852 ();
 sg13g2_decap_8 FILLER_36_1859 ();
 sg13g2_decap_4 FILLER_36_1866 ();
 sg13g2_decap_8 FILLER_36_1898 ();
 sg13g2_fill_2 FILLER_36_1905 ();
 sg13g2_decap_8 FILLER_36_1944 ();
 sg13g2_fill_2 FILLER_36_1998 ();
 sg13g2_fill_1 FILLER_36_2000 ();
 sg13g2_decap_8 FILLER_36_2017 ();
 sg13g2_fill_2 FILLER_36_2024 ();
 sg13g2_fill_2 FILLER_36_2060 ();
 sg13g2_decap_8 FILLER_36_2067 ();
 sg13g2_fill_2 FILLER_36_2078 ();
 sg13g2_fill_1 FILLER_36_2088 ();
 sg13g2_fill_1 FILLER_36_2100 ();
 sg13g2_fill_1 FILLER_36_2115 ();
 sg13g2_decap_8 FILLER_36_2128 ();
 sg13g2_decap_8 FILLER_36_2135 ();
 sg13g2_decap_8 FILLER_36_2174 ();
 sg13g2_fill_2 FILLER_36_2244 ();
 sg13g2_fill_1 FILLER_36_2246 ();
 sg13g2_decap_8 FILLER_36_2277 ();
 sg13g2_decap_4 FILLER_36_2284 ();
 sg13g2_fill_2 FILLER_36_2288 ();
 sg13g2_fill_2 FILLER_36_2304 ();
 sg13g2_fill_1 FILLER_36_2310 ();
 sg13g2_decap_8 FILLER_36_2338 ();
 sg13g2_decap_8 FILLER_36_2345 ();
 sg13g2_decap_4 FILLER_36_2352 ();
 sg13g2_decap_8 FILLER_36_2365 ();
 sg13g2_decap_8 FILLER_36_2372 ();
 sg13g2_decap_8 FILLER_36_2379 ();
 sg13g2_fill_1 FILLER_36_2386 ();
 sg13g2_decap_8 FILLER_36_2396 ();
 sg13g2_fill_1 FILLER_36_2403 ();
 sg13g2_fill_1 FILLER_36_2431 ();
 sg13g2_decap_8 FILLER_36_2449 ();
 sg13g2_decap_8 FILLER_36_2456 ();
 sg13g2_decap_8 FILLER_36_2463 ();
 sg13g2_decap_4 FILLER_36_2470 ();
 sg13g2_fill_2 FILLER_36_2474 ();
 sg13g2_decap_8 FILLER_36_2512 ();
 sg13g2_decap_8 FILLER_36_2519 ();
 sg13g2_decap_8 FILLER_36_2526 ();
 sg13g2_fill_1 FILLER_36_2533 ();
 sg13g2_fill_2 FILLER_36_2565 ();
 sg13g2_fill_1 FILLER_36_2567 ();
 sg13g2_decap_8 FILLER_36_2622 ();
 sg13g2_fill_1 FILLER_36_2629 ();
 sg13g2_decap_4 FILLER_36_2657 ();
 sg13g2_decap_8 FILLER_36_2670 ();
 sg13g2_decap_8 FILLER_36_2677 ();
 sg13g2_decap_4 FILLER_36_2684 ();
 sg13g2_fill_2 FILLER_36_2740 ();
 sg13g2_fill_1 FILLER_36_2742 ();
 sg13g2_fill_1 FILLER_36_2770 ();
 sg13g2_decap_8 FILLER_36_2808 ();
 sg13g2_decap_4 FILLER_36_2815 ();
 sg13g2_fill_2 FILLER_36_2819 ();
 sg13g2_fill_2 FILLER_36_2834 ();
 sg13g2_fill_2 FILLER_36_2863 ();
 sg13g2_fill_1 FILLER_36_2865 ();
 sg13g2_decap_4 FILLER_36_2870 ();
 sg13g2_fill_1 FILLER_36_2884 ();
 sg13g2_decap_8 FILLER_36_2922 ();
 sg13g2_decap_8 FILLER_36_2929 ();
 sg13g2_decap_8 FILLER_36_2936 ();
 sg13g2_decap_8 FILLER_36_2943 ();
 sg13g2_decap_8 FILLER_36_2981 ();
 sg13g2_decap_8 FILLER_36_2988 ();
 sg13g2_decap_8 FILLER_36_2995 ();
 sg13g2_decap_8 FILLER_36_3002 ();
 sg13g2_decap_8 FILLER_36_3009 ();
 sg13g2_decap_8 FILLER_36_3016 ();
 sg13g2_fill_2 FILLER_36_3023 ();
 sg13g2_decap_4 FILLER_36_3034 ();
 sg13g2_fill_2 FILLER_36_3038 ();
 sg13g2_decap_8 FILLER_36_3070 ();
 sg13g2_decap_8 FILLER_36_3077 ();
 sg13g2_decap_8 FILLER_36_3123 ();
 sg13g2_decap_8 FILLER_36_3130 ();
 sg13g2_fill_1 FILLER_36_3137 ();
 sg13g2_decap_4 FILLER_36_3170 ();
 sg13g2_fill_2 FILLER_36_3246 ();
 sg13g2_fill_1 FILLER_36_3248 ();
 sg13g2_fill_1 FILLER_36_3259 ();
 sg13g2_fill_2 FILLER_36_3287 ();
 sg13g2_fill_1 FILLER_36_3289 ();
 sg13g2_decap_8 FILLER_36_3303 ();
 sg13g2_decap_4 FILLER_36_3310 ();
 sg13g2_fill_2 FILLER_36_3314 ();
 sg13g2_fill_2 FILLER_36_3353 ();
 sg13g2_fill_1 FILLER_36_3355 ();
 sg13g2_decap_8 FILLER_36_3360 ();
 sg13g2_fill_2 FILLER_36_3367 ();
 sg13g2_fill_2 FILLER_36_3416 ();
 sg13g2_decap_8 FILLER_36_3428 ();
 sg13g2_decap_8 FILLER_36_3435 ();
 sg13g2_decap_8 FILLER_36_3491 ();
 sg13g2_fill_2 FILLER_36_3498 ();
 sg13g2_decap_4 FILLER_36_3544 ();
 sg13g2_fill_1 FILLER_36_3548 ();
 sg13g2_fill_1 FILLER_36_3553 ();
 sg13g2_decap_8 FILLER_36_3563 ();
 sg13g2_decap_8 FILLER_36_3570 ();
 sg13g2_fill_1 FILLER_36_3577 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_53 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_110 ();
 sg13g2_decap_4 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_4 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_decap_4 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_299 ();
 sg13g2_decap_4 FILLER_37_310 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_decap_8 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_372 ();
 sg13g2_fill_1 FILLER_37_384 ();
 sg13g2_decap_4 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_37_412 ();
 sg13g2_decap_8 FILLER_37_419 ();
 sg13g2_decap_8 FILLER_37_426 ();
 sg13g2_decap_8 FILLER_37_433 ();
 sg13g2_decap_8 FILLER_37_440 ();
 sg13g2_decap_8 FILLER_37_447 ();
 sg13g2_decap_8 FILLER_37_454 ();
 sg13g2_decap_4 FILLER_37_489 ();
 sg13g2_fill_2 FILLER_37_493 ();
 sg13g2_decap_8 FILLER_37_536 ();
 sg13g2_decap_4 FILLER_37_543 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_fill_1 FILLER_37_580 ();
 sg13g2_decap_8 FILLER_37_593 ();
 sg13g2_decap_8 FILLER_37_654 ();
 sg13g2_decap_8 FILLER_37_661 ();
 sg13g2_decap_8 FILLER_37_671 ();
 sg13g2_decap_8 FILLER_37_678 ();
 sg13g2_decap_8 FILLER_37_685 ();
 sg13g2_decap_4 FILLER_37_692 ();
 sg13g2_fill_1 FILLER_37_696 ();
 sg13g2_fill_1 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_740 ();
 sg13g2_decap_8 FILLER_37_747 ();
 sg13g2_decap_8 FILLER_37_754 ();
 sg13g2_fill_2 FILLER_37_767 ();
 sg13g2_fill_2 FILLER_37_774 ();
 sg13g2_fill_1 FILLER_37_776 ();
 sg13g2_decap_4 FILLER_37_790 ();
 sg13g2_fill_1 FILLER_37_799 ();
 sg13g2_decap_8 FILLER_37_809 ();
 sg13g2_fill_2 FILLER_37_816 ();
 sg13g2_fill_2 FILLER_37_855 ();
 sg13g2_decap_8 FILLER_37_871 ();
 sg13g2_decap_8 FILLER_37_891 ();
 sg13g2_decap_8 FILLER_37_898 ();
 sg13g2_fill_2 FILLER_37_905 ();
 sg13g2_fill_2 FILLER_37_920 ();
 sg13g2_fill_1 FILLER_37_931 ();
 sg13g2_decap_4 FILLER_37_945 ();
 sg13g2_fill_2 FILLER_37_949 ();
 sg13g2_fill_1 FILLER_37_956 ();
 sg13g2_fill_1 FILLER_37_966 ();
 sg13g2_fill_1 FILLER_37_974 ();
 sg13g2_decap_8 FILLER_37_983 ();
 sg13g2_decap_8 FILLER_37_990 ();
 sg13g2_decap_4 FILLER_37_1024 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_decap_8 FILLER_37_1033 ();
 sg13g2_decap_8 FILLER_37_1040 ();
 sg13g2_decap_8 FILLER_37_1047 ();
 sg13g2_decap_4 FILLER_37_1054 ();
 sg13g2_fill_1 FILLER_37_1058 ();
 sg13g2_fill_1 FILLER_37_1067 ();
 sg13g2_decap_8 FILLER_37_1110 ();
 sg13g2_decap_8 FILLER_37_1117 ();
 sg13g2_decap_8 FILLER_37_1124 ();
 sg13g2_decap_4 FILLER_37_1131 ();
 sg13g2_decap_8 FILLER_37_1140 ();
 sg13g2_fill_2 FILLER_37_1147 ();
 sg13g2_decap_4 FILLER_37_1154 ();
 sg13g2_fill_2 FILLER_37_1158 ();
 sg13g2_fill_1 FILLER_37_1164 ();
 sg13g2_fill_2 FILLER_37_1178 ();
 sg13g2_fill_2 FILLER_37_1189 ();
 sg13g2_decap_8 FILLER_37_1200 ();
 sg13g2_decap_8 FILLER_37_1207 ();
 sg13g2_decap_4 FILLER_37_1214 ();
 sg13g2_decap_8 FILLER_37_1227 ();
 sg13g2_fill_1 FILLER_37_1234 ();
 sg13g2_decap_8 FILLER_37_1245 ();
 sg13g2_fill_1 FILLER_37_1252 ();
 sg13g2_fill_2 FILLER_37_1268 ();
 sg13g2_fill_1 FILLER_37_1270 ();
 sg13g2_decap_4 FILLER_37_1286 ();
 sg13g2_fill_2 FILLER_37_1303 ();
 sg13g2_fill_2 FILLER_37_1310 ();
 sg13g2_fill_2 FILLER_37_1327 ();
 sg13g2_decap_8 FILLER_37_1342 ();
 sg13g2_fill_2 FILLER_37_1349 ();
 sg13g2_fill_1 FILLER_37_1351 ();
 sg13g2_fill_1 FILLER_37_1394 ();
 sg13g2_fill_2 FILLER_37_1409 ();
 sg13g2_fill_1 FILLER_37_1411 ();
 sg13g2_decap_4 FILLER_37_1420 ();
 sg13g2_fill_2 FILLER_37_1424 ();
 sg13g2_decap_8 FILLER_37_1430 ();
 sg13g2_fill_2 FILLER_37_1437 ();
 sg13g2_fill_1 FILLER_37_1439 ();
 sg13g2_fill_1 FILLER_37_1445 ();
 sg13g2_fill_2 FILLER_37_1463 ();
 sg13g2_decap_8 FILLER_37_1509 ();
 sg13g2_decap_8 FILLER_37_1516 ();
 sg13g2_decap_8 FILLER_37_1523 ();
 sg13g2_decap_8 FILLER_37_1530 ();
 sg13g2_fill_1 FILLER_37_1537 ();
 sg13g2_decap_4 FILLER_37_1546 ();
 sg13g2_fill_2 FILLER_37_1550 ();
 sg13g2_decap_4 FILLER_37_1571 ();
 sg13g2_fill_1 FILLER_37_1575 ();
 sg13g2_decap_4 FILLER_37_1586 ();
 sg13g2_fill_2 FILLER_37_1590 ();
 sg13g2_decap_8 FILLER_37_1607 ();
 sg13g2_fill_2 FILLER_37_1614 ();
 sg13g2_fill_1 FILLER_37_1616 ();
 sg13g2_fill_1 FILLER_37_1632 ();
 sg13g2_decap_8 FILLER_37_1658 ();
 sg13g2_decap_8 FILLER_37_1665 ();
 sg13g2_decap_8 FILLER_37_1672 ();
 sg13g2_fill_2 FILLER_37_1679 ();
 sg13g2_decap_4 FILLER_37_1686 ();
 sg13g2_fill_1 FILLER_37_1690 ();
 sg13g2_fill_1 FILLER_37_1718 ();
 sg13g2_decap_4 FILLER_37_1732 ();
 sg13g2_fill_2 FILLER_37_1779 ();
 sg13g2_fill_1 FILLER_37_1781 ();
 sg13g2_fill_1 FILLER_37_1790 ();
 sg13g2_fill_1 FILLER_37_1814 ();
 sg13g2_decap_4 FILLER_37_1824 ();
 sg13g2_fill_1 FILLER_37_1828 ();
 sg13g2_fill_2 FILLER_37_1837 ();
 sg13g2_fill_2 FILLER_37_1853 ();
 sg13g2_fill_1 FILLER_37_1855 ();
 sg13g2_decap_8 FILLER_37_1860 ();
 sg13g2_decap_4 FILLER_37_1867 ();
 sg13g2_fill_1 FILLER_37_1871 ();
 sg13g2_fill_1 FILLER_37_1893 ();
 sg13g2_decap_8 FILLER_37_1910 ();
 sg13g2_fill_1 FILLER_37_1917 ();
 sg13g2_decap_8 FILLER_37_1927 ();
 sg13g2_decap_8 FILLER_37_1934 ();
 sg13g2_decap_8 FILLER_37_1941 ();
 sg13g2_decap_4 FILLER_37_1948 ();
 sg13g2_fill_2 FILLER_37_1952 ();
 sg13g2_fill_1 FILLER_37_1967 ();
 sg13g2_fill_2 FILLER_37_1973 ();
 sg13g2_decap_8 FILLER_37_1983 ();
 sg13g2_decap_4 FILLER_37_1990 ();
 sg13g2_fill_2 FILLER_37_1994 ();
 sg13g2_fill_2 FILLER_37_2014 ();
 sg13g2_fill_1 FILLER_37_2016 ();
 sg13g2_decap_8 FILLER_37_2026 ();
 sg13g2_fill_2 FILLER_37_2033 ();
 sg13g2_fill_2 FILLER_37_2041 ();
 sg13g2_fill_2 FILLER_37_2051 ();
 sg13g2_fill_1 FILLER_37_2053 ();
 sg13g2_decap_8 FILLER_37_2058 ();
 sg13g2_fill_2 FILLER_37_2065 ();
 sg13g2_fill_1 FILLER_37_2067 ();
 sg13g2_decap_8 FILLER_37_2087 ();
 sg13g2_fill_2 FILLER_37_2094 ();
 sg13g2_fill_1 FILLER_37_2096 ();
 sg13g2_fill_1 FILLER_37_2119 ();
 sg13g2_decap_8 FILLER_37_2128 ();
 sg13g2_decap_4 FILLER_37_2135 ();
 sg13g2_fill_1 FILLER_37_2139 ();
 sg13g2_fill_2 FILLER_37_2153 ();
 sg13g2_fill_1 FILLER_37_2155 ();
 sg13g2_decap_8 FILLER_37_2175 ();
 sg13g2_decap_8 FILLER_37_2182 ();
 sg13g2_fill_2 FILLER_37_2189 ();
 sg13g2_fill_1 FILLER_37_2199 ();
 sg13g2_decap_8 FILLER_37_2210 ();
 sg13g2_fill_2 FILLER_37_2217 ();
 sg13g2_decap_8 FILLER_37_2275 ();
 sg13g2_decap_8 FILLER_37_2282 ();
 sg13g2_decap_8 FILLER_37_2289 ();
 sg13g2_fill_1 FILLER_37_2296 ();
 sg13g2_decap_8 FILLER_37_2338 ();
 sg13g2_decap_8 FILLER_37_2345 ();
 sg13g2_fill_2 FILLER_37_2352 ();
 sg13g2_decap_8 FILLER_37_2371 ();
 sg13g2_decap_4 FILLER_37_2378 ();
 sg13g2_fill_2 FILLER_37_2382 ();
 sg13g2_decap_8 FILLER_37_2424 ();
 sg13g2_fill_2 FILLER_37_2431 ();
 sg13g2_decap_8 FILLER_37_2460 ();
 sg13g2_fill_2 FILLER_37_2467 ();
 sg13g2_fill_1 FILLER_37_2469 ();
 sg13g2_decap_8 FILLER_37_2520 ();
 sg13g2_decap_8 FILLER_37_2527 ();
 sg13g2_decap_8 FILLER_37_2534 ();
 sg13g2_fill_2 FILLER_37_2541 ();
 sg13g2_fill_1 FILLER_37_2543 ();
 sg13g2_fill_1 FILLER_37_2557 ();
 sg13g2_fill_1 FILLER_37_2571 ();
 sg13g2_decap_8 FILLER_37_2597 ();
 sg13g2_fill_2 FILLER_37_2613 ();
 sg13g2_fill_1 FILLER_37_2615 ();
 sg13g2_decap_8 FILLER_37_2670 ();
 sg13g2_decap_4 FILLER_37_2677 ();
 sg13g2_fill_1 FILLER_37_2681 ();
 sg13g2_fill_1 FILLER_37_2740 ();
 sg13g2_fill_2 FILLER_37_2777 ();
 sg13g2_decap_8 FILLER_37_2815 ();
 sg13g2_decap_8 FILLER_37_2835 ();
 sg13g2_decap_8 FILLER_37_2842 ();
 sg13g2_decap_8 FILLER_37_2849 ();
 sg13g2_decap_8 FILLER_37_2856 ();
 sg13g2_decap_4 FILLER_37_2863 ();
 sg13g2_decap_8 FILLER_37_2931 ();
 sg13g2_decap_8 FILLER_37_2938 ();
 sg13g2_decap_4 FILLER_37_2945 ();
 sg13g2_fill_1 FILLER_37_2949 ();
 sg13g2_decap_8 FILLER_37_2977 ();
 sg13g2_decap_8 FILLER_37_2984 ();
 sg13g2_decap_8 FILLER_37_2991 ();
 sg13g2_decap_4 FILLER_37_2998 ();
 sg13g2_fill_2 FILLER_37_3002 ();
 sg13g2_fill_1 FILLER_37_3051 ();
 sg13g2_fill_2 FILLER_37_3056 ();
 sg13g2_fill_1 FILLER_37_3058 ();
 sg13g2_decap_8 FILLER_37_3068 ();
 sg13g2_decap_8 FILLER_37_3075 ();
 sg13g2_fill_2 FILLER_37_3134 ();
 sg13g2_fill_1 FILLER_37_3136 ();
 sg13g2_fill_2 FILLER_37_3150 ();
 sg13g2_fill_1 FILLER_37_3152 ();
 sg13g2_decap_8 FILLER_37_3171 ();
 sg13g2_fill_2 FILLER_37_3178 ();
 sg13g2_decap_8 FILLER_37_3184 ();
 sg13g2_decap_8 FILLER_37_3191 ();
 sg13g2_decap_4 FILLER_37_3198 ();
 sg13g2_fill_2 FILLER_37_3202 ();
 sg13g2_fill_1 FILLER_37_3287 ();
 sg13g2_decap_4 FILLER_37_3301 ();
 sg13g2_fill_1 FILLER_37_3305 ();
 sg13g2_decap_8 FILLER_37_3365 ();
 sg13g2_fill_1 FILLER_37_3372 ();
 sg13g2_fill_1 FILLER_37_3421 ();
 sg13g2_fill_1 FILLER_37_3453 ();
 sg13g2_fill_1 FILLER_37_3467 ();
 sg13g2_decap_8 FILLER_37_3481 ();
 sg13g2_decap_4 FILLER_37_3488 ();
 sg13g2_decap_8 FILLER_37_3529 ();
 sg13g2_decap_8 FILLER_37_3555 ();
 sg13g2_decap_8 FILLER_37_3562 ();
 sg13g2_decap_8 FILLER_37_3569 ();
 sg13g2_fill_2 FILLER_37_3576 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_43 ();
 sg13g2_decap_8 FILLER_38_48 ();
 sg13g2_decap_8 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_fill_2 FILLER_38_73 ();
 sg13g2_fill_1 FILLER_38_75 ();
 sg13g2_fill_1 FILLER_38_89 ();
 sg13g2_fill_2 FILLER_38_94 ();
 sg13g2_fill_1 FILLER_38_96 ();
 sg13g2_decap_4 FILLER_38_110 ();
 sg13g2_fill_1 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_146 ();
 sg13g2_decap_8 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_fill_1 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_252 ();
 sg13g2_decap_4 FILLER_38_262 ();
 sg13g2_fill_1 FILLER_38_266 ();
 sg13g2_fill_2 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_318 ();
 sg13g2_fill_1 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_353 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_362 ();
 sg13g2_fill_2 FILLER_38_416 ();
 sg13g2_decap_8 FILLER_38_423 ();
 sg13g2_decap_8 FILLER_38_430 ();
 sg13g2_decap_4 FILLER_38_437 ();
 sg13g2_decap_8 FILLER_38_469 ();
 sg13g2_decap_4 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_521 ();
 sg13g2_decap_8 FILLER_38_528 ();
 sg13g2_decap_8 FILLER_38_535 ();
 sg13g2_fill_1 FILLER_38_542 ();
 sg13g2_decap_8 FILLER_38_548 ();
 sg13g2_decap_8 FILLER_38_582 ();
 sg13g2_decap_8 FILLER_38_589 ();
 sg13g2_decap_8 FILLER_38_596 ();
 sg13g2_decap_8 FILLER_38_603 ();
 sg13g2_fill_2 FILLER_38_614 ();
 sg13g2_fill_1 FILLER_38_634 ();
 sg13g2_fill_2 FILLER_38_663 ();
 sg13g2_fill_1 FILLER_38_674 ();
 sg13g2_decap_8 FILLER_38_680 ();
 sg13g2_decap_8 FILLER_38_687 ();
 sg13g2_decap_8 FILLER_38_694 ();
 sg13g2_fill_2 FILLER_38_705 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_fill_2 FILLER_38_728 ();
 sg13g2_fill_1 FILLER_38_730 ();
 sg13g2_decap_8 FILLER_38_750 ();
 sg13g2_decap_8 FILLER_38_757 ();
 sg13g2_fill_2 FILLER_38_764 ();
 sg13g2_decap_4 FILLER_38_775 ();
 sg13g2_fill_1 FILLER_38_779 ();
 sg13g2_fill_1 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_874 ();
 sg13g2_decap_8 FILLER_38_881 ();
 sg13g2_decap_8 FILLER_38_888 ();
 sg13g2_decap_8 FILLER_38_895 ();
 sg13g2_decap_8 FILLER_38_902 ();
 sg13g2_decap_8 FILLER_38_909 ();
 sg13g2_fill_1 FILLER_38_916 ();
 sg13g2_decap_8 FILLER_38_942 ();
 sg13g2_fill_1 FILLER_38_949 ();
 sg13g2_fill_2 FILLER_38_962 ();
 sg13g2_decap_8 FILLER_38_967 ();
 sg13g2_fill_2 FILLER_38_974 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_4 FILLER_38_1049 ();
 sg13g2_fill_1 FILLER_38_1053 ();
 sg13g2_fill_1 FILLER_38_1094 ();
 sg13g2_decap_4 FILLER_38_1113 ();
 sg13g2_decap_8 FILLER_38_1123 ();
 sg13g2_decap_8 FILLER_38_1130 ();
 sg13g2_decap_8 FILLER_38_1137 ();
 sg13g2_decap_8 FILLER_38_1144 ();
 sg13g2_decap_4 FILLER_38_1151 ();
 sg13g2_fill_1 FILLER_38_1198 ();
 sg13g2_decap_8 FILLER_38_1212 ();
 sg13g2_decap_8 FILLER_38_1219 ();
 sg13g2_decap_8 FILLER_38_1226 ();
 sg13g2_decap_8 FILLER_38_1233 ();
 sg13g2_decap_8 FILLER_38_1245 ();
 sg13g2_fill_2 FILLER_38_1252 ();
 sg13g2_decap_4 FILLER_38_1294 ();
 sg13g2_fill_1 FILLER_38_1298 ();
 sg13g2_fill_2 FILLER_38_1312 ();
 sg13g2_decap_8 FILLER_38_1320 ();
 sg13g2_decap_4 FILLER_38_1327 ();
 sg13g2_fill_1 FILLER_38_1331 ();
 sg13g2_decap_8 FILLER_38_1336 ();
 sg13g2_decap_8 FILLER_38_1343 ();
 sg13g2_decap_4 FILLER_38_1350 ();
 sg13g2_fill_1 FILLER_38_1390 ();
 sg13g2_fill_1 FILLER_38_1404 ();
 sg13g2_decap_8 FILLER_38_1428 ();
 sg13g2_decap_4 FILLER_38_1435 ();
 sg13g2_fill_1 FILLER_38_1439 ();
 sg13g2_decap_4 FILLER_38_1453 ();
 sg13g2_fill_1 FILLER_38_1457 ();
 sg13g2_decap_4 FILLER_38_1471 ();
 sg13g2_fill_1 FILLER_38_1475 ();
 sg13g2_fill_2 FILLER_38_1495 ();
 sg13g2_fill_1 FILLER_38_1497 ();
 sg13g2_decap_8 FILLER_38_1508 ();
 sg13g2_decap_8 FILLER_38_1515 ();
 sg13g2_fill_2 FILLER_38_1522 ();
 sg13g2_fill_1 FILLER_38_1524 ();
 sg13g2_decap_8 FILLER_38_1534 ();
 sg13g2_fill_2 FILLER_38_1541 ();
 sg13g2_decap_8 FILLER_38_1556 ();
 sg13g2_decap_8 FILLER_38_1563 ();
 sg13g2_decap_4 FILLER_38_1570 ();
 sg13g2_fill_1 FILLER_38_1574 ();
 sg13g2_decap_4 FILLER_38_1591 ();
 sg13g2_decap_8 FILLER_38_1609 ();
 sg13g2_decap_8 FILLER_38_1616 ();
 sg13g2_decap_4 FILLER_38_1623 ();
 sg13g2_fill_2 FILLER_38_1627 ();
 sg13g2_fill_2 FILLER_38_1655 ();
 sg13g2_decap_8 FILLER_38_1665 ();
 sg13g2_decap_4 FILLER_38_1672 ();
 sg13g2_fill_2 FILLER_38_1712 ();
 sg13g2_fill_1 FILLER_38_1714 ();
 sg13g2_fill_2 FILLER_38_1730 ();
 sg13g2_fill_1 FILLER_38_1732 ();
 sg13g2_fill_2 FILLER_38_1751 ();
 sg13g2_fill_1 FILLER_38_1753 ();
 sg13g2_fill_1 FILLER_38_1809 ();
 sg13g2_fill_2 FILLER_38_1817 ();
 sg13g2_decap_8 FILLER_38_1856 ();
 sg13g2_fill_2 FILLER_38_1863 ();
 sg13g2_fill_1 FILLER_38_1877 ();
 sg13g2_decap_8 FILLER_38_1901 ();
 sg13g2_decap_8 FILLER_38_1908 ();
 sg13g2_fill_2 FILLER_38_1915 ();
 sg13g2_fill_1 FILLER_38_1917 ();
 sg13g2_decap_8 FILLER_38_1923 ();
 sg13g2_decap_8 FILLER_38_1930 ();
 sg13g2_fill_1 FILLER_38_1937 ();
 sg13g2_decap_8 FILLER_38_1946 ();
 sg13g2_decap_4 FILLER_38_1953 ();
 sg13g2_fill_2 FILLER_38_1957 ();
 sg13g2_fill_2 FILLER_38_1963 ();
 sg13g2_fill_1 FILLER_38_1965 ();
 sg13g2_decap_8 FILLER_38_1980 ();
 sg13g2_decap_8 FILLER_38_1987 ();
 sg13g2_fill_1 FILLER_38_1994 ();
 sg13g2_decap_8 FILLER_38_1999 ();
 sg13g2_decap_8 FILLER_38_2006 ();
 sg13g2_decap_8 FILLER_38_2013 ();
 sg13g2_decap_8 FILLER_38_2020 ();
 sg13g2_decap_8 FILLER_38_2027 ();
 sg13g2_decap_8 FILLER_38_2034 ();
 sg13g2_fill_1 FILLER_38_2041 ();
 sg13g2_fill_1 FILLER_38_2048 ();
 sg13g2_fill_1 FILLER_38_2066 ();
 sg13g2_fill_2 FILLER_38_2072 ();
 sg13g2_decap_8 FILLER_38_2079 ();
 sg13g2_decap_8 FILLER_38_2086 ();
 sg13g2_decap_4 FILLER_38_2093 ();
 sg13g2_fill_2 FILLER_38_2100 ();
 sg13g2_decap_8 FILLER_38_2106 ();
 sg13g2_decap_4 FILLER_38_2113 ();
 sg13g2_fill_1 FILLER_38_2117 ();
 sg13g2_decap_8 FILLER_38_2126 ();
 sg13g2_decap_8 FILLER_38_2133 ();
 sg13g2_decap_8 FILLER_38_2140 ();
 sg13g2_decap_8 FILLER_38_2147 ();
 sg13g2_decap_4 FILLER_38_2154 ();
 sg13g2_fill_2 FILLER_38_2158 ();
 sg13g2_decap_8 FILLER_38_2164 ();
 sg13g2_decap_8 FILLER_38_2171 ();
 sg13g2_decap_8 FILLER_38_2178 ();
 sg13g2_decap_8 FILLER_38_2185 ();
 sg13g2_decap_8 FILLER_38_2192 ();
 sg13g2_decap_4 FILLER_38_2203 ();
 sg13g2_decap_4 FILLER_38_2215 ();
 sg13g2_fill_1 FILLER_38_2219 ();
 sg13g2_decap_4 FILLER_38_2225 ();
 sg13g2_fill_1 FILLER_38_2229 ();
 sg13g2_decap_4 FILLER_38_2234 ();
 sg13g2_fill_1 FILLER_38_2238 ();
 sg13g2_decap_4 FILLER_38_2249 ();
 sg13g2_decap_8 FILLER_38_2269 ();
 sg13g2_decap_8 FILLER_38_2276 ();
 sg13g2_decap_8 FILLER_38_2283 ();
 sg13g2_fill_2 FILLER_38_2326 ();
 sg13g2_fill_1 FILLER_38_2328 ();
 sg13g2_decap_8 FILLER_38_2383 ();
 sg13g2_decap_8 FILLER_38_2390 ();
 sg13g2_decap_4 FILLER_38_2397 ();
 sg13g2_fill_2 FILLER_38_2463 ();
 sg13g2_fill_1 FILLER_38_2478 ();
 sg13g2_decap_8 FILLER_38_2520 ();
 sg13g2_decap_8 FILLER_38_2527 ();
 sg13g2_decap_8 FILLER_38_2534 ();
 sg13g2_fill_2 FILLER_38_2541 ();
 sg13g2_fill_1 FILLER_38_2582 ();
 sg13g2_decap_8 FILLER_38_2602 ();
 sg13g2_fill_2 FILLER_38_2680 ();
 sg13g2_decap_8 FILLER_38_2732 ();
 sg13g2_decap_4 FILLER_38_2739 ();
 sg13g2_fill_1 FILLER_38_2743 ();
 sg13g2_decap_8 FILLER_38_2801 ();
 sg13g2_fill_1 FILLER_38_2821 ();
 sg13g2_decap_8 FILLER_38_2835 ();
 sg13g2_fill_1 FILLER_38_2842 ();
 sg13g2_decap_8 FILLER_38_2856 ();
 sg13g2_decap_8 FILLER_38_2863 ();
 sg13g2_decap_4 FILLER_38_2870 ();
 sg13g2_fill_1 FILLER_38_2874 ();
 sg13g2_decap_8 FILLER_38_2924 ();
 sg13g2_decap_8 FILLER_38_2931 ();
 sg13g2_fill_2 FILLER_38_2938 ();
 sg13g2_fill_1 FILLER_38_2940 ();
 sg13g2_fill_1 FILLER_38_2967 ();
 sg13g2_decap_4 FILLER_38_2981 ();
 sg13g2_fill_2 FILLER_38_2985 ();
 sg13g2_fill_1 FILLER_38_3036 ();
 sg13g2_fill_2 FILLER_38_3064 ();
 sg13g2_fill_1 FILLER_38_3066 ();
 sg13g2_decap_8 FILLER_38_3072 ();
 sg13g2_decap_8 FILLER_38_3079 ();
 sg13g2_decap_8 FILLER_38_3160 ();
 sg13g2_decap_4 FILLER_38_3167 ();
 sg13g2_fill_1 FILLER_38_3171 ();
 sg13g2_decap_8 FILLER_38_3193 ();
 sg13g2_decap_8 FILLER_38_3200 ();
 sg13g2_decap_8 FILLER_38_3207 ();
 sg13g2_fill_1 FILLER_38_3214 ();
 sg13g2_fill_2 FILLER_38_3242 ();
 sg13g2_fill_1 FILLER_38_3244 ();
 sg13g2_decap_8 FILLER_38_3286 ();
 sg13g2_decap_8 FILLER_38_3293 ();
 sg13g2_fill_2 FILLER_38_3300 ();
 sg13g2_decap_8 FILLER_38_3374 ();
 sg13g2_fill_1 FILLER_38_3381 ();
 sg13g2_fill_2 FILLER_38_3425 ();
 sg13g2_decap_4 FILLER_38_3431 ();
 sg13g2_fill_1 FILLER_38_3435 ();
 sg13g2_decap_8 FILLER_38_3445 ();
 sg13g2_decap_8 FILLER_38_3452 ();
 sg13g2_decap_8 FILLER_38_3462 ();
 sg13g2_decap_4 FILLER_38_3469 ();
 sg13g2_fill_2 FILLER_38_3473 ();
 sg13g2_decap_8 FILLER_38_3479 ();
 sg13g2_decap_8 FILLER_38_3486 ();
 sg13g2_decap_8 FILLER_38_3493 ();
 sg13g2_decap_8 FILLER_38_3500 ();
 sg13g2_decap_4 FILLER_38_3507 ();
 sg13g2_fill_1 FILLER_38_3511 ();
 sg13g2_fill_2 FILLER_38_3531 ();
 sg13g2_decap_8 FILLER_38_3560 ();
 sg13g2_decap_8 FILLER_38_3567 ();
 sg13g2_decap_4 FILLER_38_3574 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_14 ();
 sg13g2_fill_1 FILLER_39_18 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_fill_1 FILLER_39_63 ();
 sg13g2_fill_2 FILLER_39_100 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_decap_8 FILLER_39_107 ();
 sg13g2_decap_4 FILLER_39_114 ();
 sg13g2_fill_1 FILLER_39_118 ();
 sg13g2_fill_2 FILLER_39_137 ();
 sg13g2_fill_1 FILLER_39_139 ();
 sg13g2_fill_2 FILLER_39_149 ();
 sg13g2_fill_1 FILLER_39_160 ();
 sg13g2_decap_8 FILLER_39_165 ();
 sg13g2_decap_8 FILLER_39_172 ();
 sg13g2_decap_8 FILLER_39_179 ();
 sg13g2_fill_1 FILLER_39_186 ();
 sg13g2_decap_4 FILLER_39_197 ();
 sg13g2_fill_2 FILLER_39_201 ();
 sg13g2_decap_4 FILLER_39_213 ();
 sg13g2_fill_1 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_227 ();
 sg13g2_decap_8 FILLER_39_234 ();
 sg13g2_decap_4 FILLER_39_241 ();
 sg13g2_fill_1 FILLER_39_245 ();
 sg13g2_fill_1 FILLER_39_251 ();
 sg13g2_decap_4 FILLER_39_256 ();
 sg13g2_fill_1 FILLER_39_260 ();
 sg13g2_decap_8 FILLER_39_270 ();
 sg13g2_fill_2 FILLER_39_277 ();
 sg13g2_decap_8 FILLER_39_282 ();
 sg13g2_decap_8 FILLER_39_289 ();
 sg13g2_decap_8 FILLER_39_296 ();
 sg13g2_fill_1 FILLER_39_303 ();
 sg13g2_decap_8 FILLER_39_368 ();
 sg13g2_fill_1 FILLER_39_375 ();
 sg13g2_fill_1 FILLER_39_385 ();
 sg13g2_decap_4 FILLER_39_409 ();
 sg13g2_decap_8 FILLER_39_431 ();
 sg13g2_decap_4 FILLER_39_438 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_fill_2 FILLER_39_477 ();
 sg13g2_fill_2 FILLER_39_519 ();
 sg13g2_fill_1 FILLER_39_521 ();
 sg13g2_fill_1 FILLER_39_526 ();
 sg13g2_fill_2 FILLER_39_531 ();
 sg13g2_fill_1 FILLER_39_533 ();
 sg13g2_decap_8 FILLER_39_552 ();
 sg13g2_decap_4 FILLER_39_559 ();
 sg13g2_decap_8 FILLER_39_580 ();
 sg13g2_decap_8 FILLER_39_587 ();
 sg13g2_decap_8 FILLER_39_594 ();
 sg13g2_decap_8 FILLER_39_601 ();
 sg13g2_decap_8 FILLER_39_608 ();
 sg13g2_decap_8 FILLER_39_615 ();
 sg13g2_decap_4 FILLER_39_622 ();
 sg13g2_fill_2 FILLER_39_626 ();
 sg13g2_decap_4 FILLER_39_678 ();
 sg13g2_fill_2 FILLER_39_682 ();
 sg13g2_decap_4 FILLER_39_693 ();
 sg13g2_fill_1 FILLER_39_697 ();
 sg13g2_fill_1 FILLER_39_711 ();
 sg13g2_decap_4 FILLER_39_717 ();
 sg13g2_fill_2 FILLER_39_721 ();
 sg13g2_decap_4 FILLER_39_755 ();
 sg13g2_decap_4 FILLER_39_815 ();
 sg13g2_fill_2 FILLER_39_837 ();
 sg13g2_fill_1 FILLER_39_839 ();
 sg13g2_decap_8 FILLER_39_879 ();
 sg13g2_fill_2 FILLER_39_886 ();
 sg13g2_fill_1 FILLER_39_888 ();
 sg13g2_decap_4 FILLER_39_912 ();
 sg13g2_fill_1 FILLER_39_916 ();
 sg13g2_decap_8 FILLER_39_922 ();
 sg13g2_fill_1 FILLER_39_929 ();
 sg13g2_decap_8 FILLER_39_948 ();
 sg13g2_decap_8 FILLER_39_955 ();
 sg13g2_fill_1 FILLER_39_962 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_decap_4 FILLER_39_979 ();
 sg13g2_fill_2 FILLER_39_983 ();
 sg13g2_fill_1 FILLER_39_989 ();
 sg13g2_fill_2 FILLER_39_1001 ();
 sg13g2_fill_2 FILLER_39_1017 ();
 sg13g2_fill_2 FILLER_39_1028 ();
 sg13g2_fill_2 FILLER_39_1044 ();
 sg13g2_fill_2 FILLER_39_1050 ();
 sg13g2_fill_1 FILLER_39_1052 ();
 sg13g2_fill_2 FILLER_39_1061 ();
 sg13g2_fill_1 FILLER_39_1073 ();
 sg13g2_decap_4 FILLER_39_1083 ();
 sg13g2_decap_8 FILLER_39_1135 ();
 sg13g2_decap_8 FILLER_39_1142 ();
 sg13g2_decap_8 FILLER_39_1159 ();
 sg13g2_fill_1 FILLER_39_1166 ();
 sg13g2_decap_8 FILLER_39_1217 ();
 sg13g2_decap_8 FILLER_39_1224 ();
 sg13g2_decap_4 FILLER_39_1231 ();
 sg13g2_fill_2 FILLER_39_1235 ();
 sg13g2_decap_8 FILLER_39_1278 ();
 sg13g2_decap_8 FILLER_39_1285 ();
 sg13g2_decap_8 FILLER_39_1292 ();
 sg13g2_decap_8 FILLER_39_1299 ();
 sg13g2_decap_8 FILLER_39_1306 ();
 sg13g2_decap_8 FILLER_39_1313 ();
 sg13g2_decap_8 FILLER_39_1320 ();
 sg13g2_fill_1 FILLER_39_1327 ();
 sg13g2_fill_1 FILLER_39_1332 ();
 sg13g2_fill_2 FILLER_39_1338 ();
 sg13g2_fill_1 FILLER_39_1340 ();
 sg13g2_decap_8 FILLER_39_1350 ();
 sg13g2_fill_1 FILLER_39_1357 ();
 sg13g2_fill_2 FILLER_39_1376 ();
 sg13g2_fill_1 FILLER_39_1378 ();
 sg13g2_fill_1 FILLER_39_1396 ();
 sg13g2_fill_1 FILLER_39_1413 ();
 sg13g2_decap_8 FILLER_39_1424 ();
 sg13g2_decap_8 FILLER_39_1431 ();
 sg13g2_decap_8 FILLER_39_1438 ();
 sg13g2_decap_8 FILLER_39_1463 ();
 sg13g2_decap_4 FILLER_39_1479 ();
 sg13g2_decap_8 FILLER_39_1502 ();
 sg13g2_decap_8 FILLER_39_1509 ();
 sg13g2_decap_8 FILLER_39_1516 ();
 sg13g2_decap_8 FILLER_39_1523 ();
 sg13g2_decap_8 FILLER_39_1558 ();
 sg13g2_decap_8 FILLER_39_1565 ();
 sg13g2_decap_8 FILLER_39_1572 ();
 sg13g2_decap_8 FILLER_39_1579 ();
 sg13g2_decap_8 FILLER_39_1591 ();
 sg13g2_fill_2 FILLER_39_1598 ();
 sg13g2_decap_8 FILLER_39_1604 ();
 sg13g2_decap_8 FILLER_39_1611 ();
 sg13g2_decap_8 FILLER_39_1618 ();
 sg13g2_decap_8 FILLER_39_1625 ();
 sg13g2_fill_2 FILLER_39_1632 ();
 sg13g2_fill_1 FILLER_39_1634 ();
 sg13g2_fill_1 FILLER_39_1639 ();
 sg13g2_decap_4 FILLER_39_1652 ();
 sg13g2_fill_2 FILLER_39_1671 ();
 sg13g2_fill_1 FILLER_39_1673 ();
 sg13g2_decap_4 FILLER_39_1684 ();
 sg13g2_fill_2 FILLER_39_1693 ();
 sg13g2_fill_1 FILLER_39_1695 ();
 sg13g2_decap_4 FILLER_39_1701 ();
 sg13g2_fill_2 FILLER_39_1705 ();
 sg13g2_decap_4 FILLER_39_1719 ();
 sg13g2_decap_4 FILLER_39_1727 ();
 sg13g2_fill_2 FILLER_39_1731 ();
 sg13g2_decap_8 FILLER_39_1738 ();
 sg13g2_decap_8 FILLER_39_1745 ();
 sg13g2_decap_8 FILLER_39_1752 ();
 sg13g2_fill_1 FILLER_39_1783 ();
 sg13g2_decap_8 FILLER_39_1814 ();
 sg13g2_fill_2 FILLER_39_1826 ();
 sg13g2_fill_1 FILLER_39_1828 ();
 sg13g2_decap_8 FILLER_39_1839 ();
 sg13g2_decap_8 FILLER_39_1846 ();
 sg13g2_decap_4 FILLER_39_1853 ();
 sg13g2_fill_2 FILLER_39_1863 ();
 sg13g2_fill_1 FILLER_39_1865 ();
 sg13g2_fill_2 FILLER_39_1875 ();
 sg13g2_fill_2 FILLER_39_1898 ();
 sg13g2_fill_1 FILLER_39_1900 ();
 sg13g2_fill_2 FILLER_39_1907 ();
 sg13g2_decap_8 FILLER_39_1913 ();
 sg13g2_fill_2 FILLER_39_1920 ();
 sg13g2_decap_8 FILLER_39_1942 ();
 sg13g2_fill_2 FILLER_39_1949 ();
 sg13g2_fill_1 FILLER_39_1964 ();
 sg13g2_fill_1 FILLER_39_1972 ();
 sg13g2_decap_8 FILLER_39_1989 ();
 sg13g2_decap_4 FILLER_39_1996 ();
 sg13g2_decap_8 FILLER_39_2008 ();
 sg13g2_fill_1 FILLER_39_2015 ();
 sg13g2_decap_4 FILLER_39_2029 ();
 sg13g2_decap_8 FILLER_39_2080 ();
 sg13g2_decap_4 FILLER_39_2087 ();
 sg13g2_fill_2 FILLER_39_2091 ();
 sg13g2_decap_8 FILLER_39_2097 ();
 sg13g2_decap_8 FILLER_39_2104 ();
 sg13g2_decap_4 FILLER_39_2111 ();
 sg13g2_fill_1 FILLER_39_2115 ();
 sg13g2_decap_8 FILLER_39_2135 ();
 sg13g2_fill_2 FILLER_39_2142 ();
 sg13g2_fill_1 FILLER_39_2144 ();
 sg13g2_decap_8 FILLER_39_2149 ();
 sg13g2_decap_8 FILLER_39_2156 ();
 sg13g2_decap_8 FILLER_39_2168 ();
 sg13g2_decap_8 FILLER_39_2175 ();
 sg13g2_decap_8 FILLER_39_2182 ();
 sg13g2_fill_2 FILLER_39_2189 ();
 sg13g2_fill_1 FILLER_39_2191 ();
 sg13g2_decap_4 FILLER_39_2223 ();
 sg13g2_fill_2 FILLER_39_2227 ();
 sg13g2_decap_8 FILLER_39_2233 ();
 sg13g2_decap_4 FILLER_39_2240 ();
 sg13g2_fill_1 FILLER_39_2244 ();
 sg13g2_decap_8 FILLER_39_2268 ();
 sg13g2_decap_8 FILLER_39_2275 ();
 sg13g2_decap_8 FILLER_39_2282 ();
 sg13g2_decap_8 FILLER_39_2289 ();
 sg13g2_fill_2 FILLER_39_2318 ();
 sg13g2_fill_1 FILLER_39_2360 ();
 sg13g2_decap_8 FILLER_39_2387 ();
 sg13g2_fill_1 FILLER_39_2394 ();
 sg13g2_fill_2 FILLER_39_2416 ();
 sg13g2_fill_2 FILLER_39_2456 ();
 sg13g2_fill_1 FILLER_39_2458 ();
 sg13g2_fill_1 FILLER_39_2468 ();
 sg13g2_decap_4 FILLER_39_2482 ();
 sg13g2_decap_8 FILLER_39_2527 ();
 sg13g2_decap_8 FILLER_39_2534 ();
 sg13g2_decap_8 FILLER_39_2541 ();
 sg13g2_fill_2 FILLER_39_2548 ();
 sg13g2_fill_1 FILLER_39_2550 ();
 sg13g2_fill_2 FILLER_39_2565 ();
 sg13g2_fill_1 FILLER_39_2567 ();
 sg13g2_decap_8 FILLER_39_2591 ();
 sg13g2_decap_8 FILLER_39_2598 ();
 sg13g2_decap_8 FILLER_39_2605 ();
 sg13g2_fill_1 FILLER_39_2612 ();
 sg13g2_decap_8 FILLER_39_2637 ();
 sg13g2_decap_8 FILLER_39_2674 ();
 sg13g2_decap_8 FILLER_39_2681 ();
 sg13g2_fill_2 FILLER_39_2702 ();
 sg13g2_fill_2 FILLER_39_2731 ();
 sg13g2_decap_4 FILLER_39_2742 ();
 sg13g2_fill_1 FILLER_39_2746 ();
 sg13g2_decap_4 FILLER_39_2771 ();
 sg13g2_decap_4 FILLER_39_2802 ();
 sg13g2_fill_2 FILLER_39_2832 ();
 sg13g2_fill_1 FILLER_39_2834 ();
 sg13g2_decap_8 FILLER_39_2850 ();
 sg13g2_fill_2 FILLER_39_2857 ();
 sg13g2_fill_1 FILLER_39_2859 ();
 sg13g2_decap_4 FILLER_39_2873 ();
 sg13g2_fill_2 FILLER_39_2904 ();
 sg13g2_decap_8 FILLER_39_2914 ();
 sg13g2_decap_8 FILLER_39_2921 ();
 sg13g2_decap_8 FILLER_39_2928 ();
 sg13g2_fill_2 FILLER_39_2935 ();
 sg13g2_fill_1 FILLER_39_2937 ();
 sg13g2_decap_4 FILLER_39_2951 ();
 sg13g2_fill_1 FILLER_39_2995 ();
 sg13g2_decap_8 FILLER_39_3069 ();
 sg13g2_decap_4 FILLER_39_3076 ();
 sg13g2_fill_1 FILLER_39_3080 ();
 sg13g2_decap_8 FILLER_39_3104 ();
 sg13g2_decap_4 FILLER_39_3111 ();
 sg13g2_fill_2 FILLER_39_3115 ();
 sg13g2_decap_8 FILLER_39_3156 ();
 sg13g2_decap_8 FILLER_39_3163 ();
 sg13g2_decap_8 FILLER_39_3170 ();
 sg13g2_fill_2 FILLER_39_3177 ();
 sg13g2_fill_1 FILLER_39_3179 ();
 sg13g2_decap_8 FILLER_39_3207 ();
 sg13g2_decap_4 FILLER_39_3214 ();
 sg13g2_fill_2 FILLER_39_3218 ();
 sg13g2_fill_1 FILLER_39_3234 ();
 sg13g2_decap_8 FILLER_39_3244 ();
 sg13g2_fill_2 FILLER_39_3251 ();
 sg13g2_decap_8 FILLER_39_3285 ();
 sg13g2_decap_8 FILLER_39_3292 ();
 sg13g2_decap_8 FILLER_39_3299 ();
 sg13g2_fill_2 FILLER_39_3306 ();
 sg13g2_fill_2 FILLER_39_3335 ();
 sg13g2_fill_1 FILLER_39_3337 ();
 sg13g2_decap_8 FILLER_39_3365 ();
 sg13g2_decap_8 FILLER_39_3372 ();
 sg13g2_decap_8 FILLER_39_3379 ();
 sg13g2_decap_8 FILLER_39_3386 ();
 sg13g2_decap_8 FILLER_39_3393 ();
 sg13g2_fill_2 FILLER_39_3404 ();
 sg13g2_decap_8 FILLER_39_3416 ();
 sg13g2_decap_8 FILLER_39_3423 ();
 sg13g2_decap_8 FILLER_39_3430 ();
 sg13g2_decap_8 FILLER_39_3437 ();
 sg13g2_decap_8 FILLER_39_3444 ();
 sg13g2_decap_4 FILLER_39_3451 ();
 sg13g2_decap_8 FILLER_39_3491 ();
 sg13g2_decap_8 FILLER_39_3498 ();
 sg13g2_decap_8 FILLER_39_3505 ();
 sg13g2_fill_2 FILLER_39_3512 ();
 sg13g2_fill_1 FILLER_39_3514 ();
 sg13g2_decap_4 FILLER_39_3573 ();
 sg13g2_fill_1 FILLER_39_3577 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_9 ();
 sg13g2_fill_1 FILLER_40_11 ();
 sg13g2_fill_2 FILLER_40_39 ();
 sg13g2_fill_1 FILLER_40_41 ();
 sg13g2_decap_8 FILLER_40_55 ();
 sg13g2_decap_4 FILLER_40_62 ();
 sg13g2_decap_8 FILLER_40_157 ();
 sg13g2_decap_8 FILLER_40_164 ();
 sg13g2_fill_1 FILLER_40_171 ();
 sg13g2_fill_2 FILLER_40_199 ();
 sg13g2_fill_1 FILLER_40_201 ();
 sg13g2_decap_4 FILLER_40_226 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_fill_2 FILLER_40_321 ();
 sg13g2_fill_1 FILLER_40_323 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_decap_4 FILLER_40_457 ();
 sg13g2_fill_2 FILLER_40_461 ();
 sg13g2_fill_1 FILLER_40_468 ();
 sg13g2_decap_8 FILLER_40_489 ();
 sg13g2_fill_1 FILLER_40_496 ();
 sg13g2_decap_8 FILLER_40_501 ();
 sg13g2_fill_2 FILLER_40_516 ();
 sg13g2_fill_1 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_523 ();
 sg13g2_decap_8 FILLER_40_530 ();
 sg13g2_fill_2 FILLER_40_537 ();
 sg13g2_fill_1 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_568 ();
 sg13g2_decap_4 FILLER_40_575 ();
 sg13g2_fill_2 FILLER_40_579 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_decap_8 FILLER_40_613 ();
 sg13g2_fill_1 FILLER_40_671 ();
 sg13g2_fill_2 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_715 ();
 sg13g2_decap_4 FILLER_40_722 ();
 sg13g2_fill_2 FILLER_40_726 ();
 sg13g2_fill_1 FILLER_40_746 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_fill_2 FILLER_40_862 ();
 sg13g2_decap_8 FILLER_40_884 ();
 sg13g2_fill_1 FILLER_40_891 ();
 sg13g2_fill_2 FILLER_40_899 ();
 sg13g2_decap_4 FILLER_40_915 ();
 sg13g2_fill_2 FILLER_40_919 ();
 sg13g2_fill_2 FILLER_40_947 ();
 sg13g2_decap_4 FILLER_40_955 ();
 sg13g2_decap_8 FILLER_40_972 ();
 sg13g2_decap_8 FILLER_40_979 ();
 sg13g2_decap_8 FILLER_40_986 ();
 sg13g2_decap_8 FILLER_40_993 ();
 sg13g2_decap_4 FILLER_40_1000 ();
 sg13g2_fill_1 FILLER_40_1004 ();
 sg13g2_decap_8 FILLER_40_1022 ();
 sg13g2_decap_8 FILLER_40_1029 ();
 sg13g2_decap_4 FILLER_40_1069 ();
 sg13g2_fill_2 FILLER_40_1073 ();
 sg13g2_decap_8 FILLER_40_1079 ();
 sg13g2_decap_8 FILLER_40_1086 ();
 sg13g2_fill_1 FILLER_40_1093 ();
 sg13g2_fill_1 FILLER_40_1108 ();
 sg13g2_fill_2 FILLER_40_1173 ();
 sg13g2_fill_1 FILLER_40_1175 ();
 sg13g2_decap_8 FILLER_40_1214 ();
 sg13g2_fill_2 FILLER_40_1221 ();
 sg13g2_fill_1 FILLER_40_1223 ();
 sg13g2_decap_4 FILLER_40_1251 ();
 sg13g2_decap_4 FILLER_40_1278 ();
 sg13g2_fill_2 FILLER_40_1282 ();
 sg13g2_fill_2 FILLER_40_1311 ();
 sg13g2_fill_2 FILLER_40_1322 ();
 sg13g2_fill_2 FILLER_40_1333 ();
 sg13g2_decap_8 FILLER_40_1358 ();
 sg13g2_decap_8 FILLER_40_1365 ();
 sg13g2_fill_1 FILLER_40_1372 ();
 sg13g2_decap_4 FILLER_40_1396 ();
 sg13g2_fill_2 FILLER_40_1400 ();
 sg13g2_decap_8 FILLER_40_1419 ();
 sg13g2_decap_8 FILLER_40_1426 ();
 sg13g2_decap_8 FILLER_40_1433 ();
 sg13g2_fill_1 FILLER_40_1477 ();
 sg13g2_fill_2 FILLER_40_1486 ();
 sg13g2_fill_1 FILLER_40_1488 ();
 sg13g2_decap_8 FILLER_40_1510 ();
 sg13g2_decap_8 FILLER_40_1517 ();
 sg13g2_decap_4 FILLER_40_1524 ();
 sg13g2_fill_1 FILLER_40_1528 ();
 sg13g2_decap_4 FILLER_40_1575 ();
 sg13g2_fill_1 FILLER_40_1579 ();
 sg13g2_decap_8 FILLER_40_1585 ();
 sg13g2_decap_4 FILLER_40_1592 ();
 sg13g2_fill_1 FILLER_40_1596 ();
 sg13g2_fill_2 FILLER_40_1621 ();
 sg13g2_fill_1 FILLER_40_1623 ();
 sg13g2_decap_8 FILLER_40_1630 ();
 sg13g2_decap_8 FILLER_40_1637 ();
 sg13g2_decap_4 FILLER_40_1644 ();
 sg13g2_fill_1 FILLER_40_1648 ();
 sg13g2_decap_4 FILLER_40_1670 ();
 sg13g2_decap_8 FILLER_40_1685 ();
 sg13g2_decap_8 FILLER_40_1692 ();
 sg13g2_decap_8 FILLER_40_1699 ();
 sg13g2_decap_4 FILLER_40_1706 ();
 sg13g2_fill_1 FILLER_40_1710 ();
 sg13g2_fill_2 FILLER_40_1728 ();
 sg13g2_fill_1 FILLER_40_1730 ();
 sg13g2_decap_8 FILLER_40_1740 ();
 sg13g2_decap_8 FILLER_40_1747 ();
 sg13g2_decap_8 FILLER_40_1754 ();
 sg13g2_fill_2 FILLER_40_1761 ();
 sg13g2_fill_1 FILLER_40_1763 ();
 sg13g2_decap_8 FILLER_40_1801 ();
 sg13g2_decap_8 FILLER_40_1808 ();
 sg13g2_decap_8 FILLER_40_1815 ();
 sg13g2_decap_8 FILLER_40_1822 ();
 sg13g2_decap_8 FILLER_40_1829 ();
 sg13g2_decap_4 FILLER_40_1836 ();
 sg13g2_decap_8 FILLER_40_1855 ();
 sg13g2_decap_4 FILLER_40_1862 ();
 sg13g2_fill_1 FILLER_40_1866 ();
 sg13g2_fill_2 FILLER_40_1872 ();
 sg13g2_fill_1 FILLER_40_1874 ();
 sg13g2_fill_2 FILLER_40_1888 ();
 sg13g2_fill_2 FILLER_40_1905 ();
 sg13g2_decap_8 FILLER_40_1912 ();
 sg13g2_fill_2 FILLER_40_1919 ();
 sg13g2_decap_8 FILLER_40_1936 ();
 sg13g2_fill_1 FILLER_40_1943 ();
 sg13g2_decap_4 FILLER_40_1989 ();
 sg13g2_fill_1 FILLER_40_1993 ();
 sg13g2_fill_2 FILLER_40_2001 ();
 sg13g2_fill_1 FILLER_40_2003 ();
 sg13g2_decap_8 FILLER_40_2017 ();
 sg13g2_decap_4 FILLER_40_2024 ();
 sg13g2_fill_2 FILLER_40_2028 ();
 sg13g2_fill_2 FILLER_40_2039 ();
 sg13g2_fill_1 FILLER_40_2041 ();
 sg13g2_decap_4 FILLER_40_2087 ();
 sg13g2_fill_1 FILLER_40_2091 ();
 sg13g2_fill_1 FILLER_40_2097 ();
 sg13g2_decap_4 FILLER_40_2111 ();
 sg13g2_fill_2 FILLER_40_2115 ();
 sg13g2_fill_1 FILLER_40_2123 ();
 sg13g2_decap_8 FILLER_40_2137 ();
 sg13g2_decap_8 FILLER_40_2144 ();
 sg13g2_decap_8 FILLER_40_2151 ();
 sg13g2_decap_8 FILLER_40_2158 ();
 sg13g2_decap_8 FILLER_40_2165 ();
 sg13g2_fill_2 FILLER_40_2172 ();
 sg13g2_decap_4 FILLER_40_2232 ();
 sg13g2_fill_1 FILLER_40_2236 ();
 sg13g2_decap_8 FILLER_40_2241 ();
 sg13g2_decap_8 FILLER_40_2248 ();
 sg13g2_decap_8 FILLER_40_2265 ();
 sg13g2_decap_8 FILLER_40_2272 ();
 sg13g2_decap_4 FILLER_40_2279 ();
 sg13g2_fill_1 FILLER_40_2283 ();
 sg13g2_fill_2 FILLER_40_2312 ();
 sg13g2_fill_2 FILLER_40_2341 ();
 sg13g2_fill_1 FILLER_40_2343 ();
 sg13g2_decap_8 FILLER_40_2380 ();
 sg13g2_decap_8 FILLER_40_2387 ();
 sg13g2_fill_2 FILLER_40_2394 ();
 sg13g2_decap_4 FILLER_40_2425 ();
 sg13g2_fill_1 FILLER_40_2429 ();
 sg13g2_decap_8 FILLER_40_2440 ();
 sg13g2_decap_8 FILLER_40_2447 ();
 sg13g2_decap_8 FILLER_40_2454 ();
 sg13g2_decap_8 FILLER_40_2485 ();
 sg13g2_fill_1 FILLER_40_2492 ();
 sg13g2_fill_2 FILLER_40_2527 ();
 sg13g2_fill_1 FILLER_40_2529 ();
 sg13g2_fill_1 FILLER_40_2534 ();
 sg13g2_fill_1 FILLER_40_2545 ();
 sg13g2_fill_2 FILLER_40_2555 ();
 sg13g2_decap_8 FILLER_40_2584 ();
 sg13g2_decap_8 FILLER_40_2591 ();
 sg13g2_decap_8 FILLER_40_2598 ();
 sg13g2_decap_4 FILLER_40_2605 ();
 sg13g2_fill_1 FILLER_40_2609 ();
 sg13g2_fill_2 FILLER_40_2623 ();
 sg13g2_fill_2 FILLER_40_2638 ();
 sg13g2_fill_2 FILLER_40_2653 ();
 sg13g2_fill_1 FILLER_40_2655 ();
 sg13g2_decap_8 FILLER_40_2669 ();
 sg13g2_decap_8 FILLER_40_2676 ();
 sg13g2_fill_2 FILLER_40_2683 ();
 sg13g2_decap_4 FILLER_40_2711 ();
 sg13g2_decap_8 FILLER_40_2728 ();
 sg13g2_decap_8 FILLER_40_2735 ();
 sg13g2_decap_8 FILLER_40_2755 ();
 sg13g2_decap_8 FILLER_40_2762 ();
 sg13g2_decap_8 FILLER_40_2769 ();
 sg13g2_decap_8 FILLER_40_2776 ();
 sg13g2_fill_2 FILLER_40_2783 ();
 sg13g2_decap_4 FILLER_40_2788 ();
 sg13g2_fill_1 FILLER_40_2792 ();
 sg13g2_decap_8 FILLER_40_2797 ();
 sg13g2_fill_1 FILLER_40_2804 ();
 sg13g2_fill_2 FILLER_40_2828 ();
 sg13g2_fill_2 FILLER_40_2856 ();
 sg13g2_decap_8 FILLER_40_2871 ();
 sg13g2_decap_8 FILLER_40_2878 ();
 sg13g2_decap_8 FILLER_40_2898 ();
 sg13g2_decap_8 FILLER_40_2905 ();
 sg13g2_decap_8 FILLER_40_2912 ();
 sg13g2_decap_4 FILLER_40_2919 ();
 sg13g2_fill_2 FILLER_40_2923 ();
 sg13g2_fill_2 FILLER_40_2938 ();
 sg13g2_fill_1 FILLER_40_2940 ();
 sg13g2_fill_1 FILLER_40_2954 ();
 sg13g2_fill_1 FILLER_40_2982 ();
 sg13g2_decap_4 FILLER_40_3000 ();
 sg13g2_fill_1 FILLER_40_3004 ();
 sg13g2_decap_8 FILLER_40_3069 ();
 sg13g2_decap_4 FILLER_40_3076 ();
 sg13g2_fill_2 FILLER_40_3080 ();
 sg13g2_decap_8 FILLER_40_3103 ();
 sg13g2_decap_4 FILLER_40_3110 ();
 sg13g2_fill_2 FILLER_40_3114 ();
 sg13g2_fill_1 FILLER_40_3125 ();
 sg13g2_decap_4 FILLER_40_3139 ();
 sg13g2_fill_1 FILLER_40_3143 ();
 sg13g2_decap_8 FILLER_40_3202 ();
 sg13g2_decap_8 FILLER_40_3209 ();
 sg13g2_decap_8 FILLER_40_3216 ();
 sg13g2_decap_8 FILLER_40_3223 ();
 sg13g2_decap_4 FILLER_40_3230 ();
 sg13g2_decap_4 FILLER_40_3238 ();
 sg13g2_fill_1 FILLER_40_3242 ();
 sg13g2_decap_4 FILLER_40_3256 ();
 sg13g2_fill_2 FILLER_40_3260 ();
 sg13g2_decap_8 FILLER_40_3279 ();
 sg13g2_decap_8 FILLER_40_3299 ();
 sg13g2_decap_8 FILLER_40_3306 ();
 sg13g2_decap_4 FILLER_40_3313 ();
 sg13g2_fill_2 FILLER_40_3317 ();
 sg13g2_decap_4 FILLER_40_3332 ();
 sg13g2_fill_2 FILLER_40_3336 ();
 sg13g2_decap_8 FILLER_40_3364 ();
 sg13g2_decap_4 FILLER_40_3371 ();
 sg13g2_decap_4 FILLER_40_3388 ();
 sg13g2_fill_2 FILLER_40_3392 ();
 sg13g2_fill_2 FILLER_40_3425 ();
 sg13g2_fill_1 FILLER_40_3427 ();
 sg13g2_decap_8 FILLER_40_3437 ();
 sg13g2_decap_8 FILLER_40_3444 ();
 sg13g2_decap_8 FILLER_40_3505 ();
 sg13g2_decap_8 FILLER_40_3512 ();
 sg13g2_decap_4 FILLER_40_3519 ();
 sg13g2_fill_2 FILLER_40_3554 ();
 sg13g2_decap_8 FILLER_40_3569 ();
 sg13g2_fill_2 FILLER_40_3576 ();
 sg13g2_fill_2 FILLER_41_112 ();
 sg13g2_fill_2 FILLER_41_146 ();
 sg13g2_fill_1 FILLER_41_148 ();
 sg13g2_decap_4 FILLER_41_166 ();
 sg13g2_fill_1 FILLER_41_170 ();
 sg13g2_decap_4 FILLER_41_225 ();
 sg13g2_fill_1 FILLER_41_229 ();
 sg13g2_fill_2 FILLER_41_259 ();
 sg13g2_fill_1 FILLER_41_261 ();
 sg13g2_fill_2 FILLER_41_277 ();
 sg13g2_decap_8 FILLER_41_289 ();
 sg13g2_decap_8 FILLER_41_296 ();
 sg13g2_decap_8 FILLER_41_303 ();
 sg13g2_decap_8 FILLER_41_310 ();
 sg13g2_decap_8 FILLER_41_317 ();
 sg13g2_decap_8 FILLER_41_324 ();
 sg13g2_fill_2 FILLER_41_331 ();
 sg13g2_decap_8 FILLER_41_360 ();
 sg13g2_decap_8 FILLER_41_367 ();
 sg13g2_decap_8 FILLER_41_374 ();
 sg13g2_decap_8 FILLER_41_381 ();
 sg13g2_decap_8 FILLER_41_388 ();
 sg13g2_fill_2 FILLER_41_395 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_decap_8 FILLER_41_439 ();
 sg13g2_decap_4 FILLER_41_446 ();
 sg13g2_fill_2 FILLER_41_450 ();
 sg13g2_decap_8 FILLER_41_457 ();
 sg13g2_decap_8 FILLER_41_464 ();
 sg13g2_decap_8 FILLER_41_471 ();
 sg13g2_fill_1 FILLER_41_478 ();
 sg13g2_decap_8 FILLER_41_484 ();
 sg13g2_fill_2 FILLER_41_491 ();
 sg13g2_fill_1 FILLER_41_493 ();
 sg13g2_fill_1 FILLER_41_503 ();
 sg13g2_fill_1 FILLER_41_517 ();
 sg13g2_fill_2 FILLER_41_528 ();
 sg13g2_decap_8 FILLER_41_534 ();
 sg13g2_fill_2 FILLER_41_541 ();
 sg13g2_fill_1 FILLER_41_543 ();
 sg13g2_fill_2 FILLER_41_575 ();
 sg13g2_decap_4 FILLER_41_605 ();
 sg13g2_fill_1 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_615 ();
 sg13g2_decap_8 FILLER_41_654 ();
 sg13g2_fill_2 FILLER_41_661 ();
 sg13g2_fill_1 FILLER_41_663 ();
 sg13g2_fill_1 FILLER_41_667 ();
 sg13g2_decap_8 FILLER_41_695 ();
 sg13g2_decap_8 FILLER_41_702 ();
 sg13g2_decap_8 FILLER_41_709 ();
 sg13g2_fill_2 FILLER_41_716 ();
 sg13g2_fill_1 FILLER_41_718 ();
 sg13g2_decap_8 FILLER_41_738 ();
 sg13g2_decap_8 FILLER_41_745 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_fill_2 FILLER_41_789 ();
 sg13g2_fill_2 FILLER_41_800 ();
 sg13g2_fill_1 FILLER_41_802 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_decap_8 FILLER_41_821 ();
 sg13g2_fill_1 FILLER_41_874 ();
 sg13g2_decap_8 FILLER_41_884 ();
 sg13g2_fill_2 FILLER_41_891 ();
 sg13g2_fill_1 FILLER_41_893 ();
 sg13g2_decap_8 FILLER_41_916 ();
 sg13g2_decap_8 FILLER_41_923 ();
 sg13g2_fill_2 FILLER_41_930 ();
 sg13g2_decap_8 FILLER_41_975 ();
 sg13g2_decap_8 FILLER_41_982 ();
 sg13g2_decap_8 FILLER_41_989 ();
 sg13g2_decap_4 FILLER_41_996 ();
 sg13g2_fill_2 FILLER_41_1013 ();
 sg13g2_decap_8 FILLER_41_1019 ();
 sg13g2_decap_8 FILLER_41_1026 ();
 sg13g2_decap_8 FILLER_41_1033 ();
 sg13g2_decap_8 FILLER_41_1040 ();
 sg13g2_decap_8 FILLER_41_1047 ();
 sg13g2_decap_8 FILLER_41_1054 ();
 sg13g2_fill_2 FILLER_41_1061 ();
 sg13g2_fill_1 FILLER_41_1063 ();
 sg13g2_decap_8 FILLER_41_1073 ();
 sg13g2_decap_8 FILLER_41_1080 ();
 sg13g2_decap_8 FILLER_41_1087 ();
 sg13g2_fill_1 FILLER_41_1094 ();
 sg13g2_fill_1 FILLER_41_1103 ();
 sg13g2_decap_8 FILLER_41_1127 ();
 sg13g2_decap_4 FILLER_41_1134 ();
 sg13g2_fill_1 FILLER_41_1138 ();
 sg13g2_decap_8 FILLER_41_1168 ();
 sg13g2_decap_8 FILLER_41_1175 ();
 sg13g2_fill_1 FILLER_41_1182 ();
 sg13g2_fill_1 FILLER_41_1187 ();
 sg13g2_decap_8 FILLER_41_1207 ();
 sg13g2_decap_4 FILLER_41_1214 ();
 sg13g2_fill_1 FILLER_41_1218 ();
 sg13g2_decap_8 FILLER_41_1225 ();
 sg13g2_decap_4 FILLER_41_1232 ();
 sg13g2_decap_4 FILLER_41_1264 ();
 sg13g2_fill_1 FILLER_41_1268 ();
 sg13g2_decap_8 FILLER_41_1282 ();
 sg13g2_fill_1 FILLER_41_1289 ();
 sg13g2_fill_2 FILLER_41_1300 ();
 sg13g2_fill_2 FILLER_41_1317 ();
 sg13g2_fill_1 FILLER_41_1319 ();
 sg13g2_decap_8 FILLER_41_1356 ();
 sg13g2_decap_8 FILLER_41_1363 ();
 sg13g2_decap_4 FILLER_41_1370 ();
 sg13g2_decap_4 FILLER_41_1420 ();
 sg13g2_decap_8 FILLER_41_1457 ();
 sg13g2_decap_4 FILLER_41_1464 ();
 sg13g2_decap_8 FILLER_41_1511 ();
 sg13g2_decap_4 FILLER_41_1518 ();
 sg13g2_decap_8 FILLER_41_1536 ();
 sg13g2_decap_8 FILLER_41_1543 ();
 sg13g2_fill_2 FILLER_41_1550 ();
 sg13g2_fill_1 FILLER_41_1565 ();
 sg13g2_fill_2 FILLER_41_1578 ();
 sg13g2_decap_8 FILLER_41_1588 ();
 sg13g2_decap_8 FILLER_41_1595 ();
 sg13g2_decap_8 FILLER_41_1602 ();
 sg13g2_fill_1 FILLER_41_1609 ();
 sg13g2_decap_8 FILLER_41_1633 ();
 sg13g2_decap_8 FILLER_41_1640 ();
 sg13g2_decap_8 FILLER_41_1647 ();
 sg13g2_decap_8 FILLER_41_1654 ();
 sg13g2_fill_2 FILLER_41_1661 ();
 sg13g2_fill_1 FILLER_41_1663 ();
 sg13g2_decap_8 FILLER_41_1694 ();
 sg13g2_fill_2 FILLER_41_1701 ();
 sg13g2_fill_1 FILLER_41_1703 ();
 sg13g2_decap_8 FILLER_41_1746 ();
 sg13g2_decap_8 FILLER_41_1753 ();
 sg13g2_decap_8 FILLER_41_1760 ();
 sg13g2_decap_8 FILLER_41_1767 ();
 sg13g2_decap_4 FILLER_41_1774 ();
 sg13g2_fill_2 FILLER_41_1778 ();
 sg13g2_decap_8 FILLER_41_1799 ();
 sg13g2_decap_8 FILLER_41_1806 ();
 sg13g2_decap_8 FILLER_41_1813 ();
 sg13g2_decap_8 FILLER_41_1820 ();
 sg13g2_fill_2 FILLER_41_1827 ();
 sg13g2_fill_2 FILLER_41_1838 ();
 sg13g2_fill_1 FILLER_41_1845 ();
 sg13g2_decap_8 FILLER_41_1859 ();
 sg13g2_decap_8 FILLER_41_1866 ();
 sg13g2_decap_8 FILLER_41_1873 ();
 sg13g2_fill_2 FILLER_41_1891 ();
 sg13g2_fill_1 FILLER_41_1903 ();
 sg13g2_fill_1 FILLER_41_1909 ();
 sg13g2_decap_8 FILLER_41_1916 ();
 sg13g2_decap_8 FILLER_41_1923 ();
 sg13g2_decap_8 FILLER_41_1930 ();
 sg13g2_decap_8 FILLER_41_1937 ();
 sg13g2_fill_2 FILLER_41_1944 ();
 sg13g2_decap_8 FILLER_41_1987 ();
 sg13g2_fill_1 FILLER_41_1994 ();
 sg13g2_decap_4 FILLER_41_2003 ();
 sg13g2_decap_8 FILLER_41_2015 ();
 sg13g2_fill_2 FILLER_41_2022 ();
 sg13g2_fill_1 FILLER_41_2024 ();
 sg13g2_fill_1 FILLER_41_2038 ();
 sg13g2_fill_1 FILLER_41_2065 ();
 sg13g2_decap_8 FILLER_41_2073 ();
 sg13g2_decap_8 FILLER_41_2080 ();
 sg13g2_decap_8 FILLER_41_2087 ();
 sg13g2_decap_8 FILLER_41_2094 ();
 sg13g2_fill_1 FILLER_41_2101 ();
 sg13g2_decap_8 FILLER_41_2105 ();
 sg13g2_decap_8 FILLER_41_2112 ();
 sg13g2_fill_2 FILLER_41_2119 ();
 sg13g2_fill_1 FILLER_41_2125 ();
 sg13g2_decap_8 FILLER_41_2154 ();
 sg13g2_decap_8 FILLER_41_2161 ();
 sg13g2_decap_4 FILLER_41_2176 ();
 sg13g2_decap_8 FILLER_41_2223 ();
 sg13g2_decap_8 FILLER_41_2253 ();
 sg13g2_decap_8 FILLER_41_2260 ();
 sg13g2_decap_8 FILLER_41_2267 ();
 sg13g2_decap_8 FILLER_41_2274 ();
 sg13g2_decap_4 FILLER_41_2309 ();
 sg13g2_fill_2 FILLER_41_2313 ();
 sg13g2_decap_8 FILLER_41_2319 ();
 sg13g2_decap_8 FILLER_41_2326 ();
 sg13g2_decap_4 FILLER_41_2333 ();
 sg13g2_fill_1 FILLER_41_2337 ();
 sg13g2_decap_8 FILLER_41_2368 ();
 sg13g2_decap_8 FILLER_41_2375 ();
 sg13g2_fill_1 FILLER_41_2382 ();
 sg13g2_decap_8 FILLER_41_2424 ();
 sg13g2_decap_8 FILLER_41_2431 ();
 sg13g2_decap_8 FILLER_41_2438 ();
 sg13g2_decap_8 FILLER_41_2445 ();
 sg13g2_fill_2 FILLER_41_2452 ();
 sg13g2_fill_1 FILLER_41_2454 ();
 sg13g2_fill_2 FILLER_41_2492 ();
 sg13g2_fill_2 FILLER_41_2552 ();
 sg13g2_decap_4 FILLER_41_2568 ();
 sg13g2_decap_8 FILLER_41_2599 ();
 sg13g2_decap_4 FILLER_41_2606 ();
 sg13g2_fill_2 FILLER_41_2610 ();
 sg13g2_decap_8 FILLER_41_2625 ();
 sg13g2_fill_1 FILLER_41_2632 ();
 sg13g2_fill_2 FILLER_41_2672 ();
 sg13g2_fill_1 FILLER_41_2674 ();
 sg13g2_decap_8 FILLER_41_2727 ();
 sg13g2_decap_4 FILLER_41_2734 ();
 sg13g2_fill_1 FILLER_41_2738 ();
 sg13g2_fill_2 FILLER_41_2762 ();
 sg13g2_decap_4 FILLER_41_2773 ();
 sg13g2_fill_2 FILLER_41_2777 ();
 sg13g2_decap_4 FILLER_41_2811 ();
 sg13g2_fill_2 FILLER_41_2815 ();
 sg13g2_decap_4 FILLER_41_2827 ();
 sg13g2_fill_1 FILLER_41_2883 ();
 sg13g2_decap_8 FILLER_41_2897 ();
 sg13g2_fill_2 FILLER_41_2904 ();
 sg13g2_fill_2 FILLER_41_2919 ();
 sg13g2_decap_8 FILLER_41_2934 ();
 sg13g2_decap_4 FILLER_41_3004 ();
 sg13g2_fill_2 FILLER_41_3008 ();
 sg13g2_decap_4 FILLER_41_3014 ();
 sg13g2_fill_1 FILLER_41_3018 ();
 sg13g2_decap_4 FILLER_41_3046 ();
 sg13g2_decap_4 FILLER_41_3059 ();
 sg13g2_decap_4 FILLER_41_3067 ();
 sg13g2_fill_2 FILLER_41_3148 ();
 sg13g2_decap_8 FILLER_41_3208 ();
 sg13g2_decap_8 FILLER_41_3215 ();
 sg13g2_decap_4 FILLER_41_3222 ();
 sg13g2_decap_8 FILLER_41_3276 ();
 sg13g2_fill_2 FILLER_41_3283 ();
 sg13g2_fill_1 FILLER_41_3285 ();
 sg13g2_decap_8 FILLER_41_3312 ();
 sg13g2_decap_4 FILLER_41_3319 ();
 sg13g2_decap_4 FILLER_41_3363 ();
 sg13g2_fill_1 FILLER_41_3367 ();
 sg13g2_decap_4 FILLER_41_3378 ();
 sg13g2_decap_4 FILLER_41_3446 ();
 sg13g2_fill_1 FILLER_41_3468 ();
 sg13g2_decap_8 FILLER_41_3506 ();
 sg13g2_decap_8 FILLER_41_3513 ();
 sg13g2_decap_8 FILLER_41_3520 ();
 sg13g2_decap_4 FILLER_41_3527 ();
 sg13g2_decap_4 FILLER_41_3572 ();
 sg13g2_fill_2 FILLER_41_3576 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_fill_2 FILLER_42_49 ();
 sg13g2_fill_2 FILLER_42_108 ();
 sg13g2_fill_1 FILLER_42_110 ();
 sg13g2_decap_8 FILLER_42_160 ();
 sg13g2_decap_4 FILLER_42_167 ();
 sg13g2_fill_1 FILLER_42_171 ();
 sg13g2_fill_2 FILLER_42_199 ();
 sg13g2_fill_1 FILLER_42_201 ();
 sg13g2_fill_2 FILLER_42_226 ();
 sg13g2_fill_2 FILLER_42_255 ();
 sg13g2_decap_8 FILLER_42_290 ();
 sg13g2_decap_8 FILLER_42_297 ();
 sg13g2_fill_2 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_314 ();
 sg13g2_decap_8 FILLER_42_330 ();
 sg13g2_decap_4 FILLER_42_337 ();
 sg13g2_fill_2 FILLER_42_341 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_2 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_410 ();
 sg13g2_fill_1 FILLER_42_439 ();
 sg13g2_decap_8 FILLER_42_467 ();
 sg13g2_decap_8 FILLER_42_474 ();
 sg13g2_fill_2 FILLER_42_481 ();
 sg13g2_fill_1 FILLER_42_483 ();
 sg13g2_fill_2 FILLER_42_491 ();
 sg13g2_fill_2 FILLER_42_498 ();
 sg13g2_fill_1 FILLER_42_525 ();
 sg13g2_decap_8 FILLER_42_531 ();
 sg13g2_decap_8 FILLER_42_538 ();
 sg13g2_fill_2 FILLER_42_545 ();
 sg13g2_fill_1 FILLER_42_547 ();
 sg13g2_fill_1 FILLER_42_579 ();
 sg13g2_decap_4 FILLER_42_598 ();
 sg13g2_fill_1 FILLER_42_602 ();
 sg13g2_fill_2 FILLER_42_616 ();
 sg13g2_fill_1 FILLER_42_618 ();
 sg13g2_decap_4 FILLER_42_624 ();
 sg13g2_fill_1 FILLER_42_628 ();
 sg13g2_fill_1 FILLER_42_639 ();
 sg13g2_decap_8 FILLER_42_654 ();
 sg13g2_decap_4 FILLER_42_661 ();
 sg13g2_fill_2 FILLER_42_665 ();
 sg13g2_fill_2 FILLER_42_676 ();
 sg13g2_fill_1 FILLER_42_678 ();
 sg13g2_decap_8 FILLER_42_682 ();
 sg13g2_decap_8 FILLER_42_689 ();
 sg13g2_decap_8 FILLER_42_696 ();
 sg13g2_decap_8 FILLER_42_703 ();
 sg13g2_decap_4 FILLER_42_710 ();
 sg13g2_fill_1 FILLER_42_747 ();
 sg13g2_decap_8 FILLER_42_762 ();
 sg13g2_decap_8 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_4 FILLER_42_819 ();
 sg13g2_fill_2 FILLER_42_823 ();
 sg13g2_fill_1 FILLER_42_877 ();
 sg13g2_decap_8 FILLER_42_881 ();
 sg13g2_decap_4 FILLER_42_888 ();
 sg13g2_fill_2 FILLER_42_892 ();
 sg13g2_fill_2 FILLER_42_919 ();
 sg13g2_fill_2 FILLER_42_928 ();
 sg13g2_fill_1 FILLER_42_930 ();
 sg13g2_decap_8 FILLER_42_941 ();
 sg13g2_decap_8 FILLER_42_983 ();
 sg13g2_fill_1 FILLER_42_990 ();
 sg13g2_decap_4 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_42_1041 ();
 sg13g2_decap_8 FILLER_42_1048 ();
 sg13g2_decap_8 FILLER_42_1055 ();
 sg13g2_decap_8 FILLER_42_1062 ();
 sg13g2_fill_2 FILLER_42_1069 ();
 sg13g2_fill_1 FILLER_42_1071 ();
 sg13g2_decap_8 FILLER_42_1077 ();
 sg13g2_decap_4 FILLER_42_1084 ();
 sg13g2_decap_4 FILLER_42_1092 ();
 sg13g2_fill_1 FILLER_42_1096 ();
 sg13g2_fill_2 FILLER_42_1114 ();
 sg13g2_decap_8 FILLER_42_1134 ();
 sg13g2_decap_4 FILLER_42_1141 ();
 sg13g2_fill_2 FILLER_42_1145 ();
 sg13g2_decap_8 FILLER_42_1152 ();
 sg13g2_fill_2 FILLER_42_1159 ();
 sg13g2_decap_8 FILLER_42_1165 ();
 sg13g2_fill_2 FILLER_42_1172 ();
 sg13g2_decap_8 FILLER_42_1183 ();
 sg13g2_decap_4 FILLER_42_1190 ();
 sg13g2_decap_8 FILLER_42_1213 ();
 sg13g2_decap_8 FILLER_42_1220 ();
 sg13g2_decap_4 FILLER_42_1227 ();
 sg13g2_decap_4 FILLER_42_1234 ();
 sg13g2_fill_2 FILLER_42_1248 ();
 sg13g2_fill_2 FILLER_42_1255 ();
 sg13g2_fill_1 FILLER_42_1274 ();
 sg13g2_fill_2 FILLER_42_1283 ();
 sg13g2_fill_1 FILLER_42_1285 ();
 sg13g2_fill_1 FILLER_42_1299 ();
 sg13g2_fill_2 FILLER_42_1311 ();
 sg13g2_fill_1 FILLER_42_1313 ();
 sg13g2_fill_1 FILLER_42_1319 ();
 sg13g2_decap_4 FILLER_42_1332 ();
 sg13g2_fill_2 FILLER_42_1336 ();
 sg13g2_fill_2 FILLER_42_1352 ();
 sg13g2_fill_1 FILLER_42_1354 ();
 sg13g2_decap_8 FILLER_42_1364 ();
 sg13g2_fill_2 FILLER_42_1371 ();
 sg13g2_decap_8 FILLER_42_1415 ();
 sg13g2_decap_8 FILLER_42_1422 ();
 sg13g2_decap_8 FILLER_42_1429 ();
 sg13g2_decap_8 FILLER_42_1444 ();
 sg13g2_decap_8 FILLER_42_1451 ();
 sg13g2_fill_1 FILLER_42_1458 ();
 sg13g2_fill_2 FILLER_42_1486 ();
 sg13g2_fill_1 FILLER_42_1488 ();
 sg13g2_decap_8 FILLER_42_1513 ();
 sg13g2_decap_8 FILLER_42_1520 ();
 sg13g2_decap_4 FILLER_42_1527 ();
 sg13g2_fill_2 FILLER_42_1531 ();
 sg13g2_fill_2 FILLER_42_1539 ();
 sg13g2_decap_4 FILLER_42_1548 ();
 sg13g2_fill_2 FILLER_42_1552 ();
 sg13g2_fill_2 FILLER_42_1595 ();
 sg13g2_fill_1 FILLER_42_1597 ();
 sg13g2_decap_8 FILLER_42_1606 ();
 sg13g2_fill_1 FILLER_42_1613 ();
 sg13g2_decap_8 FILLER_42_1637 ();
 sg13g2_decap_8 FILLER_42_1644 ();
 sg13g2_decap_8 FILLER_42_1651 ();
 sg13g2_decap_8 FILLER_42_1658 ();
 sg13g2_fill_2 FILLER_42_1670 ();
 sg13g2_decap_8 FILLER_42_1685 ();
 sg13g2_decap_8 FILLER_42_1692 ();
 sg13g2_decap_8 FILLER_42_1699 ();
 sg13g2_decap_8 FILLER_42_1706 ();
 sg13g2_decap_8 FILLER_42_1752 ();
 sg13g2_decap_4 FILLER_42_1759 ();
 sg13g2_fill_2 FILLER_42_1763 ();
 sg13g2_fill_1 FILLER_42_1771 ();
 sg13g2_fill_2 FILLER_42_1778 ();
 sg13g2_fill_1 FILLER_42_1780 ();
 sg13g2_decap_8 FILLER_42_1787 ();
 sg13g2_fill_1 FILLER_42_1794 ();
 sg13g2_decap_4 FILLER_42_1813 ();
 sg13g2_fill_1 FILLER_42_1817 ();
 sg13g2_decap_8 FILLER_42_1864 ();
 sg13g2_decap_8 FILLER_42_1871 ();
 sg13g2_decap_8 FILLER_42_1878 ();
 sg13g2_decap_8 FILLER_42_1885 ();
 sg13g2_decap_8 FILLER_42_1892 ();
 sg13g2_fill_1 FILLER_42_1899 ();
 sg13g2_decap_8 FILLER_42_1904 ();
 sg13g2_fill_1 FILLER_42_1927 ();
 sg13g2_decap_8 FILLER_42_1938 ();
 sg13g2_decap_8 FILLER_42_1945 ();
 sg13g2_fill_1 FILLER_42_1956 ();
 sg13g2_fill_2 FILLER_42_1967 ();
 sg13g2_fill_1 FILLER_42_1969 ();
 sg13g2_fill_2 FILLER_42_1975 ();
 sg13g2_decap_4 FILLER_42_1981 ();
 sg13g2_fill_1 FILLER_42_1985 ();
 sg13g2_decap_8 FILLER_42_2009 ();
 sg13g2_decap_8 FILLER_42_2016 ();
 sg13g2_fill_2 FILLER_42_2023 ();
 sg13g2_decap_4 FILLER_42_2038 ();
 sg13g2_fill_2 FILLER_42_2055 ();
 sg13g2_fill_2 FILLER_42_2069 ();
 sg13g2_decap_8 FILLER_42_2076 ();
 sg13g2_decap_8 FILLER_42_2083 ();
 sg13g2_decap_8 FILLER_42_2090 ();
 sg13g2_decap_8 FILLER_42_2114 ();
 sg13g2_decap_8 FILLER_42_2121 ();
 sg13g2_fill_2 FILLER_42_2128 ();
 sg13g2_fill_2 FILLER_42_2135 ();
 sg13g2_decap_8 FILLER_42_2158 ();
 sg13g2_decap_8 FILLER_42_2165 ();
 sg13g2_fill_1 FILLER_42_2172 ();
 sg13g2_fill_2 FILLER_42_2178 ();
 sg13g2_decap_8 FILLER_42_2215 ();
 sg13g2_decap_8 FILLER_42_2222 ();
 sg13g2_fill_2 FILLER_42_2229 ();
 sg13g2_fill_1 FILLER_42_2231 ();
 sg13g2_fill_1 FILLER_42_2246 ();
 sg13g2_decap_8 FILLER_42_2257 ();
 sg13g2_decap_8 FILLER_42_2264 ();
 sg13g2_fill_2 FILLER_42_2271 ();
 sg13g2_decap_8 FILLER_42_2311 ();
 sg13g2_decap_8 FILLER_42_2318 ();
 sg13g2_decap_8 FILLER_42_2325 ();
 sg13g2_fill_2 FILLER_42_2332 ();
 sg13g2_fill_1 FILLER_42_2334 ();
 sg13g2_decap_4 FILLER_42_2367 ();
 sg13g2_fill_1 FILLER_42_2371 ();
 sg13g2_fill_2 FILLER_42_2385 ();
 sg13g2_decap_8 FILLER_42_2435 ();
 sg13g2_decap_4 FILLER_42_2442 ();
 sg13g2_fill_2 FILLER_42_2522 ();
 sg13g2_fill_1 FILLER_42_2524 ();
 sg13g2_fill_1 FILLER_42_2530 ();
 sg13g2_decap_8 FILLER_42_2600 ();
 sg13g2_fill_1 FILLER_42_2607 ();
 sg13g2_fill_1 FILLER_42_2621 ();
 sg13g2_fill_2 FILLER_42_2770 ();
 sg13g2_fill_1 FILLER_42_2772 ();
 sg13g2_decap_8 FILLER_42_2819 ();
 sg13g2_fill_1 FILLER_42_2826 ();
 sg13g2_decap_8 FILLER_42_2873 ();
 sg13g2_fill_2 FILLER_42_2880 ();
 sg13g2_fill_1 FILLER_42_2882 ();
 sg13g2_decap_4 FILLER_42_2909 ();
 sg13g2_fill_2 FILLER_42_2913 ();
 sg13g2_decap_8 FILLER_42_2994 ();
 sg13g2_fill_1 FILLER_42_3001 ();
 sg13g2_fill_2 FILLER_42_3012 ();
 sg13g2_fill_1 FILLER_42_3014 ();
 sg13g2_decap_8 FILLER_42_3045 ();
 sg13g2_decap_8 FILLER_42_3052 ();
 sg13g2_decap_8 FILLER_42_3059 ();
 sg13g2_fill_1 FILLER_42_3112 ();
 sg13g2_decap_8 FILLER_42_3117 ();
 sg13g2_decap_8 FILLER_42_3124 ();
 sg13g2_fill_2 FILLER_42_3131 ();
 sg13g2_fill_1 FILLER_42_3133 ();
 sg13g2_fill_2 FILLER_42_3147 ();
 sg13g2_decap_4 FILLER_42_3153 ();
 sg13g2_fill_2 FILLER_42_3157 ();
 sg13g2_fill_1 FILLER_42_3178 ();
 sg13g2_fill_2 FILLER_42_3216 ();
 sg13g2_fill_1 FILLER_42_3218 ();
 sg13g2_fill_2 FILLER_42_3275 ();
 sg13g2_fill_1 FILLER_42_3277 ();
 sg13g2_decap_4 FILLER_42_3354 ();
 sg13g2_fill_1 FILLER_42_3417 ();
 sg13g2_decap_8 FILLER_42_3439 ();
 sg13g2_decap_8 FILLER_42_3446 ();
 sg13g2_decap_4 FILLER_42_3453 ();
 sg13g2_fill_2 FILLER_42_3457 ();
 sg13g2_fill_2 FILLER_42_3469 ();
 sg13g2_fill_1 FILLER_42_3471 ();
 sg13g2_decap_8 FILLER_42_3508 ();
 sg13g2_decap_8 FILLER_42_3515 ();
 sg13g2_decap_8 FILLER_42_3522 ();
 sg13g2_decap_8 FILLER_42_3529 ();
 sg13g2_decap_4 FILLER_42_3545 ();
 sg13g2_fill_1 FILLER_42_3549 ();
 sg13g2_fill_1 FILLER_42_3554 ();
 sg13g2_decap_8 FILLER_42_3564 ();
 sg13g2_decap_8 FILLER_42_3571 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_4 ();
 sg13g2_fill_2 FILLER_43_36 ();
 sg13g2_decap_8 FILLER_43_47 ();
 sg13g2_fill_2 FILLER_43_90 ();
 sg13g2_fill_1 FILLER_43_92 ();
 sg13g2_decap_8 FILLER_43_106 ();
 sg13g2_fill_2 FILLER_43_113 ();
 sg13g2_fill_2 FILLER_43_128 ();
 sg13g2_decap_8 FILLER_43_151 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_decap_4 FILLER_43_172 ();
 sg13g2_decap_4 FILLER_43_222 ();
 sg13g2_fill_1 FILLER_43_226 ();
 sg13g2_fill_2 FILLER_43_256 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_decap_4 FILLER_43_292 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_decap_8 FILLER_43_339 ();
 sg13g2_fill_1 FILLER_43_381 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_fill_1 FILLER_43_407 ();
 sg13g2_fill_1 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_419 ();
 sg13g2_decap_8 FILLER_43_426 ();
 sg13g2_decap_8 FILLER_43_433 ();
 sg13g2_fill_1 FILLER_43_440 ();
 sg13g2_decap_4 FILLER_43_478 ();
 sg13g2_fill_1 FILLER_43_509 ();
 sg13g2_decap_4 FILLER_43_528 ();
 sg13g2_fill_1 FILLER_43_536 ();
 sg13g2_decap_8 FILLER_43_541 ();
 sg13g2_decap_8 FILLER_43_548 ();
 sg13g2_decap_4 FILLER_43_555 ();
 sg13g2_decap_8 FILLER_43_600 ();
 sg13g2_decap_8 FILLER_43_607 ();
 sg13g2_decap_4 FILLER_43_614 ();
 sg13g2_decap_8 FILLER_43_652 ();
 sg13g2_decap_8 FILLER_43_659 ();
 sg13g2_decap_8 FILLER_43_666 ();
 sg13g2_decap_4 FILLER_43_673 ();
 sg13g2_fill_1 FILLER_43_677 ();
 sg13g2_fill_2 FILLER_43_688 ();
 sg13g2_fill_1 FILLER_43_690 ();
 sg13g2_decap_8 FILLER_43_696 ();
 sg13g2_decap_4 FILLER_43_703 ();
 sg13g2_fill_2 FILLER_43_707 ();
 sg13g2_fill_1 FILLER_43_750 ();
 sg13g2_decap_8 FILLER_43_755 ();
 sg13g2_decap_8 FILLER_43_762 ();
 sg13g2_decap_4 FILLER_43_769 ();
 sg13g2_fill_2 FILLER_43_773 ();
 sg13g2_decap_4 FILLER_43_813 ();
 sg13g2_fill_1 FILLER_43_817 ();
 sg13g2_fill_2 FILLER_43_832 ();
 sg13g2_fill_1 FILLER_43_843 ();
 sg13g2_decap_8 FILLER_43_878 ();
 sg13g2_decap_8 FILLER_43_885 ();
 sg13g2_fill_2 FILLER_43_892 ();
 sg13g2_decap_4 FILLER_43_938 ();
 sg13g2_fill_1 FILLER_43_950 ();
 sg13g2_fill_1 FILLER_43_954 ();
 sg13g2_fill_2 FILLER_43_970 ();
 sg13g2_fill_1 FILLER_43_972 ();
 sg13g2_fill_1 FILLER_43_978 ();
 sg13g2_fill_1 FILLER_43_1005 ();
 sg13g2_decap_8 FILLER_43_1044 ();
 sg13g2_decap_8 FILLER_43_1051 ();
 sg13g2_fill_1 FILLER_43_1058 ();
 sg13g2_fill_2 FILLER_43_1101 ();
 sg13g2_fill_2 FILLER_43_1114 ();
 sg13g2_fill_2 FILLER_43_1133 ();
 sg13g2_fill_1 FILLER_43_1135 ();
 sg13g2_fill_2 FILLER_43_1164 ();
 sg13g2_fill_1 FILLER_43_1174 ();
 sg13g2_fill_2 FILLER_43_1188 ();
 sg13g2_fill_1 FILLER_43_1190 ();
 sg13g2_fill_2 FILLER_43_1205 ();
 sg13g2_decap_8 FILLER_43_1235 ();
 sg13g2_fill_1 FILLER_43_1242 ();
 sg13g2_fill_2 FILLER_43_1271 ();
 sg13g2_fill_1 FILLER_43_1273 ();
 sg13g2_fill_1 FILLER_43_1299 ();
 sg13g2_fill_1 FILLER_43_1314 ();
 sg13g2_decap_8 FILLER_43_1320 ();
 sg13g2_decap_8 FILLER_43_1327 ();
 sg13g2_fill_1 FILLER_43_1334 ();
 sg13g2_fill_1 FILLER_43_1348 ();
 sg13g2_fill_2 FILLER_43_1358 ();
 sg13g2_fill_1 FILLER_43_1387 ();
 sg13g2_fill_1 FILLER_43_1405 ();
 sg13g2_decap_8 FILLER_43_1415 ();
 sg13g2_decap_8 FILLER_43_1422 ();
 sg13g2_decap_8 FILLER_43_1429 ();
 sg13g2_decap_8 FILLER_43_1436 ();
 sg13g2_decap_4 FILLER_43_1443 ();
 sg13g2_fill_1 FILLER_43_1447 ();
 sg13g2_decap_8 FILLER_43_1458 ();
 sg13g2_fill_1 FILLER_43_1465 ();
 sg13g2_decap_8 FILLER_43_1509 ();
 sg13g2_decap_8 FILLER_43_1516 ();
 sg13g2_fill_2 FILLER_43_1523 ();
 sg13g2_fill_1 FILLER_43_1525 ();
 sg13g2_fill_1 FILLER_43_1544 ();
 sg13g2_fill_1 FILLER_43_1567 ();
 sg13g2_decap_8 FILLER_43_1586 ();
 sg13g2_decap_8 FILLER_43_1593 ();
 sg13g2_decap_8 FILLER_43_1600 ();
 sg13g2_fill_1 FILLER_43_1607 ();
 sg13g2_decap_8 FILLER_43_1639 ();
 sg13g2_decap_4 FILLER_43_1646 ();
 sg13g2_decap_8 FILLER_43_1658 ();
 sg13g2_fill_1 FILLER_43_1665 ();
 sg13g2_fill_2 FILLER_43_1670 ();
 sg13g2_decap_8 FILLER_43_1692 ();
 sg13g2_decap_8 FILLER_43_1699 ();
 sg13g2_decap_8 FILLER_43_1706 ();
 sg13g2_decap_4 FILLER_43_1713 ();
 sg13g2_fill_1 FILLER_43_1717 ();
 sg13g2_fill_2 FILLER_43_1724 ();
 sg13g2_fill_1 FILLER_43_1726 ();
 sg13g2_decap_8 FILLER_43_1739 ();
 sg13g2_decap_4 FILLER_43_1746 ();
 sg13g2_fill_2 FILLER_43_1750 ();
 sg13g2_decap_8 FILLER_43_1790 ();
 sg13g2_decap_8 FILLER_43_1797 ();
 sg13g2_fill_1 FILLER_43_1817 ();
 sg13g2_fill_1 FILLER_43_1840 ();
 sg13g2_decap_8 FILLER_43_1855 ();
 sg13g2_decap_8 FILLER_43_1862 ();
 sg13g2_decap_8 FILLER_43_1869 ();
 sg13g2_decap_8 FILLER_43_1876 ();
 sg13g2_decap_8 FILLER_43_1883 ();
 sg13g2_decap_8 FILLER_43_1890 ();
 sg13g2_decap_4 FILLER_43_1897 ();
 sg13g2_fill_2 FILLER_43_1901 ();
 sg13g2_decap_8 FILLER_43_1928 ();
 sg13g2_decap_8 FILLER_43_1935 ();
 sg13g2_decap_8 FILLER_43_1942 ();
 sg13g2_fill_2 FILLER_43_1949 ();
 sg13g2_fill_1 FILLER_43_1969 ();
 sg13g2_decap_8 FILLER_43_1998 ();
 sg13g2_decap_8 FILLER_43_2005 ();
 sg13g2_fill_2 FILLER_43_2012 ();
 sg13g2_fill_1 FILLER_43_2014 ();
 sg13g2_decap_8 FILLER_43_2025 ();
 sg13g2_decap_8 FILLER_43_2032 ();
 sg13g2_decap_8 FILLER_43_2039 ();
 sg13g2_fill_1 FILLER_43_2046 ();
 sg13g2_decap_8 FILLER_43_2065 ();
 sg13g2_fill_1 FILLER_43_2072 ();
 sg13g2_fill_1 FILLER_43_2078 ();
 sg13g2_fill_1 FILLER_43_2086 ();
 sg13g2_fill_2 FILLER_43_2104 ();
 sg13g2_fill_2 FILLER_43_2119 ();
 sg13g2_fill_1 FILLER_43_2121 ();
 sg13g2_fill_1 FILLER_43_2137 ();
 sg13g2_decap_8 FILLER_43_2156 ();
 sg13g2_decap_8 FILLER_43_2163 ();
 sg13g2_decap_4 FILLER_43_2170 ();
 sg13g2_fill_2 FILLER_43_2174 ();
 sg13g2_fill_2 FILLER_43_2194 ();
 sg13g2_decap_8 FILLER_43_2209 ();
 sg13g2_fill_2 FILLER_43_2216 ();
 sg13g2_decap_8 FILLER_43_2221 ();
 sg13g2_fill_2 FILLER_43_2228 ();
 sg13g2_decap_4 FILLER_43_2271 ();
 sg13g2_fill_1 FILLER_43_2275 ();
 sg13g2_fill_1 FILLER_43_2293 ();
 sg13g2_fill_2 FILLER_43_2303 ();
 sg13g2_fill_1 FILLER_43_2305 ();
 sg13g2_decap_8 FILLER_43_2319 ();
 sg13g2_fill_2 FILLER_43_2326 ();
 sg13g2_fill_1 FILLER_43_2328 ();
 sg13g2_decap_4 FILLER_43_2380 ();
 sg13g2_fill_1 FILLER_43_2384 ();
 sg13g2_fill_2 FILLER_43_2422 ();
 sg13g2_fill_1 FILLER_43_2424 ();
 sg13g2_decap_8 FILLER_43_2438 ();
 sg13g2_decap_8 FILLER_43_2445 ();
 sg13g2_fill_2 FILLER_43_2452 ();
 sg13g2_fill_1 FILLER_43_2454 ();
 sg13g2_decap_4 FILLER_43_2504 ();
 sg13g2_fill_2 FILLER_43_2508 ();
 sg13g2_decap_4 FILLER_43_2520 ();
 sg13g2_decap_8 FILLER_43_2533 ();
 sg13g2_decap_8 FILLER_43_2565 ();
 sg13g2_decap_4 FILLER_43_2572 ();
 sg13g2_fill_1 FILLER_43_2576 ();
 sg13g2_fill_2 FILLER_43_2595 ();
 sg13g2_fill_1 FILLER_43_2597 ();
 sg13g2_decap_8 FILLER_43_2607 ();
 sg13g2_decap_8 FILLER_43_2614 ();
 sg13g2_fill_2 FILLER_43_2621 ();
 sg13g2_fill_2 FILLER_43_2675 ();
 sg13g2_fill_1 FILLER_43_2690 ();
 sg13g2_decap_8 FILLER_43_2731 ();
 sg13g2_fill_2 FILLER_43_2738 ();
 sg13g2_fill_1 FILLER_43_2740 ();
 sg13g2_fill_2 FILLER_43_2764 ();
 sg13g2_fill_2 FILLER_43_2776 ();
 sg13g2_fill_1 FILLER_43_2778 ();
 sg13g2_decap_8 FILLER_43_2810 ();
 sg13g2_decap_4 FILLER_43_2817 ();
 sg13g2_fill_2 FILLER_43_2834 ();
 sg13g2_fill_1 FILLER_43_2836 ();
 sg13g2_fill_1 FILLER_43_2855 ();
 sg13g2_decap_4 FILLER_43_2908 ();
 sg13g2_fill_2 FILLER_43_2912 ();
 sg13g2_decap_8 FILLER_43_2940 ();
 sg13g2_decap_8 FILLER_43_2947 ();
 sg13g2_fill_1 FILLER_43_2954 ();
 sg13g2_decap_8 FILLER_43_3003 ();
 sg13g2_fill_2 FILLER_43_3010 ();
 sg13g2_decap_4 FILLER_43_3049 ();
 sg13g2_fill_1 FILLER_43_3053 ();
 sg13g2_decap_8 FILLER_43_3063 ();
 sg13g2_fill_1 FILLER_43_3070 ();
 sg13g2_fill_1 FILLER_43_3075 ();
 sg13g2_decap_8 FILLER_43_3107 ();
 sg13g2_decap_8 FILLER_43_3114 ();
 sg13g2_decap_8 FILLER_43_3121 ();
 sg13g2_decap_4 FILLER_43_3128 ();
 sg13g2_fill_2 FILLER_43_3132 ();
 sg13g2_decap_8 FILLER_43_3147 ();
 sg13g2_decap_8 FILLER_43_3154 ();
 sg13g2_decap_8 FILLER_43_3161 ();
 sg13g2_fill_2 FILLER_43_3168 ();
 sg13g2_fill_2 FILLER_43_3180 ();
 sg13g2_decap_8 FILLER_43_3208 ();
 sg13g2_fill_1 FILLER_43_3215 ();
 sg13g2_fill_1 FILLER_43_3243 ();
 sg13g2_decap_8 FILLER_43_3280 ();
 sg13g2_fill_2 FILLER_43_3287 ();
 sg13g2_decap_8 FILLER_43_3360 ();
 sg13g2_decap_8 FILLER_43_3367 ();
 sg13g2_fill_2 FILLER_43_3374 ();
 sg13g2_decap_4 FILLER_43_3380 ();
 sg13g2_fill_1 FILLER_43_3384 ();
 sg13g2_decap_8 FILLER_43_3394 ();
 sg13g2_decap_4 FILLER_43_3401 ();
 sg13g2_fill_2 FILLER_43_3405 ();
 sg13g2_decap_8 FILLER_43_3424 ();
 sg13g2_decap_4 FILLER_43_3431 ();
 sg13g2_fill_2 FILLER_43_3435 ();
 sg13g2_fill_2 FILLER_43_3445 ();
 sg13g2_fill_2 FILLER_43_3462 ();
 sg13g2_fill_1 FILLER_43_3464 ();
 sg13g2_decap_8 FILLER_43_3508 ();
 sg13g2_decap_8 FILLER_43_3515 ();
 sg13g2_decap_4 FILLER_43_3522 ();
 sg13g2_decap_4 FILLER_43_3539 ();
 sg13g2_fill_2 FILLER_43_3543 ();
 sg13g2_decap_8 FILLER_43_3558 ();
 sg13g2_decap_8 FILLER_43_3565 ();
 sg13g2_decap_4 FILLER_43_3572 ();
 sg13g2_fill_2 FILLER_43_3576 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_11 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_fill_2 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_58 ();
 sg13g2_fill_2 FILLER_44_63 ();
 sg13g2_fill_1 FILLER_44_65 ();
 sg13g2_decap_8 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_decap_8 FILLER_44_116 ();
 sg13g2_fill_2 FILLER_44_123 ();
 sg13g2_fill_1 FILLER_44_125 ();
 sg13g2_decap_8 FILLER_44_153 ();
 sg13g2_decap_8 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_167 ();
 sg13g2_fill_2 FILLER_44_220 ();
 sg13g2_fill_1 FILLER_44_222 ();
 sg13g2_decap_8 FILLER_44_254 ();
 sg13g2_decap_8 FILLER_44_261 ();
 sg13g2_fill_2 FILLER_44_268 ();
 sg13g2_fill_1 FILLER_44_270 ();
 sg13g2_decap_4 FILLER_44_275 ();
 sg13g2_decap_8 FILLER_44_288 ();
 sg13g2_decap_4 FILLER_44_295 ();
 sg13g2_fill_2 FILLER_44_299 ();
 sg13g2_fill_2 FILLER_44_373 ();
 sg13g2_fill_1 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_423 ();
 sg13g2_decap_8 FILLER_44_430 ();
 sg13g2_decap_8 FILLER_44_437 ();
 sg13g2_decap_8 FILLER_44_444 ();
 sg13g2_decap_8 FILLER_44_451 ();
 sg13g2_decap_8 FILLER_44_458 ();
 sg13g2_decap_8 FILLER_44_465 ();
 sg13g2_decap_8 FILLER_44_472 ();
 sg13g2_decap_8 FILLER_44_479 ();
 sg13g2_fill_1 FILLER_44_486 ();
 sg13g2_fill_2 FILLER_44_496 ();
 sg13g2_decap_4 FILLER_44_503 ();
 sg13g2_fill_1 FILLER_44_507 ();
 sg13g2_fill_2 FILLER_44_512 ();
 sg13g2_decap_4 FILLER_44_522 ();
 sg13g2_fill_1 FILLER_44_526 ();
 sg13g2_fill_1 FILLER_44_531 ();
 sg13g2_decap_8 FILLER_44_536 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_557 ();
 sg13g2_decap_4 FILLER_44_564 ();
 sg13g2_decap_8 FILLER_44_572 ();
 sg13g2_decap_4 FILLER_44_579 ();
 sg13g2_fill_2 FILLER_44_583 ();
 sg13g2_decap_8 FILLER_44_589 ();
 sg13g2_fill_1 FILLER_44_596 ();
 sg13g2_decap_8 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_609 ();
 sg13g2_decap_8 FILLER_44_650 ();
 sg13g2_decap_8 FILLER_44_657 ();
 sg13g2_fill_2 FILLER_44_664 ();
 sg13g2_decap_8 FILLER_44_702 ();
 sg13g2_fill_2 FILLER_44_709 ();
 sg13g2_fill_1 FILLER_44_721 ();
 sg13g2_decap_8 FILLER_44_762 ();
 sg13g2_decap_4 FILLER_44_769 ();
 sg13g2_fill_1 FILLER_44_773 ();
 sg13g2_fill_2 FILLER_44_801 ();
 sg13g2_fill_1 FILLER_44_849 ();
 sg13g2_decap_8 FILLER_44_877 ();
 sg13g2_fill_2 FILLER_44_884 ();
 sg13g2_fill_1 FILLER_44_886 ();
 sg13g2_fill_2 FILLER_44_896 ();
 sg13g2_fill_1 FILLER_44_898 ();
 sg13g2_fill_1 FILLER_44_915 ();
 sg13g2_fill_1 FILLER_44_924 ();
 sg13g2_fill_2 FILLER_44_931 ();
 sg13g2_decap_8 FILLER_44_951 ();
 sg13g2_decap_8 FILLER_44_958 ();
 sg13g2_decap_4 FILLER_44_985 ();
 sg13g2_fill_1 FILLER_44_989 ();
 sg13g2_decap_8 FILLER_44_1040 ();
 sg13g2_decap_8 FILLER_44_1047 ();
 sg13g2_fill_1 FILLER_44_1054 ();
 sg13g2_fill_2 FILLER_44_1083 ();
 sg13g2_fill_1 FILLER_44_1085 ();
 sg13g2_fill_2 FILLER_44_1104 ();
 sg13g2_fill_1 FILLER_44_1121 ();
 sg13g2_fill_2 FILLER_44_1132 ();
 sg13g2_fill_1 FILLER_44_1134 ();
 sg13g2_decap_4 FILLER_44_1148 ();
 sg13g2_fill_1 FILLER_44_1152 ();
 sg13g2_fill_1 FILLER_44_1159 ();
 sg13g2_fill_2 FILLER_44_1178 ();
 sg13g2_decap_4 FILLER_44_1255 ();
 sg13g2_fill_1 FILLER_44_1259 ();
 sg13g2_fill_1 FILLER_44_1278 ();
 sg13g2_decap_4 FILLER_44_1315 ();
 sg13g2_fill_1 FILLER_44_1319 ();
 sg13g2_fill_2 FILLER_44_1352 ();
 sg13g2_fill_2 FILLER_44_1426 ();
 sg13g2_fill_1 FILLER_44_1428 ();
 sg13g2_decap_8 FILLER_44_1447 ();
 sg13g2_decap_8 FILLER_44_1454 ();
 sg13g2_decap_4 FILLER_44_1461 ();
 sg13g2_fill_2 FILLER_44_1481 ();
 sg13g2_decap_8 FILLER_44_1507 ();
 sg13g2_decap_8 FILLER_44_1514 ();
 sg13g2_decap_8 FILLER_44_1521 ();
 sg13g2_decap_4 FILLER_44_1528 ();
 sg13g2_fill_1 FILLER_44_1532 ();
 sg13g2_fill_1 FILLER_44_1537 ();
 sg13g2_decap_4 FILLER_44_1549 ();
 sg13g2_decap_4 FILLER_44_1558 ();
 sg13g2_fill_2 FILLER_44_1562 ();
 sg13g2_fill_1 FILLER_44_1572 ();
 sg13g2_fill_2 FILLER_44_1581 ();
 sg13g2_fill_1 FILLER_44_1583 ();
 sg13g2_fill_2 FILLER_44_1589 ();
 sg13g2_decap_8 FILLER_44_1597 ();
 sg13g2_decap_4 FILLER_44_1604 ();
 sg13g2_fill_2 FILLER_44_1608 ();
 sg13g2_fill_2 FILLER_44_1631 ();
 sg13g2_decap_8 FILLER_44_1649 ();
 sg13g2_decap_8 FILLER_44_1656 ();
 sg13g2_fill_2 FILLER_44_1663 ();
 sg13g2_fill_1 FILLER_44_1665 ();
 sg13g2_decap_8 FILLER_44_1699 ();
 sg13g2_decap_8 FILLER_44_1706 ();
 sg13g2_decap_8 FILLER_44_1713 ();
 sg13g2_decap_8 FILLER_44_1720 ();
 sg13g2_decap_8 FILLER_44_1727 ();
 sg13g2_decap_8 FILLER_44_1734 ();
 sg13g2_fill_2 FILLER_44_1741 ();
 sg13g2_fill_1 FILLER_44_1743 ();
 sg13g2_fill_2 FILLER_44_1771 ();
 sg13g2_fill_1 FILLER_44_1773 ();
 sg13g2_decap_8 FILLER_44_1791 ();
 sg13g2_decap_8 FILLER_44_1798 ();
 sg13g2_fill_2 FILLER_44_1814 ();
 sg13g2_decap_8 FILLER_44_1841 ();
 sg13g2_decap_8 FILLER_44_1848 ();
 sg13g2_decap_8 FILLER_44_1855 ();
 sg13g2_decap_8 FILLER_44_1862 ();
 sg13g2_fill_2 FILLER_44_1869 ();
 sg13g2_decap_8 FILLER_44_1879 ();
 sg13g2_decap_8 FILLER_44_1886 ();
 sg13g2_fill_1 FILLER_44_1893 ();
 sg13g2_decap_8 FILLER_44_1938 ();
 sg13g2_decap_8 FILLER_44_1945 ();
 sg13g2_decap_8 FILLER_44_1952 ();
 sg13g2_decap_8 FILLER_44_1964 ();
 sg13g2_decap_8 FILLER_44_1971 ();
 sg13g2_decap_8 FILLER_44_1978 ();
 sg13g2_decap_4 FILLER_44_1989 ();
 sg13g2_fill_2 FILLER_44_1993 ();
 sg13g2_decap_8 FILLER_44_2007 ();
 sg13g2_fill_2 FILLER_44_2014 ();
 sg13g2_decap_8 FILLER_44_2021 ();
 sg13g2_fill_1 FILLER_44_2028 ();
 sg13g2_decap_8 FILLER_44_2034 ();
 sg13g2_decap_8 FILLER_44_2041 ();
 sg13g2_decap_4 FILLER_44_2048 ();
 sg13g2_decap_8 FILLER_44_2068 ();
 sg13g2_fill_2 FILLER_44_2083 ();
 sg13g2_fill_2 FILLER_44_2097 ();
 sg13g2_decap_8 FILLER_44_2122 ();
 sg13g2_fill_2 FILLER_44_2129 ();
 sg13g2_decap_8 FILLER_44_2153 ();
 sg13g2_decap_8 FILLER_44_2160 ();
 sg13g2_decap_8 FILLER_44_2167 ();
 sg13g2_fill_2 FILLER_44_2174 ();
 sg13g2_decap_8 FILLER_44_2199 ();
 sg13g2_decap_8 FILLER_44_2206 ();
 sg13g2_decap_8 FILLER_44_2213 ();
 sg13g2_decap_4 FILLER_44_2220 ();
 sg13g2_decap_8 FILLER_44_2264 ();
 sg13g2_decap_8 FILLER_44_2271 ();
 sg13g2_decap_8 FILLER_44_2278 ();
 sg13g2_fill_1 FILLER_44_2285 ();
 sg13g2_decap_4 FILLER_44_2314 ();
 sg13g2_fill_2 FILLER_44_2318 ();
 sg13g2_decap_8 FILLER_44_2361 ();
 sg13g2_decap_8 FILLER_44_2368 ();
 sg13g2_decap_8 FILLER_44_2375 ();
 sg13g2_decap_8 FILLER_44_2382 ();
 sg13g2_decap_4 FILLER_44_2389 ();
 sg13g2_fill_1 FILLER_44_2393 ();
 sg13g2_decap_8 FILLER_44_2434 ();
 sg13g2_decap_8 FILLER_44_2441 ();
 sg13g2_decap_8 FILLER_44_2448 ();
 sg13g2_decap_4 FILLER_44_2455 ();
 sg13g2_decap_8 FILLER_44_2490 ();
 sg13g2_decap_8 FILLER_44_2497 ();
 sg13g2_fill_2 FILLER_44_2504 ();
 sg13g2_fill_1 FILLER_44_2506 ();
 sg13g2_decap_8 FILLER_44_2534 ();
 sg13g2_fill_2 FILLER_44_2541 ();
 sg13g2_fill_1 FILLER_44_2543 ();
 sg13g2_decap_8 FILLER_44_2566 ();
 sg13g2_decap_8 FILLER_44_2610 ();
 sg13g2_decap_8 FILLER_44_2617 ();
 sg13g2_fill_1 FILLER_44_2624 ();
 sg13g2_decap_8 FILLER_44_2664 ();
 sg13g2_decap_8 FILLER_44_2671 ();
 sg13g2_fill_1 FILLER_44_2678 ();
 sg13g2_fill_2 FILLER_44_2706 ();
 sg13g2_fill_1 FILLER_44_2708 ();
 sg13g2_decap_8 FILLER_44_2722 ();
 sg13g2_decap_8 FILLER_44_2729 ();
 sg13g2_decap_8 FILLER_44_2736 ();
 sg13g2_decap_8 FILLER_44_2760 ();
 sg13g2_decap_4 FILLER_44_2767 ();
 sg13g2_decap_8 FILLER_44_2776 ();
 sg13g2_decap_4 FILLER_44_2783 ();
 sg13g2_fill_1 FILLER_44_2787 ();
 sg13g2_fill_2 FILLER_44_2791 ();
 sg13g2_fill_1 FILLER_44_2793 ();
 sg13g2_decap_4 FILLER_44_2799 ();
 sg13g2_decap_8 FILLER_44_2808 ();
 sg13g2_decap_8 FILLER_44_2815 ();
 sg13g2_decap_8 FILLER_44_2822 ();
 sg13g2_decap_8 FILLER_44_2829 ();
 sg13g2_fill_1 FILLER_44_2836 ();
 sg13g2_fill_1 FILLER_44_2855 ();
 sg13g2_decap_8 FILLER_44_2869 ();
 sg13g2_decap_4 FILLER_44_2876 ();
 sg13g2_fill_2 FILLER_44_2880 ();
 sg13g2_fill_2 FILLER_44_2921 ();
 sg13g2_decap_8 FILLER_44_2949 ();
 sg13g2_decap_8 FILLER_44_2956 ();
 sg13g2_fill_2 FILLER_44_2963 ();
 sg13g2_fill_1 FILLER_44_2965 ();
 sg13g2_decap_8 FILLER_44_2989 ();
 sg13g2_decap_4 FILLER_44_3033 ();
 sg13g2_decap_8 FILLER_44_3064 ();
 sg13g2_decap_8 FILLER_44_3071 ();
 sg13g2_fill_2 FILLER_44_3078 ();
 sg13g2_decap_8 FILLER_44_3108 ();
 sg13g2_decap_8 FILLER_44_3115 ();
 sg13g2_decap_8 FILLER_44_3122 ();
 sg13g2_fill_2 FILLER_44_3129 ();
 sg13g2_decap_8 FILLER_44_3157 ();
 sg13g2_fill_2 FILLER_44_3164 ();
 sg13g2_decap_8 FILLER_44_3193 ();
 sg13g2_decap_8 FILLER_44_3200 ();
 sg13g2_decap_8 FILLER_44_3207 ();
 sg13g2_decap_8 FILLER_44_3214 ();
 sg13g2_fill_2 FILLER_44_3225 ();
 sg13g2_fill_2 FILLER_44_3246 ();
 sg13g2_fill_1 FILLER_44_3248 ();
 sg13g2_decap_8 FILLER_44_3270 ();
 sg13g2_decap_8 FILLER_44_3277 ();
 sg13g2_decap_8 FILLER_44_3284 ();
 sg13g2_fill_2 FILLER_44_3291 ();
 sg13g2_fill_1 FILLER_44_3293 ();
 sg13g2_decap_8 FILLER_44_3357 ();
 sg13g2_decap_8 FILLER_44_3364 ();
 sg13g2_fill_2 FILLER_44_3371 ();
 sg13g2_fill_2 FILLER_44_3408 ();
 sg13g2_fill_1 FILLER_44_3410 ();
 sg13g2_decap_8 FILLER_44_3429 ();
 sg13g2_decap_8 FILLER_44_3436 ();
 sg13g2_decap_8 FILLER_44_3448 ();
 sg13g2_decap_4 FILLER_44_3455 ();
 sg13g2_fill_2 FILLER_44_3459 ();
 sg13g2_fill_2 FILLER_44_3469 ();
 sg13g2_fill_1 FILLER_44_3523 ();
 sg13g2_decap_4 FILLER_44_3572 ();
 sg13g2_fill_2 FILLER_44_3576 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_decap_4 FILLER_45_22 ();
 sg13g2_fill_1 FILLER_45_26 ();
 sg13g2_decap_8 FILLER_45_37 ();
 sg13g2_decap_8 FILLER_45_44 ();
 sg13g2_decap_8 FILLER_45_51 ();
 sg13g2_decap_8 FILLER_45_58 ();
 sg13g2_decap_4 FILLER_45_65 ();
 sg13g2_fill_2 FILLER_45_69 ();
 sg13g2_fill_2 FILLER_45_75 ();
 sg13g2_fill_1 FILLER_45_96 ();
 sg13g2_decap_4 FILLER_45_124 ();
 sg13g2_fill_1 FILLER_45_128 ();
 sg13g2_fill_2 FILLER_45_143 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_4 FILLER_45_182 ();
 sg13g2_fill_2 FILLER_45_186 ();
 sg13g2_fill_2 FILLER_45_206 ();
 sg13g2_fill_2 FILLER_45_217 ();
 sg13g2_fill_2 FILLER_45_224 ();
 sg13g2_fill_1 FILLER_45_226 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_fill_1 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_247 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_2 FILLER_45_260 ();
 sg13g2_fill_1 FILLER_45_262 ();
 sg13g2_decap_8 FILLER_45_282 ();
 sg13g2_decap_8 FILLER_45_289 ();
 sg13g2_decap_8 FILLER_45_296 ();
 sg13g2_decap_4 FILLER_45_303 ();
 sg13g2_fill_1 FILLER_45_307 ();
 sg13g2_decap_4 FILLER_45_312 ();
 sg13g2_fill_2 FILLER_45_333 ();
 sg13g2_fill_1 FILLER_45_335 ();
 sg13g2_fill_2 FILLER_45_363 ();
 sg13g2_fill_1 FILLER_45_365 ();
 sg13g2_fill_2 FILLER_45_376 ();
 sg13g2_fill_1 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_419 ();
 sg13g2_decap_8 FILLER_45_426 ();
 sg13g2_decap_8 FILLER_45_433 ();
 sg13g2_decap_8 FILLER_45_440 ();
 sg13g2_decap_8 FILLER_45_447 ();
 sg13g2_decap_8 FILLER_45_454 ();
 sg13g2_fill_2 FILLER_45_461 ();
 sg13g2_fill_1 FILLER_45_463 ();
 sg13g2_decap_8 FILLER_45_507 ();
 sg13g2_decap_4 FILLER_45_514 ();
 sg13g2_fill_2 FILLER_45_518 ();
 sg13g2_fill_2 FILLER_45_532 ();
 sg13g2_decap_8 FILLER_45_561 ();
 sg13g2_decap_4 FILLER_45_568 ();
 sg13g2_fill_2 FILLER_45_572 ();
 sg13g2_fill_1 FILLER_45_602 ();
 sg13g2_decap_8 FILLER_45_608 ();
 sg13g2_decap_4 FILLER_45_615 ();
 sg13g2_fill_1 FILLER_45_619 ();
 sg13g2_fill_1 FILLER_45_633 ();
 sg13g2_decap_8 FILLER_45_646 ();
 sg13g2_decap_4 FILLER_45_653 ();
 sg13g2_fill_2 FILLER_45_657 ();
 sg13g2_decap_8 FILLER_45_693 ();
 sg13g2_decap_8 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_707 ();
 sg13g2_decap_8 FILLER_45_714 ();
 sg13g2_fill_2 FILLER_45_721 ();
 sg13g2_fill_2 FILLER_45_733 ();
 sg13g2_fill_1 FILLER_45_748 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_fill_1 FILLER_45_807 ();
 sg13g2_fill_1 FILLER_45_864 ();
 sg13g2_decap_8 FILLER_45_874 ();
 sg13g2_decap_8 FILLER_45_881 ();
 sg13g2_decap_4 FILLER_45_888 ();
 sg13g2_fill_1 FILLER_45_892 ();
 sg13g2_decap_8 FILLER_45_898 ();
 sg13g2_decap_4 FILLER_45_905 ();
 sg13g2_fill_1 FILLER_45_922 ();
 sg13g2_fill_1 FILLER_45_928 ();
 sg13g2_fill_1 FILLER_45_934 ();
 sg13g2_decap_8 FILLER_45_946 ();
 sg13g2_decap_8 FILLER_45_953 ();
 sg13g2_decap_8 FILLER_45_960 ();
 sg13g2_fill_2 FILLER_45_967 ();
 sg13g2_fill_1 FILLER_45_969 ();
 sg13g2_decap_8 FILLER_45_974 ();
 sg13g2_decap_8 FILLER_45_981 ();
 sg13g2_decap_8 FILLER_45_988 ();
 sg13g2_fill_2 FILLER_45_995 ();
 sg13g2_fill_1 FILLER_45_997 ();
 sg13g2_decap_8 FILLER_45_1039 ();
 sg13g2_decap_8 FILLER_45_1046 ();
 sg13g2_decap_8 FILLER_45_1053 ();
 sg13g2_decap_8 FILLER_45_1060 ();
 sg13g2_decap_8 FILLER_45_1067 ();
 sg13g2_decap_8 FILLER_45_1074 ();
 sg13g2_fill_1 FILLER_45_1145 ();
 sg13g2_decap_8 FILLER_45_1149 ();
 sg13g2_fill_2 FILLER_45_1156 ();
 sg13g2_fill_2 FILLER_45_1161 ();
 sg13g2_fill_1 FILLER_45_1163 ();
 sg13g2_fill_2 FILLER_45_1181 ();
 sg13g2_fill_1 FILLER_45_1183 ();
 sg13g2_fill_2 FILLER_45_1202 ();
 sg13g2_fill_1 FILLER_45_1211 ();
 sg13g2_decap_8 FILLER_45_1231 ();
 sg13g2_decap_8 FILLER_45_1238 ();
 sg13g2_decap_8 FILLER_45_1245 ();
 sg13g2_fill_2 FILLER_45_1252 ();
 sg13g2_fill_1 FILLER_45_1254 ();
 sg13g2_fill_1 FILLER_45_1308 ();
 sg13g2_decap_8 FILLER_45_1318 ();
 sg13g2_fill_1 FILLER_45_1325 ();
 sg13g2_decap_4 FILLER_45_1330 ();
 sg13g2_fill_2 FILLER_45_1338 ();
 sg13g2_fill_2 FILLER_45_1358 ();
 sg13g2_fill_1 FILLER_45_1391 ();
 sg13g2_fill_2 FILLER_45_1405 ();
 sg13g2_decap_4 FILLER_45_1416 ();
 sg13g2_fill_1 FILLER_45_1430 ();
 sg13g2_decap_8 FILLER_45_1437 ();
 sg13g2_fill_2 FILLER_45_1444 ();
 sg13g2_decap_8 FILLER_45_1451 ();
 sg13g2_decap_8 FILLER_45_1458 ();
 sg13g2_decap_8 FILLER_45_1465 ();
 sg13g2_fill_2 FILLER_45_1472 ();
 sg13g2_fill_1 FILLER_45_1489 ();
 sg13g2_decap_4 FILLER_45_1507 ();
 sg13g2_fill_1 FILLER_45_1511 ();
 sg13g2_decap_4 FILLER_45_1518 ();
 sg13g2_decap_8 FILLER_45_1527 ();
 sg13g2_decap_8 FILLER_45_1534 ();
 sg13g2_decap_8 FILLER_45_1541 ();
 sg13g2_decap_8 FILLER_45_1548 ();
 sg13g2_decap_8 FILLER_45_1555 ();
 sg13g2_decap_4 FILLER_45_1562 ();
 sg13g2_fill_2 FILLER_45_1600 ();
 sg13g2_fill_1 FILLER_45_1607 ();
 sg13g2_decap_8 FILLER_45_1613 ();
 sg13g2_decap_8 FILLER_45_1620 ();
 sg13g2_decap_8 FILLER_45_1627 ();
 sg13g2_decap_8 FILLER_45_1634 ();
 sg13g2_decap_8 FILLER_45_1653 ();
 sg13g2_decap_8 FILLER_45_1660 ();
 sg13g2_decap_8 FILLER_45_1667 ();
 sg13g2_decap_8 FILLER_45_1697 ();
 sg13g2_fill_2 FILLER_45_1704 ();
 sg13g2_fill_1 FILLER_45_1706 ();
 sg13g2_decap_8 FILLER_45_1711 ();
 sg13g2_decap_8 FILLER_45_1718 ();
 sg13g2_decap_8 FILLER_45_1725 ();
 sg13g2_decap_8 FILLER_45_1732 ();
 sg13g2_decap_4 FILLER_45_1739 ();
 sg13g2_fill_2 FILLER_45_1743 ();
 sg13g2_decap_4 FILLER_45_1766 ();
 sg13g2_fill_2 FILLER_45_1770 ();
 sg13g2_decap_8 FILLER_45_1776 ();
 sg13g2_decap_8 FILLER_45_1783 ();
 sg13g2_decap_8 FILLER_45_1790 ();
 sg13g2_decap_8 FILLER_45_1797 ();
 sg13g2_decap_8 FILLER_45_1804 ();
 sg13g2_decap_8 FILLER_45_1836 ();
 sg13g2_decap_8 FILLER_45_1843 ();
 sg13g2_decap_8 FILLER_45_1850 ();
 sg13g2_fill_2 FILLER_45_1857 ();
 sg13g2_fill_2 FILLER_45_1881 ();
 sg13g2_fill_1 FILLER_45_1883 ();
 sg13g2_fill_2 FILLER_45_1913 ();
 sg13g2_decap_8 FILLER_45_1939 ();
 sg13g2_decap_8 FILLER_45_1946 ();
 sg13g2_decap_8 FILLER_45_1953 ();
 sg13g2_fill_2 FILLER_45_1960 ();
 sg13g2_decap_8 FILLER_45_1975 ();
 sg13g2_decap_8 FILLER_45_1982 ();
 sg13g2_fill_2 FILLER_45_1989 ();
 sg13g2_decap_4 FILLER_45_2017 ();
 sg13g2_decap_8 FILLER_45_2046 ();
 sg13g2_decap_8 FILLER_45_2053 ();
 sg13g2_fill_1 FILLER_45_2060 ();
 sg13g2_decap_8 FILLER_45_2066 ();
 sg13g2_decap_8 FILLER_45_2073 ();
 sg13g2_fill_2 FILLER_45_2088 ();
 sg13g2_fill_1 FILLER_45_2090 ();
 sg13g2_decap_8 FILLER_45_2095 ();
 sg13g2_fill_1 FILLER_45_2114 ();
 sg13g2_decap_8 FILLER_45_2125 ();
 sg13g2_fill_2 FILLER_45_2132 ();
 sg13g2_fill_1 FILLER_45_2143 ();
 sg13g2_decap_8 FILLER_45_2149 ();
 sg13g2_fill_2 FILLER_45_2156 ();
 sg13g2_fill_1 FILLER_45_2158 ();
 sg13g2_fill_1 FILLER_45_2163 ();
 sg13g2_decap_8 FILLER_45_2199 ();
 sg13g2_fill_1 FILLER_45_2206 ();
 sg13g2_decap_8 FILLER_45_2210 ();
 sg13g2_fill_2 FILLER_45_2217 ();
 sg13g2_decap_8 FILLER_45_2268 ();
 sg13g2_decap_8 FILLER_45_2275 ();
 sg13g2_fill_2 FILLER_45_2291 ();
 sg13g2_decap_8 FILLER_45_2320 ();
 sg13g2_decap_4 FILLER_45_2327 ();
 sg13g2_fill_2 FILLER_45_2331 ();
 sg13g2_fill_2 FILLER_45_2350 ();
 sg13g2_fill_1 FILLER_45_2352 ();
 sg13g2_decap_8 FILLER_45_2366 ();
 sg13g2_decap_8 FILLER_45_2373 ();
 sg13g2_decap_8 FILLER_45_2380 ();
 sg13g2_fill_1 FILLER_45_2387 ();
 sg13g2_decap_8 FILLER_45_2424 ();
 sg13g2_decap_8 FILLER_45_2431 ();
 sg13g2_fill_2 FILLER_45_2447 ();
 sg13g2_fill_1 FILLER_45_2449 ();
 sg13g2_decap_4 FILLER_45_2460 ();
 sg13g2_fill_2 FILLER_45_2464 ();
 sg13g2_decap_8 FILLER_45_2479 ();
 sg13g2_decap_8 FILLER_45_2486 ();
 sg13g2_decap_8 FILLER_45_2493 ();
 sg13g2_decap_8 FILLER_45_2541 ();
 sg13g2_decap_8 FILLER_45_2548 ();
 sg13g2_decap_8 FILLER_45_2555 ();
 sg13g2_decap_4 FILLER_45_2562 ();
 sg13g2_fill_1 FILLER_45_2570 ();
 sg13g2_decap_8 FILLER_45_2607 ();
 sg13g2_decap_8 FILLER_45_2614 ();
 sg13g2_decap_8 FILLER_45_2621 ();
 sg13g2_fill_1 FILLER_45_2650 ();
 sg13g2_fill_1 FILLER_45_2655 ();
 sg13g2_fill_2 FILLER_45_2669 ();
 sg13g2_decap_8 FILLER_45_2737 ();
 sg13g2_fill_2 FILLER_45_2744 ();
 sg13g2_decap_8 FILLER_45_2751 ();
 sg13g2_decap_8 FILLER_45_2758 ();
 sg13g2_decap_8 FILLER_45_2765 ();
 sg13g2_decap_8 FILLER_45_2772 ();
 sg13g2_decap_8 FILLER_45_2779 ();
 sg13g2_decap_4 FILLER_45_2786 ();
 sg13g2_decap_8 FILLER_45_2812 ();
 sg13g2_decap_8 FILLER_45_2819 ();
 sg13g2_decap_8 FILLER_45_2826 ();
 sg13g2_decap_4 FILLER_45_2833 ();
 sg13g2_fill_1 FILLER_45_2861 ();
 sg13g2_decap_8 FILLER_45_2880 ();
 sg13g2_decap_4 FILLER_45_2887 ();
 sg13g2_decap_8 FILLER_45_2917 ();
 sg13g2_decap_8 FILLER_45_2955 ();
 sg13g2_decap_8 FILLER_45_2962 ();
 sg13g2_decap_8 FILLER_45_2969 ();
 sg13g2_decap_4 FILLER_45_2976 ();
 sg13g2_decap_8 FILLER_45_2989 ();
 sg13g2_decap_4 FILLER_45_2996 ();
 sg13g2_fill_1 FILLER_45_3000 ();
 sg13g2_decap_4 FILLER_45_3005 ();
 sg13g2_fill_2 FILLER_45_3009 ();
 sg13g2_decap_8 FILLER_45_3046 ();
 sg13g2_decap_8 FILLER_45_3053 ();
 sg13g2_decap_8 FILLER_45_3060 ();
 sg13g2_decap_8 FILLER_45_3067 ();
 sg13g2_decap_8 FILLER_45_3074 ();
 sg13g2_decap_8 FILLER_45_3081 ();
 sg13g2_fill_2 FILLER_45_3088 ();
 sg13g2_decap_8 FILLER_45_3094 ();
 sg13g2_decap_8 FILLER_45_3101 ();
 sg13g2_fill_2 FILLER_45_3108 ();
 sg13g2_fill_1 FILLER_45_3110 ();
 sg13g2_fill_2 FILLER_45_3138 ();
 sg13g2_fill_1 FILLER_45_3140 ();
 sg13g2_decap_8 FILLER_45_3154 ();
 sg13g2_fill_2 FILLER_45_3161 ();
 sg13g2_decap_8 FILLER_45_3203 ();
 sg13g2_decap_8 FILLER_45_3210 ();
 sg13g2_decap_8 FILLER_45_3217 ();
 sg13g2_decap_4 FILLER_45_3224 ();
 sg13g2_fill_1 FILLER_45_3228 ();
 sg13g2_decap_4 FILLER_45_3243 ();
 sg13g2_fill_1 FILLER_45_3247 ();
 sg13g2_decap_8 FILLER_45_3261 ();
 sg13g2_decap_8 FILLER_45_3268 ();
 sg13g2_decap_8 FILLER_45_3275 ();
 sg13g2_fill_2 FILLER_45_3282 ();
 sg13g2_fill_1 FILLER_45_3284 ();
 sg13g2_decap_4 FILLER_45_3308 ();
 sg13g2_fill_1 FILLER_45_3312 ();
 sg13g2_fill_1 FILLER_45_3336 ();
 sg13g2_decap_8 FILLER_45_3350 ();
 sg13g2_decap_8 FILLER_45_3357 ();
 sg13g2_decap_8 FILLER_45_3364 ();
 sg13g2_fill_2 FILLER_45_3371 ();
 sg13g2_decap_8 FILLER_45_3383 ();
 sg13g2_fill_1 FILLER_45_3390 ();
 sg13g2_fill_2 FILLER_45_3458 ();
 sg13g2_decap_4 FILLER_45_3511 ();
 sg13g2_fill_2 FILLER_45_3515 ();
 sg13g2_decap_8 FILLER_45_3567 ();
 sg13g2_decap_4 FILLER_45_3574 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_11 ();
 sg13g2_fill_2 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_55 ();
 sg13g2_decap_8 FILLER_46_62 ();
 sg13g2_decap_8 FILLER_46_69 ();
 sg13g2_decap_4 FILLER_46_76 ();
 sg13g2_fill_1 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_125 ();
 sg13g2_decap_8 FILLER_46_132 ();
 sg13g2_fill_2 FILLER_46_139 ();
 sg13g2_fill_1 FILLER_46_141 ();
 sg13g2_fill_2 FILLER_46_155 ();
 sg13g2_decap_8 FILLER_46_166 ();
 sg13g2_decap_8 FILLER_46_173 ();
 sg13g2_fill_1 FILLER_46_180 ();
 sg13g2_fill_1 FILLER_46_208 ();
 sg13g2_decap_8 FILLER_46_228 ();
 sg13g2_decap_8 FILLER_46_235 ();
 sg13g2_decap_8 FILLER_46_242 ();
 sg13g2_fill_2 FILLER_46_249 ();
 sg13g2_decap_8 FILLER_46_283 ();
 sg13g2_decap_8 FILLER_46_290 ();
 sg13g2_decap_8 FILLER_46_297 ();
 sg13g2_decap_8 FILLER_46_304 ();
 sg13g2_decap_4 FILLER_46_311 ();
 sg13g2_fill_1 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_339 ();
 sg13g2_decap_4 FILLER_46_346 ();
 sg13g2_fill_2 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_419 ();
 sg13g2_decap_8 FILLER_46_426 ();
 sg13g2_decap_8 FILLER_46_433 ();
 sg13g2_decap_8 FILLER_46_440 ();
 sg13g2_fill_1 FILLER_46_447 ();
 sg13g2_decap_8 FILLER_46_461 ();
 sg13g2_decap_8 FILLER_46_468 ();
 sg13g2_decap_8 FILLER_46_475 ();
 sg13g2_decap_8 FILLER_46_482 ();
 sg13g2_decap_8 FILLER_46_489 ();
 sg13g2_decap_8 FILLER_46_496 ();
 sg13g2_decap_8 FILLER_46_503 ();
 sg13g2_decap_8 FILLER_46_510 ();
 sg13g2_decap_8 FILLER_46_517 ();
 sg13g2_decap_8 FILLER_46_524 ();
 sg13g2_fill_2 FILLER_46_531 ();
 sg13g2_decap_8 FILLER_46_561 ();
 sg13g2_decap_8 FILLER_46_568 ();
 sg13g2_decap_8 FILLER_46_575 ();
 sg13g2_decap_8 FILLER_46_582 ();
 sg13g2_fill_2 FILLER_46_589 ();
 sg13g2_fill_1 FILLER_46_591 ();
 sg13g2_fill_2 FILLER_46_633 ();
 sg13g2_decap_4 FILLER_46_645 ();
 sg13g2_fill_1 FILLER_46_649 ();
 sg13g2_decap_4 FILLER_46_655 ();
 sg13g2_fill_1 FILLER_46_672 ();
 sg13g2_fill_2 FILLER_46_686 ();
 sg13g2_fill_1 FILLER_46_688 ();
 sg13g2_decap_8 FILLER_46_713 ();
 sg13g2_decap_8 FILLER_46_720 ();
 sg13g2_decap_4 FILLER_46_727 ();
 sg13g2_decap_4 FILLER_46_776 ();
 sg13g2_fill_1 FILLER_46_780 ();
 sg13g2_decap_4 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_795 ();
 sg13g2_decap_8 FILLER_46_802 ();
 sg13g2_decap_8 FILLER_46_809 ();
 sg13g2_fill_2 FILLER_46_816 ();
 sg13g2_fill_1 FILLER_46_818 ();
 sg13g2_decap_8 FILLER_46_823 ();
 sg13g2_fill_1 FILLER_46_830 ();
 sg13g2_decap_4 FILLER_46_845 ();
 sg13g2_decap_4 FILLER_46_859 ();
 sg13g2_fill_1 FILLER_46_863 ();
 sg13g2_decap_4 FILLER_46_873 ();
 sg13g2_fill_2 FILLER_46_877 ();
 sg13g2_decap_8 FILLER_46_883 ();
 sg13g2_decap_4 FILLER_46_890 ();
 sg13g2_fill_1 FILLER_46_894 ();
 sg13g2_decap_4 FILLER_46_900 ();
 sg13g2_fill_2 FILLER_46_904 ();
 sg13g2_fill_2 FILLER_46_910 ();
 sg13g2_fill_1 FILLER_46_912 ();
 sg13g2_decap_8 FILLER_46_922 ();
 sg13g2_decap_8 FILLER_46_934 ();
 sg13g2_fill_2 FILLER_46_953 ();
 sg13g2_fill_1 FILLER_46_955 ();
 sg13g2_decap_8 FILLER_46_960 ();
 sg13g2_decap_8 FILLER_46_967 ();
 sg13g2_decap_8 FILLER_46_974 ();
 sg13g2_fill_1 FILLER_46_981 ();
 sg13g2_decap_8 FILLER_46_991 ();
 sg13g2_decap_4 FILLER_46_998 ();
 sg13g2_fill_2 FILLER_46_1002 ();
 sg13g2_decap_8 FILLER_46_1017 ();
 sg13g2_decap_8 FILLER_46_1024 ();
 sg13g2_decap_8 FILLER_46_1031 ();
 sg13g2_decap_8 FILLER_46_1038 ();
 sg13g2_fill_1 FILLER_46_1045 ();
 sg13g2_decap_8 FILLER_46_1055 ();
 sg13g2_fill_2 FILLER_46_1062 ();
 sg13g2_fill_2 FILLER_46_1077 ();
 sg13g2_fill_1 FILLER_46_1079 ();
 sg13g2_fill_2 FILLER_46_1086 ();
 sg13g2_fill_1 FILLER_46_1100 ();
 sg13g2_fill_1 FILLER_46_1147 ();
 sg13g2_fill_2 FILLER_46_1163 ();
 sg13g2_fill_2 FILLER_46_1178 ();
 sg13g2_fill_2 FILLER_46_1209 ();
 sg13g2_fill_2 FILLER_46_1239 ();
 sg13g2_fill_1 FILLER_46_1241 ();
 sg13g2_fill_2 FILLER_46_1256 ();
 sg13g2_fill_2 FILLER_46_1273 ();
 sg13g2_decap_4 FILLER_46_1297 ();
 sg13g2_decap_4 FILLER_46_1315 ();
 sg13g2_fill_1 FILLER_46_1324 ();
 sg13g2_decap_8 FILLER_46_1330 ();
 sg13g2_fill_2 FILLER_46_1337 ();
 sg13g2_fill_1 FILLER_46_1339 ();
 sg13g2_fill_1 FILLER_46_1353 ();
 sg13g2_decap_4 FILLER_46_1400 ();
 sg13g2_fill_2 FILLER_46_1404 ();
 sg13g2_fill_1 FILLER_46_1453 ();
 sg13g2_decap_8 FILLER_46_1467 ();
 sg13g2_fill_2 FILLER_46_1474 ();
 sg13g2_fill_1 FILLER_46_1476 ();
 sg13g2_fill_2 FILLER_46_1486 ();
 sg13g2_fill_1 FILLER_46_1488 ();
 sg13g2_decap_8 FILLER_46_1499 ();
 sg13g2_fill_1 FILLER_46_1506 ();
 sg13g2_decap_4 FILLER_46_1512 ();
 sg13g2_fill_2 FILLER_46_1516 ();
 sg13g2_fill_2 FILLER_46_1535 ();
 sg13g2_fill_1 FILLER_46_1537 ();
 sg13g2_decap_8 FILLER_46_1546 ();
 sg13g2_decap_4 FILLER_46_1553 ();
 sg13g2_fill_1 FILLER_46_1557 ();
 sg13g2_decap_4 FILLER_46_1603 ();
 sg13g2_decap_8 FILLER_46_1624 ();
 sg13g2_decap_8 FILLER_46_1631 ();
 sg13g2_decap_8 FILLER_46_1638 ();
 sg13g2_fill_2 FILLER_46_1645 ();
 sg13g2_fill_1 FILLER_46_1647 ();
 sg13g2_decap_8 FILLER_46_1658 ();
 sg13g2_fill_2 FILLER_46_1665 ();
 sg13g2_fill_1 FILLER_46_1667 ();
 sg13g2_fill_1 FILLER_46_1685 ();
 sg13g2_decap_4 FILLER_46_1698 ();
 sg13g2_fill_1 FILLER_46_1702 ();
 sg13g2_decap_8 FILLER_46_1711 ();
 sg13g2_decap_8 FILLER_46_1718 ();
 sg13g2_decap_8 FILLER_46_1725 ();
 sg13g2_fill_2 FILLER_46_1732 ();
 sg13g2_fill_2 FILLER_46_1747 ();
 sg13g2_fill_1 FILLER_46_1749 ();
 sg13g2_decap_8 FILLER_46_1771 ();
 sg13g2_decap_8 FILLER_46_1778 ();
 sg13g2_decap_8 FILLER_46_1785 ();
 sg13g2_decap_8 FILLER_46_1792 ();
 sg13g2_decap_8 FILLER_46_1799 ();
 sg13g2_fill_2 FILLER_46_1806 ();
 sg13g2_fill_1 FILLER_46_1808 ();
 sg13g2_fill_1 FILLER_46_1827 ();
 sg13g2_decap_4 FILLER_46_1836 ();
 sg13g2_fill_1 FILLER_46_1840 ();
 sg13g2_decap_8 FILLER_46_1854 ();
 sg13g2_decap_8 FILLER_46_1861 ();
 sg13g2_fill_2 FILLER_46_1868 ();
 sg13g2_fill_1 FILLER_46_1870 ();
 sg13g2_decap_8 FILLER_46_1876 ();
 sg13g2_decap_8 FILLER_46_1883 ();
 sg13g2_fill_2 FILLER_46_1890 ();
 sg13g2_fill_1 FILLER_46_1892 ();
 sg13g2_fill_2 FILLER_46_1897 ();
 sg13g2_fill_1 FILLER_46_1904 ();
 sg13g2_decap_8 FILLER_46_1931 ();
 sg13g2_decap_8 FILLER_46_1938 ();
 sg13g2_decap_8 FILLER_46_1945 ();
 sg13g2_fill_1 FILLER_46_1952 ();
 sg13g2_fill_2 FILLER_46_1971 ();
 sg13g2_fill_2 FILLER_46_2007 ();
 sg13g2_fill_2 FILLER_46_2030 ();
 sg13g2_decap_8 FILLER_46_2049 ();
 sg13g2_fill_1 FILLER_46_2061 ();
 sg13g2_decap_8 FILLER_46_2084 ();
 sg13g2_decap_8 FILLER_46_2091 ();
 sg13g2_decap_8 FILLER_46_2098 ();
 sg13g2_decap_8 FILLER_46_2105 ();
 sg13g2_decap_8 FILLER_46_2112 ();
 sg13g2_fill_1 FILLER_46_2119 ();
 sg13g2_decap_8 FILLER_46_2137 ();
 sg13g2_decap_4 FILLER_46_2144 ();
 sg13g2_fill_2 FILLER_46_2148 ();
 sg13g2_fill_1 FILLER_46_2227 ();
 sg13g2_decap_8 FILLER_46_2250 ();
 sg13g2_decap_8 FILLER_46_2257 ();
 sg13g2_decap_8 FILLER_46_2264 ();
 sg13g2_decap_8 FILLER_46_2271 ();
 sg13g2_decap_8 FILLER_46_2278 ();
 sg13g2_fill_2 FILLER_46_2349 ();
 sg13g2_fill_1 FILLER_46_2351 ();
 sg13g2_decap_8 FILLER_46_2379 ();
 sg13g2_fill_2 FILLER_46_2386 ();
 sg13g2_fill_2 FILLER_46_2415 ();
 sg13g2_fill_1 FILLER_46_2417 ();
 sg13g2_decap_8 FILLER_46_2491 ();
 sg13g2_decap_4 FILLER_46_2498 ();
 sg13g2_decap_4 FILLER_46_2552 ();
 sg13g2_fill_1 FILLER_46_2556 ();
 sg13g2_decap_8 FILLER_46_2609 ();
 sg13g2_decap_8 FILLER_46_2616 ();
 sg13g2_decap_4 FILLER_46_2623 ();
 sg13g2_fill_2 FILLER_46_2627 ();
 sg13g2_decap_4 FILLER_46_2639 ();
 sg13g2_fill_2 FILLER_46_2643 ();
 sg13g2_decap_8 FILLER_46_2666 ();
 sg13g2_decap_8 FILLER_46_2673 ();
 sg13g2_decap_8 FILLER_46_2707 ();
 sg13g2_fill_2 FILLER_46_2714 ();
 sg13g2_decap_8 FILLER_46_2764 ();
 sg13g2_decap_8 FILLER_46_2771 ();
 sg13g2_decap_8 FILLER_46_2815 ();
 sg13g2_decap_8 FILLER_46_2886 ();
 sg13g2_decap_8 FILLER_46_2893 ();
 sg13g2_decap_8 FILLER_46_2900 ();
 sg13g2_decap_8 FILLER_46_2907 ();
 sg13g2_fill_2 FILLER_46_2914 ();
 sg13g2_fill_1 FILLER_46_2916 ();
 sg13g2_fill_2 FILLER_46_2957 ();
 sg13g2_fill_1 FILLER_46_2959 ();
 sg13g2_decap_8 FILLER_46_2965 ();
 sg13g2_decap_4 FILLER_46_2972 ();
 sg13g2_fill_1 FILLER_46_2976 ();
 sg13g2_fill_2 FILLER_46_2991 ();
 sg13g2_decap_8 FILLER_46_3002 ();
 sg13g2_decap_8 FILLER_46_3009 ();
 sg13g2_decap_8 FILLER_46_3042 ();
 sg13g2_fill_2 FILLER_46_3049 ();
 sg13g2_decap_8 FILLER_46_3088 ();
 sg13g2_decap_8 FILLER_46_3095 ();
 sg13g2_decap_8 FILLER_46_3133 ();
 sg13g2_decap_4 FILLER_46_3140 ();
 sg13g2_fill_2 FILLER_46_3157 ();
 sg13g2_decap_8 FILLER_46_3205 ();
 sg13g2_decap_8 FILLER_46_3212 ();
 sg13g2_decap_8 FILLER_46_3219 ();
 sg13g2_decap_4 FILLER_46_3226 ();
 sg13g2_fill_1 FILLER_46_3230 ();
 sg13g2_fill_2 FILLER_46_3284 ();
 sg13g2_decap_8 FILLER_46_3352 ();
 sg13g2_decap_8 FILLER_46_3359 ();
 sg13g2_fill_2 FILLER_46_3366 ();
 sg13g2_fill_1 FILLER_46_3368 ();
 sg13g2_fill_2 FILLER_46_3396 ();
 sg13g2_decap_8 FILLER_46_3425 ();
 sg13g2_decap_8 FILLER_46_3432 ();
 sg13g2_decap_8 FILLER_46_3439 ();
 sg13g2_decap_4 FILLER_46_3446 ();
 sg13g2_fill_1 FILLER_46_3450 ();
 sg13g2_fill_2 FILLER_46_3482 ();
 sg13g2_fill_1 FILLER_46_3484 ();
 sg13g2_fill_1 FILLER_46_3498 ();
 sg13g2_decap_4 FILLER_46_3572 ();
 sg13g2_fill_2 FILLER_46_3576 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_42 ();
 sg13g2_fill_1 FILLER_47_73 ();
 sg13g2_decap_8 FILLER_47_128 ();
 sg13g2_decap_8 FILLER_47_135 ();
 sg13g2_fill_1 FILLER_47_142 ();
 sg13g2_decap_8 FILLER_47_170 ();
 sg13g2_decap_8 FILLER_47_177 ();
 sg13g2_decap_4 FILLER_47_184 ();
 sg13g2_fill_1 FILLER_47_188 ();
 sg13g2_fill_1 FILLER_47_223 ();
 sg13g2_fill_1 FILLER_47_237 ();
 sg13g2_decap_8 FILLER_47_242 ();
 sg13g2_fill_2 FILLER_47_249 ();
 sg13g2_fill_2 FILLER_47_259 ();
 sg13g2_fill_1 FILLER_47_275 ();
 sg13g2_decap_4 FILLER_47_317 ();
 sg13g2_fill_1 FILLER_47_321 ();
 sg13g2_decap_8 FILLER_47_335 ();
 sg13g2_decap_8 FILLER_47_342 ();
 sg13g2_decap_8 FILLER_47_389 ();
 sg13g2_fill_2 FILLER_47_396 ();
 sg13g2_decap_8 FILLER_47_415 ();
 sg13g2_decap_8 FILLER_47_422 ();
 sg13g2_decap_8 FILLER_47_429 ();
 sg13g2_fill_1 FILLER_47_468 ();
 sg13g2_decap_8 FILLER_47_496 ();
 sg13g2_decap_8 FILLER_47_503 ();
 sg13g2_decap_8 FILLER_47_510 ();
 sg13g2_fill_1 FILLER_47_517 ();
 sg13g2_decap_8 FILLER_47_559 ();
 sg13g2_decap_4 FILLER_47_566 ();
 sg13g2_fill_2 FILLER_47_570 ();
 sg13g2_decap_8 FILLER_47_576 ();
 sg13g2_fill_2 FILLER_47_583 ();
 sg13g2_decap_8 FILLER_47_618 ();
 sg13g2_decap_4 FILLER_47_625 ();
 sg13g2_fill_2 FILLER_47_634 ();
 sg13g2_fill_2 FILLER_47_660 ();
 sg13g2_decap_8 FILLER_47_671 ();
 sg13g2_decap_8 FILLER_47_678 ();
 sg13g2_decap_4 FILLER_47_711 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_766 ();
 sg13g2_decap_8 FILLER_47_799 ();
 sg13g2_fill_2 FILLER_47_806 ();
 sg13g2_fill_1 FILLER_47_808 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_fill_1 FILLER_47_843 ();
 sg13g2_decap_8 FILLER_47_849 ();
 sg13g2_fill_2 FILLER_47_856 ();
 sg13g2_fill_1 FILLER_47_858 ();
 sg13g2_decap_4 FILLER_47_868 ();
 sg13g2_fill_1 FILLER_47_872 ();
 sg13g2_fill_1 FILLER_47_882 ();
 sg13g2_fill_1 FILLER_47_892 ();
 sg13g2_fill_1 FILLER_47_921 ();
 sg13g2_fill_1 FILLER_47_931 ();
 sg13g2_fill_1 FILLER_47_954 ();
 sg13g2_fill_1 FILLER_47_982 ();
 sg13g2_fill_2 FILLER_47_1025 ();
 sg13g2_fill_1 FILLER_47_1027 ();
 sg13g2_fill_1 FILLER_47_1033 ();
 sg13g2_decap_8 FILLER_47_1040 ();
 sg13g2_decap_4 FILLER_47_1047 ();
 sg13g2_fill_2 FILLER_47_1051 ();
 sg13g2_fill_2 FILLER_47_1094 ();
 sg13g2_fill_1 FILLER_47_1096 ();
 sg13g2_fill_1 FILLER_47_1134 ();
 sg13g2_fill_1 FILLER_47_1150 ();
 sg13g2_fill_2 FILLER_47_1160 ();
 sg13g2_fill_1 FILLER_47_1162 ();
 sg13g2_fill_1 FILLER_47_1192 ();
 sg13g2_decap_4 FILLER_47_1227 ();
 sg13g2_fill_2 FILLER_47_1231 ();
 sg13g2_fill_2 FILLER_47_1254 ();
 sg13g2_fill_1 FILLER_47_1283 ();
 sg13g2_decap_8 FILLER_47_1322 ();
 sg13g2_decap_4 FILLER_47_1329 ();
 sg13g2_fill_2 FILLER_47_1333 ();
 sg13g2_decap_8 FILLER_47_1402 ();
 sg13g2_fill_1 FILLER_47_1409 ();
 sg13g2_decap_8 FILLER_47_1431 ();
 sg13g2_decap_8 FILLER_47_1438 ();
 sg13g2_decap_8 FILLER_47_1445 ();
 sg13g2_decap_8 FILLER_47_1452 ();
 sg13g2_decap_8 FILLER_47_1459 ();
 sg13g2_decap_4 FILLER_47_1466 ();
 sg13g2_fill_1 FILLER_47_1470 ();
 sg13g2_fill_2 FILLER_47_1476 ();
 sg13g2_fill_2 FILLER_47_1483 ();
 sg13g2_fill_2 FILLER_47_1507 ();
 sg13g2_fill_1 FILLER_47_1533 ();
 sg13g2_decap_4 FILLER_47_1540 ();
 sg13g2_fill_1 FILLER_47_1544 ();
 sg13g2_fill_1 FILLER_47_1555 ();
 sg13g2_fill_2 FILLER_47_1572 ();
 sg13g2_fill_1 FILLER_47_1574 ();
 sg13g2_fill_2 FILLER_47_1590 ();
 sg13g2_fill_1 FILLER_47_1592 ();
 sg13g2_fill_1 FILLER_47_1606 ();
 sg13g2_decap_8 FILLER_47_1625 ();
 sg13g2_decap_8 FILLER_47_1632 ();
 sg13g2_decap_4 FILLER_47_1639 ();
 sg13g2_decap_4 FILLER_47_1664 ();
 sg13g2_decap_8 FILLER_47_1704 ();
 sg13g2_decap_8 FILLER_47_1711 ();
 sg13g2_decap_4 FILLER_47_1718 ();
 sg13g2_fill_2 FILLER_47_1740 ();
 sg13g2_fill_1 FILLER_47_1742 ();
 sg13g2_decap_8 FILLER_47_1764 ();
 sg13g2_decap_8 FILLER_47_1771 ();
 sg13g2_decap_4 FILLER_47_1778 ();
 sg13g2_fill_2 FILLER_47_1782 ();
 sg13g2_decap_4 FILLER_47_1792 ();
 sg13g2_fill_1 FILLER_47_1796 ();
 sg13g2_decap_4 FILLER_47_1807 ();
 sg13g2_fill_1 FILLER_47_1816 ();
 sg13g2_decap_8 FILLER_47_1827 ();
 sg13g2_decap_8 FILLER_47_1834 ();
 sg13g2_fill_2 FILLER_47_1841 ();
 sg13g2_fill_2 FILLER_47_1859 ();
 sg13g2_fill_1 FILLER_47_1861 ();
 sg13g2_decap_8 FILLER_47_1866 ();
 sg13g2_decap_8 FILLER_47_1873 ();
 sg13g2_fill_2 FILLER_47_1880 ();
 sg13g2_fill_1 FILLER_47_1882 ();
 sg13g2_fill_2 FILLER_47_1888 ();
 sg13g2_fill_1 FILLER_47_1904 ();
 sg13g2_decap_8 FILLER_47_1921 ();
 sg13g2_decap_8 FILLER_47_1928 ();
 sg13g2_decap_8 FILLER_47_1935 ();
 sg13g2_fill_2 FILLER_47_1942 ();
 sg13g2_fill_1 FILLER_47_1944 ();
 sg13g2_fill_1 FILLER_47_1980 ();
 sg13g2_decap_4 FILLER_47_1986 ();
 sg13g2_fill_1 FILLER_47_1990 ();
 sg13g2_fill_2 FILLER_47_2004 ();
 sg13g2_fill_1 FILLER_47_2006 ();
 sg13g2_fill_1 FILLER_47_2020 ();
 sg13g2_fill_1 FILLER_47_2030 ();
 sg13g2_fill_1 FILLER_47_2039 ();
 sg13g2_decap_8 FILLER_47_2044 ();
 sg13g2_decap_8 FILLER_47_2055 ();
 sg13g2_decap_4 FILLER_47_2062 ();
 sg13g2_decap_8 FILLER_47_2109 ();
 sg13g2_decap_8 FILLER_47_2116 ();
 sg13g2_fill_1 FILLER_47_2123 ();
 sg13g2_decap_8 FILLER_47_2129 ();
 sg13g2_decap_8 FILLER_47_2136 ();
 sg13g2_decap_4 FILLER_47_2143 ();
 sg13g2_fill_2 FILLER_47_2174 ();
 sg13g2_fill_2 FILLER_47_2185 ();
 sg13g2_fill_1 FILLER_47_2187 ();
 sg13g2_decap_8 FILLER_47_2251 ();
 sg13g2_fill_2 FILLER_47_2262 ();
 sg13g2_fill_1 FILLER_47_2264 ();
 sg13g2_decap_4 FILLER_47_2270 ();
 sg13g2_fill_2 FILLER_47_2274 ();
 sg13g2_fill_2 FILLER_47_2304 ();
 sg13g2_fill_2 FILLER_47_2319 ();
 sg13g2_fill_1 FILLER_47_2321 ();
 sg13g2_decap_4 FILLER_47_2327 ();
 sg13g2_fill_1 FILLER_47_2331 ();
 sg13g2_fill_2 FILLER_47_2354 ();
 sg13g2_fill_1 FILLER_47_2356 ();
 sg13g2_decap_8 FILLER_47_2361 ();
 sg13g2_decap_8 FILLER_47_2368 ();
 sg13g2_decap_4 FILLER_47_2375 ();
 sg13g2_decap_8 FILLER_47_2441 ();
 sg13g2_fill_1 FILLER_47_2448 ();
 sg13g2_decap_8 FILLER_47_2490 ();
 sg13g2_fill_2 FILLER_47_2497 ();
 sg13g2_fill_1 FILLER_47_2499 ();
 sg13g2_fill_2 FILLER_47_2509 ();
 sg13g2_decap_8 FILLER_47_2549 ();
 sg13g2_decap_8 FILLER_47_2556 ();
 sg13g2_fill_2 FILLER_47_2563 ();
 sg13g2_fill_1 FILLER_47_2575 ();
 sg13g2_fill_2 FILLER_47_2603 ();
 sg13g2_fill_1 FILLER_47_2605 ();
 sg13g2_decap_4 FILLER_47_2673 ();
 sg13g2_fill_2 FILLER_47_2687 ();
 sg13g2_decap_8 FILLER_47_2702 ();
 sg13g2_decap_8 FILLER_47_2709 ();
 sg13g2_decap_8 FILLER_47_2716 ();
 sg13g2_decap_4 FILLER_47_2723 ();
 sg13g2_decap_8 FILLER_47_2764 ();
 sg13g2_decap_4 FILLER_47_2771 ();
 sg13g2_decap_8 FILLER_47_2820 ();
 sg13g2_decap_8 FILLER_47_2827 ();
 sg13g2_fill_2 FILLER_47_2834 ();
 sg13g2_fill_1 FILLER_47_2836 ();
 sg13g2_decap_8 FILLER_47_2841 ();
 sg13g2_fill_2 FILLER_47_2862 ();
 sg13g2_fill_1 FILLER_47_2864 ();
 sg13g2_decap_8 FILLER_47_2895 ();
 sg13g2_decap_8 FILLER_47_2902 ();
 sg13g2_decap_8 FILLER_47_2909 ();
 sg13g2_decap_8 FILLER_47_2966 ();
 sg13g2_fill_1 FILLER_47_2973 ();
 sg13g2_decap_8 FILLER_47_3005 ();
 sg13g2_fill_2 FILLER_47_3012 ();
 sg13g2_decap_4 FILLER_47_3024 ();
 sg13g2_fill_2 FILLER_47_3028 ();
 sg13g2_decap_8 FILLER_47_3039 ();
 sg13g2_fill_1 FILLER_47_3046 ();
 sg13g2_decap_4 FILLER_47_3093 ();
 sg13g2_fill_1 FILLER_47_3097 ();
 sg13g2_decap_8 FILLER_47_3134 ();
 sg13g2_decap_4 FILLER_47_3141 ();
 sg13g2_fill_1 FILLER_47_3163 ();
 sg13g2_fill_1 FILLER_47_3184 ();
 sg13g2_decap_8 FILLER_47_3206 ();
 sg13g2_decap_8 FILLER_47_3213 ();
 sg13g2_decap_8 FILLER_47_3220 ();
 sg13g2_fill_1 FILLER_47_3264 ();
 sg13g2_decap_8 FILLER_47_3278 ();
 sg13g2_fill_2 FILLER_47_3285 ();
 sg13g2_decap_4 FILLER_47_3336 ();
 sg13g2_decap_4 FILLER_47_3353 ();
 sg13g2_fill_1 FILLER_47_3357 ();
 sg13g2_fill_2 FILLER_47_3410 ();
 sg13g2_decap_8 FILLER_47_3425 ();
 sg13g2_decap_8 FILLER_47_3432 ();
 sg13g2_decap_8 FILLER_47_3439 ();
 sg13g2_decap_8 FILLER_47_3446 ();
 sg13g2_fill_2 FILLER_47_3453 ();
 sg13g2_fill_1 FILLER_47_3455 ();
 sg13g2_decap_8 FILLER_47_3502 ();
 sg13g2_decap_8 FILLER_47_3509 ();
 sg13g2_decap_8 FILLER_47_3558 ();
 sg13g2_decap_8 FILLER_47_3565 ();
 sg13g2_decap_4 FILLER_47_3572 ();
 sg13g2_fill_2 FILLER_47_3576 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_4 FILLER_48_14 ();
 sg13g2_fill_2 FILLER_48_18 ();
 sg13g2_decap_4 FILLER_48_24 ();
 sg13g2_fill_1 FILLER_48_28 ();
 sg13g2_decap_4 FILLER_48_58 ();
 sg13g2_fill_1 FILLER_48_62 ();
 sg13g2_decap_8 FILLER_48_72 ();
 sg13g2_decap_4 FILLER_48_79 ();
 sg13g2_fill_1 FILLER_48_83 ();
 sg13g2_decap_4 FILLER_48_94 ();
 sg13g2_fill_2 FILLER_48_98 ();
 sg13g2_fill_1 FILLER_48_119 ();
 sg13g2_decap_4 FILLER_48_135 ();
 sg13g2_decap_4 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_180 ();
 sg13g2_decap_8 FILLER_48_240 ();
 sg13g2_decap_8 FILLER_48_247 ();
 sg13g2_decap_4 FILLER_48_254 ();
 sg13g2_fill_2 FILLER_48_258 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_4 FILLER_48_287 ();
 sg13g2_fill_1 FILLER_48_291 ();
 sg13g2_decap_4 FILLER_48_319 ();
 sg13g2_fill_2 FILLER_48_351 ();
 sg13g2_decap_4 FILLER_48_384 ();
 sg13g2_decap_8 FILLER_48_424 ();
 sg13g2_decap_4 FILLER_48_431 ();
 sg13g2_fill_1 FILLER_48_435 ();
 sg13g2_fill_1 FILLER_48_475 ();
 sg13g2_decap_4 FILLER_48_494 ();
 sg13g2_decap_8 FILLER_48_526 ();
 sg13g2_fill_2 FILLER_48_533 ();
 sg13g2_decap_4 FILLER_48_563 ();
 sg13g2_fill_1 FILLER_48_575 ();
 sg13g2_decap_8 FILLER_48_606 ();
 sg13g2_decap_4 FILLER_48_613 ();
 sg13g2_fill_1 FILLER_48_617 ();
 sg13g2_fill_2 FILLER_48_631 ();
 sg13g2_fill_2 FILLER_48_645 ();
 sg13g2_decap_4 FILLER_48_675 ();
 sg13g2_fill_2 FILLER_48_712 ();
 sg13g2_fill_2 FILLER_48_760 ();
 sg13g2_decap_4 FILLER_48_766 ();
 sg13g2_fill_1 FILLER_48_834 ();
 sg13g2_decap_8 FILLER_48_845 ();
 sg13g2_fill_2 FILLER_48_880 ();
 sg13g2_fill_1 FILLER_48_909 ();
 sg13g2_decap_4 FILLER_48_916 ();
 sg13g2_decap_8 FILLER_48_1009 ();
 sg13g2_fill_1 FILLER_48_1016 ();
 sg13g2_fill_2 FILLER_48_1022 ();
 sg13g2_fill_1 FILLER_48_1024 ();
 sg13g2_fill_1 FILLER_48_1033 ();
 sg13g2_fill_2 FILLER_48_1092 ();
 sg13g2_decap_8 FILLER_48_1109 ();
 sg13g2_decap_8 FILLER_48_1116 ();
 sg13g2_fill_1 FILLER_48_1123 ();
 sg13g2_fill_2 FILLER_48_1186 ();
 sg13g2_fill_1 FILLER_48_1188 ();
 sg13g2_decap_8 FILLER_48_1194 ();
 sg13g2_fill_1 FILLER_48_1201 ();
 sg13g2_fill_2 FILLER_48_1207 ();
 sg13g2_fill_2 FILLER_48_1247 ();
 sg13g2_fill_2 FILLER_48_1253 ();
 sg13g2_fill_1 FILLER_48_1255 ();
 sg13g2_decap_8 FILLER_48_1261 ();
 sg13g2_decap_8 FILLER_48_1268 ();
 sg13g2_fill_2 FILLER_48_1275 ();
 sg13g2_decap_8 FILLER_48_1327 ();
 sg13g2_decap_8 FILLER_48_1334 ();
 sg13g2_fill_1 FILLER_48_1372 ();
 sg13g2_decap_8 FILLER_48_1395 ();
 sg13g2_decap_8 FILLER_48_1402 ();
 sg13g2_fill_2 FILLER_48_1409 ();
 sg13g2_decap_4 FILLER_48_1416 ();
 sg13g2_fill_2 FILLER_48_1420 ();
 sg13g2_decap_8 FILLER_48_1430 ();
 sg13g2_decap_8 FILLER_48_1437 ();
 sg13g2_decap_8 FILLER_48_1444 ();
 sg13g2_decap_8 FILLER_48_1451 ();
 sg13g2_decap_8 FILLER_48_1458 ();
 sg13g2_decap_4 FILLER_48_1465 ();
 sg13g2_fill_1 FILLER_48_1469 ();
 sg13g2_fill_2 FILLER_48_1496 ();
 sg13g2_decap_8 FILLER_48_1515 ();
 sg13g2_decap_8 FILLER_48_1522 ();
 sg13g2_decap_8 FILLER_48_1529 ();
 sg13g2_decap_8 FILLER_48_1536 ();
 sg13g2_decap_8 FILLER_48_1543 ();
 sg13g2_decap_4 FILLER_48_1550 ();
 sg13g2_fill_2 FILLER_48_1572 ();
 sg13g2_fill_1 FILLER_48_1574 ();
 sg13g2_decap_4 FILLER_48_1608 ();
 sg13g2_fill_2 FILLER_48_1612 ();
 sg13g2_decap_8 FILLER_48_1622 ();
 sg13g2_decap_8 FILLER_48_1629 ();
 sg13g2_decap_8 FILLER_48_1636 ();
 sg13g2_decap_8 FILLER_48_1643 ();
 sg13g2_decap_8 FILLER_48_1650 ();
 sg13g2_decap_8 FILLER_48_1657 ();
 sg13g2_decap_8 FILLER_48_1664 ();
 sg13g2_fill_2 FILLER_48_1671 ();
 sg13g2_decap_8 FILLER_48_1700 ();
 sg13g2_decap_8 FILLER_48_1707 ();
 sg13g2_fill_2 FILLER_48_1714 ();
 sg13g2_decap_8 FILLER_48_1747 ();
 sg13g2_fill_1 FILLER_48_1754 ();
 sg13g2_decap_8 FILLER_48_1759 ();
 sg13g2_decap_4 FILLER_48_1766 ();
 sg13g2_fill_1 FILLER_48_1770 ();
 sg13g2_fill_2 FILLER_48_1778 ();
 sg13g2_fill_1 FILLER_48_1780 ();
 sg13g2_decap_8 FILLER_48_1802 ();
 sg13g2_decap_8 FILLER_48_1827 ();
 sg13g2_decap_8 FILLER_48_1834 ();
 sg13g2_fill_2 FILLER_48_1841 ();
 sg13g2_fill_2 FILLER_48_1888 ();
 sg13g2_fill_1 FILLER_48_1890 ();
 sg13g2_decap_8 FILLER_48_1910 ();
 sg13g2_decap_8 FILLER_48_1917 ();
 sg13g2_decap_8 FILLER_48_1924 ();
 sg13g2_fill_2 FILLER_48_1931 ();
 sg13g2_decap_8 FILLER_48_1937 ();
 sg13g2_fill_2 FILLER_48_1944 ();
 sg13g2_decap_4 FILLER_48_1970 ();
 sg13g2_fill_1 FILLER_48_1974 ();
 sg13g2_fill_1 FILLER_48_1999 ();
 sg13g2_fill_2 FILLER_48_2010 ();
 sg13g2_decap_8 FILLER_48_2020 ();
 sg13g2_fill_1 FILLER_48_2027 ();
 sg13g2_fill_2 FILLER_48_2035 ();
 sg13g2_fill_1 FILLER_48_2037 ();
 sg13g2_fill_1 FILLER_48_2051 ();
 sg13g2_decap_8 FILLER_48_2066 ();
 sg13g2_fill_1 FILLER_48_2073 ();
 sg13g2_decap_8 FILLER_48_2083 ();
 sg13g2_decap_4 FILLER_48_2090 ();
 sg13g2_decap_8 FILLER_48_2121 ();
 sg13g2_decap_8 FILLER_48_2128 ();
 sg13g2_decap_8 FILLER_48_2135 ();
 sg13g2_fill_2 FILLER_48_2142 ();
 sg13g2_fill_1 FILLER_48_2144 ();
 sg13g2_decap_4 FILLER_48_2220 ();
 sg13g2_fill_2 FILLER_48_2224 ();
 sg13g2_decap_8 FILLER_48_2280 ();
 sg13g2_decap_8 FILLER_48_2287 ();
 sg13g2_decap_4 FILLER_48_2294 ();
 sg13g2_fill_1 FILLER_48_2302 ();
 sg13g2_decap_8 FILLER_48_2338 ();
 sg13g2_decap_8 FILLER_48_2345 ();
 sg13g2_fill_1 FILLER_48_2352 ();
 sg13g2_decap_8 FILLER_48_2367 ();
 sg13g2_decap_8 FILLER_48_2374 ();
 sg13g2_fill_1 FILLER_48_2381 ();
 sg13g2_fill_2 FILLER_48_2422 ();
 sg13g2_decap_8 FILLER_48_2437 ();
 sg13g2_decap_8 FILLER_48_2444 ();
 sg13g2_fill_1 FILLER_48_2451 ();
 sg13g2_decap_4 FILLER_48_2478 ();
 sg13g2_fill_2 FILLER_48_2482 ();
 sg13g2_decap_8 FILLER_48_2504 ();
 sg13g2_fill_1 FILLER_48_2511 ();
 sg13g2_decap_8 FILLER_48_2534 ();
 sg13g2_decap_8 FILLER_48_2541 ();
 sg13g2_fill_1 FILLER_48_2548 ();
 sg13g2_fill_1 FILLER_48_2575 ();
 sg13g2_decap_8 FILLER_48_2604 ();
 sg13g2_decap_4 FILLER_48_2611 ();
 sg13g2_fill_1 FILLER_48_2615 ();
 sg13g2_fill_2 FILLER_48_2663 ();
 sg13g2_decap_4 FILLER_48_2726 ();
 sg13g2_fill_1 FILLER_48_2740 ();
 sg13g2_decap_8 FILLER_48_2767 ();
 sg13g2_decap_4 FILLER_48_2774 ();
 sg13g2_decap_8 FILLER_48_2819 ();
 sg13g2_decap_8 FILLER_48_2826 ();
 sg13g2_decap_8 FILLER_48_2833 ();
 sg13g2_decap_4 FILLER_48_2840 ();
 sg13g2_fill_1 FILLER_48_2844 ();
 sg13g2_decap_8 FILLER_48_2896 ();
 sg13g2_decap_8 FILLER_48_2903 ();
 sg13g2_decap_8 FILLER_48_2910 ();
 sg13g2_fill_1 FILLER_48_2917 ();
 sg13g2_decap_8 FILLER_48_2960 ();
 sg13g2_fill_2 FILLER_48_2967 ();
 sg13g2_fill_1 FILLER_48_2969 ();
 sg13g2_decap_8 FILLER_48_3016 ();
 sg13g2_decap_8 FILLER_48_3023 ();
 sg13g2_decap_8 FILLER_48_3030 ();
 sg13g2_decap_4 FILLER_48_3037 ();
 sg13g2_fill_1 FILLER_48_3041 ();
 sg13g2_decap_8 FILLER_48_3086 ();
 sg13g2_decap_8 FILLER_48_3093 ();
 sg13g2_decap_4 FILLER_48_3100 ();
 sg13g2_fill_2 FILLER_48_3104 ();
 sg13g2_decap_4 FILLER_48_3116 ();
 sg13g2_fill_2 FILLER_48_3120 ();
 sg13g2_decap_8 FILLER_48_3131 ();
 sg13g2_decap_4 FILLER_48_3138 ();
 sg13g2_fill_1 FILLER_48_3142 ();
 sg13g2_decap_8 FILLER_48_3156 ();
 sg13g2_decap_4 FILLER_48_3163 ();
 sg13g2_decap_8 FILLER_48_3207 ();
 sg13g2_decap_4 FILLER_48_3214 ();
 sg13g2_decap_4 FILLER_48_3276 ();
 sg13g2_fill_2 FILLER_48_3280 ();
 sg13g2_fill_2 FILLER_48_3326 ();
 sg13g2_fill_2 FILLER_48_3365 ();
 sg13g2_fill_2 FILLER_48_3381 ();
 sg13g2_fill_1 FILLER_48_3383 ();
 sg13g2_decap_8 FILLER_48_3416 ();
 sg13g2_decap_8 FILLER_48_3423 ();
 sg13g2_decap_8 FILLER_48_3430 ();
 sg13g2_decap_8 FILLER_48_3437 ();
 sg13g2_decap_8 FILLER_48_3444 ();
 sg13g2_decap_8 FILLER_48_3451 ();
 sg13g2_decap_8 FILLER_48_3458 ();
 sg13g2_decap_8 FILLER_48_3493 ();
 sg13g2_decap_8 FILLER_48_3500 ();
 sg13g2_decap_8 FILLER_48_3507 ();
 sg13g2_decap_8 FILLER_48_3514 ();
 sg13g2_decap_8 FILLER_48_3521 ();
 sg13g2_fill_1 FILLER_48_3549 ();
 sg13g2_decap_8 FILLER_48_3554 ();
 sg13g2_decap_8 FILLER_48_3561 ();
 sg13g2_decap_8 FILLER_48_3568 ();
 sg13g2_fill_2 FILLER_48_3575 ();
 sg13g2_fill_1 FILLER_48_3577 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_50 ();
 sg13g2_decap_8 FILLER_49_57 ();
 sg13g2_decap_8 FILLER_49_64 ();
 sg13g2_decap_4 FILLER_49_71 ();
 sg13g2_decap_4 FILLER_49_121 ();
 sg13g2_fill_1 FILLER_49_125 ();
 sg13g2_decap_4 FILLER_49_163 ();
 sg13g2_decap_8 FILLER_49_176 ();
 sg13g2_decap_8 FILLER_49_183 ();
 sg13g2_decap_4 FILLER_49_190 ();
 sg13g2_fill_1 FILLER_49_194 ();
 sg13g2_decap_8 FILLER_49_198 ();
 sg13g2_fill_1 FILLER_49_205 ();
 sg13g2_fill_2 FILLER_49_221 ();
 sg13g2_fill_1 FILLER_49_223 ();
 sg13g2_fill_1 FILLER_49_233 ();
 sg13g2_fill_1 FILLER_49_244 ();
 sg13g2_decap_4 FILLER_49_300 ();
 sg13g2_fill_2 FILLER_49_304 ();
 sg13g2_decap_8 FILLER_49_334 ();
 sg13g2_decap_8 FILLER_49_341 ();
 sg13g2_decap_8 FILLER_49_348 ();
 sg13g2_decap_8 FILLER_49_422 ();
 sg13g2_decap_8 FILLER_49_429 ();
 sg13g2_decap_4 FILLER_49_436 ();
 sg13g2_fill_2 FILLER_49_440 ();
 sg13g2_decap_8 FILLER_49_484 ();
 sg13g2_decap_8 FILLER_49_491 ();
 sg13g2_decap_8 FILLER_49_498 ();
 sg13g2_decap_8 FILLER_49_505 ();
 sg13g2_decap_8 FILLER_49_512 ();
 sg13g2_decap_8 FILLER_49_519 ();
 sg13g2_decap_8 FILLER_49_526 ();
 sg13g2_decap_8 FILLER_49_533 ();
 sg13g2_fill_1 FILLER_49_540 ();
 sg13g2_fill_1 FILLER_49_576 ();
 sg13g2_decap_8 FILLER_49_596 ();
 sg13g2_decap_8 FILLER_49_603 ();
 sg13g2_decap_8 FILLER_49_610 ();
 sg13g2_decap_8 FILLER_49_617 ();
 sg13g2_decap_4 FILLER_49_624 ();
 sg13g2_fill_1 FILLER_49_628 ();
 sg13g2_decap_4 FILLER_49_643 ();
 sg13g2_fill_2 FILLER_49_647 ();
 sg13g2_decap_8 FILLER_49_654 ();
 sg13g2_decap_8 FILLER_49_661 ();
 sg13g2_decap_8 FILLER_49_668 ();
 sg13g2_decap_8 FILLER_49_675 ();
 sg13g2_decap_8 FILLER_49_715 ();
 sg13g2_fill_1 FILLER_49_722 ();
 sg13g2_decap_8 FILLER_49_745 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_decap_8 FILLER_49_759 ();
 sg13g2_decap_8 FILLER_49_766 ();
 sg13g2_decap_4 FILLER_49_773 ();
 sg13g2_decap_8 FILLER_49_785 ();
 sg13g2_fill_1 FILLER_49_792 ();
 sg13g2_fill_1 FILLER_49_797 ();
 sg13g2_fill_2 FILLER_49_835 ();
 sg13g2_fill_1 FILLER_49_837 ();
 sg13g2_fill_2 FILLER_49_847 ();
 sg13g2_fill_1 FILLER_49_849 ();
 sg13g2_decap_8 FILLER_49_858 ();
 sg13g2_fill_2 FILLER_49_865 ();
 sg13g2_decap_8 FILLER_49_871 ();
 sg13g2_decap_4 FILLER_49_878 ();
 sg13g2_fill_2 FILLER_49_886 ();
 sg13g2_fill_1 FILLER_49_888 ();
 sg13g2_fill_2 FILLER_49_893 ();
 sg13g2_fill_2 FILLER_49_909 ();
 sg13g2_fill_1 FILLER_49_937 ();
 sg13g2_decap_8 FILLER_49_1006 ();
 sg13g2_decap_8 FILLER_49_1013 ();
 sg13g2_fill_2 FILLER_49_1020 ();
 sg13g2_fill_1 FILLER_49_1033 ();
 sg13g2_decap_8 FILLER_49_1041 ();
 sg13g2_decap_8 FILLER_49_1048 ();
 sg13g2_fill_2 FILLER_49_1088 ();
 sg13g2_decap_8 FILLER_49_1100 ();
 sg13g2_decap_8 FILLER_49_1107 ();
 sg13g2_decap_8 FILLER_49_1114 ();
 sg13g2_decap_8 FILLER_49_1121 ();
 sg13g2_decap_8 FILLER_49_1137 ();
 sg13g2_decap_4 FILLER_49_1144 ();
 sg13g2_fill_2 FILLER_49_1148 ();
 sg13g2_decap_8 FILLER_49_1192 ();
 sg13g2_decap_8 FILLER_49_1199 ();
 sg13g2_decap_4 FILLER_49_1206 ();
 sg13g2_fill_1 FILLER_49_1210 ();
 sg13g2_decap_8 FILLER_49_1220 ();
 sg13g2_decap_8 FILLER_49_1227 ();
 sg13g2_fill_2 FILLER_49_1234 ();
 sg13g2_decap_4 FILLER_49_1280 ();
 sg13g2_decap_8 FILLER_49_1341 ();
 sg13g2_decap_4 FILLER_49_1348 ();
 sg13g2_fill_2 FILLER_49_1362 ();
 sg13g2_fill_1 FILLER_49_1364 ();
 sg13g2_fill_1 FILLER_49_1374 ();
 sg13g2_decap_8 FILLER_49_1388 ();
 sg13g2_decap_8 FILLER_49_1395 ();
 sg13g2_fill_1 FILLER_49_1402 ();
 sg13g2_fill_2 FILLER_49_1408 ();
 sg13g2_decap_8 FILLER_49_1437 ();
 sg13g2_decap_8 FILLER_49_1444 ();
 sg13g2_decap_8 FILLER_49_1451 ();
 sg13g2_decap_8 FILLER_49_1458 ();
 sg13g2_decap_8 FILLER_49_1465 ();
 sg13g2_fill_1 FILLER_49_1472 ();
 sg13g2_fill_2 FILLER_49_1489 ();
 sg13g2_decap_8 FILLER_49_1517 ();
 sg13g2_decap_8 FILLER_49_1524 ();
 sg13g2_decap_8 FILLER_49_1531 ();
 sg13g2_fill_2 FILLER_49_1538 ();
 sg13g2_fill_1 FILLER_49_1576 ();
 sg13g2_fill_1 FILLER_49_1588 ();
 sg13g2_decap_8 FILLER_49_1593 ();
 sg13g2_decap_8 FILLER_49_1600 ();
 sg13g2_fill_1 FILLER_49_1607 ();
 sg13g2_decap_8 FILLER_49_1616 ();
 sg13g2_fill_2 FILLER_49_1623 ();
 sg13g2_decap_8 FILLER_49_1654 ();
 sg13g2_decap_8 FILLER_49_1661 ();
 sg13g2_decap_8 FILLER_49_1668 ();
 sg13g2_decap_4 FILLER_49_1675 ();
 sg13g2_fill_2 FILLER_49_1679 ();
 sg13g2_decap_8 FILLER_49_1696 ();
 sg13g2_decap_8 FILLER_49_1703 ();
 sg13g2_decap_8 FILLER_49_1710 ();
 sg13g2_fill_2 FILLER_49_1717 ();
 sg13g2_decap_8 FILLER_49_1738 ();
 sg13g2_decap_8 FILLER_49_1745 ();
 sg13g2_decap_8 FILLER_49_1752 ();
 sg13g2_fill_2 FILLER_49_1759 ();
 sg13g2_fill_1 FILLER_49_1761 ();
 sg13g2_fill_2 FILLER_49_1783 ();
 sg13g2_decap_8 FILLER_49_1804 ();
 sg13g2_decap_8 FILLER_49_1811 ();
 sg13g2_decap_8 FILLER_49_1818 ();
 sg13g2_decap_8 FILLER_49_1825 ();
 sg13g2_decap_8 FILLER_49_1832 ();
 sg13g2_fill_2 FILLER_49_1839 ();
 sg13g2_fill_2 FILLER_49_1870 ();
 sg13g2_fill_2 FILLER_49_1890 ();
 sg13g2_decap_8 FILLER_49_1901 ();
 sg13g2_decap_8 FILLER_49_1908 ();
 sg13g2_decap_8 FILLER_49_1915 ();
 sg13g2_decap_8 FILLER_49_1922 ();
 sg13g2_decap_8 FILLER_49_1929 ();
 sg13g2_decap_4 FILLER_49_1936 ();
 sg13g2_fill_2 FILLER_49_1940 ();
 sg13g2_fill_2 FILLER_49_1951 ();
 sg13g2_fill_1 FILLER_49_1953 ();
 sg13g2_decap_8 FILLER_49_1968 ();
 sg13g2_decap_8 FILLER_49_1975 ();
 sg13g2_decap_8 FILLER_49_1982 ();
 sg13g2_decap_4 FILLER_49_1989 ();
 sg13g2_decap_8 FILLER_49_1997 ();
 sg13g2_decap_4 FILLER_49_2004 ();
 sg13g2_fill_1 FILLER_49_2008 ();
 sg13g2_decap_8 FILLER_49_2017 ();
 sg13g2_fill_2 FILLER_49_2024 ();
 sg13g2_fill_1 FILLER_49_2058 ();
 sg13g2_decap_8 FILLER_49_2069 ();
 sg13g2_decap_8 FILLER_49_2076 ();
 sg13g2_decap_8 FILLER_49_2128 ();
 sg13g2_decap_8 FILLER_49_2135 ();
 sg13g2_decap_4 FILLER_49_2142 ();
 sg13g2_fill_2 FILLER_49_2183 ();
 sg13g2_decap_8 FILLER_49_2199 ();
 sg13g2_decap_8 FILLER_49_2206 ();
 sg13g2_decap_4 FILLER_49_2213 ();
 sg13g2_fill_1 FILLER_49_2244 ();
 sg13g2_fill_2 FILLER_49_2296 ();
 sg13g2_fill_1 FILLER_49_2298 ();
 sg13g2_fill_2 FILLER_49_2304 ();
 sg13g2_fill_1 FILLER_49_2306 ();
 sg13g2_decap_8 FILLER_49_2335 ();
 sg13g2_decap_8 FILLER_49_2342 ();
 sg13g2_fill_2 FILLER_49_2349 ();
 sg13g2_fill_1 FILLER_49_2351 ();
 sg13g2_decap_4 FILLER_49_2389 ();
 sg13g2_decap_4 FILLER_49_2425 ();
 sg13g2_fill_1 FILLER_49_2429 ();
 sg13g2_decap_8 FILLER_49_2440 ();
 sg13g2_decap_8 FILLER_49_2447 ();
 sg13g2_decap_8 FILLER_49_2454 ();
 sg13g2_fill_1 FILLER_49_2461 ();
 sg13g2_decap_8 FILLER_49_2528 ();
 sg13g2_decap_8 FILLER_49_2535 ();
 sg13g2_decap_8 FILLER_49_2542 ();
 sg13g2_fill_2 FILLER_49_2549 ();
 sg13g2_decap_4 FILLER_49_2555 ();
 sg13g2_decap_8 FILLER_49_2563 ();
 sg13g2_decap_8 FILLER_49_2570 ();
 sg13g2_decap_4 FILLER_49_2577 ();
 sg13g2_fill_1 FILLER_49_2581 ();
 sg13g2_fill_2 FILLER_49_2590 ();
 sg13g2_fill_1 FILLER_49_2592 ();
 sg13g2_decap_8 FILLER_49_2598 ();
 sg13g2_decap_8 FILLER_49_2605 ();
 sg13g2_decap_4 FILLER_49_2612 ();
 sg13g2_fill_1 FILLER_49_2616 ();
 sg13g2_decap_4 FILLER_49_2670 ();
 sg13g2_fill_2 FILLER_49_2711 ();
 sg13g2_fill_1 FILLER_49_2713 ();
 sg13g2_decap_4 FILLER_49_2741 ();
 sg13g2_decap_8 FILLER_49_2758 ();
 sg13g2_decap_8 FILLER_49_2765 ();
 sg13g2_decap_4 FILLER_49_2772 ();
 sg13g2_fill_1 FILLER_49_2776 ();
 sg13g2_decap_8 FILLER_49_2811 ();
 sg13g2_decap_4 FILLER_49_2818 ();
 sg13g2_fill_1 FILLER_49_2822 ();
 sg13g2_decap_8 FILLER_49_2842 ();
 sg13g2_decap_8 FILLER_49_2899 ();
 sg13g2_decap_4 FILLER_49_2906 ();
 sg13g2_fill_2 FILLER_49_2910 ();
 sg13g2_fill_1 FILLER_49_2939 ();
 sg13g2_decap_8 FILLER_49_2953 ();
 sg13g2_decap_4 FILLER_49_2960 ();
 sg13g2_fill_1 FILLER_49_2964 ();
 sg13g2_decap_8 FILLER_49_3015 ();
 sg13g2_decap_8 FILLER_49_3022 ();
 sg13g2_fill_2 FILLER_49_3066 ();
 sg13g2_fill_1 FILLER_49_3158 ();
 sg13g2_decap_4 FILLER_49_3168 ();
 sg13g2_fill_2 FILLER_49_3172 ();
 sg13g2_fill_1 FILLER_49_3201 ();
 sg13g2_decap_8 FILLER_49_3264 ();
 sg13g2_decap_4 FILLER_49_3271 ();
 sg13g2_fill_1 FILLER_49_3275 ();
 sg13g2_decap_8 FILLER_49_3281 ();
 sg13g2_decap_4 FILLER_49_3288 ();
 sg13g2_fill_2 FILLER_49_3306 ();
 sg13g2_fill_1 FILLER_49_3308 ();
 sg13g2_decap_8 FILLER_49_3330 ();
 sg13g2_fill_1 FILLER_49_3347 ();
 sg13g2_decap_8 FILLER_49_3357 ();
 sg13g2_decap_8 FILLER_49_3364 ();
 sg13g2_decap_8 FILLER_49_3371 ();
 sg13g2_fill_2 FILLER_49_3378 ();
 sg13g2_decap_8 FILLER_49_3389 ();
 sg13g2_decap_4 FILLER_49_3396 ();
 sg13g2_fill_2 FILLER_49_3400 ();
 sg13g2_decap_8 FILLER_49_3415 ();
 sg13g2_fill_1 FILLER_49_3422 ();
 sg13g2_decap_8 FILLER_49_3436 ();
 sg13g2_fill_1 FILLER_49_3443 ();
 sg13g2_decap_4 FILLER_49_3475 ();
 sg13g2_decap_4 FILLER_49_3506 ();
 sg13g2_fill_1 FILLER_49_3510 ();
 sg13g2_decap_8 FILLER_49_3521 ();
 sg13g2_decap_8 FILLER_49_3565 ();
 sg13g2_decap_4 FILLER_49_3572 ();
 sg13g2_fill_2 FILLER_49_3576 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_53 ();
 sg13g2_decap_8 FILLER_50_60 ();
 sg13g2_fill_2 FILLER_50_67 ();
 sg13g2_fill_1 FILLER_50_69 ();
 sg13g2_fill_2 FILLER_50_74 ();
 sg13g2_decap_4 FILLER_50_114 ();
 sg13g2_decap_8 FILLER_50_123 ();
 sg13g2_fill_1 FILLER_50_130 ();
 sg13g2_fill_1 FILLER_50_135 ();
 sg13g2_decap_8 FILLER_50_186 ();
 sg13g2_decap_8 FILLER_50_193 ();
 sg13g2_decap_8 FILLER_50_200 ();
 sg13g2_decap_4 FILLER_50_207 ();
 sg13g2_fill_2 FILLER_50_211 ();
 sg13g2_fill_2 FILLER_50_249 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_decap_8 FILLER_50_265 ();
 sg13g2_decap_8 FILLER_50_281 ();
 sg13g2_decap_8 FILLER_50_288 ();
 sg13g2_decap_8 FILLER_50_295 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_fill_1 FILLER_50_304 ();
 sg13g2_decap_4 FILLER_50_336 ();
 sg13g2_fill_1 FILLER_50_353 ();
 sg13g2_decap_8 FILLER_50_367 ();
 sg13g2_decap_4 FILLER_50_374 ();
 sg13g2_decap_8 FILLER_50_383 ();
 sg13g2_decap_4 FILLER_50_390 ();
 sg13g2_fill_2 FILLER_50_394 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_50_409 ();
 sg13g2_decap_4 FILLER_50_416 ();
 sg13g2_fill_2 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_428 ();
 sg13g2_decap_4 FILLER_50_435 ();
 sg13g2_fill_2 FILLER_50_443 ();
 sg13g2_fill_1 FILLER_50_445 ();
 sg13g2_decap_8 FILLER_50_488 ();
 sg13g2_decap_8 FILLER_50_495 ();
 sg13g2_decap_8 FILLER_50_502 ();
 sg13g2_fill_1 FILLER_50_509 ();
 sg13g2_fill_2 FILLER_50_538 ();
 sg13g2_fill_1 FILLER_50_543 ();
 sg13g2_fill_1 FILLER_50_557 ();
 sg13g2_fill_1 FILLER_50_562 ();
 sg13g2_fill_1 FILLER_50_572 ();
 sg13g2_decap_4 FILLER_50_623 ();
 sg13g2_fill_2 FILLER_50_627 ();
 sg13g2_decap_8 FILLER_50_672 ();
 sg13g2_decap_8 FILLER_50_679 ();
 sg13g2_fill_2 FILLER_50_686 ();
 sg13g2_fill_1 FILLER_50_688 ();
 sg13g2_fill_1 FILLER_50_694 ();
 sg13g2_decap_8 FILLER_50_713 ();
 sg13g2_decap_8 FILLER_50_720 ();
 sg13g2_decap_8 FILLER_50_727 ();
 sg13g2_decap_8 FILLER_50_734 ();
 sg13g2_decap_8 FILLER_50_741 ();
 sg13g2_fill_2 FILLER_50_748 ();
 sg13g2_decap_8 FILLER_50_771 ();
 sg13g2_decap_4 FILLER_50_778 ();
 sg13g2_fill_2 FILLER_50_782 ();
 sg13g2_decap_8 FILLER_50_791 ();
 sg13g2_decap_8 FILLER_50_798 ();
 sg13g2_fill_1 FILLER_50_805 ();
 sg13g2_decap_8 FILLER_50_809 ();
 sg13g2_fill_1 FILLER_50_825 ();
 sg13g2_decap_4 FILLER_50_854 ();
 sg13g2_fill_2 FILLER_50_858 ();
 sg13g2_fill_2 FILLER_50_868 ();
 sg13g2_fill_1 FILLER_50_870 ();
 sg13g2_decap_8 FILLER_50_880 ();
 sg13g2_fill_2 FILLER_50_887 ();
 sg13g2_fill_2 FILLER_50_898 ();
 sg13g2_fill_1 FILLER_50_906 ();
 sg13g2_fill_2 FILLER_50_921 ();
 sg13g2_fill_2 FILLER_50_928 ();
 sg13g2_fill_1 FILLER_50_930 ();
 sg13g2_fill_1 FILLER_50_969 ();
 sg13g2_decap_4 FILLER_50_978 ();
 sg13g2_fill_2 FILLER_50_982 ();
 sg13g2_decap_8 FILLER_50_1006 ();
 sg13g2_decap_8 FILLER_50_1013 ();
 sg13g2_decap_8 FILLER_50_1020 ();
 sg13g2_fill_1 FILLER_50_1027 ();
 sg13g2_decap_8 FILLER_50_1037 ();
 sg13g2_decap_8 FILLER_50_1044 ();
 sg13g2_decap_8 FILLER_50_1051 ();
 sg13g2_decap_4 FILLER_50_1058 ();
 sg13g2_fill_1 FILLER_50_1062 ();
 sg13g2_fill_2 FILLER_50_1079 ();
 sg13g2_fill_1 FILLER_50_1086 ();
 sg13g2_decap_8 FILLER_50_1096 ();
 sg13g2_decap_8 FILLER_50_1103 ();
 sg13g2_decap_4 FILLER_50_1110 ();
 sg13g2_fill_2 FILLER_50_1119 ();
 sg13g2_fill_1 FILLER_50_1121 ();
 sg13g2_fill_1 FILLER_50_1131 ();
 sg13g2_decap_8 FILLER_50_1143 ();
 sg13g2_decap_8 FILLER_50_1150 ();
 sg13g2_decap_4 FILLER_50_1170 ();
 sg13g2_decap_8 FILLER_50_1188 ();
 sg13g2_decap_4 FILLER_50_1195 ();
 sg13g2_fill_2 FILLER_50_1199 ();
 sg13g2_fill_2 FILLER_50_1218 ();
 sg13g2_fill_2 FILLER_50_1229 ();
 sg13g2_fill_2 FILLER_50_1235 ();
 sg13g2_fill_1 FILLER_50_1237 ();
 sg13g2_decap_8 FILLER_50_1244 ();
 sg13g2_decap_8 FILLER_50_1251 ();
 sg13g2_decap_8 FILLER_50_1258 ();
 sg13g2_fill_2 FILLER_50_1265 ();
 sg13g2_decap_8 FILLER_50_1283 ();
 sg13g2_decap_8 FILLER_50_1290 ();
 sg13g2_fill_2 FILLER_50_1297 ();
 sg13g2_fill_1 FILLER_50_1308 ();
 sg13g2_decap_8 FILLER_50_1336 ();
 sg13g2_decap_4 FILLER_50_1343 ();
 sg13g2_decap_8 FILLER_50_1379 ();
 sg13g2_decap_8 FILLER_50_1386 ();
 sg13g2_fill_1 FILLER_50_1393 ();
 sg13g2_decap_4 FILLER_50_1427 ();
 sg13g2_fill_2 FILLER_50_1431 ();
 sg13g2_decap_8 FILLER_50_1442 ();
 sg13g2_decap_8 FILLER_50_1449 ();
 sg13g2_decap_8 FILLER_50_1456 ();
 sg13g2_fill_2 FILLER_50_1463 ();
 sg13g2_fill_2 FILLER_50_1485 ();
 sg13g2_fill_1 FILLER_50_1487 ();
 sg13g2_fill_2 FILLER_50_1492 ();
 sg13g2_decap_8 FILLER_50_1503 ();
 sg13g2_decap_8 FILLER_50_1510 ();
 sg13g2_decap_8 FILLER_50_1517 ();
 sg13g2_decap_8 FILLER_50_1524 ();
 sg13g2_decap_8 FILLER_50_1531 ();
 sg13g2_decap_8 FILLER_50_1538 ();
 sg13g2_decap_8 FILLER_50_1545 ();
 sg13g2_decap_8 FILLER_50_1552 ();
 sg13g2_fill_2 FILLER_50_1559 ();
 sg13g2_fill_1 FILLER_50_1561 ();
 sg13g2_decap_8 FILLER_50_1579 ();
 sg13g2_decap_8 FILLER_50_1586 ();
 sg13g2_decap_8 FILLER_50_1593 ();
 sg13g2_decap_4 FILLER_50_1600 ();
 sg13g2_decap_8 FILLER_50_1628 ();
 sg13g2_decap_8 FILLER_50_1635 ();
 sg13g2_decap_8 FILLER_50_1642 ();
 sg13g2_decap_8 FILLER_50_1649 ();
 sg13g2_decap_8 FILLER_50_1656 ();
 sg13g2_fill_1 FILLER_50_1663 ();
 sg13g2_decap_8 FILLER_50_1668 ();
 sg13g2_decap_4 FILLER_50_1675 ();
 sg13g2_decap_8 FILLER_50_1684 ();
 sg13g2_decap_8 FILLER_50_1691 ();
 sg13g2_decap_8 FILLER_50_1698 ();
 sg13g2_decap_4 FILLER_50_1705 ();
 sg13g2_fill_2 FILLER_50_1709 ();
 sg13g2_decap_8 FILLER_50_1715 ();
 sg13g2_decap_8 FILLER_50_1722 ();
 sg13g2_fill_1 FILLER_50_1729 ();
 sg13g2_fill_2 FILLER_50_1735 ();
 sg13g2_decap_4 FILLER_50_1745 ();
 sg13g2_decap_8 FILLER_50_1755 ();
 sg13g2_decap_8 FILLER_50_1762 ();
 sg13g2_decap_8 FILLER_50_1799 ();
 sg13g2_decap_4 FILLER_50_1806 ();
 sg13g2_fill_2 FILLER_50_1823 ();
 sg13g2_decap_8 FILLER_50_1838 ();
 sg13g2_decap_4 FILLER_50_1845 ();
 sg13g2_fill_1 FILLER_50_1849 ();
 sg13g2_decap_8 FILLER_50_1867 ();
 sg13g2_decap_8 FILLER_50_1874 ();
 sg13g2_fill_2 FILLER_50_1881 ();
 sg13g2_fill_1 FILLER_50_1883 ();
 sg13g2_fill_2 FILLER_50_1889 ();
 sg13g2_fill_1 FILLER_50_1891 ();
 sg13g2_fill_2 FILLER_50_1897 ();
 sg13g2_fill_1 FILLER_50_1899 ();
 sg13g2_decap_4 FILLER_50_1914 ();
 sg13g2_fill_1 FILLER_50_1922 ();
 sg13g2_decap_8 FILLER_50_1968 ();
 sg13g2_fill_2 FILLER_50_1988 ();
 sg13g2_fill_1 FILLER_50_1990 ();
 sg13g2_fill_2 FILLER_50_1996 ();
 sg13g2_fill_1 FILLER_50_2002 ();
 sg13g2_fill_2 FILLER_50_2006 ();
 sg13g2_decap_8 FILLER_50_2017 ();
 sg13g2_fill_2 FILLER_50_2024 ();
 sg13g2_decap_4 FILLER_50_2052 ();
 sg13g2_fill_2 FILLER_50_2069 ();
 sg13g2_decap_4 FILLER_50_2075 ();
 sg13g2_fill_1 FILLER_50_2079 ();
 sg13g2_decap_4 FILLER_50_2089 ();
 sg13g2_decap_4 FILLER_50_2129 ();
 sg13g2_fill_1 FILLER_50_2143 ();
 sg13g2_fill_2 FILLER_50_2162 ();
 sg13g2_decap_8 FILLER_50_2191 ();
 sg13g2_decap_8 FILLER_50_2198 ();
 sg13g2_decap_8 FILLER_50_2205 ();
 sg13g2_decap_4 FILLER_50_2212 ();
 sg13g2_decap_8 FILLER_50_2225 ();
 sg13g2_decap_8 FILLER_50_2232 ();
 sg13g2_decap_8 FILLER_50_2239 ();
 sg13g2_decap_8 FILLER_50_2246 ();
 sg13g2_decap_4 FILLER_50_2253 ();
 sg13g2_fill_2 FILLER_50_2289 ();
 sg13g2_fill_1 FILLER_50_2291 ();
 sg13g2_decap_8 FILLER_50_2348 ();
 sg13g2_fill_1 FILLER_50_2355 ();
 sg13g2_fill_1 FILLER_50_2361 ();
 sg13g2_decap_8 FILLER_50_2392 ();
 sg13g2_decap_8 FILLER_50_2399 ();
 sg13g2_fill_1 FILLER_50_2406 ();
 sg13g2_decap_8 FILLER_50_2412 ();
 sg13g2_decap_8 FILLER_50_2465 ();
 sg13g2_fill_2 FILLER_50_2472 ();
 sg13g2_decap_8 FILLER_50_2529 ();
 sg13g2_decap_8 FILLER_50_2536 ();
 sg13g2_fill_2 FILLER_50_2543 ();
 sg13g2_fill_1 FILLER_50_2545 ();
 sg13g2_decap_8 FILLER_50_2594 ();
 sg13g2_decap_8 FILLER_50_2601 ();
 sg13g2_decap_8 FILLER_50_2608 ();
 sg13g2_decap_8 FILLER_50_2615 ();
 sg13g2_decap_4 FILLER_50_2622 ();
 sg13g2_fill_2 FILLER_50_2626 ();
 sg13g2_decap_8 FILLER_50_2642 ();
 sg13g2_decap_8 FILLER_50_2662 ();
 sg13g2_decap_8 FILLER_50_2669 ();
 sg13g2_fill_2 FILLER_50_2676 ();
 sg13g2_fill_1 FILLER_50_2678 ();
 sg13g2_decap_4 FILLER_50_2723 ();
 sg13g2_decap_8 FILLER_50_2736 ();
 sg13g2_decap_8 FILLER_50_2743 ();
 sg13g2_fill_2 FILLER_50_2750 ();
 sg13g2_decap_4 FILLER_50_2762 ();
 sg13g2_fill_2 FILLER_50_2766 ();
 sg13g2_decap_4 FILLER_50_2782 ();
 sg13g2_decap_8 FILLER_50_2804 ();
 sg13g2_decap_8 FILLER_50_2811 ();
 sg13g2_fill_1 FILLER_50_2818 ();
 sg13g2_decap_4 FILLER_50_2850 ();
 sg13g2_fill_1 FILLER_50_2854 ();
 sg13g2_decap_8 FILLER_50_2891 ();
 sg13g2_decap_4 FILLER_50_2898 ();
 sg13g2_fill_1 FILLER_50_2902 ();
 sg13g2_fill_2 FILLER_50_2930 ();
 sg13g2_decap_8 FILLER_50_2953 ();
 sg13g2_decap_8 FILLER_50_2960 ();
 sg13g2_decap_8 FILLER_50_2967 ();
 sg13g2_decap_8 FILLER_50_3011 ();
 sg13g2_decap_8 FILLER_50_3018 ();
 sg13g2_decap_8 FILLER_50_3025 ();
 sg13g2_decap_4 FILLER_50_3032 ();
 sg13g2_fill_2 FILLER_50_3036 ();
 sg13g2_fill_2 FILLER_50_3052 ();
 sg13g2_fill_1 FILLER_50_3054 ();
 sg13g2_decap_8 FILLER_50_3068 ();
 sg13g2_decap_4 FILLER_50_3075 ();
 sg13g2_fill_1 FILLER_50_3079 ();
 sg13g2_decap_8 FILLER_50_3115 ();
 sg13g2_fill_2 FILLER_50_3122 ();
 sg13g2_fill_2 FILLER_50_3128 ();
 sg13g2_fill_1 FILLER_50_3140 ();
 sg13g2_decap_8 FILLER_50_3172 ();
 sg13g2_decap_4 FILLER_50_3179 ();
 sg13g2_fill_2 FILLER_50_3183 ();
 sg13g2_decap_4 FILLER_50_3189 ();
 sg13g2_fill_2 FILLER_50_3193 ();
 sg13g2_decap_8 FILLER_50_3204 ();
 sg13g2_decap_8 FILLER_50_3211 ();
 sg13g2_fill_2 FILLER_50_3218 ();
 sg13g2_decap_4 FILLER_50_3224 ();
 sg13g2_decap_8 FILLER_50_3242 ();
 sg13g2_fill_1 FILLER_50_3249 ();
 sg13g2_decap_8 FILLER_50_3263 ();
 sg13g2_decap_4 FILLER_50_3270 ();
 sg13g2_fill_2 FILLER_50_3274 ();
 sg13g2_decap_8 FILLER_50_3325 ();
 sg13g2_decap_8 FILLER_50_3332 ();
 sg13g2_decap_8 FILLER_50_3339 ();
 sg13g2_fill_1 FILLER_50_3346 ();
 sg13g2_decap_4 FILLER_50_3351 ();
 sg13g2_decap_8 FILLER_50_3419 ();
 sg13g2_decap_8 FILLER_50_3426 ();
 sg13g2_fill_2 FILLER_50_3433 ();
 sg13g2_fill_2 FILLER_50_3462 ();
 sg13g2_fill_1 FILLER_50_3464 ();
 sg13g2_decap_8 FILLER_50_3502 ();
 sg13g2_fill_1 FILLER_50_3509 ();
 sg13g2_decap_8 FILLER_50_3564 ();
 sg13g2_decap_8 FILLER_50_3571 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_50 ();
 sg13g2_fill_2 FILLER_51_63 ();
 sg13g2_decap_4 FILLER_51_92 ();
 sg13g2_decap_4 FILLER_51_111 ();
 sg13g2_decap_8 FILLER_51_129 ();
 sg13g2_fill_1 FILLER_51_164 ();
 sg13g2_decap_8 FILLER_51_192 ();
 sg13g2_fill_2 FILLER_51_199 ();
 sg13g2_fill_1 FILLER_51_205 ();
 sg13g2_fill_1 FILLER_51_215 ();
 sg13g2_fill_2 FILLER_51_221 ();
 sg13g2_fill_1 FILLER_51_223 ();
 sg13g2_decap_8 FILLER_51_229 ();
 sg13g2_decap_8 FILLER_51_236 ();
 sg13g2_decap_8 FILLER_51_243 ();
 sg13g2_decap_4 FILLER_51_250 ();
 sg13g2_fill_2 FILLER_51_254 ();
 sg13g2_decap_8 FILLER_51_283 ();
 sg13g2_decap_4 FILLER_51_290 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_331 ();
 sg13g2_decap_8 FILLER_51_338 ();
 sg13g2_decap_8 FILLER_51_345 ();
 sg13g2_decap_8 FILLER_51_352 ();
 sg13g2_fill_1 FILLER_51_359 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_decap_8 FILLER_51_406 ();
 sg13g2_decap_8 FILLER_51_413 ();
 sg13g2_decap_8 FILLER_51_433 ();
 sg13g2_fill_2 FILLER_51_440 ();
 sg13g2_fill_2 FILLER_51_475 ();
 sg13g2_fill_1 FILLER_51_477 ();
 sg13g2_decap_8 FILLER_51_506 ();
 sg13g2_decap_4 FILLER_51_549 ();
 sg13g2_fill_2 FILLER_51_553 ();
 sg13g2_decap_4 FILLER_51_573 ();
 sg13g2_fill_1 FILLER_51_577 ();
 sg13g2_fill_2 FILLER_51_586 ();
 sg13g2_fill_1 FILLER_51_588 ();
 sg13g2_decap_8 FILLER_51_617 ();
 sg13g2_decap_4 FILLER_51_624 ();
 sg13g2_fill_1 FILLER_51_628 ();
 sg13g2_decap_8 FILLER_51_696 ();
 sg13g2_fill_1 FILLER_51_703 ();
 sg13g2_fill_2 FILLER_51_731 ();
 sg13g2_fill_1 FILLER_51_733 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_decap_4 FILLER_51_786 ();
 sg13g2_fill_2 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_813 ();
 sg13g2_fill_2 FILLER_51_820 ();
 sg13g2_decap_4 FILLER_51_826 ();
 sg13g2_decap_8 FILLER_51_844 ();
 sg13g2_fill_2 FILLER_51_851 ();
 sg13g2_decap_4 FILLER_51_862 ();
 sg13g2_fill_1 FILLER_51_866 ();
 sg13g2_decap_8 FILLER_51_900 ();
 sg13g2_fill_1 FILLER_51_907 ();
 sg13g2_fill_2 FILLER_51_936 ();
 sg13g2_fill_1 FILLER_51_938 ();
 sg13g2_decap_8 FILLER_51_967 ();
 sg13g2_decap_8 FILLER_51_974 ();
 sg13g2_decap_8 FILLER_51_981 ();
 sg13g2_decap_8 FILLER_51_988 ();
 sg13g2_decap_8 FILLER_51_995 ();
 sg13g2_decap_4 FILLER_51_1002 ();
 sg13g2_fill_1 FILLER_51_1019 ();
 sg13g2_fill_1 FILLER_51_1032 ();
 sg13g2_fill_1 FILLER_51_1079 ();
 sg13g2_fill_1 FILLER_51_1095 ();
 sg13g2_fill_2 FILLER_51_1105 ();
 sg13g2_fill_1 FILLER_51_1137 ();
 sg13g2_decap_4 FILLER_51_1160 ();
 sg13g2_fill_2 FILLER_51_1182 ();
 sg13g2_decap_4 FILLER_51_1197 ();
 sg13g2_fill_2 FILLER_51_1201 ();
 sg13g2_fill_1 FILLER_51_1207 ();
 sg13g2_decap_8 FILLER_51_1222 ();
 sg13g2_decap_8 FILLER_51_1229 ();
 sg13g2_decap_8 FILLER_51_1236 ();
 sg13g2_decap_8 FILLER_51_1243 ();
 sg13g2_fill_2 FILLER_51_1250 ();
 sg13g2_decap_8 FILLER_51_1293 ();
 sg13g2_decap_4 FILLER_51_1300 ();
 sg13g2_decap_4 FILLER_51_1344 ();
 sg13g2_fill_2 FILLER_51_1348 ();
 sg13g2_decap_8 FILLER_51_1359 ();
 sg13g2_decap_4 FILLER_51_1366 ();
 sg13g2_fill_2 FILLER_51_1375 ();
 sg13g2_decap_8 FILLER_51_1386 ();
 sg13g2_fill_2 FILLER_51_1402 ();
 sg13g2_fill_1 FILLER_51_1404 ();
 sg13g2_fill_2 FILLER_51_1417 ();
 sg13g2_decap_8 FILLER_51_1431 ();
 sg13g2_decap_8 FILLER_51_1438 ();
 sg13g2_decap_8 FILLER_51_1445 ();
 sg13g2_decap_8 FILLER_51_1452 ();
 sg13g2_fill_1 FILLER_51_1459 ();
 sg13g2_fill_2 FILLER_51_1468 ();
 sg13g2_fill_1 FILLER_51_1470 ();
 sg13g2_fill_1 FILLER_51_1498 ();
 sg13g2_decap_8 FILLER_51_1512 ();
 sg13g2_decap_8 FILLER_51_1519 ();
 sg13g2_decap_8 FILLER_51_1526 ();
 sg13g2_fill_2 FILLER_51_1533 ();
 sg13g2_fill_1 FILLER_51_1535 ();
 sg13g2_decap_8 FILLER_51_1576 ();
 sg13g2_decap_8 FILLER_51_1583 ();
 sg13g2_decap_8 FILLER_51_1590 ();
 sg13g2_fill_1 FILLER_51_1618 ();
 sg13g2_fill_2 FILLER_51_1624 ();
 sg13g2_fill_1 FILLER_51_1626 ();
 sg13g2_decap_8 FILLER_51_1636 ();
 sg13g2_fill_2 FILLER_51_1643 ();
 sg13g2_fill_1 FILLER_51_1645 ();
 sg13g2_fill_2 FILLER_51_1691 ();
 sg13g2_decap_4 FILLER_51_1734 ();
 sg13g2_fill_2 FILLER_51_1738 ();
 sg13g2_decap_8 FILLER_51_1749 ();
 sg13g2_decap_8 FILLER_51_1756 ();
 sg13g2_fill_2 FILLER_51_1763 ();
 sg13g2_decap_8 FILLER_51_1770 ();
 sg13g2_decap_4 FILLER_51_1777 ();
 sg13g2_fill_1 FILLER_51_1781 ();
 sg13g2_fill_1 FILLER_51_1822 ();
 sg13g2_decap_4 FILLER_51_1835 ();
 sg13g2_fill_2 FILLER_51_1848 ();
 sg13g2_decap_8 FILLER_51_1868 ();
 sg13g2_decap_8 FILLER_51_1875 ();
 sg13g2_decap_4 FILLER_51_1882 ();
 sg13g2_fill_2 FILLER_51_1886 ();
 sg13g2_fill_2 FILLER_51_1933 ();
 sg13g2_fill_1 FILLER_51_1935 ();
 sg13g2_fill_2 FILLER_51_1963 ();
 sg13g2_fill_2 FILLER_51_1978 ();
 sg13g2_decap_4 FILLER_51_2011 ();
 sg13g2_decap_4 FILLER_51_2028 ();
 sg13g2_fill_2 FILLER_51_2081 ();
 sg13g2_fill_1 FILLER_51_2083 ();
 sg13g2_fill_2 FILLER_51_2094 ();
 sg13g2_fill_1 FILLER_51_2114 ();
 sg13g2_decap_8 FILLER_51_2127 ();
 sg13g2_decap_8 FILLER_51_2134 ();
 sg13g2_decap_8 FILLER_51_2141 ();
 sg13g2_decap_4 FILLER_51_2148 ();
 sg13g2_decap_4 FILLER_51_2165 ();
 sg13g2_decap_8 FILLER_51_2183 ();
 sg13g2_decap_8 FILLER_51_2190 ();
 sg13g2_decap_8 FILLER_51_2197 ();
 sg13g2_decap_8 FILLER_51_2204 ();
 sg13g2_decap_4 FILLER_51_2211 ();
 sg13g2_fill_2 FILLER_51_2215 ();
 sg13g2_decap_8 FILLER_51_2222 ();
 sg13g2_fill_1 FILLER_51_2229 ();
 sg13g2_decap_8 FILLER_51_2258 ();
 sg13g2_fill_1 FILLER_51_2265 ();
 sg13g2_decap_4 FILLER_51_2279 ();
 sg13g2_fill_2 FILLER_51_2283 ();
 sg13g2_decap_8 FILLER_51_2303 ();
 sg13g2_decap_8 FILLER_51_2323 ();
 sg13g2_decap_4 FILLER_51_2330 ();
 sg13g2_decap_8 FILLER_51_2343 ();
 sg13g2_decap_8 FILLER_51_2350 ();
 sg13g2_decap_8 FILLER_51_2357 ();
 sg13g2_fill_1 FILLER_51_2364 ();
 sg13g2_fill_1 FILLER_51_2370 ();
 sg13g2_decap_4 FILLER_51_2406 ();
 sg13g2_fill_1 FILLER_51_2410 ();
 sg13g2_decap_8 FILLER_51_2469 ();
 sg13g2_decap_4 FILLER_51_2476 ();
 sg13g2_fill_1 FILLER_51_2480 ();
 sg13g2_decap_4 FILLER_51_2529 ();
 sg13g2_fill_2 FILLER_51_2533 ();
 sg13g2_decap_4 FILLER_51_2576 ();
 sg13g2_decap_8 FILLER_51_2611 ();
 sg13g2_decap_8 FILLER_51_2618 ();
 sg13g2_decap_4 FILLER_51_2625 ();
 sg13g2_fill_2 FILLER_51_2629 ();
 sg13g2_decap_8 FILLER_51_2662 ();
 sg13g2_decap_4 FILLER_51_2679 ();
 sg13g2_fill_2 FILLER_51_2683 ();
 sg13g2_fill_1 FILLER_51_2708 ();
 sg13g2_decap_4 FILLER_51_2719 ();
 sg13g2_fill_1 FILLER_51_2723 ();
 sg13g2_fill_1 FILLER_51_2737 ();
 sg13g2_decap_8 FILLER_51_2801 ();
 sg13g2_decap_4 FILLER_51_2854 ();
 sg13g2_fill_2 FILLER_51_2858 ();
 sg13g2_fill_1 FILLER_51_2864 ();
 sg13g2_decap_8 FILLER_51_2891 ();
 sg13g2_decap_8 FILLER_51_2898 ();
 sg13g2_fill_1 FILLER_51_2905 ();
 sg13g2_decap_4 FILLER_51_2943 ();
 sg13g2_fill_2 FILLER_51_2947 ();
 sg13g2_fill_2 FILLER_51_2975 ();
 sg13g2_fill_1 FILLER_51_2977 ();
 sg13g2_decap_8 FILLER_51_3003 ();
 sg13g2_decap_8 FILLER_51_3010 ();
 sg13g2_decap_4 FILLER_51_3017 ();
 sg13g2_fill_1 FILLER_51_3048 ();
 sg13g2_decap_8 FILLER_51_3067 ();
 sg13g2_decap_8 FILLER_51_3074 ();
 sg13g2_decap_4 FILLER_51_3081 ();
 sg13g2_fill_2 FILLER_51_3085 ();
 sg13g2_fill_2 FILLER_51_3116 ();
 sg13g2_fill_1 FILLER_51_3118 ();
 sg13g2_decap_8 FILLER_51_3187 ();
 sg13g2_decap_8 FILLER_51_3194 ();
 sg13g2_decap_8 FILLER_51_3201 ();
 sg13g2_fill_2 FILLER_51_3208 ();
 sg13g2_decap_8 FILLER_51_3223 ();
 sg13g2_fill_2 FILLER_51_3230 ();
 sg13g2_decap_8 FILLER_51_3241 ();
 sg13g2_decap_8 FILLER_51_3248 ();
 sg13g2_decap_8 FILLER_51_3255 ();
 sg13g2_fill_1 FILLER_51_3299 ();
 sg13g2_fill_2 FILLER_51_3314 ();
 sg13g2_decap_8 FILLER_51_3338 ();
 sg13g2_decap_4 FILLER_51_3426 ();
 sg13g2_decap_4 FILLER_51_3466 ();
 sg13g2_decap_8 FILLER_51_3504 ();
 sg13g2_decap_4 FILLER_51_3572 ();
 sg13g2_fill_2 FILLER_51_3576 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_11 ();
 sg13g2_fill_2 FILLER_52_66 ();
 sg13g2_decap_4 FILLER_52_78 ();
 sg13g2_fill_2 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_125 ();
 sg13g2_decap_8 FILLER_52_132 ();
 sg13g2_decap_8 FILLER_52_139 ();
 sg13g2_decap_4 FILLER_52_146 ();
 sg13g2_decap_4 FILLER_52_181 ();
 sg13g2_fill_1 FILLER_52_185 ();
 sg13g2_decap_8 FILLER_52_228 ();
 sg13g2_decap_4 FILLER_52_235 ();
 sg13g2_decap_8 FILLER_52_342 ();
 sg13g2_decap_8 FILLER_52_349 ();
 sg13g2_decap_8 FILLER_52_356 ();
 sg13g2_fill_1 FILLER_52_390 ();
 sg13g2_decap_4 FILLER_52_404 ();
 sg13g2_fill_2 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_52_423 ();
 sg13g2_decap_4 FILLER_52_430 ();
 sg13g2_fill_1 FILLER_52_434 ();
 sg13g2_fill_2 FILLER_52_468 ();
 sg13g2_fill_1 FILLER_52_470 ();
 sg13g2_fill_2 FILLER_52_476 ();
 sg13g2_fill_1 FILLER_52_478 ();
 sg13g2_decap_8 FILLER_52_482 ();
 sg13g2_decap_8 FILLER_52_489 ();
 sg13g2_decap_8 FILLER_52_496 ();
 sg13g2_decap_8 FILLER_52_503 ();
 sg13g2_fill_1 FILLER_52_510 ();
 sg13g2_fill_2 FILLER_52_538 ();
 sg13g2_fill_2 FILLER_52_545 ();
 sg13g2_fill_1 FILLER_52_547 ();
 sg13g2_fill_1 FILLER_52_590 ();
 sg13g2_decap_8 FILLER_52_609 ();
 sg13g2_decap_8 FILLER_52_616 ();
 sg13g2_decap_4 FILLER_52_694 ();
 sg13g2_decap_4 FILLER_52_711 ();
 sg13g2_decap_4 FILLER_52_755 ();
 sg13g2_fill_2 FILLER_52_759 ();
 sg13g2_decap_8 FILLER_52_815 ();
 sg13g2_decap_8 FILLER_52_822 ();
 sg13g2_decap_8 FILLER_52_829 ();
 sg13g2_fill_2 FILLER_52_836 ();
 sg13g2_fill_1 FILLER_52_838 ();
 sg13g2_decap_8 FILLER_52_891 ();
 sg13g2_decap_8 FILLER_52_898 ();
 sg13g2_decap_8 FILLER_52_905 ();
 sg13g2_decap_4 FILLER_52_912 ();
 sg13g2_decap_8 FILLER_52_948 ();
 sg13g2_decap_8 FILLER_52_955 ();
 sg13g2_fill_1 FILLER_52_962 ();
 sg13g2_decap_8 FILLER_52_968 ();
 sg13g2_decap_8 FILLER_52_975 ();
 sg13g2_fill_2 FILLER_52_1072 ();
 sg13g2_fill_1 FILLER_52_1074 ();
 sg13g2_fill_2 FILLER_52_1103 ();
 sg13g2_decap_4 FILLER_52_1159 ();
 sg13g2_fill_1 FILLER_52_1163 ();
 sg13g2_decap_8 FILLER_52_1213 ();
 sg13g2_decap_8 FILLER_52_1220 ();
 sg13g2_decap_8 FILLER_52_1227 ();
 sg13g2_decap_8 FILLER_52_1234 ();
 sg13g2_decap_8 FILLER_52_1241 ();
 sg13g2_decap_4 FILLER_52_1248 ();
 sg13g2_fill_1 FILLER_52_1252 ();
 sg13g2_fill_2 FILLER_52_1269 ();
 sg13g2_fill_2 FILLER_52_1301 ();
 sg13g2_fill_1 FILLER_52_1303 ();
 sg13g2_fill_1 FILLER_52_1335 ();
 sg13g2_decap_8 FILLER_52_1341 ();
 sg13g2_decap_8 FILLER_52_1348 ();
 sg13g2_decap_8 FILLER_52_1355 ();
 sg13g2_decap_8 FILLER_52_1362 ();
 sg13g2_fill_2 FILLER_52_1369 ();
 sg13g2_fill_1 FILLER_52_1398 ();
 sg13g2_fill_2 FILLER_52_1425 ();
 sg13g2_decap_4 FILLER_52_1437 ();
 sg13g2_fill_2 FILLER_52_1477 ();
 sg13g2_fill_1 FILLER_52_1479 ();
 sg13g2_fill_2 FILLER_52_1488 ();
 sg13g2_fill_1 FILLER_52_1490 ();
 sg13g2_fill_2 FILLER_52_1501 ();
 sg13g2_fill_1 FILLER_52_1503 ();
 sg13g2_decap_8 FILLER_52_1517 ();
 sg13g2_fill_2 FILLER_52_1551 ();
 sg13g2_decap_8 FILLER_52_1580 ();
 sg13g2_decap_8 FILLER_52_1587 ();
 sg13g2_fill_2 FILLER_52_1594 ();
 sg13g2_fill_2 FILLER_52_1612 ();
 sg13g2_fill_1 FILLER_52_1614 ();
 sg13g2_fill_2 FILLER_52_1649 ();
 sg13g2_fill_1 FILLER_52_1678 ();
 sg13g2_decap_4 FILLER_52_1694 ();
 sg13g2_fill_2 FILLER_52_1712 ();
 sg13g2_fill_1 FILLER_52_1714 ();
 sg13g2_fill_2 FILLER_52_1718 ();
 sg13g2_decap_8 FILLER_52_1743 ();
 sg13g2_decap_4 FILLER_52_1750 ();
 sg13g2_fill_1 FILLER_52_1754 ();
 sg13g2_fill_1 FILLER_52_1773 ();
 sg13g2_decap_8 FILLER_52_1787 ();
 sg13g2_fill_2 FILLER_52_1807 ();
 sg13g2_fill_1 FILLER_52_1809 ();
 sg13g2_fill_1 FILLER_52_1841 ();
 sg13g2_decap_4 FILLER_52_1875 ();
 sg13g2_fill_2 FILLER_52_1879 ();
 sg13g2_fill_2 FILLER_52_1951 ();
 sg13g2_fill_1 FILLER_52_1953 ();
 sg13g2_fill_2 FILLER_52_1968 ();
 sg13g2_decap_8 FILLER_52_1983 ();
 sg13g2_fill_1 FILLER_52_1990 ();
 sg13g2_fill_1 FILLER_52_1996 ();
 sg13g2_fill_2 FILLER_52_2002 ();
 sg13g2_fill_2 FILLER_52_2024 ();
 sg13g2_fill_2 FILLER_52_2029 ();
 sg13g2_fill_1 FILLER_52_2031 ();
 sg13g2_decap_4 FILLER_52_2037 ();
 sg13g2_fill_1 FILLER_52_2041 ();
 sg13g2_fill_2 FILLER_52_2050 ();
 sg13g2_decap_8 FILLER_52_2067 ();
 sg13g2_decap_4 FILLER_52_2074 ();
 sg13g2_fill_1 FILLER_52_2078 ();
 sg13g2_decap_4 FILLER_52_2089 ();
 sg13g2_fill_1 FILLER_52_2093 ();
 sg13g2_decap_4 FILLER_52_2099 ();
 sg13g2_fill_1 FILLER_52_2103 ();
 sg13g2_decap_4 FILLER_52_2108 ();
 sg13g2_decap_8 FILLER_52_2124 ();
 sg13g2_decap_8 FILLER_52_2131 ();
 sg13g2_fill_1 FILLER_52_2138 ();
 sg13g2_decap_8 FILLER_52_2157 ();
 sg13g2_decap_8 FILLER_52_2164 ();
 sg13g2_decap_8 FILLER_52_2171 ();
 sg13g2_fill_2 FILLER_52_2178 ();
 sg13g2_fill_1 FILLER_52_2180 ();
 sg13g2_decap_4 FILLER_52_2193 ();
 sg13g2_fill_2 FILLER_52_2197 ();
 sg13g2_decap_8 FILLER_52_2204 ();
 sg13g2_fill_2 FILLER_52_2211 ();
 sg13g2_fill_1 FILLER_52_2213 ();
 sg13g2_decap_8 FILLER_52_2217 ();
 sg13g2_decap_4 FILLER_52_2224 ();
 sg13g2_fill_1 FILLER_52_2228 ();
 sg13g2_fill_1 FILLER_52_2247 ();
 sg13g2_decap_8 FILLER_52_2281 ();
 sg13g2_decap_4 FILLER_52_2288 ();
 sg13g2_decap_8 FILLER_52_2296 ();
 sg13g2_decap_4 FILLER_52_2303 ();
 sg13g2_fill_1 FILLER_52_2307 ();
 sg13g2_decap_8 FILLER_52_2313 ();
 sg13g2_decap_8 FILLER_52_2320 ();
 sg13g2_fill_1 FILLER_52_2327 ();
 sg13g2_fill_1 FILLER_52_2369 ();
 sg13g2_decap_8 FILLER_52_2398 ();
 sg13g2_decap_4 FILLER_52_2405 ();
 sg13g2_fill_1 FILLER_52_2409 ();
 sg13g2_decap_8 FILLER_52_2464 ();
 sg13g2_decap_8 FILLER_52_2471 ();
 sg13g2_decap_8 FILLER_52_2478 ();
 sg13g2_fill_1 FILLER_52_2485 ();
 sg13g2_decap_4 FILLER_52_2515 ();
 sg13g2_fill_2 FILLER_52_2519 ();
 sg13g2_decap_8 FILLER_52_2534 ();
 sg13g2_fill_2 FILLER_52_2541 ();
 sg13g2_fill_1 FILLER_52_2543 ();
 sg13g2_decap_8 FILLER_52_2609 ();
 sg13g2_decap_4 FILLER_52_2616 ();
 sg13g2_fill_1 FILLER_52_2620 ();
 sg13g2_fill_2 FILLER_52_2648 ();
 sg13g2_fill_1 FILLER_52_2650 ();
 sg13g2_decap_4 FILLER_52_2705 ();
 sg13g2_fill_2 FILLER_52_2709 ();
 sg13g2_decap_8 FILLER_52_2720 ();
 sg13g2_decap_8 FILLER_52_2727 ();
 sg13g2_decap_8 FILLER_52_2793 ();
 sg13g2_decap_4 FILLER_52_2800 ();
 sg13g2_fill_1 FILLER_52_2804 ();
 sg13g2_decap_8 FILLER_52_2855 ();
 sg13g2_decap_8 FILLER_52_2862 ();
 sg13g2_fill_2 FILLER_52_2869 ();
 sg13g2_fill_1 FILLER_52_2871 ();
 sg13g2_decap_8 FILLER_52_2881 ();
 sg13g2_decap_8 FILLER_52_2888 ();
 sg13g2_decap_8 FILLER_52_2895 ();
 sg13g2_decap_8 FILLER_52_2902 ();
 sg13g2_decap_4 FILLER_52_2909 ();
 sg13g2_fill_1 FILLER_52_2913 ();
 sg13g2_decap_8 FILLER_52_2924 ();
 sg13g2_decap_8 FILLER_52_2952 ();
 sg13g2_decap_8 FILLER_52_2959 ();
 sg13g2_decap_8 FILLER_52_2966 ();
 sg13g2_decap_4 FILLER_52_2973 ();
 sg13g2_fill_2 FILLER_52_2977 ();
 sg13g2_fill_2 FILLER_52_2983 ();
 sg13g2_decap_8 FILLER_52_3007 ();
 sg13g2_fill_2 FILLER_52_3014 ();
 sg13g2_fill_1 FILLER_52_3016 ();
 sg13g2_decap_8 FILLER_52_3057 ();
 sg13g2_decap_8 FILLER_52_3064 ();
 sg13g2_decap_8 FILLER_52_3071 ();
 sg13g2_decap_8 FILLER_52_3078 ();
 sg13g2_decap_8 FILLER_52_3085 ();
 sg13g2_fill_2 FILLER_52_3092 ();
 sg13g2_fill_1 FILLER_52_3094 ();
 sg13g2_fill_1 FILLER_52_3108 ();
 sg13g2_decap_8 FILLER_52_3118 ();
 sg13g2_decap_8 FILLER_52_3125 ();
 sg13g2_fill_2 FILLER_52_3132 ();
 sg13g2_fill_1 FILLER_52_3134 ();
 sg13g2_fill_2 FILLER_52_3175 ();
 sg13g2_fill_1 FILLER_52_3177 ();
 sg13g2_decap_8 FILLER_52_3187 ();
 sg13g2_decap_4 FILLER_52_3194 ();
 sg13g2_fill_2 FILLER_52_3198 ();
 sg13g2_decap_4 FILLER_52_3231 ();
 sg13g2_decap_8 FILLER_52_3244 ();
 sg13g2_decap_4 FILLER_52_3251 ();
 sg13g2_decap_8 FILLER_52_3334 ();
 sg13g2_fill_1 FILLER_52_3341 ();
 sg13g2_decap_8 FILLER_52_3347 ();
 sg13g2_fill_1 FILLER_52_3377 ();
 sg13g2_decap_8 FILLER_52_3422 ();
 sg13g2_decap_8 FILLER_52_3429 ();
 sg13g2_decap_4 FILLER_52_3436 ();
 sg13g2_fill_1 FILLER_52_3440 ();
 sg13g2_fill_2 FILLER_52_3445 ();
 sg13g2_fill_1 FILLER_52_3447 ();
 sg13g2_decap_8 FILLER_52_3513 ();
 sg13g2_fill_1 FILLER_52_3520 ();
 sg13g2_fill_2 FILLER_52_3575 ();
 sg13g2_fill_1 FILLER_52_3577 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_11 ();
 sg13g2_fill_2 FILLER_53_48 ();
 sg13g2_fill_1 FILLER_53_50 ();
 sg13g2_fill_2 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_80 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_decap_8 FILLER_53_146 ();
 sg13g2_decap_8 FILLER_53_163 ();
 sg13g2_decap_8 FILLER_53_179 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_2 FILLER_53_275 ();
 sg13g2_fill_1 FILLER_53_277 ();
 sg13g2_decap_8 FILLER_53_335 ();
 sg13g2_decap_8 FILLER_53_342 ();
 sg13g2_fill_1 FILLER_53_349 ();
 sg13g2_fill_1 FILLER_53_378 ();
 sg13g2_fill_1 FILLER_53_388 ();
 sg13g2_decap_8 FILLER_53_424 ();
 sg13g2_decap_8 FILLER_53_431 ();
 sg13g2_decap_8 FILLER_53_438 ();
 sg13g2_fill_1 FILLER_53_445 ();
 sg13g2_decap_4 FILLER_53_502 ();
 sg13g2_fill_1 FILLER_53_506 ();
 sg13g2_fill_2 FILLER_53_516 ();
 sg13g2_fill_1 FILLER_53_518 ();
 sg13g2_decap_8 FILLER_53_594 ();
 sg13g2_decap_8 FILLER_53_601 ();
 sg13g2_decap_8 FILLER_53_608 ();
 sg13g2_fill_1 FILLER_53_615 ();
 sg13g2_fill_2 FILLER_53_650 ();
 sg13g2_fill_2 FILLER_53_675 ();
 sg13g2_fill_1 FILLER_53_677 ();
 sg13g2_decap_4 FILLER_53_692 ();
 sg13g2_decap_8 FILLER_53_705 ();
 sg13g2_fill_1 FILLER_53_712 ();
 sg13g2_fill_1 FILLER_53_821 ();
 sg13g2_fill_1 FILLER_53_858 ();
 sg13g2_decap_8 FILLER_53_886 ();
 sg13g2_decap_8 FILLER_53_902 ();
 sg13g2_decap_8 FILLER_53_909 ();
 sg13g2_fill_2 FILLER_53_916 ();
 sg13g2_fill_1 FILLER_53_918 ();
 sg13g2_fill_1 FILLER_53_932 ();
 sg13g2_decap_4 FILLER_53_946 ();
 sg13g2_fill_2 FILLER_53_959 ();
 sg13g2_fill_1 FILLER_53_967 ();
 sg13g2_decap_4 FILLER_53_1001 ();
 sg13g2_decap_4 FILLER_53_1018 ();
 sg13g2_decap_4 FILLER_53_1095 ();
 sg13g2_fill_2 FILLER_53_1099 ();
 sg13g2_decap_8 FILLER_53_1148 ();
 sg13g2_decap_8 FILLER_53_1155 ();
 sg13g2_decap_4 FILLER_53_1162 ();
 sg13g2_fill_2 FILLER_53_1166 ();
 sg13g2_decap_4 FILLER_53_1218 ();
 sg13g2_fill_2 FILLER_53_1222 ();
 sg13g2_decap_8 FILLER_53_1229 ();
 sg13g2_decap_8 FILLER_53_1236 ();
 sg13g2_fill_1 FILLER_53_1243 ();
 sg13g2_decap_8 FILLER_53_1251 ();
 sg13g2_fill_2 FILLER_53_1258 ();
 sg13g2_fill_2 FILLER_53_1273 ();
 sg13g2_fill_1 FILLER_53_1275 ();
 sg13g2_decap_8 FILLER_53_1297 ();
 sg13g2_fill_1 FILLER_53_1315 ();
 sg13g2_decap_8 FILLER_53_1334 ();
 sg13g2_fill_1 FILLER_53_1341 ();
 sg13g2_fill_2 FILLER_53_1355 ();
 sg13g2_fill_1 FILLER_53_1357 ();
 sg13g2_decap_8 FILLER_53_1435 ();
 sg13g2_decap_4 FILLER_53_1442 ();
 sg13g2_fill_2 FILLER_53_1492 ();
 sg13g2_decap_4 FILLER_53_1509 ();
 sg13g2_fill_2 FILLER_53_1513 ();
 sg13g2_fill_2 FILLER_53_1528 ();
 sg13g2_fill_1 FILLER_53_1530 ();
 sg13g2_decap_4 FILLER_53_1540 ();
 sg13g2_fill_1 FILLER_53_1556 ();
 sg13g2_fill_1 FILLER_53_1560 ();
 sg13g2_decap_8 FILLER_53_1576 ();
 sg13g2_decap_8 FILLER_53_1583 ();
 sg13g2_decap_8 FILLER_53_1590 ();
 sg13g2_fill_2 FILLER_53_1597 ();
 sg13g2_fill_2 FILLER_53_1615 ();
 sg13g2_decap_8 FILLER_53_1621 ();
 sg13g2_decap_8 FILLER_53_1628 ();
 sg13g2_fill_2 FILLER_53_1635 ();
 sg13g2_fill_1 FILLER_53_1684 ();
 sg13g2_fill_1 FILLER_53_1737 ();
 sg13g2_decap_8 FILLER_53_1751 ();
 sg13g2_decap_8 FILLER_53_1781 ();
 sg13g2_decap_8 FILLER_53_1788 ();
 sg13g2_decap_8 FILLER_53_1795 ();
 sg13g2_decap_8 FILLER_53_1802 ();
 sg13g2_fill_2 FILLER_53_1809 ();
 sg13g2_fill_1 FILLER_53_1811 ();
 sg13g2_fill_2 FILLER_53_1822 ();
 sg13g2_decap_4 FILLER_53_1873 ();
 sg13g2_fill_1 FILLER_53_1877 ();
 sg13g2_decap_8 FILLER_53_1914 ();
 sg13g2_decap_8 FILLER_53_1921 ();
 sg13g2_fill_2 FILLER_53_1928 ();
 sg13g2_fill_1 FILLER_53_1930 ();
 sg13g2_decap_4 FILLER_53_1936 ();
 sg13g2_fill_1 FILLER_53_1940 ();
 sg13g2_decap_8 FILLER_53_1963 ();
 sg13g2_decap_8 FILLER_53_1970 ();
 sg13g2_decap_8 FILLER_53_1977 ();
 sg13g2_decap_8 FILLER_53_1984 ();
 sg13g2_fill_2 FILLER_53_1991 ();
 sg13g2_fill_1 FILLER_53_1993 ();
 sg13g2_decap_8 FILLER_53_2043 ();
 sg13g2_decap_8 FILLER_53_2050 ();
 sg13g2_decap_8 FILLER_53_2057 ();
 sg13g2_decap_8 FILLER_53_2064 ();
 sg13g2_decap_8 FILLER_53_2071 ();
 sg13g2_decap_4 FILLER_53_2078 ();
 sg13g2_fill_1 FILLER_53_2082 ();
 sg13g2_decap_8 FILLER_53_2087 ();
 sg13g2_decap_8 FILLER_53_2094 ();
 sg13g2_decap_8 FILLER_53_2101 ();
 sg13g2_decap_8 FILLER_53_2108 ();
 sg13g2_decap_8 FILLER_53_2115 ();
 sg13g2_decap_8 FILLER_53_2122 ();
 sg13g2_decap_8 FILLER_53_2145 ();
 sg13g2_decap_8 FILLER_53_2152 ();
 sg13g2_decap_8 FILLER_53_2159 ();
 sg13g2_decap_8 FILLER_53_2166 ();
 sg13g2_decap_4 FILLER_53_2173 ();
 sg13g2_fill_1 FILLER_53_2177 ();
 sg13g2_fill_1 FILLER_53_2212 ();
 sg13g2_decap_8 FILLER_53_2226 ();
 sg13g2_fill_2 FILLER_53_2233 ();
 sg13g2_decap_8 FILLER_53_2257 ();
 sg13g2_fill_2 FILLER_53_2264 ();
 sg13g2_fill_1 FILLER_53_2303 ();
 sg13g2_fill_2 FILLER_53_2336 ();
 sg13g2_decap_4 FILLER_53_2366 ();
 sg13g2_fill_1 FILLER_53_2370 ();
 sg13g2_decap_8 FILLER_53_2384 ();
 sg13g2_decap_4 FILLER_53_2391 ();
 sg13g2_decap_8 FILLER_53_2408 ();
 sg13g2_decap_4 FILLER_53_2419 ();
 sg13g2_decap_8 FILLER_53_2455 ();
 sg13g2_decap_8 FILLER_53_2462 ();
 sg13g2_decap_8 FILLER_53_2469 ();
 sg13g2_decap_4 FILLER_53_2476 ();
 sg13g2_fill_2 FILLER_53_2489 ();
 sg13g2_fill_1 FILLER_53_2491 ();
 sg13g2_decap_8 FILLER_53_2505 ();
 sg13g2_decap_8 FILLER_53_2512 ();
 sg13g2_decap_8 FILLER_53_2519 ();
 sg13g2_decap_8 FILLER_53_2526 ();
 sg13g2_decap_8 FILLER_53_2533 ();
 sg13g2_decap_8 FILLER_53_2540 ();
 sg13g2_fill_2 FILLER_53_2547 ();
 sg13g2_fill_1 FILLER_53_2549 ();
 sg13g2_fill_1 FILLER_53_2593 ();
 sg13g2_decap_8 FILLER_53_2599 ();
 sg13g2_decap_4 FILLER_53_2606 ();
 sg13g2_fill_1 FILLER_53_2610 ();
 sg13g2_decap_4 FILLER_53_2642 ();
 sg13g2_decap_4 FILLER_53_2678 ();
 sg13g2_fill_1 FILLER_53_2682 ();
 sg13g2_decap_8 FILLER_53_2687 ();
 sg13g2_decap_8 FILLER_53_2694 ();
 sg13g2_decap_4 FILLER_53_2701 ();
 sg13g2_fill_1 FILLER_53_2705 ();
 sg13g2_decap_8 FILLER_53_2719 ();
 sg13g2_decap_8 FILLER_53_2726 ();
 sg13g2_fill_2 FILLER_53_2750 ();
 sg13g2_fill_1 FILLER_53_2752 ();
 sg13g2_fill_2 FILLER_53_2788 ();
 sg13g2_decap_8 FILLER_53_2857 ();
 sg13g2_fill_1 FILLER_53_2864 ();
 sg13g2_fill_1 FILLER_53_2879 ();
 sg13g2_decap_8 FILLER_53_2889 ();
 sg13g2_decap_8 FILLER_53_2896 ();
 sg13g2_fill_1 FILLER_53_2903 ();
 sg13g2_decap_8 FILLER_53_2959 ();
 sg13g2_decap_4 FILLER_53_2966 ();
 sg13g2_decap_8 FILLER_53_3001 ();
 sg13g2_fill_2 FILLER_53_3008 ();
 sg13g2_fill_1 FILLER_53_3010 ();
 sg13g2_decap_8 FILLER_53_3073 ();
 sg13g2_decap_8 FILLER_53_3080 ();
 sg13g2_decap_8 FILLER_53_3087 ();
 sg13g2_fill_2 FILLER_53_3094 ();
 sg13g2_fill_1 FILLER_53_3096 ();
 sg13g2_decap_8 FILLER_53_3110 ();
 sg13g2_decap_4 FILLER_53_3117 ();
 sg13g2_fill_2 FILLER_53_3121 ();
 sg13g2_fill_2 FILLER_53_3133 ();
 sg13g2_fill_1 FILLER_53_3135 ();
 sg13g2_fill_2 FILLER_53_3145 ();
 sg13g2_fill_1 FILLER_53_3147 ();
 sg13g2_decap_8 FILLER_53_3175 ();
 sg13g2_fill_2 FILLER_53_3182 ();
 sg13g2_fill_2 FILLER_53_3211 ();
 sg13g2_decap_8 FILLER_53_3244 ();
 sg13g2_decap_8 FILLER_53_3251 ();
 sg13g2_fill_2 FILLER_53_3258 ();
 sg13g2_decap_8 FILLER_53_3297 ();
 sg13g2_decap_4 FILLER_53_3304 ();
 sg13g2_fill_2 FILLER_53_3308 ();
 sg13g2_decap_8 FILLER_53_3324 ();
 sg13g2_decap_8 FILLER_53_3331 ();
 sg13g2_decap_8 FILLER_53_3338 ();
 sg13g2_decap_8 FILLER_53_3345 ();
 sg13g2_decap_8 FILLER_53_3352 ();
 sg13g2_fill_1 FILLER_53_3359 ();
 sg13g2_decap_8 FILLER_53_3364 ();
 sg13g2_fill_1 FILLER_53_3371 ();
 sg13g2_decap_8 FILLER_53_3381 ();
 sg13g2_fill_1 FILLER_53_3388 ();
 sg13g2_decap_4 FILLER_53_3399 ();
 sg13g2_fill_2 FILLER_53_3403 ();
 sg13g2_decap_8 FILLER_53_3414 ();
 sg13g2_decap_8 FILLER_53_3421 ();
 sg13g2_fill_2 FILLER_53_3428 ();
 sg13g2_fill_1 FILLER_53_3430 ();
 sg13g2_decap_8 FILLER_53_3436 ();
 sg13g2_decap_8 FILLER_53_3443 ();
 sg13g2_fill_2 FILLER_53_3450 ();
 sg13g2_fill_1 FILLER_53_3452 ();
 sg13g2_fill_2 FILLER_53_3475 ();
 sg13g2_fill_2 FILLER_53_3503 ();
 sg13g2_fill_1 FILLER_53_3505 ();
 sg13g2_decap_8 FILLER_53_3519 ();
 sg13g2_decap_8 FILLER_53_3526 ();
 sg13g2_decap_8 FILLER_53_3570 ();
 sg13g2_fill_1 FILLER_53_3577 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_32 ();
 sg13g2_fill_1 FILLER_54_34 ();
 sg13g2_fill_1 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_4 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_136 ();
 sg13g2_fill_1 FILLER_54_138 ();
 sg13g2_decap_8 FILLER_54_179 ();
 sg13g2_decap_8 FILLER_54_186 ();
 sg13g2_decap_4 FILLER_54_193 ();
 sg13g2_fill_2 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_236 ();
 sg13g2_decap_4 FILLER_54_263 ();
 sg13g2_decap_4 FILLER_54_288 ();
 sg13g2_fill_2 FILLER_54_292 ();
 sg13g2_decap_4 FILLER_54_303 ();
 sg13g2_fill_2 FILLER_54_307 ();
 sg13g2_decap_8 FILLER_54_318 ();
 sg13g2_decap_8 FILLER_54_338 ();
 sg13g2_decap_8 FILLER_54_345 ();
 sg13g2_decap_4 FILLER_54_352 ();
 sg13g2_fill_1 FILLER_54_356 ();
 sg13g2_fill_2 FILLER_54_384 ();
 sg13g2_fill_1 FILLER_54_386 ();
 sg13g2_fill_1 FILLER_54_410 ();
 sg13g2_decap_8 FILLER_54_419 ();
 sg13g2_decap_8 FILLER_54_426 ();
 sg13g2_decap_8 FILLER_54_433 ();
 sg13g2_decap_8 FILLER_54_440 ();
 sg13g2_decap_8 FILLER_54_478 ();
 sg13g2_decap_8 FILLER_54_485 ();
 sg13g2_decap_8 FILLER_54_492 ();
 sg13g2_decap_8 FILLER_54_503 ();
 sg13g2_decap_8 FILLER_54_510 ();
 sg13g2_fill_1 FILLER_54_558 ();
 sg13g2_decap_8 FILLER_54_598 ();
 sg13g2_decap_8 FILLER_54_605 ();
 sg13g2_decap_8 FILLER_54_612 ();
 sg13g2_decap_8 FILLER_54_619 ();
 sg13g2_fill_1 FILLER_54_626 ();
 sg13g2_fill_2 FILLER_54_632 ();
 sg13g2_fill_1 FILLER_54_634 ();
 sg13g2_decap_4 FILLER_54_641 ();
 sg13g2_fill_2 FILLER_54_645 ();
 sg13g2_decap_4 FILLER_54_654 ();
 sg13g2_decap_8 FILLER_54_711 ();
 sg13g2_decap_8 FILLER_54_718 ();
 sg13g2_decap_4 FILLER_54_725 ();
 sg13g2_fill_1 FILLER_54_729 ();
 sg13g2_decap_4 FILLER_54_739 ();
 sg13g2_fill_2 FILLER_54_743 ();
 sg13g2_fill_2 FILLER_54_758 ();
 sg13g2_fill_1 FILLER_54_781 ();
 sg13g2_decap_8 FILLER_54_818 ();
 sg13g2_decap_8 FILLER_54_825 ();
 sg13g2_decap_8 FILLER_54_832 ();
 sg13g2_decap_4 FILLER_54_839 ();
 sg13g2_decap_4 FILLER_54_870 ();
 sg13g2_fill_1 FILLER_54_874 ();
 sg13g2_decap_8 FILLER_54_902 ();
 sg13g2_decap_8 FILLER_54_909 ();
 sg13g2_decap_8 FILLER_54_916 ();
 sg13g2_fill_1 FILLER_54_923 ();
 sg13g2_decap_8 FILLER_54_937 ();
 sg13g2_decap_8 FILLER_54_944 ();
 sg13g2_fill_2 FILLER_54_951 ();
 sg13g2_fill_2 FILLER_54_995 ();
 sg13g2_fill_1 FILLER_54_997 ();
 sg13g2_fill_1 FILLER_54_1044 ();
 sg13g2_decap_4 FILLER_54_1063 ();
 sg13g2_fill_1 FILLER_54_1082 ();
 sg13g2_decap_4 FILLER_54_1101 ();
 sg13g2_fill_1 FILLER_54_1105 ();
 sg13g2_fill_2 FILLER_54_1119 ();
 sg13g2_fill_1 FILLER_54_1121 ();
 sg13g2_fill_2 FILLER_54_1140 ();
 sg13g2_decap_4 FILLER_54_1155 ();
 sg13g2_fill_1 FILLER_54_1159 ();
 sg13g2_fill_2 FILLER_54_1213 ();
 sg13g2_fill_2 FILLER_54_1223 ();
 sg13g2_fill_1 FILLER_54_1230 ();
 sg13g2_decap_8 FILLER_54_1243 ();
 sg13g2_decap_4 FILLER_54_1250 ();
 sg13g2_fill_1 FILLER_54_1254 ();
 sg13g2_fill_1 FILLER_54_1272 ();
 sg13g2_fill_2 FILLER_54_1283 ();
 sg13g2_decap_8 FILLER_54_1290 ();
 sg13g2_fill_2 FILLER_54_1297 ();
 sg13g2_fill_1 FILLER_54_1299 ();
 sg13g2_fill_2 FILLER_54_1313 ();
 sg13g2_decap_8 FILLER_54_1328 ();
 sg13g2_decap_8 FILLER_54_1335 ();
 sg13g2_fill_2 FILLER_54_1342 ();
 sg13g2_fill_1 FILLER_54_1414 ();
 sg13g2_decap_8 FILLER_54_1430 ();
 sg13g2_fill_2 FILLER_54_1437 ();
 sg13g2_fill_2 FILLER_54_1462 ();
 sg13g2_fill_1 FILLER_54_1464 ();
 sg13g2_fill_2 FILLER_54_1485 ();
 sg13g2_decap_8 FILLER_54_1498 ();
 sg13g2_decap_8 FILLER_54_1505 ();
 sg13g2_decap_8 FILLER_54_1512 ();
 sg13g2_decap_8 FILLER_54_1519 ();
 sg13g2_decap_8 FILLER_54_1567 ();
 sg13g2_decap_8 FILLER_54_1574 ();
 sg13g2_decap_8 FILLER_54_1581 ();
 sg13g2_fill_2 FILLER_54_1588 ();
 sg13g2_fill_2 FILLER_54_1617 ();
 sg13g2_decap_8 FILLER_54_1647 ();
 sg13g2_decap_8 FILLER_54_1654 ();
 sg13g2_decap_4 FILLER_54_1661 ();
 sg13g2_fill_1 FILLER_54_1665 ();
 sg13g2_fill_2 FILLER_54_1714 ();
 sg13g2_fill_1 FILLER_54_1716 ();
 sg13g2_decap_8 FILLER_54_1745 ();
 sg13g2_decap_8 FILLER_54_1792 ();
 sg13g2_decap_8 FILLER_54_1799 ();
 sg13g2_fill_2 FILLER_54_1806 ();
 sg13g2_fill_1 FILLER_54_1808 ();
 sg13g2_fill_2 FILLER_54_1816 ();
 sg13g2_fill_2 FILLER_54_1823 ();
 sg13g2_decap_8 FILLER_54_1830 ();
 sg13g2_fill_2 FILLER_54_1837 ();
 sg13g2_fill_1 FILLER_54_1839 ();
 sg13g2_decap_8 FILLER_54_1867 ();
 sg13g2_decap_4 FILLER_54_1874 ();
 sg13g2_fill_2 FILLER_54_1878 ();
 sg13g2_decap_8 FILLER_54_1884 ();
 sg13g2_decap_8 FILLER_54_1918 ();
 sg13g2_decap_8 FILLER_54_1925 ();
 sg13g2_decap_8 FILLER_54_1932 ();
 sg13g2_decap_8 FILLER_54_1939 ();
 sg13g2_decap_8 FILLER_54_1959 ();
 sg13g2_decap_8 FILLER_54_1966 ();
 sg13g2_decap_8 FILLER_54_1973 ();
 sg13g2_fill_2 FILLER_54_1980 ();
 sg13g2_decap_8 FILLER_54_2023 ();
 sg13g2_decap_8 FILLER_54_2030 ();
 sg13g2_fill_1 FILLER_54_2037 ();
 sg13g2_decap_8 FILLER_54_2048 ();
 sg13g2_decap_8 FILLER_54_2055 ();
 sg13g2_decap_8 FILLER_54_2072 ();
 sg13g2_decap_8 FILLER_54_2079 ();
 sg13g2_decap_4 FILLER_54_2086 ();
 sg13g2_decap_8 FILLER_54_2098 ();
 sg13g2_fill_2 FILLER_54_2105 ();
 sg13g2_fill_1 FILLER_54_2107 ();
 sg13g2_decap_4 FILLER_54_2113 ();
 sg13g2_fill_1 FILLER_54_2125 ();
 sg13g2_decap_4 FILLER_54_2131 ();
 sg13g2_fill_2 FILLER_54_2135 ();
 sg13g2_fill_2 FILLER_54_2153 ();
 sg13g2_fill_1 FILLER_54_2155 ();
 sg13g2_fill_2 FILLER_54_2169 ();
 sg13g2_fill_2 FILLER_54_2176 ();
 sg13g2_fill_2 FILLER_54_2182 ();
 sg13g2_fill_1 FILLER_54_2191 ();
 sg13g2_decap_4 FILLER_54_2207 ();
 sg13g2_decap_4 FILLER_54_2234 ();
 sg13g2_fill_2 FILLER_54_2238 ();
 sg13g2_decap_8 FILLER_54_2245 ();
 sg13g2_decap_8 FILLER_54_2252 ();
 sg13g2_fill_1 FILLER_54_2259 ();
 sg13g2_decap_8 FILLER_54_2297 ();
 sg13g2_decap_8 FILLER_54_2304 ();
 sg13g2_decap_4 FILLER_54_2311 ();
 sg13g2_fill_2 FILLER_54_2315 ();
 sg13g2_fill_2 FILLER_54_2343 ();
 sg13g2_fill_1 FILLER_54_2345 ();
 sg13g2_decap_4 FILLER_54_2359 ();
 sg13g2_decap_8 FILLER_54_2390 ();
 sg13g2_decap_8 FILLER_54_2397 ();
 sg13g2_decap_8 FILLER_54_2404 ();
 sg13g2_decap_8 FILLER_54_2411 ();
 sg13g2_decap_8 FILLER_54_2418 ();
 sg13g2_fill_1 FILLER_54_2425 ();
 sg13g2_fill_2 FILLER_54_2435 ();
 sg13g2_fill_1 FILLER_54_2445 ();
 sg13g2_decap_8 FILLER_54_2456 ();
 sg13g2_decap_8 FILLER_54_2473 ();
 sg13g2_decap_8 FILLER_54_2507 ();
 sg13g2_decap_8 FILLER_54_2514 ();
 sg13g2_decap_8 FILLER_54_2521 ();
 sg13g2_decap_8 FILLER_54_2528 ();
 sg13g2_decap_8 FILLER_54_2535 ();
 sg13g2_fill_1 FILLER_54_2542 ();
 sg13g2_fill_1 FILLER_54_2584 ();
 sg13g2_decap_4 FILLER_54_2598 ();
 sg13g2_fill_2 FILLER_54_2602 ();
 sg13g2_decap_4 FILLER_54_2609 ();
 sg13g2_fill_2 FILLER_54_2613 ();
 sg13g2_decap_8 FILLER_54_2648 ();
 sg13g2_fill_1 FILLER_54_2655 ();
 sg13g2_fill_2 FILLER_54_2691 ();
 sg13g2_decap_4 FILLER_54_2702 ();
 sg13g2_fill_1 FILLER_54_2706 ();
 sg13g2_decap_8 FILLER_54_2720 ();
 sg13g2_fill_2 FILLER_54_2727 ();
 sg13g2_fill_1 FILLER_54_2729 ();
 sg13g2_decap_4 FILLER_54_2747 ();
 sg13g2_fill_1 FILLER_54_2751 ();
 sg13g2_decap_8 FILLER_54_2775 ();
 sg13g2_decap_4 FILLER_54_2782 ();
 sg13g2_decap_8 FILLER_54_2795 ();
 sg13g2_decap_8 FILLER_54_2802 ();
 sg13g2_decap_4 FILLER_54_2809 ();
 sg13g2_fill_1 FILLER_54_2817 ();
 sg13g2_decap_8 FILLER_54_2848 ();
 sg13g2_decap_8 FILLER_54_2855 ();
 sg13g2_fill_1 FILLER_54_2862 ();
 sg13g2_fill_1 FILLER_54_2890 ();
 sg13g2_decap_4 FILLER_54_2896 ();
 sg13g2_fill_1 FILLER_54_2900 ();
 sg13g2_decap_8 FILLER_54_2947 ();
 sg13g2_decap_8 FILLER_54_2954 ();
 sg13g2_fill_2 FILLER_54_3016 ();
 sg13g2_fill_2 FILLER_54_3028 ();
 sg13g2_fill_2 FILLER_54_3049 ();
 sg13g2_fill_1 FILLER_54_3051 ();
 sg13g2_fill_2 FILLER_54_3084 ();
 sg13g2_decap_8 FILLER_54_3099 ();
 sg13g2_fill_2 FILLER_54_3106 ();
 sg13g2_decap_4 FILLER_54_3144 ();
 sg13g2_fill_2 FILLER_54_3162 ();
 sg13g2_decap_4 FILLER_54_3173 ();
 sg13g2_fill_2 FILLER_54_3177 ();
 sg13g2_decap_8 FILLER_54_3237 ();
 sg13g2_decap_8 FILLER_54_3244 ();
 sg13g2_decap_8 FILLER_54_3251 ();
 sg13g2_decap_8 FILLER_54_3258 ();
 sg13g2_decap_4 FILLER_54_3265 ();
 sg13g2_fill_1 FILLER_54_3269 ();
 sg13g2_decap_8 FILLER_54_3289 ();
 sg13g2_decap_8 FILLER_54_3296 ();
 sg13g2_decap_8 FILLER_54_3303 ();
 sg13g2_decap_8 FILLER_54_3310 ();
 sg13g2_decap_8 FILLER_54_3317 ();
 sg13g2_decap_4 FILLER_54_3324 ();
 sg13g2_decap_4 FILLER_54_3338 ();
 sg13g2_decap_8 FILLER_54_3355 ();
 sg13g2_decap_4 FILLER_54_3362 ();
 sg13g2_decap_8 FILLER_54_3403 ();
 sg13g2_fill_1 FILLER_54_3410 ();
 sg13g2_decap_4 FILLER_54_3421 ();
 sg13g2_fill_2 FILLER_54_3425 ();
 sg13g2_fill_1 FILLER_54_3463 ();
 sg13g2_decap_4 FILLER_54_3518 ();
 sg13g2_decap_8 FILLER_54_3568 ();
 sg13g2_fill_2 FILLER_54_3575 ();
 sg13g2_fill_1 FILLER_54_3577 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_54 ();
 sg13g2_decap_8 FILLER_55_60 ();
 sg13g2_decap_4 FILLER_55_67 ();
 sg13g2_fill_2 FILLER_55_71 ();
 sg13g2_decap_4 FILLER_55_100 ();
 sg13g2_fill_2 FILLER_55_113 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_fill_2 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_198 ();
 sg13g2_fill_2 FILLER_55_205 ();
 sg13g2_fill_1 FILLER_55_207 ();
 sg13g2_decap_8 FILLER_55_235 ();
 sg13g2_decap_4 FILLER_55_242 ();
 sg13g2_fill_1 FILLER_55_246 ();
 sg13g2_fill_2 FILLER_55_252 ();
 sg13g2_fill_1 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_fill_1 FILLER_55_294 ();
 sg13g2_decap_8 FILLER_55_334 ();
 sg13g2_decap_8 FILLER_55_341 ();
 sg13g2_fill_1 FILLER_55_348 ();
 sg13g2_decap_8 FILLER_55_423 ();
 sg13g2_decap_4 FILLER_55_430 ();
 sg13g2_decap_4 FILLER_55_447 ();
 sg13g2_fill_1 FILLER_55_451 ();
 sg13g2_fill_1 FILLER_55_465 ();
 sg13g2_decap_8 FILLER_55_488 ();
 sg13g2_decap_8 FILLER_55_495 ();
 sg13g2_fill_2 FILLER_55_529 ();
 sg13g2_fill_1 FILLER_55_577 ();
 sg13g2_fill_2 FILLER_55_583 ();
 sg13g2_decap_8 FILLER_55_590 ();
 sg13g2_decap_8 FILLER_55_597 ();
 sg13g2_fill_2 FILLER_55_604 ();
 sg13g2_fill_1 FILLER_55_606 ();
 sg13g2_decap_8 FILLER_55_620 ();
 sg13g2_decap_4 FILLER_55_627 ();
 sg13g2_fill_1 FILLER_55_631 ();
 sg13g2_fill_2 FILLER_55_659 ();
 sg13g2_fill_1 FILLER_55_661 ();
 sg13g2_decap_4 FILLER_55_682 ();
 sg13g2_fill_2 FILLER_55_686 ();
 sg13g2_fill_2 FILLER_55_693 ();
 sg13g2_fill_1 FILLER_55_695 ();
 sg13g2_decap_8 FILLER_55_724 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_decap_4 FILLER_55_762 ();
 sg13g2_fill_1 FILLER_55_766 ();
 sg13g2_fill_2 FILLER_55_782 ();
 sg13g2_fill_1 FILLER_55_784 ();
 sg13g2_decap_4 FILLER_55_794 ();
 sg13g2_fill_1 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_829 ();
 sg13g2_fill_2 FILLER_55_836 ();
 sg13g2_decap_8 FILLER_55_842 ();
 sg13g2_fill_2 FILLER_55_849 ();
 sg13g2_fill_1 FILLER_55_864 ();
 sg13g2_decap_8 FILLER_55_874 ();
 sg13g2_decap_8 FILLER_55_881 ();
 sg13g2_decap_8 FILLER_55_888 ();
 sg13g2_decap_8 FILLER_55_895 ();
 sg13g2_decap_8 FILLER_55_902 ();
 sg13g2_decap_8 FILLER_55_909 ();
 sg13g2_decap_4 FILLER_55_916 ();
 sg13g2_fill_2 FILLER_55_920 ();
 sg13g2_decap_8 FILLER_55_925 ();
 sg13g2_decap_8 FILLER_55_932 ();
 sg13g2_fill_2 FILLER_55_939 ();
 sg13g2_fill_1 FILLER_55_941 ();
 sg13g2_fill_2 FILLER_55_954 ();
 sg13g2_fill_1 FILLER_55_1013 ();
 sg13g2_decap_4 FILLER_55_1052 ();
 sg13g2_fill_1 FILLER_55_1108 ();
 sg13g2_fill_1 FILLER_55_1122 ();
 sg13g2_fill_2 FILLER_55_1129 ();
 sg13g2_decap_8 FILLER_55_1155 ();
 sg13g2_decap_4 FILLER_55_1162 ();
 sg13g2_fill_1 FILLER_55_1166 ();
 sg13g2_fill_2 FILLER_55_1232 ();
 sg13g2_fill_1 FILLER_55_1234 ();
 sg13g2_fill_1 FILLER_55_1290 ();
 sg13g2_fill_1 FILLER_55_1304 ();
 sg13g2_decap_8 FILLER_55_1338 ();
 sg13g2_fill_1 FILLER_55_1345 ();
 sg13g2_fill_1 FILLER_55_1359 ();
 sg13g2_decap_4 FILLER_55_1389 ();
 sg13g2_fill_2 FILLER_55_1393 ();
 sg13g2_fill_2 FILLER_55_1405 ();
 sg13g2_decap_8 FILLER_55_1428 ();
 sg13g2_fill_2 FILLER_55_1435 ();
 sg13g2_fill_1 FILLER_55_1464 ();
 sg13g2_decap_4 FILLER_55_1486 ();
 sg13g2_decap_8 FILLER_55_1495 ();
 sg13g2_decap_4 FILLER_55_1502 ();
 sg13g2_fill_1 FILLER_55_1506 ();
 sg13g2_decap_4 FILLER_55_1512 ();
 sg13g2_fill_1 FILLER_55_1516 ();
 sg13g2_fill_1 FILLER_55_1521 ();
 sg13g2_decap_8 FILLER_55_1571 ();
 sg13g2_fill_2 FILLER_55_1617 ();
 sg13g2_decap_8 FILLER_55_1633 ();
 sg13g2_decap_8 FILLER_55_1640 ();
 sg13g2_decap_8 FILLER_55_1647 ();
 sg13g2_decap_8 FILLER_55_1654 ();
 sg13g2_decap_4 FILLER_55_1661 ();
 sg13g2_fill_2 FILLER_55_1665 ();
 sg13g2_fill_1 FILLER_55_1676 ();
 sg13g2_fill_1 FILLER_55_1682 ();
 sg13g2_decap_4 FILLER_55_1725 ();
 sg13g2_decap_8 FILLER_55_1734 ();
 sg13g2_decap_8 FILLER_55_1741 ();
 sg13g2_decap_8 FILLER_55_1748 ();
 sg13g2_decap_8 FILLER_55_1755 ();
 sg13g2_fill_2 FILLER_55_1798 ();
 sg13g2_fill_1 FILLER_55_1800 ();
 sg13g2_fill_1 FILLER_55_1813 ();
 sg13g2_decap_8 FILLER_55_1830 ();
 sg13g2_decap_8 FILLER_55_1837 ();
 sg13g2_decap_8 FILLER_55_1844 ();
 sg13g2_fill_2 FILLER_55_1860 ();
 sg13g2_fill_1 FILLER_55_1862 ();
 sg13g2_fill_2 FILLER_55_1878 ();
 sg13g2_fill_1 FILLER_55_1880 ();
 sg13g2_decap_8 FILLER_55_1914 ();
 sg13g2_decap_8 FILLER_55_1921 ();
 sg13g2_decap_8 FILLER_55_1928 ();
 sg13g2_fill_2 FILLER_55_1975 ();
 sg13g2_decap_4 FILLER_55_2010 ();
 sg13g2_decap_4 FILLER_55_2023 ();
 sg13g2_decap_8 FILLER_55_2060 ();
 sg13g2_fill_2 FILLER_55_2076 ();
 sg13g2_decap_4 FILLER_55_2104 ();
 sg13g2_fill_1 FILLER_55_2117 ();
 sg13g2_decap_8 FILLER_55_2137 ();
 sg13g2_decap_8 FILLER_55_2144 ();
 sg13g2_decap_4 FILLER_55_2151 ();
 sg13g2_fill_1 FILLER_55_2155 ();
 sg13g2_decap_8 FILLER_55_2167 ();
 sg13g2_decap_8 FILLER_55_2174 ();
 sg13g2_fill_2 FILLER_55_2181 ();
 sg13g2_decap_8 FILLER_55_2191 ();
 sg13g2_decap_8 FILLER_55_2198 ();
 sg13g2_fill_2 FILLER_55_2213 ();
 sg13g2_fill_1 FILLER_55_2215 ();
 sg13g2_decap_8 FILLER_55_2231 ();
 sg13g2_decap_8 FILLER_55_2238 ();
 sg13g2_decap_8 FILLER_55_2245 ();
 sg13g2_decap_8 FILLER_55_2252 ();
 sg13g2_decap_8 FILLER_55_2259 ();
 sg13g2_fill_2 FILLER_55_2266 ();
 sg13g2_fill_1 FILLER_55_2286 ();
 sg13g2_decap_8 FILLER_55_2296 ();
 sg13g2_decap_8 FILLER_55_2303 ();
 sg13g2_decap_8 FILLER_55_2310 ();
 sg13g2_fill_2 FILLER_55_2317 ();
 sg13g2_fill_1 FILLER_55_2350 ();
 sg13g2_decap_8 FILLER_55_2419 ();
 sg13g2_decap_8 FILLER_55_2426 ();
 sg13g2_decap_4 FILLER_55_2433 ();
 sg13g2_fill_1 FILLER_55_2437 ();
 sg13g2_decap_8 FILLER_55_2513 ();
 sg13g2_decap_4 FILLER_55_2520 ();
 sg13g2_fill_1 FILLER_55_2524 ();
 sg13g2_fill_1 FILLER_55_2530 ();
 sg13g2_fill_2 FILLER_55_2612 ();
 sg13g2_fill_1 FILLER_55_2614 ();
 sg13g2_fill_2 FILLER_55_2620 ();
 sg13g2_decap_4 FILLER_55_2666 ();
 sg13g2_decap_8 FILLER_55_2707 ();
 sg13g2_decap_4 FILLER_55_2714 ();
 sg13g2_fill_1 FILLER_55_2718 ();
 sg13g2_decap_4 FILLER_55_2729 ();
 sg13g2_decap_4 FILLER_55_2742 ();
 sg13g2_fill_2 FILLER_55_2746 ();
 sg13g2_fill_2 FILLER_55_2758 ();
 sg13g2_fill_1 FILLER_55_2760 ();
 sg13g2_decap_8 FILLER_55_2780 ();
 sg13g2_decap_8 FILLER_55_2800 ();
 sg13g2_decap_4 FILLER_55_2807 ();
 sg13g2_decap_8 FILLER_55_2841 ();
 sg13g2_decap_8 FILLER_55_2848 ();
 sg13g2_decap_4 FILLER_55_2855 ();
 sg13g2_fill_1 FILLER_55_2859 ();
 sg13g2_decap_8 FILLER_55_2891 ();
 sg13g2_decap_8 FILLER_55_2898 ();
 sg13g2_decap_4 FILLER_55_2905 ();
 sg13g2_decap_8 FILLER_55_2940 ();
 sg13g2_decap_8 FILLER_55_2947 ();
 sg13g2_decap_4 FILLER_55_2954 ();
 sg13g2_decap_4 FILLER_55_3010 ();
 sg13g2_fill_1 FILLER_55_3014 ();
 sg13g2_decap_4 FILLER_55_3032 ();
 sg13g2_fill_1 FILLER_55_3036 ();
 sg13g2_decap_8 FILLER_55_3076 ();
 sg13g2_decap_8 FILLER_55_3083 ();
 sg13g2_decap_8 FILLER_55_3090 ();
 sg13g2_decap_8 FILLER_55_3097 ();
 sg13g2_fill_2 FILLER_55_3104 ();
 sg13g2_decap_8 FILLER_55_3143 ();
 sg13g2_decap_8 FILLER_55_3177 ();
 sg13g2_decap_8 FILLER_55_3246 ();
 sg13g2_decap_8 FILLER_55_3253 ();
 sg13g2_fill_2 FILLER_55_3260 ();
 sg13g2_fill_2 FILLER_55_3303 ();
 sg13g2_fill_1 FILLER_55_3305 ();
 sg13g2_decap_8 FILLER_55_3310 ();
 sg13g2_fill_2 FILLER_55_3317 ();
 sg13g2_fill_1 FILLER_55_3319 ();
 sg13g2_fill_2 FILLER_55_3351 ();
 sg13g2_fill_1 FILLER_55_3353 ();
 sg13g2_decap_4 FILLER_55_3417 ();
 sg13g2_fill_1 FILLER_55_3467 ();
 sg13g2_decap_4 FILLER_55_3505 ();
 sg13g2_decap_4 FILLER_55_3513 ();
 sg13g2_decap_4 FILLER_55_3527 ();
 sg13g2_fill_2 FILLER_55_3531 ();
 sg13g2_decap_8 FILLER_55_3571 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_68 ();
 sg13g2_fill_2 FILLER_56_75 ();
 sg13g2_decap_4 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_117 ();
 sg13g2_fill_2 FILLER_56_133 ();
 sg13g2_fill_2 FILLER_56_145 ();
 sg13g2_fill_1 FILLER_56_152 ();
 sg13g2_fill_2 FILLER_56_159 ();
 sg13g2_fill_2 FILLER_56_174 ();
 sg13g2_fill_1 FILLER_56_176 ();
 sg13g2_decap_4 FILLER_56_213 ();
 sg13g2_fill_1 FILLER_56_217 ();
 sg13g2_fill_1 FILLER_56_245 ();
 sg13g2_decap_4 FILLER_56_255 ();
 sg13g2_decap_4 FILLER_56_286 ();
 sg13g2_fill_2 FILLER_56_290 ();
 sg13g2_fill_1 FILLER_56_305 ();
 sg13g2_decap_4 FILLER_56_310 ();
 sg13g2_fill_1 FILLER_56_314 ();
 sg13g2_decap_8 FILLER_56_328 ();
 sg13g2_decap_8 FILLER_56_335 ();
 sg13g2_fill_2 FILLER_56_342 ();
 sg13g2_fill_1 FILLER_56_344 ();
 sg13g2_decap_4 FILLER_56_372 ();
 sg13g2_fill_2 FILLER_56_398 ();
 sg13g2_decap_4 FILLER_56_449 ();
 sg13g2_fill_2 FILLER_56_453 ();
 sg13g2_fill_2 FILLER_56_488 ();
 sg13g2_fill_1 FILLER_56_490 ();
 sg13g2_fill_2 FILLER_56_532 ();
 sg13g2_fill_1 FILLER_56_567 ();
 sg13g2_fill_2 FILLER_56_586 ();
 sg13g2_fill_2 FILLER_56_615 ();
 sg13g2_fill_2 FILLER_56_622 ();
 sg13g2_fill_1 FILLER_56_624 ();
 sg13g2_fill_1 FILLER_56_641 ();
 sg13g2_decap_4 FILLER_56_673 ();
 sg13g2_fill_1 FILLER_56_677 ();
 sg13g2_decap_8 FILLER_56_690 ();
 sg13g2_decap_8 FILLER_56_697 ();
 sg13g2_fill_2 FILLER_56_704 ();
 sg13g2_decap_8 FILLER_56_715 ();
 sg13g2_decap_8 FILLER_56_722 ();
 sg13g2_decap_8 FILLER_56_729 ();
 sg13g2_fill_1 FILLER_56_741 ();
 sg13g2_fill_1 FILLER_56_778 ();
 sg13g2_fill_1 FILLER_56_825 ();
 sg13g2_fill_2 FILLER_56_832 ();
 sg13g2_decap_4 FILLER_56_849 ();
 sg13g2_decap_8 FILLER_56_867 ();
 sg13g2_decap_8 FILLER_56_874 ();
 sg13g2_decap_8 FILLER_56_881 ();
 sg13g2_fill_2 FILLER_56_888 ();
 sg13g2_decap_4 FILLER_56_894 ();
 sg13g2_fill_1 FILLER_56_956 ();
 sg13g2_fill_2 FILLER_56_980 ();
 sg13g2_fill_1 FILLER_56_996 ();
 sg13g2_fill_1 FILLER_56_1033 ();
 sg13g2_fill_1 FILLER_56_1054 ();
 sg13g2_fill_2 FILLER_56_1085 ();
 sg13g2_decap_4 FILLER_56_1120 ();
 sg13g2_fill_2 FILLER_56_1166 ();
 sg13g2_fill_1 FILLER_56_1168 ();
 sg13g2_fill_2 FILLER_56_1187 ();
 sg13g2_fill_1 FILLER_56_1189 ();
 sg13g2_fill_1 FILLER_56_1247 ();
 sg13g2_decap_8 FILLER_56_1253 ();
 sg13g2_fill_2 FILLER_56_1260 ();
 sg13g2_decap_8 FILLER_56_1292 ();
 sg13g2_fill_1 FILLER_56_1299 ();
 sg13g2_fill_2 FILLER_56_1323 ();
 sg13g2_decap_8 FILLER_56_1334 ();
 sg13g2_decap_8 FILLER_56_1341 ();
 sg13g2_decap_8 FILLER_56_1348 ();
 sg13g2_fill_1 FILLER_56_1355 ();
 sg13g2_fill_1 FILLER_56_1383 ();
 sg13g2_decap_4 FILLER_56_1398 ();
 sg13g2_decap_8 FILLER_56_1425 ();
 sg13g2_decap_8 FILLER_56_1432 ();
 sg13g2_decap_8 FILLER_56_1439 ();
 sg13g2_decap_8 FILLER_56_1446 ();
 sg13g2_decap_4 FILLER_56_1453 ();
 sg13g2_fill_2 FILLER_56_1474 ();
 sg13g2_fill_1 FILLER_56_1476 ();
 sg13g2_decap_4 FILLER_56_1483 ();
 sg13g2_fill_2 FILLER_56_1496 ();
 sg13g2_fill_1 FILLER_56_1506 ();
 sg13g2_decap_8 FILLER_56_1549 ();
 sg13g2_decap_8 FILLER_56_1556 ();
 sg13g2_decap_4 FILLER_56_1563 ();
 sg13g2_fill_2 FILLER_56_1567 ();
 sg13g2_fill_1 FILLER_56_1579 ();
 sg13g2_fill_2 FILLER_56_1585 ();
 sg13g2_fill_1 FILLER_56_1587 ();
 sg13g2_decap_4 FILLER_56_1617 ();
 sg13g2_fill_2 FILLER_56_1631 ();
 sg13g2_fill_1 FILLER_56_1633 ();
 sg13g2_decap_8 FILLER_56_1647 ();
 sg13g2_decap_8 FILLER_56_1654 ();
 sg13g2_decap_8 FILLER_56_1661 ();
 sg13g2_fill_2 FILLER_56_1668 ();
 sg13g2_fill_1 FILLER_56_1670 ();
 sg13g2_decap_8 FILLER_56_1681 ();
 sg13g2_fill_1 FILLER_56_1688 ();
 sg13g2_decap_4 FILLER_56_1699 ();
 sg13g2_decap_8 FILLER_56_1717 ();
 sg13g2_decap_8 FILLER_56_1724 ();
 sg13g2_decap_8 FILLER_56_1731 ();
 sg13g2_decap_8 FILLER_56_1738 ();
 sg13g2_fill_2 FILLER_56_1745 ();
 sg13g2_decap_8 FILLER_56_1756 ();
 sg13g2_decap_8 FILLER_56_1782 ();
 sg13g2_fill_1 FILLER_56_1789 ();
 sg13g2_fill_2 FILLER_56_1794 ();
 sg13g2_decap_4 FILLER_56_1819 ();
 sg13g2_fill_1 FILLER_56_1823 ();
 sg13g2_decap_8 FILLER_56_1830 ();
 sg13g2_fill_1 FILLER_56_1837 ();
 sg13g2_decap_8 FILLER_56_1851 ();
 sg13g2_decap_8 FILLER_56_1858 ();
 sg13g2_fill_2 FILLER_56_1865 ();
 sg13g2_fill_2 FILLER_56_1881 ();
 sg13g2_fill_1 FILLER_56_1883 ();
 sg13g2_decap_8 FILLER_56_1914 ();
 sg13g2_fill_2 FILLER_56_1921 ();
 sg13g2_fill_1 FILLER_56_1923 ();
 sg13g2_fill_1 FILLER_56_1938 ();
 sg13g2_fill_2 FILLER_56_1980 ();
 sg13g2_decap_4 FILLER_56_1986 ();
 sg13g2_fill_2 FILLER_56_2017 ();
 sg13g2_fill_2 FILLER_56_2027 ();
 sg13g2_fill_1 FILLER_56_2029 ();
 sg13g2_decap_4 FILLER_56_2095 ();
 sg13g2_fill_2 FILLER_56_2099 ();
 sg13g2_decap_4 FILLER_56_2147 ();
 sg13g2_fill_1 FILLER_56_2151 ();
 sg13g2_fill_2 FILLER_56_2174 ();
 sg13g2_decap_8 FILLER_56_2192 ();
 sg13g2_decap_8 FILLER_56_2199 ();
 sg13g2_fill_1 FILLER_56_2206 ();
 sg13g2_fill_1 FILLER_56_2216 ();
 sg13g2_decap_8 FILLER_56_2225 ();
 sg13g2_decap_8 FILLER_56_2232 ();
 sg13g2_decap_8 FILLER_56_2239 ();
 sg13g2_decap_8 FILLER_56_2246 ();
 sg13g2_decap_8 FILLER_56_2253 ();
 sg13g2_decap_4 FILLER_56_2260 ();
 sg13g2_decap_8 FILLER_56_2307 ();
 sg13g2_decap_8 FILLER_56_2314 ();
 sg13g2_decap_4 FILLER_56_2321 ();
 sg13g2_fill_2 FILLER_56_2364 ();
 sg13g2_fill_1 FILLER_56_2366 ();
 sg13g2_decap_8 FILLER_56_2403 ();
 sg13g2_decap_8 FILLER_56_2410 ();
 sg13g2_decap_8 FILLER_56_2417 ();
 sg13g2_decap_8 FILLER_56_2424 ();
 sg13g2_decap_8 FILLER_56_2431 ();
 sg13g2_decap_4 FILLER_56_2438 ();
 sg13g2_fill_2 FILLER_56_2442 ();
 sg13g2_decap_4 FILLER_56_2448 ();
 sg13g2_fill_1 FILLER_56_2452 ();
 sg13g2_fill_2 FILLER_56_2470 ();
 sg13g2_fill_1 FILLER_56_2472 ();
 sg13g2_decap_8 FILLER_56_2510 ();
 sg13g2_decap_8 FILLER_56_2517 ();
 sg13g2_decap_8 FILLER_56_2524 ();
 sg13g2_decap_8 FILLER_56_2604 ();
 sg13g2_fill_1 FILLER_56_2611 ();
 sg13g2_decap_8 FILLER_56_2616 ();
 sg13g2_decap_8 FILLER_56_2623 ();
 sg13g2_fill_1 FILLER_56_2630 ();
 sg13g2_decap_8 FILLER_56_2704 ();
 sg13g2_decap_4 FILLER_56_2711 ();
 sg13g2_decap_4 FILLER_56_2742 ();
 sg13g2_decap_8 FILLER_56_2777 ();
 sg13g2_decap_8 FILLER_56_2784 ();
 sg13g2_decap_8 FILLER_56_2791 ();
 sg13g2_fill_2 FILLER_56_2798 ();
 sg13g2_decap_4 FILLER_56_2846 ();
 sg13g2_fill_2 FILLER_56_2850 ();
 sg13g2_fill_1 FILLER_56_2902 ();
 sg13g2_decap_8 FILLER_56_2943 ();
 sg13g2_decap_8 FILLER_56_2950 ();
 sg13g2_decap_8 FILLER_56_2957 ();
 sg13g2_decap_4 FILLER_56_2964 ();
 sg13g2_decap_8 FILLER_56_2988 ();
 sg13g2_fill_1 FILLER_56_2995 ();
 sg13g2_decap_4 FILLER_56_3009 ();
 sg13g2_fill_1 FILLER_56_3013 ();
 sg13g2_fill_1 FILLER_56_3027 ();
 sg13g2_decap_8 FILLER_56_3032 ();
 sg13g2_decap_8 FILLER_56_3039 ();
 sg13g2_fill_1 FILLER_56_3046 ();
 sg13g2_fill_1 FILLER_56_3057 ();
 sg13g2_decap_8 FILLER_56_3066 ();
 sg13g2_fill_2 FILLER_56_3073 ();
 sg13g2_fill_2 FILLER_56_3079 ();
 sg13g2_fill_1 FILLER_56_3081 ();
 sg13g2_decap_8 FILLER_56_3095 ();
 sg13g2_decap_4 FILLER_56_3102 ();
 sg13g2_fill_1 FILLER_56_3106 ();
 sg13g2_fill_2 FILLER_56_3142 ();
 sg13g2_decap_8 FILLER_56_3180 ();
 sg13g2_fill_1 FILLER_56_3187 ();
 sg13g2_decap_4 FILLER_56_3198 ();
 sg13g2_decap_8 FILLER_56_3231 ();
 sg13g2_decap_8 FILLER_56_3238 ();
 sg13g2_decap_8 FILLER_56_3245 ();
 sg13g2_decap_4 FILLER_56_3252 ();
 sg13g2_fill_1 FILLER_56_3256 ();
 sg13g2_decap_8 FILLER_56_3314 ();
 sg13g2_decap_8 FILLER_56_3321 ();
 sg13g2_fill_2 FILLER_56_3328 ();
 sg13g2_fill_1 FILLER_56_3330 ();
 sg13g2_fill_2 FILLER_56_3341 ();
 sg13g2_fill_1 FILLER_56_3343 ();
 sg13g2_fill_1 FILLER_56_3353 ();
 sg13g2_fill_1 FILLER_56_3383 ();
 sg13g2_fill_2 FILLER_56_3425 ();
 sg13g2_fill_2 FILLER_56_3431 ();
 sg13g2_fill_1 FILLER_56_3433 ();
 sg13g2_decap_8 FILLER_56_3451 ();
 sg13g2_decap_8 FILLER_56_3458 ();
 sg13g2_decap_4 FILLER_56_3465 ();
 sg13g2_fill_2 FILLER_56_3469 ();
 sg13g2_decap_8 FILLER_56_3511 ();
 sg13g2_decap_4 FILLER_56_3572 ();
 sg13g2_fill_2 FILLER_56_3576 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_15 ();
 sg13g2_fill_1 FILLER_57_56 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_fill_2 FILLER_57_95 ();
 sg13g2_fill_1 FILLER_57_97 ();
 sg13g2_fill_1 FILLER_57_120 ();
 sg13g2_fill_2 FILLER_57_148 ();
 sg13g2_fill_1 FILLER_57_163 ();
 sg13g2_decap_4 FILLER_57_209 ();
 sg13g2_fill_1 FILLER_57_244 ();
 sg13g2_decap_4 FILLER_57_272 ();
 sg13g2_decap_8 FILLER_57_294 ();
 sg13g2_fill_1 FILLER_57_301 ();
 sg13g2_fill_1 FILLER_57_307 ();
 sg13g2_decap_8 FILLER_57_321 ();
 sg13g2_decap_8 FILLER_57_328 ();
 sg13g2_fill_2 FILLER_57_335 ();
 sg13g2_fill_1 FILLER_57_337 ();
 sg13g2_fill_2 FILLER_57_402 ();
 sg13g2_fill_2 FILLER_57_417 ();
 sg13g2_fill_1 FILLER_57_419 ();
 sg13g2_decap_8 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_57_436 ();
 sg13g2_decap_4 FILLER_57_443 ();
 sg13g2_fill_2 FILLER_57_484 ();
 sg13g2_decap_8 FILLER_57_512 ();
 sg13g2_decap_8 FILLER_57_519 ();
 sg13g2_decap_4 FILLER_57_526 ();
 sg13g2_fill_1 FILLER_57_530 ();
 sg13g2_decap_8 FILLER_57_599 ();
 sg13g2_fill_2 FILLER_57_606 ();
 sg13g2_fill_2 FILLER_57_628 ();
 sg13g2_fill_1 FILLER_57_630 ();
 sg13g2_fill_1 FILLER_57_641 ();
 sg13g2_decap_8 FILLER_57_655 ();
 sg13g2_decap_4 FILLER_57_662 ();
 sg13g2_fill_2 FILLER_57_666 ();
 sg13g2_decap_8 FILLER_57_719 ();
 sg13g2_decap_8 FILLER_57_726 ();
 sg13g2_decap_8 FILLER_57_733 ();
 sg13g2_decap_4 FILLER_57_740 ();
 sg13g2_fill_2 FILLER_57_744 ();
 sg13g2_fill_2 FILLER_57_773 ();
 sg13g2_fill_1 FILLER_57_775 ();
 sg13g2_fill_2 FILLER_57_830 ();
 sg13g2_fill_2 FILLER_57_887 ();
 sg13g2_decap_8 FILLER_57_993 ();
 sg13g2_fill_1 FILLER_57_1000 ();
 sg13g2_decap_8 FILLER_57_1046 ();
 sg13g2_decap_4 FILLER_57_1053 ();
 sg13g2_fill_2 FILLER_57_1085 ();
 sg13g2_decap_4 FILLER_57_1114 ();
 sg13g2_decap_8 FILLER_57_1159 ();
 sg13g2_fill_1 FILLER_57_1166 ();
 sg13g2_fill_2 FILLER_57_1194 ();
 sg13g2_fill_1 FILLER_57_1218 ();
 sg13g2_fill_1 FILLER_57_1228 ();
 sg13g2_fill_2 FILLER_57_1248 ();
 sg13g2_decap_8 FILLER_57_1281 ();
 sg13g2_decap_8 FILLER_57_1288 ();
 sg13g2_decap_8 FILLER_57_1330 ();
 sg13g2_decap_8 FILLER_57_1337 ();
 sg13g2_decap_8 FILLER_57_1380 ();
 sg13g2_fill_1 FILLER_57_1387 ();
 sg13g2_decap_4 FILLER_57_1398 ();
 sg13g2_fill_2 FILLER_57_1423 ();
 sg13g2_decap_8 FILLER_57_1438 ();
 sg13g2_fill_2 FILLER_57_1445 ();
 sg13g2_fill_2 FILLER_57_1482 ();
 sg13g2_decap_4 FILLER_57_1499 ();
 sg13g2_decap_8 FILLER_57_1508 ();
 sg13g2_decap_4 FILLER_57_1515 ();
 sg13g2_decap_8 FILLER_57_1538 ();
 sg13g2_decap_8 FILLER_57_1545 ();
 sg13g2_decap_4 FILLER_57_1552 ();
 sg13g2_decap_4 FILLER_57_1561 ();
 sg13g2_decap_8 FILLER_57_1574 ();
 sg13g2_decap_8 FILLER_57_1581 ();
 sg13g2_decap_4 FILLER_57_1598 ();
 sg13g2_fill_1 FILLER_57_1602 ();
 sg13g2_fill_1 FILLER_57_1616 ();
 sg13g2_decap_8 FILLER_57_1627 ();
 sg13g2_decap_8 FILLER_57_1634 ();
 sg13g2_fill_1 FILLER_57_1641 ();
 sg13g2_fill_2 FILLER_57_1678 ();
 sg13g2_fill_1 FILLER_57_1680 ();
 sg13g2_decap_8 FILLER_57_1713 ();
 sg13g2_fill_2 FILLER_57_1720 ();
 sg13g2_fill_1 FILLER_57_1722 ();
 sg13g2_decap_8 FILLER_57_1766 ();
 sg13g2_decap_8 FILLER_57_1773 ();
 sg13g2_fill_1 FILLER_57_1780 ();
 sg13g2_decap_4 FILLER_57_1787 ();
 sg13g2_decap_8 FILLER_57_1810 ();
 sg13g2_decap_8 FILLER_57_1817 ();
 sg13g2_decap_4 FILLER_57_1824 ();
 sg13g2_fill_2 FILLER_57_1828 ();
 sg13g2_decap_4 FILLER_57_1856 ();
 sg13g2_fill_2 FILLER_57_1874 ();
 sg13g2_fill_1 FILLER_57_1876 ();
 sg13g2_fill_1 FILLER_57_1914 ();
 sg13g2_fill_2 FILLER_57_1928 ();
 sg13g2_decap_8 FILLER_57_1973 ();
 sg13g2_decap_4 FILLER_57_1980 ();
 sg13g2_fill_1 FILLER_57_2002 ();
 sg13g2_decap_8 FILLER_57_2011 ();
 sg13g2_fill_1 FILLER_57_2018 ();
 sg13g2_decap_4 FILLER_57_2028 ();
 sg13g2_fill_2 FILLER_57_2032 ();
 sg13g2_fill_1 FILLER_57_2047 ();
 sg13g2_decap_8 FILLER_57_2057 ();
 sg13g2_decap_8 FILLER_57_2064 ();
 sg13g2_fill_2 FILLER_57_2071 ();
 sg13g2_decap_4 FILLER_57_2086 ();
 sg13g2_fill_2 FILLER_57_2098 ();
 sg13g2_decap_8 FILLER_57_2146 ();
 sg13g2_decap_8 FILLER_57_2153 ();
 sg13g2_decap_8 FILLER_57_2160 ();
 sg13g2_decap_4 FILLER_57_2167 ();
 sg13g2_fill_1 FILLER_57_2171 ();
 sg13g2_decap_8 FILLER_57_2196 ();
 sg13g2_decap_8 FILLER_57_2234 ();
 sg13g2_decap_8 FILLER_57_2241 ();
 sg13g2_decap_8 FILLER_57_2248 ();
 sg13g2_fill_1 FILLER_57_2281 ();
 sg13g2_decap_4 FILLER_57_2308 ();
 sg13g2_fill_1 FILLER_57_2312 ();
 sg13g2_decap_8 FILLER_57_2361 ();
 sg13g2_decap_4 FILLER_57_2368 ();
 sg13g2_fill_2 FILLER_57_2372 ();
 sg13g2_decap_8 FILLER_57_2432 ();
 sg13g2_decap_4 FILLER_57_2439 ();
 sg13g2_fill_1 FILLER_57_2457 ();
 sg13g2_decap_8 FILLER_57_2467 ();
 sg13g2_decap_4 FILLER_57_2474 ();
 sg13g2_fill_1 FILLER_57_2478 ();
 sg13g2_fill_2 FILLER_57_2497 ();
 sg13g2_decap_8 FILLER_57_2533 ();
 sg13g2_fill_2 FILLER_57_2540 ();
 sg13g2_fill_1 FILLER_57_2599 ();
 sg13g2_decap_8 FILLER_57_2609 ();
 sg13g2_decap_8 FILLER_57_2616 ();
 sg13g2_fill_2 FILLER_57_2623 ();
 sg13g2_fill_1 FILLER_57_2625 ();
 sg13g2_fill_2 FILLER_57_2639 ();
 sg13g2_fill_1 FILLER_57_2641 ();
 sg13g2_decap_8 FILLER_57_2659 ();
 sg13g2_decap_4 FILLER_57_2666 ();
 sg13g2_fill_2 FILLER_57_2687 ();
 sg13g2_fill_1 FILLER_57_2689 ();
 sg13g2_decap_4 FILLER_57_2699 ();
 sg13g2_fill_1 FILLER_57_2703 ();
 sg13g2_decap_8 FILLER_57_2772 ();
 sg13g2_decap_8 FILLER_57_2779 ();
 sg13g2_decap_8 FILLER_57_2786 ();
 sg13g2_fill_2 FILLER_57_2793 ();
 sg13g2_fill_1 FILLER_57_2795 ();
 sg13g2_decap_8 FILLER_57_2844 ();
 sg13g2_decap_4 FILLER_57_2851 ();
 sg13g2_decap_8 FILLER_57_2899 ();
 sg13g2_fill_1 FILLER_57_2906 ();
 sg13g2_fill_2 FILLER_57_2920 ();
 sg13g2_fill_1 FILLER_57_2922 ();
 sg13g2_decap_8 FILLER_57_2953 ();
 sg13g2_decap_4 FILLER_57_2960 ();
 sg13g2_fill_2 FILLER_57_2964 ();
 sg13g2_fill_1 FILLER_57_2998 ();
 sg13g2_decap_8 FILLER_57_3012 ();
 sg13g2_fill_2 FILLER_57_3033 ();
 sg13g2_fill_1 FILLER_57_3035 ();
 sg13g2_decap_8 FILLER_57_3063 ();
 sg13g2_decap_8 FILLER_57_3106 ();
 sg13g2_fill_2 FILLER_57_3113 ();
 sg13g2_decap_4 FILLER_57_3129 ();
 sg13g2_fill_2 FILLER_57_3154 ();
 sg13g2_fill_1 FILLER_57_3156 ();
 sg13g2_decap_8 FILLER_57_3191 ();
 sg13g2_fill_1 FILLER_57_3198 ();
 sg13g2_decap_8 FILLER_57_3242 ();
 sg13g2_decap_4 FILLER_57_3249 ();
 sg13g2_fill_2 FILLER_57_3284 ();
 sg13g2_decap_8 FILLER_57_3318 ();
 sg13g2_decap_4 FILLER_57_3325 ();
 sg13g2_fill_1 FILLER_57_3381 ();
 sg13g2_fill_1 FILLER_57_3390 ();
 sg13g2_decap_8 FILLER_57_3412 ();
 sg13g2_fill_2 FILLER_57_3419 ();
 sg13g2_decap_8 FILLER_57_3434 ();
 sg13g2_decap_8 FILLER_57_3441 ();
 sg13g2_decap_8 FILLER_57_3448 ();
 sg13g2_decap_8 FILLER_57_3455 ();
 sg13g2_decap_8 FILLER_57_3462 ();
 sg13g2_fill_2 FILLER_57_3469 ();
 sg13g2_fill_1 FILLER_57_3498 ();
 sg13g2_decap_8 FILLER_57_3508 ();
 sg13g2_decap_8 FILLER_57_3515 ();
 sg13g2_fill_2 FILLER_57_3545 ();
 sg13g2_fill_1 FILLER_57_3547 ();
 sg13g2_fill_2 FILLER_57_3552 ();
 sg13g2_fill_1 FILLER_57_3554 ();
 sg13g2_decap_8 FILLER_57_3564 ();
 sg13g2_decap_8 FILLER_57_3571 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_11 ();
 sg13g2_fill_2 FILLER_58_43 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_4 FILLER_58_77 ();
 sg13g2_fill_2 FILLER_58_85 ();
 sg13g2_fill_1 FILLER_58_116 ();
 sg13g2_decap_4 FILLER_58_121 ();
 sg13g2_fill_1 FILLER_58_125 ();
 sg13g2_decap_4 FILLER_58_130 ();
 sg13g2_fill_2 FILLER_58_134 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_4 FILLER_58_203 ();
 sg13g2_fill_1 FILLER_58_207 ();
 sg13g2_decap_8 FILLER_58_213 ();
 sg13g2_fill_2 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_257 ();
 sg13g2_fill_1 FILLER_58_288 ();
 sg13g2_decap_4 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_330 ();
 sg13g2_fill_1 FILLER_58_414 ();
 sg13g2_fill_1 FILLER_58_420 ();
 sg13g2_decap_4 FILLER_58_430 ();
 sg13g2_decap_8 FILLER_58_443 ();
 sg13g2_fill_2 FILLER_58_450 ();
 sg13g2_fill_1 FILLER_58_452 ();
 sg13g2_decap_8 FILLER_58_490 ();
 sg13g2_decap_8 FILLER_58_497 ();
 sg13g2_decap_8 FILLER_58_504 ();
 sg13g2_decap_8 FILLER_58_511 ();
 sg13g2_decap_8 FILLER_58_518 ();
 sg13g2_decap_8 FILLER_58_525 ();
 sg13g2_decap_8 FILLER_58_532 ();
 sg13g2_decap_8 FILLER_58_539 ();
 sg13g2_fill_2 FILLER_58_546 ();
 sg13g2_fill_1 FILLER_58_548 ();
 sg13g2_fill_2 FILLER_58_575 ();
 sg13g2_fill_1 FILLER_58_577 ();
 sg13g2_fill_2 FILLER_58_583 ();
 sg13g2_fill_1 FILLER_58_585 ();
 sg13g2_decap_8 FILLER_58_596 ();
 sg13g2_decap_8 FILLER_58_649 ();
 sg13g2_decap_8 FILLER_58_656 ();
 sg13g2_decap_8 FILLER_58_663 ();
 sg13g2_decap_8 FILLER_58_670 ();
 sg13g2_fill_2 FILLER_58_677 ();
 sg13g2_decap_8 FILLER_58_725 ();
 sg13g2_decap_8 FILLER_58_732 ();
 sg13g2_fill_1 FILLER_58_770 ();
 sg13g2_decap_8 FILLER_58_780 ();
 sg13g2_decap_4 FILLER_58_787 ();
 sg13g2_fill_1 FILLER_58_808 ();
 sg13g2_fill_1 FILLER_58_850 ();
 sg13g2_fill_2 FILLER_58_865 ();
 sg13g2_decap_8 FILLER_58_923 ();
 sg13g2_decap_4 FILLER_58_930 ();
 sg13g2_fill_1 FILLER_58_934 ();
 sg13g2_fill_2 FILLER_58_979 ();
 sg13g2_decap_8 FILLER_58_994 ();
 sg13g2_decap_4 FILLER_58_1001 ();
 sg13g2_fill_1 FILLER_58_1032 ();
 sg13g2_decap_8 FILLER_58_1042 ();
 sg13g2_decap_8 FILLER_58_1049 ();
 sg13g2_fill_2 FILLER_58_1056 ();
 sg13g2_fill_1 FILLER_58_1058 ();
 sg13g2_fill_2 FILLER_58_1105 ();
 sg13g2_decap_4 FILLER_58_1142 ();
 sg13g2_decap_8 FILLER_58_1155 ();
 sg13g2_decap_8 FILLER_58_1162 ();
 sg13g2_fill_2 FILLER_58_1169 ();
 sg13g2_fill_1 FILLER_58_1171 ();
 sg13g2_fill_1 FILLER_58_1242 ();
 sg13g2_decap_4 FILLER_58_1277 ();
 sg13g2_fill_2 FILLER_58_1281 ();
 sg13g2_fill_2 FILLER_58_1296 ();
 sg13g2_decap_8 FILLER_58_1339 ();
 sg13g2_decap_8 FILLER_58_1346 ();
 sg13g2_decap_4 FILLER_58_1353 ();
 sg13g2_fill_2 FILLER_58_1357 ();
 sg13g2_decap_4 FILLER_58_1413 ();
 sg13g2_fill_2 FILLER_58_1426 ();
 sg13g2_fill_2 FILLER_58_1446 ();
 sg13g2_fill_1 FILLER_58_1448 ();
 sg13g2_decap_4 FILLER_58_1481 ();
 sg13g2_fill_1 FILLER_58_1489 ();
 sg13g2_fill_1 FILLER_58_1495 ();
 sg13g2_decap_8 FILLER_58_1504 ();
 sg13g2_decap_8 FILLER_58_1518 ();
 sg13g2_decap_4 FILLER_58_1525 ();
 sg13g2_decap_8 FILLER_58_1533 ();
 sg13g2_decap_8 FILLER_58_1540 ();
 sg13g2_decap_8 FILLER_58_1547 ();
 sg13g2_fill_2 FILLER_58_1554 ();
 sg13g2_fill_2 FILLER_58_1574 ();
 sg13g2_fill_1 FILLER_58_1576 ();
 sg13g2_decap_8 FILLER_58_1587 ();
 sg13g2_decap_8 FILLER_58_1594 ();
 sg13g2_decap_8 FILLER_58_1601 ();
 sg13g2_fill_2 FILLER_58_1608 ();
 sg13g2_decap_4 FILLER_58_1615 ();
 sg13g2_decap_8 FILLER_58_1623 ();
 sg13g2_decap_8 FILLER_58_1630 ();
 sg13g2_decap_4 FILLER_58_1637 ();
 sg13g2_decap_4 FILLER_58_1699 ();
 sg13g2_decap_8 FILLER_58_1712 ();
 sg13g2_fill_2 FILLER_58_1719 ();
 sg13g2_fill_1 FILLER_58_1721 ();
 sg13g2_decap_4 FILLER_58_1764 ();
 sg13g2_fill_1 FILLER_58_1768 ();
 sg13g2_decap_4 FILLER_58_1792 ();
 sg13g2_fill_1 FILLER_58_1796 ();
 sg13g2_decap_8 FILLER_58_1801 ();
 sg13g2_decap_8 FILLER_58_1808 ();
 sg13g2_fill_1 FILLER_58_1815 ();
 sg13g2_decap_4 FILLER_58_1821 ();
 sg13g2_fill_1 FILLER_58_1825 ();
 sg13g2_fill_2 FILLER_58_1835 ();
 sg13g2_decap_8 FILLER_58_1858 ();
 sg13g2_fill_2 FILLER_58_1865 ();
 sg13g2_fill_2 FILLER_58_1871 ();
 sg13g2_decap_4 FILLER_58_1905 ();
 sg13g2_fill_1 FILLER_58_1909 ();
 sg13g2_fill_1 FILLER_58_1990 ();
 sg13g2_decap_8 FILLER_58_2037 ();
 sg13g2_decap_8 FILLER_58_2044 ();
 sg13g2_decap_8 FILLER_58_2051 ();
 sg13g2_decap_4 FILLER_58_2058 ();
 sg13g2_decap_4 FILLER_58_2098 ();
 sg13g2_fill_1 FILLER_58_2102 ();
 sg13g2_decap_8 FILLER_58_2108 ();
 sg13g2_fill_1 FILLER_58_2119 ();
 sg13g2_fill_1 FILLER_58_2128 ();
 sg13g2_decap_8 FILLER_58_2145 ();
 sg13g2_decap_8 FILLER_58_2152 ();
 sg13g2_decap_4 FILLER_58_2159 ();
 sg13g2_fill_2 FILLER_58_2163 ();
 sg13g2_decap_4 FILLER_58_2198 ();
 sg13g2_decap_4 FILLER_58_2236 ();
 sg13g2_fill_2 FILLER_58_2240 ();
 sg13g2_fill_1 FILLER_58_2255 ();
 sg13g2_fill_2 FILLER_58_2262 ();
 sg13g2_fill_1 FILLER_58_2300 ();
 sg13g2_decap_8 FILLER_58_2315 ();
 sg13g2_fill_2 FILLER_58_2327 ();
 sg13g2_fill_1 FILLER_58_2329 ();
 sg13g2_fill_1 FILLER_58_2387 ();
 sg13g2_decap_8 FILLER_58_2424 ();
 sg13g2_decap_8 FILLER_58_2431 ();
 sg13g2_fill_1 FILLER_58_2438 ();
 sg13g2_decap_8 FILLER_58_2475 ();
 sg13g2_decap_8 FILLER_58_2482 ();
 sg13g2_decap_8 FILLER_58_2489 ();
 sg13g2_fill_2 FILLER_58_2496 ();
 sg13g2_fill_1 FILLER_58_2498 ();
 sg13g2_decap_8 FILLER_58_2508 ();
 sg13g2_decap_8 FILLER_58_2515 ();
 sg13g2_fill_1 FILLER_58_2522 ();
 sg13g2_fill_2 FILLER_58_2560 ();
 sg13g2_fill_2 FILLER_58_2588 ();
 sg13g2_decap_8 FILLER_58_2622 ();
 sg13g2_decap_8 FILLER_58_2629 ();
 sg13g2_decap_8 FILLER_58_2636 ();
 sg13g2_decap_8 FILLER_58_2643 ();
 sg13g2_fill_2 FILLER_58_2650 ();
 sg13g2_decap_8 FILLER_58_2656 ();
 sg13g2_decap_8 FILLER_58_2663 ();
 sg13g2_decap_4 FILLER_58_2684 ();
 sg13g2_decap_4 FILLER_58_2697 ();
 sg13g2_fill_1 FILLER_58_2701 ();
 sg13g2_fill_1 FILLER_58_2708 ();
 sg13g2_decap_4 FILLER_58_2743 ();
 sg13g2_decap_8 FILLER_58_2778 ();
 sg13g2_decap_8 FILLER_58_2785 ();
 sg13g2_fill_1 FILLER_58_2792 ();
 sg13g2_fill_2 FILLER_58_2797 ();
 sg13g2_fill_1 FILLER_58_2799 ();
 sg13g2_fill_1 FILLER_58_2810 ();
 sg13g2_decap_8 FILLER_58_2843 ();
 sg13g2_fill_2 FILLER_58_2850 ();
 sg13g2_decap_8 FILLER_58_2889 ();
 sg13g2_decap_8 FILLER_58_2896 ();
 sg13g2_decap_8 FILLER_58_2903 ();
 sg13g2_fill_1 FILLER_58_2910 ();
 sg13g2_fill_2 FILLER_58_2942 ();
 sg13g2_decap_8 FILLER_58_2957 ();
 sg13g2_fill_1 FILLER_58_2964 ();
 sg13g2_fill_1 FILLER_58_2992 ();
 sg13g2_decap_8 FILLER_58_3066 ();
 sg13g2_fill_2 FILLER_58_3073 ();
 sg13g2_decap_8 FILLER_58_3106 ();
 sg13g2_decap_8 FILLER_58_3113 ();
 sg13g2_decap_8 FILLER_58_3120 ();
 sg13g2_fill_1 FILLER_58_3127 ();
 sg13g2_decap_8 FILLER_58_3137 ();
 sg13g2_fill_2 FILLER_58_3144 ();
 sg13g2_fill_1 FILLER_58_3146 ();
 sg13g2_decap_8 FILLER_58_3157 ();
 sg13g2_decap_8 FILLER_58_3164 ();
 sg13g2_decap_8 FILLER_58_3171 ();
 sg13g2_decap_8 FILLER_58_3178 ();
 sg13g2_fill_2 FILLER_58_3212 ();
 sg13g2_decap_8 FILLER_58_3241 ();
 sg13g2_decap_8 FILLER_58_3248 ();
 sg13g2_decap_4 FILLER_58_3255 ();
 sg13g2_fill_1 FILLER_58_3277 ();
 sg13g2_fill_1 FILLER_58_3301 ();
 sg13g2_decap_8 FILLER_58_3315 ();
 sg13g2_decap_8 FILLER_58_3353 ();
 sg13g2_decap_8 FILLER_58_3360 ();
 sg13g2_fill_2 FILLER_58_3367 ();
 sg13g2_fill_1 FILLER_58_3369 ();
 sg13g2_fill_1 FILLER_58_3379 ();
 sg13g2_decap_8 FILLER_58_3393 ();
 sg13g2_decap_8 FILLER_58_3405 ();
 sg13g2_decap_8 FILLER_58_3412 ();
 sg13g2_decap_4 FILLER_58_3419 ();
 sg13g2_fill_1 FILLER_58_3423 ();
 sg13g2_decap_8 FILLER_58_3450 ();
 sg13g2_decap_8 FILLER_58_3457 ();
 sg13g2_decap_8 FILLER_58_3464 ();
 sg13g2_decap_4 FILLER_58_3471 ();
 sg13g2_fill_1 FILLER_58_3475 ();
 sg13g2_decap_8 FILLER_58_3503 ();
 sg13g2_decap_8 FILLER_58_3510 ();
 sg13g2_decap_8 FILLER_58_3517 ();
 sg13g2_decap_4 FILLER_58_3524 ();
 sg13g2_fill_1 FILLER_58_3528 ();
 sg13g2_decap_8 FILLER_58_3538 ();
 sg13g2_decap_8 FILLER_58_3545 ();
 sg13g2_decap_8 FILLER_58_3552 ();
 sg13g2_decap_8 FILLER_58_3559 ();
 sg13g2_decap_8 FILLER_58_3566 ();
 sg13g2_decap_4 FILLER_58_3573 ();
 sg13g2_fill_1 FILLER_58_3577 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_4 FILLER_59_39 ();
 sg13g2_decap_8 FILLER_59_74 ();
 sg13g2_decap_8 FILLER_59_81 ();
 sg13g2_fill_1 FILLER_59_88 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_4 FILLER_59_133 ();
 sg13g2_fill_2 FILLER_59_143 ();
 sg13g2_fill_2 FILLER_59_153 ();
 sg13g2_fill_2 FILLER_59_165 ();
 sg13g2_fill_1 FILLER_59_167 ();
 sg13g2_fill_2 FILLER_59_177 ();
 sg13g2_fill_1 FILLER_59_194 ();
 sg13g2_fill_1 FILLER_59_205 ();
 sg13g2_fill_1 FILLER_59_213 ();
 sg13g2_decap_8 FILLER_59_227 ();
 sg13g2_decap_4 FILLER_59_234 ();
 sg13g2_fill_1 FILLER_59_238 ();
 sg13g2_decap_8 FILLER_59_276 ();
 sg13g2_decap_8 FILLER_59_283 ();
 sg13g2_decap_4 FILLER_59_299 ();
 sg13g2_fill_2 FILLER_59_310 ();
 sg13g2_fill_1 FILLER_59_410 ();
 sg13g2_fill_2 FILLER_59_444 ();
 sg13g2_fill_1 FILLER_59_446 ();
 sg13g2_decap_8 FILLER_59_451 ();
 sg13g2_fill_1 FILLER_59_467 ();
 sg13g2_fill_2 FILLER_59_486 ();
 sg13g2_decap_8 FILLER_59_493 ();
 sg13g2_decap_4 FILLER_59_500 ();
 sg13g2_decap_8 FILLER_59_508 ();
 sg13g2_fill_2 FILLER_59_515 ();
 sg13g2_decap_8 FILLER_59_544 ();
 sg13g2_decap_4 FILLER_59_551 ();
 sg13g2_decap_8 FILLER_59_570 ();
 sg13g2_decap_8 FILLER_59_577 ();
 sg13g2_decap_8 FILLER_59_584 ();
 sg13g2_decap_4 FILLER_59_591 ();
 sg13g2_fill_2 FILLER_59_595 ();
 sg13g2_fill_1 FILLER_59_634 ();
 sg13g2_decap_8 FILLER_59_645 ();
 sg13g2_decap_8 FILLER_59_652 ();
 sg13g2_decap_8 FILLER_59_659 ();
 sg13g2_decap_8 FILLER_59_666 ();
 sg13g2_fill_2 FILLER_59_673 ();
 sg13g2_fill_1 FILLER_59_675 ();
 sg13g2_fill_2 FILLER_59_721 ();
 sg13g2_decap_8 FILLER_59_757 ();
 sg13g2_decap_8 FILLER_59_764 ();
 sg13g2_decap_8 FILLER_59_771 ();
 sg13g2_decap_8 FILLER_59_787 ();
 sg13g2_decap_4 FILLER_59_794 ();
 sg13g2_fill_2 FILLER_59_798 ();
 sg13g2_fill_2 FILLER_59_818 ();
 sg13g2_fill_1 FILLER_59_820 ();
 sg13g2_decap_8 FILLER_59_826 ();
 sg13g2_fill_2 FILLER_59_833 ();
 sg13g2_decap_4 FILLER_59_857 ();
 sg13g2_fill_1 FILLER_59_892 ();
 sg13g2_fill_2 FILLER_59_907 ();
 sg13g2_decap_8 FILLER_59_931 ();
 sg13g2_fill_2 FILLER_59_938 ();
 sg13g2_fill_1 FILLER_59_940 ();
 sg13g2_fill_2 FILLER_59_945 ();
 sg13g2_fill_1 FILLER_59_965 ();
 sg13g2_decap_8 FILLER_59_975 ();
 sg13g2_decap_8 FILLER_59_982 ();
 sg13g2_decap_8 FILLER_59_989 ();
 sg13g2_decap_8 FILLER_59_996 ();
 sg13g2_decap_8 FILLER_59_1003 ();
 sg13g2_fill_1 FILLER_59_1010 ();
 sg13g2_fill_2 FILLER_59_1017 ();
 sg13g2_fill_1 FILLER_59_1019 ();
 sg13g2_fill_2 FILLER_59_1029 ();
 sg13g2_fill_1 FILLER_59_1031 ();
 sg13g2_decap_8 FILLER_59_1036 ();
 sg13g2_fill_2 FILLER_59_1043 ();
 sg13g2_fill_1 FILLER_59_1045 ();
 sg13g2_fill_1 FILLER_59_1090 ();
 sg13g2_decap_8 FILLER_59_1094 ();
 sg13g2_decap_8 FILLER_59_1101 ();
 sg13g2_decap_8 FILLER_59_1108 ();
 sg13g2_decap_4 FILLER_59_1115 ();
 sg13g2_fill_1 FILLER_59_1119 ();
 sg13g2_fill_2 FILLER_59_1128 ();
 sg13g2_fill_1 FILLER_59_1130 ();
 sg13g2_fill_1 FILLER_59_1150 ();
 sg13g2_decap_8 FILLER_59_1155 ();
 sg13g2_decap_8 FILLER_59_1162 ();
 sg13g2_decap_8 FILLER_59_1169 ();
 sg13g2_decap_4 FILLER_59_1176 ();
 sg13g2_fill_1 FILLER_59_1180 ();
 sg13g2_fill_2 FILLER_59_1236 ();
 sg13g2_decap_8 FILLER_59_1281 ();
 sg13g2_decap_4 FILLER_59_1288 ();
 sg13g2_decap_8 FILLER_59_1336 ();
 sg13g2_decap_8 FILLER_59_1343 ();
 sg13g2_decap_8 FILLER_59_1350 ();
 sg13g2_decap_4 FILLER_59_1357 ();
 sg13g2_fill_1 FILLER_59_1361 ();
 sg13g2_fill_2 FILLER_59_1375 ();
 sg13g2_fill_1 FILLER_59_1386 ();
 sg13g2_fill_2 FILLER_59_1405 ();
 sg13g2_decap_8 FILLER_59_1442 ();
 sg13g2_decap_4 FILLER_59_1449 ();
 sg13g2_decap_8 FILLER_59_1480 ();
 sg13g2_decap_4 FILLER_59_1487 ();
 sg13g2_fill_2 FILLER_59_1491 ();
 sg13g2_fill_1 FILLER_59_1522 ();
 sg13g2_decap_4 FILLER_59_1541 ();
 sg13g2_fill_1 FILLER_59_1545 ();
 sg13g2_fill_1 FILLER_59_1569 ();
 sg13g2_decap_8 FILLER_59_1584 ();
 sg13g2_decap_8 FILLER_59_1591 ();
 sg13g2_decap_8 FILLER_59_1598 ();
 sg13g2_decap_8 FILLER_59_1605 ();
 sg13g2_decap_8 FILLER_59_1612 ();
 sg13g2_decap_4 FILLER_59_1619 ();
 sg13g2_fill_2 FILLER_59_1623 ();
 sg13g2_decap_8 FILLER_59_1657 ();
 sg13g2_fill_2 FILLER_59_1664 ();
 sg13g2_fill_1 FILLER_59_1666 ();
 sg13g2_fill_2 FILLER_59_1700 ();
 sg13g2_decap_8 FILLER_59_1708 ();
 sg13g2_decap_4 FILLER_59_1715 ();
 sg13g2_fill_1 FILLER_59_1719 ();
 sg13g2_decap_8 FILLER_59_1768 ();
 sg13g2_decap_8 FILLER_59_1775 ();
 sg13g2_fill_2 FILLER_59_1782 ();
 sg13g2_decap_8 FILLER_59_1818 ();
 sg13g2_fill_2 FILLER_59_1825 ();
 sg13g2_fill_1 FILLER_59_1827 ();
 sg13g2_fill_2 FILLER_59_1860 ();
 sg13g2_fill_1 FILLER_59_1862 ();
 sg13g2_fill_2 FILLER_59_1876 ();
 sg13g2_fill_1 FILLER_59_1878 ();
 sg13g2_decap_8 FILLER_59_1907 ();
 sg13g2_fill_1 FILLER_59_1936 ();
 sg13g2_fill_2 FILLER_59_1959 ();
 sg13g2_decap_8 FILLER_59_2006 ();
 sg13g2_decap_8 FILLER_59_2013 ();
 sg13g2_fill_2 FILLER_59_2020 ();
 sg13g2_decap_8 FILLER_59_2032 ();
 sg13g2_decap_8 FILLER_59_2039 ();
 sg13g2_decap_8 FILLER_59_2046 ();
 sg13g2_decap_8 FILLER_59_2053 ();
 sg13g2_decap_8 FILLER_59_2060 ();
 sg13g2_decap_8 FILLER_59_2083 ();
 sg13g2_decap_8 FILLER_59_2090 ();
 sg13g2_decap_8 FILLER_59_2097 ();
 sg13g2_decap_8 FILLER_59_2104 ();
 sg13g2_decap_8 FILLER_59_2111 ();
 sg13g2_decap_8 FILLER_59_2118 ();
 sg13g2_decap_4 FILLER_59_2125 ();
 sg13g2_decap_8 FILLER_59_2134 ();
 sg13g2_decap_8 FILLER_59_2141 ();
 sg13g2_decap_8 FILLER_59_2148 ();
 sg13g2_decap_8 FILLER_59_2155 ();
 sg13g2_decap_8 FILLER_59_2162 ();
 sg13g2_fill_2 FILLER_59_2169 ();
 sg13g2_fill_1 FILLER_59_2171 ();
 sg13g2_decap_8 FILLER_59_2193 ();
 sg13g2_decap_8 FILLER_59_2200 ();
 sg13g2_fill_2 FILLER_59_2207 ();
 sg13g2_decap_8 FILLER_59_2234 ();
 sg13g2_decap_8 FILLER_59_2241 ();
 sg13g2_decap_4 FILLER_59_2248 ();
 sg13g2_fill_2 FILLER_59_2252 ();
 sg13g2_decap_4 FILLER_59_2267 ();
 sg13g2_fill_1 FILLER_59_2271 ();
 sg13g2_fill_2 FILLER_59_2281 ();
 sg13g2_fill_1 FILLER_59_2283 ();
 sg13g2_fill_2 FILLER_59_2297 ();
 sg13g2_fill_1 FILLER_59_2299 ();
 sg13g2_fill_1 FILLER_59_2309 ();
 sg13g2_decap_8 FILLER_59_2323 ();
 sg13g2_fill_1 FILLER_59_2330 ();
 sg13g2_decap_8 FILLER_59_2381 ();
 sg13g2_fill_2 FILLER_59_2388 ();
 sg13g2_fill_1 FILLER_59_2394 ();
 sg13g2_decap_4 FILLER_59_2408 ();
 sg13g2_decap_4 FILLER_59_2426 ();
 sg13g2_fill_2 FILLER_59_2430 ();
 sg13g2_decap_8 FILLER_59_2468 ();
 sg13g2_decap_8 FILLER_59_2475 ();
 sg13g2_decap_8 FILLER_59_2482 ();
 sg13g2_decap_8 FILLER_59_2489 ();
 sg13g2_decap_8 FILLER_59_2496 ();
 sg13g2_fill_2 FILLER_59_2523 ();
 sg13g2_fill_1 FILLER_59_2525 ();
 sg13g2_decap_8 FILLER_59_2539 ();
 sg13g2_fill_1 FILLER_59_2546 ();
 sg13g2_decap_8 FILLER_59_2593 ();
 sg13g2_decap_8 FILLER_59_2600 ();
 sg13g2_decap_4 FILLER_59_2607 ();
 sg13g2_fill_2 FILLER_59_2611 ();
 sg13g2_decap_8 FILLER_59_2622 ();
 sg13g2_decap_8 FILLER_59_2629 ();
 sg13g2_fill_1 FILLER_59_2636 ();
 sg13g2_decap_8 FILLER_59_2701 ();
 sg13g2_fill_2 FILLER_59_2708 ();
 sg13g2_fill_1 FILLER_59_2710 ();
 sg13g2_fill_2 FILLER_59_2724 ();
 sg13g2_fill_2 FILLER_59_2748 ();
 sg13g2_fill_1 FILLER_59_2750 ();
 sg13g2_fill_2 FILLER_59_2786 ();
 sg13g2_decap_4 FILLER_59_2855 ();
 sg13g2_decap_8 FILLER_59_2885 ();
 sg13g2_decap_8 FILLER_59_2892 ();
 sg13g2_decap_4 FILLER_59_2899 ();
 sg13g2_decap_8 FILLER_59_2961 ();
 sg13g2_fill_1 FILLER_59_2968 ();
 sg13g2_fill_2 FILLER_59_3019 ();
 sg13g2_fill_1 FILLER_59_3021 ();
 sg13g2_decap_8 FILLER_59_3052 ();
 sg13g2_fill_2 FILLER_59_3059 ();
 sg13g2_fill_1 FILLER_59_3061 ();
 sg13g2_decap_8 FILLER_59_3099 ();
 sg13g2_decap_8 FILLER_59_3106 ();
 sg13g2_decap_8 FILLER_59_3113 ();
 sg13g2_decap_8 FILLER_59_3177 ();
 sg13g2_decap_4 FILLER_59_3184 ();
 sg13g2_fill_2 FILLER_59_3188 ();
 sg13g2_fill_2 FILLER_59_3194 ();
 sg13g2_fill_1 FILLER_59_3196 ();
 sg13g2_decap_8 FILLER_59_3238 ();
 sg13g2_decap_8 FILLER_59_3245 ();
 sg13g2_decap_8 FILLER_59_3252 ();
 sg13g2_decap_8 FILLER_59_3259 ();
 sg13g2_decap_4 FILLER_59_3266 ();
 sg13g2_fill_1 FILLER_59_3270 ();
 sg13g2_decap_8 FILLER_59_3307 ();
 sg13g2_decap_8 FILLER_59_3314 ();
 sg13g2_decap_8 FILLER_59_3321 ();
 sg13g2_fill_2 FILLER_59_3328 ();
 sg13g2_fill_1 FILLER_59_3330 ();
 sg13g2_fill_2 FILLER_59_3345 ();
 sg13g2_fill_1 FILLER_59_3347 ();
 sg13g2_decap_8 FILLER_59_3357 ();
 sg13g2_fill_2 FILLER_59_3364 ();
 sg13g2_decap_4 FILLER_59_3396 ();
 sg13g2_fill_2 FILLER_59_3400 ();
 sg13g2_decap_8 FILLER_59_3415 ();
 sg13g2_decap_4 FILLER_59_3453 ();
 sg13g2_decap_8 FILLER_59_3503 ();
 sg13g2_fill_2 FILLER_59_3510 ();
 sg13g2_fill_1 FILLER_59_3512 ();
 sg13g2_decap_8 FILLER_59_3549 ();
 sg13g2_decap_8 FILLER_59_3556 ();
 sg13g2_decap_8 FILLER_59_3563 ();
 sg13g2_decap_8 FILLER_59_3570 ();
 sg13g2_fill_1 FILLER_59_3577 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_11 ();
 sg13g2_fill_1 FILLER_60_48 ();
 sg13g2_decap_8 FILLER_60_80 ();
 sg13g2_fill_2 FILLER_60_87 ();
 sg13g2_decap_8 FILLER_60_130 ();
 sg13g2_decap_8 FILLER_60_137 ();
 sg13g2_decap_8 FILLER_60_144 ();
 sg13g2_decap_4 FILLER_60_151 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_fill_1 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_221 ();
 sg13g2_decap_4 FILLER_60_228 ();
 sg13g2_fill_1 FILLER_60_232 ();
 sg13g2_decap_8 FILLER_60_279 ();
 sg13g2_decap_4 FILLER_60_286 ();
 sg13g2_fill_1 FILLER_60_309 ();
 sg13g2_fill_2 FILLER_60_318 ();
 sg13g2_fill_1 FILLER_60_343 ();
 sg13g2_fill_1 FILLER_60_372 ();
 sg13g2_fill_1 FILLER_60_398 ();
 sg13g2_fill_1 FILLER_60_460 ();
 sg13g2_decap_4 FILLER_60_464 ();
 sg13g2_fill_1 FILLER_60_468 ();
 sg13g2_fill_1 FILLER_60_473 ();
 sg13g2_decap_8 FILLER_60_504 ();
 sg13g2_fill_1 FILLER_60_511 ();
 sg13g2_decap_8 FILLER_60_576 ();
 sg13g2_decap_4 FILLER_60_595 ();
 sg13g2_decap_8 FILLER_60_640 ();
 sg13g2_decap_8 FILLER_60_647 ();
 sg13g2_decap_8 FILLER_60_654 ();
 sg13g2_decap_8 FILLER_60_665 ();
 sg13g2_fill_1 FILLER_60_672 ();
 sg13g2_fill_2 FILLER_60_683 ();
 sg13g2_fill_1 FILLER_60_694 ();
 sg13g2_fill_1 FILLER_60_704 ();
 sg13g2_fill_1 FILLER_60_715 ();
 sg13g2_decap_4 FILLER_60_753 ();
 sg13g2_fill_1 FILLER_60_757 ();
 sg13g2_decap_8 FILLER_60_796 ();
 sg13g2_decap_8 FILLER_60_803 ();
 sg13g2_decap_8 FILLER_60_810 ();
 sg13g2_decap_8 FILLER_60_821 ();
 sg13g2_decap_8 FILLER_60_828 ();
 sg13g2_fill_2 FILLER_60_835 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_8 FILLER_60_925 ();
 sg13g2_decap_8 FILLER_60_932 ();
 sg13g2_decap_8 FILLER_60_939 ();
 sg13g2_fill_2 FILLER_60_946 ();
 sg13g2_fill_1 FILLER_60_948 ();
 sg13g2_fill_1 FILLER_60_952 ();
 sg13g2_fill_2 FILLER_60_958 ();
 sg13g2_decap_8 FILLER_60_984 ();
 sg13g2_decap_8 FILLER_60_991 ();
 sg13g2_decap_4 FILLER_60_998 ();
 sg13g2_fill_2 FILLER_60_1002 ();
 sg13g2_decap_8 FILLER_60_1008 ();
 sg13g2_decap_8 FILLER_60_1015 ();
 sg13g2_decap_8 FILLER_60_1028 ();
 sg13g2_fill_2 FILLER_60_1035 ();
 sg13g2_fill_1 FILLER_60_1037 ();
 sg13g2_fill_2 FILLER_60_1043 ();
 sg13g2_fill_1 FILLER_60_1045 ();
 sg13g2_fill_1 FILLER_60_1061 ();
 sg13g2_fill_2 FILLER_60_1075 ();
 sg13g2_decap_4 FILLER_60_1080 ();
 sg13g2_fill_2 FILLER_60_1084 ();
 sg13g2_fill_2 FILLER_60_1091 ();
 sg13g2_decap_8 FILLER_60_1101 ();
 sg13g2_fill_1 FILLER_60_1108 ();
 sg13g2_decap_8 FILLER_60_1118 ();
 sg13g2_fill_2 FILLER_60_1143 ();
 sg13g2_fill_1 FILLER_60_1145 ();
 sg13g2_fill_1 FILLER_60_1156 ();
 sg13g2_decap_8 FILLER_60_1162 ();
 sg13g2_decap_8 FILLER_60_1169 ();
 sg13g2_fill_2 FILLER_60_1176 ();
 sg13g2_fill_1 FILLER_60_1206 ();
 sg13g2_fill_1 FILLER_60_1216 ();
 sg13g2_decap_8 FILLER_60_1277 ();
 sg13g2_decap_8 FILLER_60_1284 ();
 sg13g2_decap_8 FILLER_60_1291 ();
 sg13g2_fill_2 FILLER_60_1298 ();
 sg13g2_fill_1 FILLER_60_1300 ();
 sg13g2_decap_8 FILLER_60_1329 ();
 sg13g2_decap_8 FILLER_60_1336 ();
 sg13g2_decap_8 FILLER_60_1343 ();
 sg13g2_decap_8 FILLER_60_1350 ();
 sg13g2_fill_2 FILLER_60_1357 ();
 sg13g2_fill_1 FILLER_60_1359 ();
 sg13g2_decap_8 FILLER_60_1363 ();
 sg13g2_fill_2 FILLER_60_1370 ();
 sg13g2_fill_1 FILLER_60_1372 ();
 sg13g2_decap_8 FILLER_60_1404 ();
 sg13g2_fill_2 FILLER_60_1447 ();
 sg13g2_fill_2 FILLER_60_1458 ();
 sg13g2_decap_4 FILLER_60_1464 ();
 sg13g2_fill_1 FILLER_60_1474 ();
 sg13g2_fill_2 FILLER_60_1487 ();
 sg13g2_fill_1 FILLER_60_1489 ();
 sg13g2_fill_2 FILLER_60_1521 ();
 sg13g2_fill_1 FILLER_60_1523 ();
 sg13g2_fill_1 FILLER_60_1529 ();
 sg13g2_fill_1 FILLER_60_1543 ();
 sg13g2_fill_2 FILLER_60_1557 ();
 sg13g2_fill_1 FILLER_60_1559 ();
 sg13g2_fill_2 FILLER_60_1601 ();
 sg13g2_decap_4 FILLER_60_1608 ();
 sg13g2_decap_8 FILLER_60_1664 ();
 sg13g2_fill_2 FILLER_60_1671 ();
 sg13g2_decap_4 FILLER_60_1692 ();
 sg13g2_fill_2 FILLER_60_1701 ();
 sg13g2_fill_2 FILLER_60_1709 ();
 sg13g2_fill_1 FILLER_60_1711 ();
 sg13g2_fill_1 FILLER_60_1716 ();
 sg13g2_fill_2 FILLER_60_1722 ();
 sg13g2_fill_1 FILLER_60_1742 ();
 sg13g2_decap_4 FILLER_60_1771 ();
 sg13g2_fill_2 FILLER_60_1775 ();
 sg13g2_fill_1 FILLER_60_1793 ();
 sg13g2_fill_2 FILLER_60_1807 ();
 sg13g2_fill_1 FILLER_60_1809 ();
 sg13g2_decap_8 FILLER_60_1821 ();
 sg13g2_decap_8 FILLER_60_1828 ();
 sg13g2_decap_8 FILLER_60_1835 ();
 sg13g2_decap_8 FILLER_60_1842 ();
 sg13g2_fill_2 FILLER_60_1849 ();
 sg13g2_fill_1 FILLER_60_1851 ();
 sg13g2_decap_8 FILLER_60_1858 ();
 sg13g2_fill_1 FILLER_60_1865 ();
 sg13g2_fill_1 FILLER_60_1875 ();
 sg13g2_decap_8 FILLER_60_1898 ();
 sg13g2_fill_2 FILLER_60_1905 ();
 sg13g2_decap_4 FILLER_60_1916 ();
 sg13g2_fill_2 FILLER_60_1920 ();
 sg13g2_decap_8 FILLER_60_1935 ();
 sg13g2_fill_2 FILLER_60_1942 ();
 sg13g2_decap_8 FILLER_60_1977 ();
 sg13g2_decap_8 FILLER_60_1984 ();
 sg13g2_fill_2 FILLER_60_1991 ();
 sg13g2_fill_1 FILLER_60_1993 ();
 sg13g2_decap_8 FILLER_60_2003 ();
 sg13g2_fill_2 FILLER_60_2010 ();
 sg13g2_decap_8 FILLER_60_2043 ();
 sg13g2_decap_8 FILLER_60_2050 ();
 sg13g2_decap_8 FILLER_60_2057 ();
 sg13g2_fill_1 FILLER_60_2064 ();
 sg13g2_decap_8 FILLER_60_2070 ();
 sg13g2_decap_8 FILLER_60_2077 ();
 sg13g2_decap_4 FILLER_60_2084 ();
 sg13g2_fill_2 FILLER_60_2088 ();
 sg13g2_decap_8 FILLER_60_2095 ();
 sg13g2_decap_8 FILLER_60_2102 ();
 sg13g2_decap_8 FILLER_60_2109 ();
 sg13g2_fill_1 FILLER_60_2116 ();
 sg13g2_decap_8 FILLER_60_2139 ();
 sg13g2_decap_4 FILLER_60_2146 ();
 sg13g2_decap_8 FILLER_60_2158 ();
 sg13g2_fill_2 FILLER_60_2165 ();
 sg13g2_decap_8 FILLER_60_2175 ();
 sg13g2_decap_8 FILLER_60_2182 ();
 sg13g2_decap_8 FILLER_60_2189 ();
 sg13g2_decap_8 FILLER_60_2196 ();
 sg13g2_fill_1 FILLER_60_2203 ();
 sg13g2_decap_4 FILLER_60_2223 ();
 sg13g2_decap_8 FILLER_60_2240 ();
 sg13g2_decap_8 FILLER_60_2247 ();
 sg13g2_decap_8 FILLER_60_2254 ();
 sg13g2_decap_8 FILLER_60_2261 ();
 sg13g2_decap_8 FILLER_60_2268 ();
 sg13g2_decap_8 FILLER_60_2275 ();
 sg13g2_fill_2 FILLER_60_2282 ();
 sg13g2_fill_1 FILLER_60_2284 ();
 sg13g2_decap_8 FILLER_60_2289 ();
 sg13g2_decap_8 FILLER_60_2296 ();
 sg13g2_decap_4 FILLER_60_2303 ();
 sg13g2_fill_1 FILLER_60_2307 ();
 sg13g2_decap_8 FILLER_60_2325 ();
 sg13g2_decap_8 FILLER_60_2332 ();
 sg13g2_decap_4 FILLER_60_2339 ();
 sg13g2_fill_1 FILLER_60_2343 ();
 sg13g2_fill_2 FILLER_60_2349 ();
 sg13g2_decap_8 FILLER_60_2355 ();
 sg13g2_fill_1 FILLER_60_2362 ();
 sg13g2_decap_4 FILLER_60_2376 ();
 sg13g2_decap_4 FILLER_60_2393 ();
 sg13g2_fill_2 FILLER_60_2397 ();
 sg13g2_decap_8 FILLER_60_2408 ();
 sg13g2_decap_8 FILLER_60_2415 ();
 sg13g2_fill_2 FILLER_60_2422 ();
 sg13g2_decap_8 FILLER_60_2482 ();
 sg13g2_decap_4 FILLER_60_2489 ();
 sg13g2_fill_2 FILLER_60_2493 ();
 sg13g2_decap_4 FILLER_60_2545 ();
 sg13g2_fill_1 FILLER_60_2549 ();
 sg13g2_decap_8 FILLER_60_2592 ();
 sg13g2_decap_8 FILLER_60_2599 ();
 sg13g2_decap_8 FILLER_60_2627 ();
 sg13g2_decap_8 FILLER_60_2634 ();
 sg13g2_decap_8 FILLER_60_2641 ();
 sg13g2_decap_8 FILLER_60_2648 ();
 sg13g2_fill_2 FILLER_60_2655 ();
 sg13g2_decap_4 FILLER_60_2666 ();
 sg13g2_decap_8 FILLER_60_2691 ();
 sg13g2_decap_8 FILLER_60_2698 ();
 sg13g2_decap_8 FILLER_60_2705 ();
 sg13g2_decap_8 FILLER_60_2712 ();
 sg13g2_decap_4 FILLER_60_2719 ();
 sg13g2_decap_8 FILLER_60_2744 ();
 sg13g2_decap_4 FILLER_60_2751 ();
 sg13g2_fill_1 FILLER_60_2768 ();
 sg13g2_decap_4 FILLER_60_2795 ();
 sg13g2_fill_1 FILLER_60_2822 ();
 sg13g2_decap_8 FILLER_60_2841 ();
 sg13g2_decap_4 FILLER_60_2848 ();
 sg13g2_fill_2 FILLER_60_2852 ();
 sg13g2_decap_8 FILLER_60_2881 ();
 sg13g2_decap_8 FILLER_60_2888 ();
 sg13g2_decap_8 FILLER_60_2895 ();
 sg13g2_decap_8 FILLER_60_2902 ();
 sg13g2_decap_8 FILLER_60_2960 ();
 sg13g2_decap_8 FILLER_60_2967 ();
 sg13g2_decap_8 FILLER_60_2974 ();
 sg13g2_fill_2 FILLER_60_2981 ();
 sg13g2_decap_8 FILLER_60_3023 ();
 sg13g2_decap_8 FILLER_60_3030 ();
 sg13g2_decap_4 FILLER_60_3037 ();
 sg13g2_fill_2 FILLER_60_3041 ();
 sg13g2_decap_8 FILLER_60_3047 ();
 sg13g2_decap_8 FILLER_60_3054 ();
 sg13g2_fill_2 FILLER_60_3061 ();
 sg13g2_decap_8 FILLER_60_3104 ();
 sg13g2_fill_1 FILLER_60_3111 ();
 sg13g2_fill_2 FILLER_60_3149 ();
 sg13g2_decap_8 FILLER_60_3182 ();
 sg13g2_decap_8 FILLER_60_3235 ();
 sg13g2_decap_8 FILLER_60_3242 ();
 sg13g2_decap_8 FILLER_60_3249 ();
 sg13g2_fill_2 FILLER_60_3275 ();
 sg13g2_decap_8 FILLER_60_3299 ();
 sg13g2_decap_8 FILLER_60_3306 ();
 sg13g2_decap_8 FILLER_60_3313 ();
 sg13g2_fill_1 FILLER_60_3320 ();
 sg13g2_fill_2 FILLER_60_3334 ();
 sg13g2_fill_1 FILLER_60_3336 ();
 sg13g2_decap_4 FILLER_60_3347 ();
 sg13g2_fill_2 FILLER_60_3351 ();
 sg13g2_decap_4 FILLER_60_3363 ();
 sg13g2_decap_8 FILLER_60_3398 ();
 sg13g2_decap_8 FILLER_60_3405 ();
 sg13g2_fill_1 FILLER_60_3412 ();
 sg13g2_fill_2 FILLER_60_3469 ();
 sg13g2_decap_8 FILLER_60_3494 ();
 sg13g2_decap_8 FILLER_60_3501 ();
 sg13g2_decap_4 FILLER_60_3508 ();
 sg13g2_fill_2 FILLER_60_3512 ();
 sg13g2_fill_2 FILLER_60_3528 ();
 sg13g2_decap_8 FILLER_60_3567 ();
 sg13g2_decap_4 FILLER_60_3574 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_decap_4 FILLER_61_62 ();
 sg13g2_fill_2 FILLER_61_66 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_fill_1 FILLER_61_101 ();
 sg13g2_decap_4 FILLER_61_117 ();
 sg13g2_decap_8 FILLER_61_130 ();
 sg13g2_decap_4 FILLER_61_137 ();
 sg13g2_fill_2 FILLER_61_141 ();
 sg13g2_fill_1 FILLER_61_179 ();
 sg13g2_decap_8 FILLER_61_216 ();
 sg13g2_fill_2 FILLER_61_223 ();
 sg13g2_fill_1 FILLER_61_283 ();
 sg13g2_decap_8 FILLER_61_332 ();
 sg13g2_decap_8 FILLER_61_339 ();
 sg13g2_fill_1 FILLER_61_346 ();
 sg13g2_fill_2 FILLER_61_405 ();
 sg13g2_fill_1 FILLER_61_453 ();
 sg13g2_fill_2 FILLER_61_503 ();
 sg13g2_fill_1 FILLER_61_505 ();
 sg13g2_fill_1 FILLER_61_524 ();
 sg13g2_fill_1 FILLER_61_559 ();
 sg13g2_fill_1 FILLER_61_590 ();
 sg13g2_decap_8 FILLER_61_635 ();
 sg13g2_decap_8 FILLER_61_642 ();
 sg13g2_fill_2 FILLER_61_694 ();
 sg13g2_fill_1 FILLER_61_696 ();
 sg13g2_fill_2 FILLER_61_707 ();
 sg13g2_fill_1 FILLER_61_709 ();
 sg13g2_fill_1 FILLER_61_718 ();
 sg13g2_fill_2 FILLER_61_737 ();
 sg13g2_decap_8 FILLER_61_744 ();
 sg13g2_decap_8 FILLER_61_751 ();
 sg13g2_decap_8 FILLER_61_796 ();
 sg13g2_decap_8 FILLER_61_803 ();
 sg13g2_decap_8 FILLER_61_810 ();
 sg13g2_decap_4 FILLER_61_817 ();
 sg13g2_fill_2 FILLER_61_821 ();
 sg13g2_fill_1 FILLER_61_842 ();
 sg13g2_fill_1 FILLER_61_875 ();
 sg13g2_decap_8 FILLER_61_942 ();
 sg13g2_decap_8 FILLER_61_949 ();
 sg13g2_decap_4 FILLER_61_956 ();
 sg13g2_fill_1 FILLER_61_964 ();
 sg13g2_decap_8 FILLER_61_1014 ();
 sg13g2_fill_2 FILLER_61_1021 ();
 sg13g2_decap_4 FILLER_61_1036 ();
 sg13g2_fill_1 FILLER_61_1040 ();
 sg13g2_fill_1 FILLER_61_1069 ();
 sg13g2_fill_2 FILLER_61_1086 ();
 sg13g2_fill_1 FILLER_61_1088 ();
 sg13g2_decap_8 FILLER_61_1109 ();
 sg13g2_decap_4 FILLER_61_1116 ();
 sg13g2_fill_1 FILLER_61_1120 ();
 sg13g2_fill_2 FILLER_61_1147 ();
 sg13g2_fill_1 FILLER_61_1149 ();
 sg13g2_decap_8 FILLER_61_1163 ();
 sg13g2_decap_8 FILLER_61_1170 ();
 sg13g2_decap_8 FILLER_61_1177 ();
 sg13g2_fill_2 FILLER_61_1238 ();
 sg13g2_decap_8 FILLER_61_1276 ();
 sg13g2_decap_8 FILLER_61_1283 ();
 sg13g2_decap_8 FILLER_61_1290 ();
 sg13g2_decap_4 FILLER_61_1297 ();
 sg13g2_fill_2 FILLER_61_1324 ();
 sg13g2_decap_8 FILLER_61_1336 ();
 sg13g2_decap_8 FILLER_61_1343 ();
 sg13g2_fill_2 FILLER_61_1350 ();
 sg13g2_decap_8 FILLER_61_1411 ();
 sg13g2_decap_8 FILLER_61_1418 ();
 sg13g2_decap_4 FILLER_61_1425 ();
 sg13g2_fill_1 FILLER_61_1438 ();
 sg13g2_fill_2 FILLER_61_1447 ();
 sg13g2_fill_2 FILLER_61_1475 ();
 sg13g2_decap_8 FILLER_61_1491 ();
 sg13g2_fill_1 FILLER_61_1498 ();
 sg13g2_fill_2 FILLER_61_1505 ();
 sg13g2_fill_1 FILLER_61_1507 ();
 sg13g2_fill_1 FILLER_61_1513 ();
 sg13g2_decap_8 FILLER_61_1521 ();
 sg13g2_fill_2 FILLER_61_1528 ();
 sg13g2_fill_1 FILLER_61_1530 ();
 sg13g2_fill_2 FILLER_61_1549 ();
 sg13g2_fill_1 FILLER_61_1551 ();
 sg13g2_decap_4 FILLER_61_1557 ();
 sg13g2_fill_1 FILLER_61_1561 ();
 sg13g2_fill_1 FILLER_61_1633 ();
 sg13g2_decap_8 FILLER_61_1656 ();
 sg13g2_decap_8 FILLER_61_1663 ();
 sg13g2_decap_4 FILLER_61_1670 ();
 sg13g2_decap_4 FILLER_61_1702 ();
 sg13g2_fill_1 FILLER_61_1706 ();
 sg13g2_decap_4 FILLER_61_1725 ();
 sg13g2_fill_1 FILLER_61_1729 ();
 sg13g2_decap_8 FILLER_61_1743 ();
 sg13g2_decap_4 FILLER_61_1750 ();
 sg13g2_fill_2 FILLER_61_1763 ();
 sg13g2_fill_2 FILLER_61_1775 ();
 sg13g2_fill_1 FILLER_61_1777 ();
 sg13g2_fill_2 FILLER_61_1788 ();
 sg13g2_fill_1 FILLER_61_1790 ();
 sg13g2_fill_2 FILLER_61_1806 ();
 sg13g2_fill_1 FILLER_61_1808 ();
 sg13g2_decap_8 FILLER_61_1827 ();
 sg13g2_decap_8 FILLER_61_1834 ();
 sg13g2_decap_8 FILLER_61_1841 ();
 sg13g2_decap_8 FILLER_61_1848 ();
 sg13g2_decap_4 FILLER_61_1855 ();
 sg13g2_decap_8 FILLER_61_1895 ();
 sg13g2_fill_2 FILLER_61_1902 ();
 sg13g2_decap_8 FILLER_61_1912 ();
 sg13g2_fill_2 FILLER_61_1919 ();
 sg13g2_fill_1 FILLER_61_1921 ();
 sg13g2_decap_8 FILLER_61_1943 ();
 sg13g2_fill_1 FILLER_61_1950 ();
 sg13g2_fill_1 FILLER_61_1959 ();
 sg13g2_decap_8 FILLER_61_1964 ();
 sg13g2_decap_8 FILLER_61_1971 ();
 sg13g2_decap_8 FILLER_61_1978 ();
 sg13g2_decap_8 FILLER_61_1985 ();
 sg13g2_decap_8 FILLER_61_1992 ();
 sg13g2_fill_1 FILLER_61_1999 ();
 sg13g2_fill_1 FILLER_61_2007 ();
 sg13g2_decap_8 FILLER_61_2054 ();
 sg13g2_decap_8 FILLER_61_2061 ();
 sg13g2_decap_8 FILLER_61_2068 ();
 sg13g2_decap_4 FILLER_61_2075 ();
 sg13g2_fill_2 FILLER_61_2079 ();
 sg13g2_fill_2 FILLER_61_2091 ();
 sg13g2_fill_1 FILLER_61_2093 ();
 sg13g2_decap_4 FILLER_61_2102 ();
 sg13g2_fill_2 FILLER_61_2106 ();
 sg13g2_fill_2 FILLER_61_2113 ();
 sg13g2_fill_1 FILLER_61_2115 ();
 sg13g2_fill_1 FILLER_61_2132 ();
 sg13g2_decap_8 FILLER_61_2146 ();
 sg13g2_decap_8 FILLER_61_2153 ();
 sg13g2_decap_8 FILLER_61_2160 ();
 sg13g2_decap_8 FILLER_61_2167 ();
 sg13g2_decap_8 FILLER_61_2174 ();
 sg13g2_decap_8 FILLER_61_2181 ();
 sg13g2_decap_4 FILLER_61_2188 ();
 sg13g2_fill_2 FILLER_61_2205 ();
 sg13g2_decap_8 FILLER_61_2225 ();
 sg13g2_fill_1 FILLER_61_2232 ();
 sg13g2_decap_8 FILLER_61_2246 ();
 sg13g2_decap_8 FILLER_61_2253 ();
 sg13g2_fill_2 FILLER_61_2260 ();
 sg13g2_fill_1 FILLER_61_2262 ();
 sg13g2_fill_1 FILLER_61_2267 ();
 sg13g2_decap_4 FILLER_61_2281 ();
 sg13g2_fill_1 FILLER_61_2285 ();
 sg13g2_decap_4 FILLER_61_2299 ();
 sg13g2_decap_8 FILLER_61_2316 ();
 sg13g2_decap_8 FILLER_61_2323 ();
 sg13g2_decap_8 FILLER_61_2330 ();
 sg13g2_decap_8 FILLER_61_2337 ();
 sg13g2_decap_8 FILLER_61_2344 ();
 sg13g2_decap_8 FILLER_61_2351 ();
 sg13g2_decap_4 FILLER_61_2358 ();
 sg13g2_decap_8 FILLER_61_2405 ();
 sg13g2_decap_8 FILLER_61_2412 ();
 sg13g2_decap_8 FILLER_61_2419 ();
 sg13g2_fill_2 FILLER_61_2426 ();
 sg13g2_fill_1 FILLER_61_2428 ();
 sg13g2_fill_2 FILLER_61_2460 ();
 sg13g2_decap_4 FILLER_61_2475 ();
 sg13g2_fill_2 FILLER_61_2479 ();
 sg13g2_fill_2 FILLER_61_2508 ();
 sg13g2_decap_8 FILLER_61_2540 ();
 sg13g2_decap_8 FILLER_61_2547 ();
 sg13g2_fill_1 FILLER_61_2554 ();
 sg13g2_fill_1 FILLER_61_2559 ();
 sg13g2_fill_2 FILLER_61_2570 ();
 sg13g2_decap_8 FILLER_61_2581 ();
 sg13g2_decap_8 FILLER_61_2588 ();
 sg13g2_fill_2 FILLER_61_2599 ();
 sg13g2_decap_8 FILLER_61_2638 ();
 sg13g2_decap_8 FILLER_61_2645 ();
 sg13g2_decap_8 FILLER_61_2652 ();
 sg13g2_decap_8 FILLER_61_2686 ();
 sg13g2_decap_8 FILLER_61_2693 ();
 sg13g2_decap_8 FILLER_61_2700 ();
 sg13g2_fill_2 FILLER_61_2707 ();
 sg13g2_fill_1 FILLER_61_2709 ();
 sg13g2_decap_8 FILLER_61_2741 ();
 sg13g2_fill_2 FILLER_61_2748 ();
 sg13g2_fill_1 FILLER_61_2750 ();
 sg13g2_decap_8 FILLER_61_2759 ();
 sg13g2_decap_4 FILLER_61_2771 ();
 sg13g2_fill_2 FILLER_61_2775 ();
 sg13g2_decap_8 FILLER_61_2782 ();
 sg13g2_decap_8 FILLER_61_2789 ();
 sg13g2_fill_2 FILLER_61_2796 ();
 sg13g2_fill_1 FILLER_61_2798 ();
 sg13g2_fill_2 FILLER_61_2820 ();
 sg13g2_decap_8 FILLER_61_2826 ();
 sg13g2_decap_8 FILLER_61_2833 ();
 sg13g2_decap_4 FILLER_61_2840 ();
 sg13g2_fill_1 FILLER_61_2844 ();
 sg13g2_decap_8 FILLER_61_2849 ();
 sg13g2_decap_8 FILLER_61_2887 ();
 sg13g2_decap_8 FILLER_61_2894 ();
 sg13g2_decap_8 FILLER_61_2901 ();
 sg13g2_decap_4 FILLER_61_2908 ();
 sg13g2_fill_2 FILLER_61_2912 ();
 sg13g2_decap_8 FILLER_61_2960 ();
 sg13g2_decap_8 FILLER_61_2967 ();
 sg13g2_decap_8 FILLER_61_2974 ();
 sg13g2_decap_4 FILLER_61_2981 ();
 sg13g2_fill_2 FILLER_61_2985 ();
 sg13g2_fill_2 FILLER_61_2992 ();
 sg13g2_fill_1 FILLER_61_2994 ();
 sg13g2_fill_2 FILLER_61_3014 ();
 sg13g2_decap_8 FILLER_61_3050 ();
 sg13g2_decap_8 FILLER_61_3057 ();
 sg13g2_fill_1 FILLER_61_3064 ();
 sg13g2_fill_2 FILLER_61_3115 ();
 sg13g2_fill_1 FILLER_61_3117 ();
 sg13g2_decap_8 FILLER_61_3167 ();
 sg13g2_decap_8 FILLER_61_3174 ();
 sg13g2_decap_8 FILLER_61_3181 ();
 sg13g2_decap_8 FILLER_61_3188 ();
 sg13g2_decap_4 FILLER_61_3195 ();
 sg13g2_fill_1 FILLER_61_3199 ();
 sg13g2_decap_8 FILLER_61_3231 ();
 sg13g2_fill_1 FILLER_61_3238 ();
 sg13g2_fill_2 FILLER_61_3276 ();
 sg13g2_decap_4 FILLER_61_3295 ();
 sg13g2_fill_1 FILLER_61_3299 ();
 sg13g2_fill_1 FILLER_61_3327 ();
 sg13g2_fill_2 FILLER_61_3387 ();
 sg13g2_decap_8 FILLER_61_3416 ();
 sg13g2_fill_2 FILLER_61_3423 ();
 sg13g2_fill_1 FILLER_61_3425 ();
 sg13g2_fill_2 FILLER_61_3439 ();
 sg13g2_fill_1 FILLER_61_3466 ();
 sg13g2_fill_2 FILLER_61_3471 ();
 sg13g2_decap_4 FILLER_61_3477 ();
 sg13g2_fill_2 FILLER_61_3481 ();
 sg13g2_decap_4 FILLER_61_3497 ();
 sg13g2_decap_8 FILLER_61_3510 ();
 sg13g2_decap_8 FILLER_61_3517 ();
 sg13g2_fill_2 FILLER_61_3524 ();
 sg13g2_decap_8 FILLER_61_3563 ();
 sg13g2_decap_8 FILLER_61_3570 ();
 sg13g2_fill_1 FILLER_61_3577 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_43 ();
 sg13g2_fill_1 FILLER_62_59 ();
 sg13g2_decap_8 FILLER_62_69 ();
 sg13g2_fill_2 FILLER_62_76 ();
 sg13g2_fill_1 FILLER_62_78 ();
 sg13g2_fill_1 FILLER_62_102 ();
 sg13g2_fill_2 FILLER_62_116 ();
 sg13g2_fill_1 FILLER_62_118 ();
 sg13g2_decap_4 FILLER_62_129 ();
 sg13g2_fill_2 FILLER_62_142 ();
 sg13g2_fill_1 FILLER_62_201 ();
 sg13g2_decap_8 FILLER_62_211 ();
 sg13g2_decap_8 FILLER_62_218 ();
 sg13g2_decap_8 FILLER_62_225 ();
 sg13g2_fill_1 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_262 ();
 sg13g2_decap_4 FILLER_62_283 ();
 sg13g2_fill_2 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_fill_1 FILLER_62_343 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_2 FILLER_62_382 ();
 sg13g2_fill_2 FILLER_62_414 ();
 sg13g2_fill_1 FILLER_62_416 ();
 sg13g2_fill_2 FILLER_62_449 ();
 sg13g2_decap_4 FILLER_62_460 ();
 sg13g2_fill_1 FILLER_62_478 ();
 sg13g2_decap_4 FILLER_62_510 ();
 sg13g2_fill_1 FILLER_62_545 ();
 sg13g2_fill_2 FILLER_62_565 ();
 sg13g2_decap_8 FILLER_62_598 ();
 sg13g2_fill_1 FILLER_62_614 ();
 sg13g2_decap_4 FILLER_62_697 ();
 sg13g2_fill_2 FILLER_62_701 ();
 sg13g2_decap_4 FILLER_62_708 ();
 sg13g2_fill_1 FILLER_62_712 ();
 sg13g2_fill_1 FILLER_62_723 ();
 sg13g2_decap_4 FILLER_62_750 ();
 sg13g2_fill_2 FILLER_62_754 ();
 sg13g2_decap_8 FILLER_62_761 ();
 sg13g2_fill_1 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_790 ();
 sg13g2_fill_1 FILLER_62_797 ();
 sg13g2_decap_8 FILLER_62_811 ();
 sg13g2_decap_4 FILLER_62_818 ();
 sg13g2_fill_1 FILLER_62_854 ();
 sg13g2_fill_1 FILLER_62_915 ();
 sg13g2_fill_2 FILLER_62_922 ();
 sg13g2_fill_1 FILLER_62_944 ();
 sg13g2_fill_2 FILLER_62_958 ();
 sg13g2_fill_1 FILLER_62_960 ();
 sg13g2_decap_8 FILLER_62_966 ();
 sg13g2_decap_8 FILLER_62_973 ();
 sg13g2_fill_2 FILLER_62_980 ();
 sg13g2_fill_2 FILLER_62_1007 ();
 sg13g2_decap_4 FILLER_62_1022 ();
 sg13g2_fill_1 FILLER_62_1026 ();
 sg13g2_fill_1 FILLER_62_1057 ();
 sg13g2_fill_1 FILLER_62_1064 ();
 sg13g2_fill_2 FILLER_62_1075 ();
 sg13g2_fill_2 FILLER_62_1105 ();
 sg13g2_decap_4 FILLER_62_1110 ();
 sg13g2_fill_1 FILLER_62_1114 ();
 sg13g2_fill_1 FILLER_62_1166 ();
 sg13g2_decap_8 FILLER_62_1175 ();
 sg13g2_decap_4 FILLER_62_1182 ();
 sg13g2_fill_1 FILLER_62_1225 ();
 sg13g2_decap_4 FILLER_62_1281 ();
 sg13g2_fill_2 FILLER_62_1285 ();
 sg13g2_decap_8 FILLER_62_1344 ();
 sg13g2_fill_1 FILLER_62_1351 ();
 sg13g2_fill_2 FILLER_62_1379 ();
 sg13g2_fill_1 FILLER_62_1381 ();
 sg13g2_decap_8 FILLER_62_1417 ();
 sg13g2_decap_4 FILLER_62_1424 ();
 sg13g2_fill_1 FILLER_62_1428 ();
 sg13g2_fill_2 FILLER_62_1486 ();
 sg13g2_fill_1 FILLER_62_1488 ();
 sg13g2_decap_8 FILLER_62_1494 ();
 sg13g2_fill_2 FILLER_62_1501 ();
 sg13g2_decap_8 FILLER_62_1512 ();
 sg13g2_decap_8 FILLER_62_1519 ();
 sg13g2_decap_4 FILLER_62_1544 ();
 sg13g2_decap_8 FILLER_62_1561 ();
 sg13g2_fill_2 FILLER_62_1568 ();
 sg13g2_decap_8 FILLER_62_1601 ();
 sg13g2_decap_8 FILLER_62_1608 ();
 sg13g2_decap_4 FILLER_62_1619 ();
 sg13g2_fill_2 FILLER_62_1623 ();
 sg13g2_decap_8 FILLER_62_1634 ();
 sg13g2_decap_8 FILLER_62_1641 ();
 sg13g2_decap_8 FILLER_62_1648 ();
 sg13g2_fill_2 FILLER_62_1655 ();
 sg13g2_fill_1 FILLER_62_1657 ();
 sg13g2_decap_4 FILLER_62_1662 ();
 sg13g2_fill_2 FILLER_62_1666 ();
 sg13g2_decap_8 FILLER_62_1677 ();
 sg13g2_decap_8 FILLER_62_1684 ();
 sg13g2_fill_2 FILLER_62_1691 ();
 sg13g2_decap_4 FILLER_62_1706 ();
 sg13g2_fill_2 FILLER_62_1710 ();
 sg13g2_decap_8 FILLER_62_1746 ();
 sg13g2_decap_8 FILLER_62_1753 ();
 sg13g2_decap_8 FILLER_62_1760 ();
 sg13g2_decap_8 FILLER_62_1767 ();
 sg13g2_decap_8 FILLER_62_1774 ();
 sg13g2_fill_1 FILLER_62_1781 ();
 sg13g2_decap_4 FILLER_62_1795 ();
 sg13g2_decap_4 FILLER_62_1808 ();
 sg13g2_decap_8 FILLER_62_1830 ();
 sg13g2_fill_2 FILLER_62_1837 ();
 sg13g2_decap_4 FILLER_62_1865 ();
 sg13g2_fill_2 FILLER_62_1874 ();
 sg13g2_fill_2 FILLER_62_1895 ();
 sg13g2_decap_8 FILLER_62_1903 ();
 sg13g2_fill_1 FILLER_62_1918 ();
 sg13g2_decap_8 FILLER_62_1928 ();
 sg13g2_decap_8 FILLER_62_1943 ();
 sg13g2_fill_1 FILLER_62_1950 ();
 sg13g2_decap_8 FILLER_62_1959 ();
 sg13g2_decap_8 FILLER_62_1966 ();
 sg13g2_decap_8 FILLER_62_1973 ();
 sg13g2_decap_8 FILLER_62_1980 ();
 sg13g2_decap_4 FILLER_62_1987 ();
 sg13g2_fill_2 FILLER_62_2012 ();
 sg13g2_fill_2 FILLER_62_2019 ();
 sg13g2_decap_8 FILLER_62_2043 ();
 sg13g2_decap_8 FILLER_62_2050 ();
 sg13g2_decap_8 FILLER_62_2057 ();
 sg13g2_decap_8 FILLER_62_2064 ();
 sg13g2_decap_8 FILLER_62_2071 ();
 sg13g2_decap_4 FILLER_62_2078 ();
 sg13g2_decap_4 FILLER_62_2087 ();
 sg13g2_fill_2 FILLER_62_2091 ();
 sg13g2_decap_4 FILLER_62_2097 ();
 sg13g2_fill_1 FILLER_62_2101 ();
 sg13g2_fill_2 FILLER_62_2107 ();
 sg13g2_fill_2 FILLER_62_2140 ();
 sg13g2_fill_2 FILLER_62_2153 ();
 sg13g2_decap_8 FILLER_62_2159 ();
 sg13g2_decap_8 FILLER_62_2166 ();
 sg13g2_fill_1 FILLER_62_2173 ();
 sg13g2_decap_8 FILLER_62_2177 ();
 sg13g2_decap_8 FILLER_62_2217 ();
 sg13g2_decap_8 FILLER_62_2224 ();
 sg13g2_decap_8 FILLER_62_2231 ();
 sg13g2_decap_8 FILLER_62_2238 ();
 sg13g2_decap_8 FILLER_62_2245 ();
 sg13g2_decap_4 FILLER_62_2252 ();
 sg13g2_fill_1 FILLER_62_2256 ();
 sg13g2_decap_8 FILLER_62_2272 ();
 sg13g2_fill_1 FILLER_62_2279 ();
 sg13g2_decap_8 FILLER_62_2285 ();
 sg13g2_decap_8 FILLER_62_2292 ();
 sg13g2_decap_4 FILLER_62_2299 ();
 sg13g2_fill_1 FILLER_62_2303 ();
 sg13g2_fill_2 FILLER_62_2317 ();
 sg13g2_decap_8 FILLER_62_2350 ();
 sg13g2_decap_8 FILLER_62_2357 ();
 sg13g2_decap_8 FILLER_62_2364 ();
 sg13g2_decap_8 FILLER_62_2371 ();
 sg13g2_decap_4 FILLER_62_2378 ();
 sg13g2_decap_8 FILLER_62_2403 ();
 sg13g2_decap_8 FILLER_62_2410 ();
 sg13g2_decap_8 FILLER_62_2417 ();
 sg13g2_decap_8 FILLER_62_2424 ();
 sg13g2_decap_4 FILLER_62_2431 ();
 sg13g2_fill_2 FILLER_62_2435 ();
 sg13g2_fill_1 FILLER_62_2470 ();
 sg13g2_fill_2 FILLER_62_2529 ();
 sg13g2_fill_2 FILLER_62_2535 ();
 sg13g2_fill_1 FILLER_62_2537 ();
 sg13g2_decap_4 FILLER_62_2562 ();
 sg13g2_fill_1 FILLER_62_2566 ();
 sg13g2_decap_8 FILLER_62_2580 ();
 sg13g2_fill_2 FILLER_62_2587 ();
 sg13g2_fill_1 FILLER_62_2589 ();
 sg13g2_decap_8 FILLER_62_2684 ();
 sg13g2_decap_8 FILLER_62_2691 ();
 sg13g2_decap_4 FILLER_62_2698 ();
 sg13g2_decap_8 FILLER_62_2758 ();
 sg13g2_decap_8 FILLER_62_2765 ();
 sg13g2_fill_2 FILLER_62_2772 ();
 sg13g2_fill_1 FILLER_62_2774 ();
 sg13g2_decap_4 FILLER_62_2790 ();
 sg13g2_fill_1 FILLER_62_2794 ();
 sg13g2_decap_8 FILLER_62_2816 ();
 sg13g2_decap_8 FILLER_62_2823 ();
 sg13g2_decap_8 FILLER_62_2830 ();
 sg13g2_fill_2 FILLER_62_2837 ();
 sg13g2_fill_1 FILLER_62_2839 ();
 sg13g2_fill_1 FILLER_62_2867 ();
 sg13g2_decap_8 FILLER_62_2895 ();
 sg13g2_decap_8 FILLER_62_2915 ();
 sg13g2_decap_8 FILLER_62_2922 ();
 sg13g2_decap_4 FILLER_62_2929 ();
 sg13g2_fill_1 FILLER_62_2933 ();
 sg13g2_decap_4 FILLER_62_2944 ();
 sg13g2_decap_8 FILLER_62_2962 ();
 sg13g2_decap_8 FILLER_62_2969 ();
 sg13g2_decap_8 FILLER_62_2976 ();
 sg13g2_decap_4 FILLER_62_2983 ();
 sg13g2_decap_4 FILLER_62_3014 ();
 sg13g2_fill_1 FILLER_62_3028 ();
 sg13g2_decap_8 FILLER_62_3056 ();
 sg13g2_decap_8 FILLER_62_3063 ();
 sg13g2_decap_8 FILLER_62_3070 ();
 sg13g2_fill_1 FILLER_62_3077 ();
 sg13g2_decap_8 FILLER_62_3109 ();
 sg13g2_decap_8 FILLER_62_3116 ();
 sg13g2_decap_8 FILLER_62_3123 ();
 sg13g2_decap_4 FILLER_62_3149 ();
 sg13g2_fill_2 FILLER_62_3153 ();
 sg13g2_decap_4 FILLER_62_3164 ();
 sg13g2_fill_2 FILLER_62_3168 ();
 sg13g2_decap_4 FILLER_62_3175 ();
 sg13g2_fill_2 FILLER_62_3179 ();
 sg13g2_decap_8 FILLER_62_3186 ();
 sg13g2_decap_8 FILLER_62_3193 ();
 sg13g2_decap_4 FILLER_62_3200 ();
 sg13g2_fill_1 FILLER_62_3204 ();
 sg13g2_decap_8 FILLER_62_3223 ();
 sg13g2_fill_2 FILLER_62_3230 ();
 sg13g2_fill_1 FILLER_62_3296 ();
 sg13g2_fill_2 FILLER_62_3311 ();
 sg13g2_fill_1 FILLER_62_3313 ();
 sg13g2_decap_8 FILLER_62_3327 ();
 sg13g2_decap_8 FILLER_62_3338 ();
 sg13g2_fill_2 FILLER_62_3345 ();
 sg13g2_fill_1 FILLER_62_3347 ();
 sg13g2_decap_4 FILLER_62_3361 ();
 sg13g2_decap_8 FILLER_62_3412 ();
 sg13g2_decap_8 FILLER_62_3419 ();
 sg13g2_fill_1 FILLER_62_3426 ();
 sg13g2_decap_8 FILLER_62_3440 ();
 sg13g2_decap_8 FILLER_62_3457 ();
 sg13g2_fill_2 FILLER_62_3464 ();
 sg13g2_fill_1 FILLER_62_3466 ();
 sg13g2_decap_8 FILLER_62_3514 ();
 sg13g2_decap_8 FILLER_62_3571 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_4 FILLER_63_14 ();
 sg13g2_fill_1 FILLER_63_18 ();
 sg13g2_fill_2 FILLER_63_24 ();
 sg13g2_decap_8 FILLER_63_62 ();
 sg13g2_decap_4 FILLER_63_69 ();
 sg13g2_fill_2 FILLER_63_73 ();
 sg13g2_fill_2 FILLER_63_102 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_decap_4 FILLER_63_110 ();
 sg13g2_fill_2 FILLER_63_114 ();
 sg13g2_decap_8 FILLER_63_143 ();
 sg13g2_fill_2 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_152 ();
 sg13g2_fill_2 FILLER_63_162 ();
 sg13g2_fill_2 FILLER_63_188 ();
 sg13g2_decap_8 FILLER_63_199 ();
 sg13g2_decap_8 FILLER_63_206 ();
 sg13g2_decap_8 FILLER_63_213 ();
 sg13g2_decap_8 FILLER_63_220 ();
 sg13g2_decap_8 FILLER_63_227 ();
 sg13g2_decap_4 FILLER_63_234 ();
 sg13g2_fill_1 FILLER_63_238 ();
 sg13g2_fill_1 FILLER_63_266 ();
 sg13g2_decap_4 FILLER_63_280 ();
 sg13g2_fill_1 FILLER_63_284 ();
 sg13g2_decap_8 FILLER_63_335 ();
 sg13g2_decap_4 FILLER_63_342 ();
 sg13g2_decap_8 FILLER_63_418 ();
 sg13g2_decap_8 FILLER_63_425 ();
 sg13g2_fill_1 FILLER_63_432 ();
 sg13g2_decap_4 FILLER_63_437 ();
 sg13g2_fill_1 FILLER_63_441 ();
 sg13g2_fill_2 FILLER_63_470 ();
 sg13g2_decap_8 FILLER_63_494 ();
 sg13g2_decap_4 FILLER_63_501 ();
 sg13g2_fill_2 FILLER_63_530 ();
 sg13g2_fill_1 FILLER_63_532 ();
 sg13g2_decap_8 FILLER_63_585 ();
 sg13g2_fill_2 FILLER_63_605 ();
 sg13g2_fill_1 FILLER_63_649 ();
 sg13g2_decap_4 FILLER_63_677 ();
 sg13g2_decap_8 FILLER_63_690 ();
 sg13g2_decap_8 FILLER_63_697 ();
 sg13g2_decap_8 FILLER_63_704 ();
 sg13g2_decap_4 FILLER_63_711 ();
 sg13g2_decap_8 FILLER_63_755 ();
 sg13g2_decap_4 FILLER_63_762 ();
 sg13g2_decap_8 FILLER_63_793 ();
 sg13g2_decap_8 FILLER_63_800 ();
 sg13g2_fill_2 FILLER_63_807 ();
 sg13g2_fill_1 FILLER_63_809 ();
 sg13g2_fill_2 FILLER_63_823 ();
 sg13g2_fill_1 FILLER_63_862 ();
 sg13g2_fill_2 FILLER_63_905 ();
 sg13g2_decap_4 FILLER_63_925 ();
 sg13g2_fill_1 FILLER_63_971 ();
 sg13g2_fill_2 FILLER_63_1030 ();
 sg13g2_decap_4 FILLER_63_1041 ();
 sg13g2_decap_8 FILLER_63_1073 ();
 sg13g2_fill_2 FILLER_63_1080 ();
 sg13g2_fill_1 FILLER_63_1082 ();
 sg13g2_fill_1 FILLER_63_1088 ();
 sg13g2_decap_4 FILLER_63_1098 ();
 sg13g2_fill_2 FILLER_63_1102 ();
 sg13g2_fill_1 FILLER_63_1134 ();
 sg13g2_fill_2 FILLER_63_1146 ();
 sg13g2_fill_2 FILLER_63_1164 ();
 sg13g2_fill_1 FILLER_63_1166 ();
 sg13g2_fill_2 FILLER_63_1180 ();
 sg13g2_fill_1 FILLER_63_1182 ();
 sg13g2_fill_2 FILLER_63_1186 ();
 sg13g2_fill_1 FILLER_63_1188 ();
 sg13g2_fill_2 FILLER_63_1228 ();
 sg13g2_decap_4 FILLER_63_1256 ();
 sg13g2_decap_8 FILLER_63_1269 ();
 sg13g2_decap_8 FILLER_63_1276 ();
 sg13g2_decap_8 FILLER_63_1283 ();
 sg13g2_decap_8 FILLER_63_1327 ();
 sg13g2_decap_8 FILLER_63_1334 ();
 sg13g2_decap_8 FILLER_63_1341 ();
 sg13g2_decap_4 FILLER_63_1348 ();
 sg13g2_fill_2 FILLER_63_1352 ();
 sg13g2_fill_1 FILLER_63_1381 ();
 sg13g2_fill_2 FILLER_63_1398 ();
 sg13g2_decap_8 FILLER_63_1422 ();
 sg13g2_decap_8 FILLER_63_1429 ();
 sg13g2_decap_8 FILLER_63_1436 ();
 sg13g2_fill_2 FILLER_63_1447 ();
 sg13g2_fill_1 FILLER_63_1449 ();
 sg13g2_decap_4 FILLER_63_1454 ();
 sg13g2_decap_4 FILLER_63_1482 ();
 sg13g2_fill_2 FILLER_63_1490 ();
 sg13g2_fill_1 FILLER_63_1492 ();
 sg13g2_decap_4 FILLER_63_1498 ();
 sg13g2_decap_4 FILLER_63_1506 ();
 sg13g2_fill_2 FILLER_63_1510 ();
 sg13g2_fill_2 FILLER_63_1518 ();
 sg13g2_fill_1 FILLER_63_1520 ();
 sg13g2_fill_1 FILLER_63_1560 ();
 sg13g2_decap_8 FILLER_63_1569 ();
 sg13g2_decap_8 FILLER_63_1576 ();
 sg13g2_decap_8 FILLER_63_1583 ();
 sg13g2_decap_8 FILLER_63_1590 ();
 sg13g2_decap_4 FILLER_63_1597 ();
 sg13g2_fill_1 FILLER_63_1601 ();
 sg13g2_decap_8 FILLER_63_1606 ();
 sg13g2_decap_8 FILLER_63_1623 ();
 sg13g2_fill_1 FILLER_63_1630 ();
 sg13g2_fill_2 FILLER_63_1640 ();
 sg13g2_fill_1 FILLER_63_1642 ();
 sg13g2_fill_1 FILLER_63_1682 ();
 sg13g2_decap_8 FILLER_63_1696 ();
 sg13g2_decap_8 FILLER_63_1703 ();
 sg13g2_decap_8 FILLER_63_1710 ();
 sg13g2_decap_8 FILLER_63_1754 ();
 sg13g2_decap_8 FILLER_63_1761 ();
 sg13g2_decap_8 FILLER_63_1768 ();
 sg13g2_decap_4 FILLER_63_1775 ();
 sg13g2_fill_2 FILLER_63_1779 ();
 sg13g2_decap_4 FILLER_63_1803 ();
 sg13g2_decap_4 FILLER_63_1815 ();
 sg13g2_fill_1 FILLER_63_1826 ();
 sg13g2_decap_8 FILLER_63_1833 ();
 sg13g2_decap_8 FILLER_63_1840 ();
 sg13g2_decap_8 FILLER_63_1847 ();
 sg13g2_fill_2 FILLER_63_1854 ();
 sg13g2_fill_1 FILLER_63_1856 ();
 sg13g2_decap_8 FILLER_63_1891 ();
 sg13g2_decap_8 FILLER_63_1898 ();
 sg13g2_decap_8 FILLER_63_1905 ();
 sg13g2_decap_4 FILLER_63_1912 ();
 sg13g2_fill_1 FILLER_63_1916 ();
 sg13g2_decap_4 FILLER_63_1922 ();
 sg13g2_fill_1 FILLER_63_1926 ();
 sg13g2_decap_8 FILLER_63_1940 ();
 sg13g2_fill_2 FILLER_63_1947 ();
 sg13g2_decap_4 FILLER_63_1957 ();
 sg13g2_decap_8 FILLER_63_1969 ();
 sg13g2_decap_8 FILLER_63_1976 ();
 sg13g2_fill_2 FILLER_63_1991 ();
 sg13g2_decap_4 FILLER_63_2021 ();
 sg13g2_fill_2 FILLER_63_2029 ();
 sg13g2_decap_8 FILLER_63_2036 ();
 sg13g2_decap_8 FILLER_63_2049 ();
 sg13g2_decap_8 FILLER_63_2056 ();
 sg13g2_fill_2 FILLER_63_2063 ();
 sg13g2_decap_8 FILLER_63_2068 ();
 sg13g2_fill_2 FILLER_63_2075 ();
 sg13g2_fill_2 FILLER_63_2085 ();
 sg13g2_fill_1 FILLER_63_2087 ();
 sg13g2_decap_4 FILLER_63_2115 ();
 sg13g2_fill_2 FILLER_63_2128 ();
 sg13g2_decap_8 FILLER_63_2138 ();
 sg13g2_decap_8 FILLER_63_2150 ();
 sg13g2_decap_4 FILLER_63_2157 ();
 sg13g2_fill_1 FILLER_63_2161 ();
 sg13g2_decap_8 FILLER_63_2222 ();
 sg13g2_decap_8 FILLER_63_2229 ();
 sg13g2_decap_8 FILLER_63_2245 ();
 sg13g2_fill_1 FILLER_63_2252 ();
 sg13g2_fill_2 FILLER_63_2300 ();
 sg13g2_fill_1 FILLER_63_2302 ();
 sg13g2_fill_2 FILLER_63_2355 ();
 sg13g2_decap_8 FILLER_63_2412 ();
 sg13g2_decap_8 FILLER_63_2419 ();
 sg13g2_fill_2 FILLER_63_2426 ();
 sg13g2_decap_8 FILLER_63_2432 ();
 sg13g2_decap_8 FILLER_63_2439 ();
 sg13g2_fill_2 FILLER_63_2446 ();
 sg13g2_fill_1 FILLER_63_2448 ();
 sg13g2_decap_8 FILLER_63_2459 ();
 sg13g2_decap_8 FILLER_63_2466 ();
 sg13g2_fill_2 FILLER_63_2473 ();
 sg13g2_fill_1 FILLER_63_2475 ();
 sg13g2_decap_4 FILLER_63_2516 ();
 sg13g2_fill_1 FILLER_63_2520 ();
 sg13g2_decap_8 FILLER_63_2530 ();
 sg13g2_fill_1 FILLER_63_2564 ();
 sg13g2_decap_8 FILLER_63_2575 ();
 sg13g2_decap_8 FILLER_63_2582 ();
 sg13g2_decap_8 FILLER_63_2589 ();
 sg13g2_decap_4 FILLER_63_2596 ();
 sg13g2_decap_4 FILLER_63_2652 ();
 sg13g2_fill_1 FILLER_63_2656 ();
 sg13g2_fill_2 FILLER_63_2671 ();
 sg13g2_decap_8 FILLER_63_2682 ();
 sg13g2_decap_8 FILLER_63_2689 ();
 sg13g2_fill_2 FILLER_63_2696 ();
 sg13g2_fill_1 FILLER_63_2698 ();
 sg13g2_decap_8 FILLER_63_2740 ();
 sg13g2_decap_8 FILLER_63_2747 ();
 sg13g2_decap_8 FILLER_63_2754 ();
 sg13g2_fill_2 FILLER_63_2761 ();
 sg13g2_fill_2 FILLER_63_2768 ();
 sg13g2_fill_1 FILLER_63_2770 ();
 sg13g2_decap_8 FILLER_63_2834 ();
 sg13g2_decap_8 FILLER_63_2841 ();
 sg13g2_fill_1 FILLER_63_2848 ();
 sg13g2_fill_2 FILLER_63_2880 ();
 sg13g2_fill_1 FILLER_63_2882 ();
 sg13g2_decap_8 FILLER_63_2910 ();
 sg13g2_decap_8 FILLER_63_2917 ();
 sg13g2_fill_1 FILLER_63_2924 ();
 sg13g2_fill_1 FILLER_63_2965 ();
 sg13g2_decap_4 FILLER_63_2975 ();
 sg13g2_fill_2 FILLER_63_2979 ();
 sg13g2_decap_8 FILLER_63_3070 ();
 sg13g2_decap_4 FILLER_63_3077 ();
 sg13g2_fill_1 FILLER_63_3085 ();
 sg13g2_decap_8 FILLER_63_3109 ();
 sg13g2_decap_8 FILLER_63_3116 ();
 sg13g2_decap_8 FILLER_63_3123 ();
 sg13g2_fill_1 FILLER_63_3130 ();
 sg13g2_fill_2 FILLER_63_3159 ();
 sg13g2_decap_8 FILLER_63_3198 ();
 sg13g2_decap_8 FILLER_63_3205 ();
 sg13g2_decap_8 FILLER_63_3212 ();
 sg13g2_decap_8 FILLER_63_3219 ();
 sg13g2_fill_2 FILLER_63_3226 ();
 sg13g2_fill_1 FILLER_63_3228 ();
 sg13g2_fill_2 FILLER_63_3285 ();
 sg13g2_fill_2 FILLER_63_3311 ();
 sg13g2_fill_1 FILLER_63_3313 ();
 sg13g2_decap_8 FILLER_63_3333 ();
 sg13g2_decap_8 FILLER_63_3340 ();
 sg13g2_decap_8 FILLER_63_3347 ();
 sg13g2_decap_8 FILLER_63_3354 ();
 sg13g2_decap_4 FILLER_63_3361 ();
 sg13g2_fill_2 FILLER_63_3365 ();
 sg13g2_fill_2 FILLER_63_3401 ();
 sg13g2_decap_8 FILLER_63_3412 ();
 sg13g2_decap_8 FILLER_63_3419 ();
 sg13g2_decap_8 FILLER_63_3447 ();
 sg13g2_fill_2 FILLER_63_3454 ();
 sg13g2_fill_1 FILLER_63_3456 ();
 sg13g2_decap_8 FILLER_63_3516 ();
 sg13g2_decap_8 FILLER_63_3523 ();
 sg13g2_fill_1 FILLER_63_3530 ();
 sg13g2_decap_8 FILLER_63_3569 ();
 sg13g2_fill_2 FILLER_63_3576 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_fill_2 FILLER_64_18 ();
 sg13g2_fill_2 FILLER_64_55 ();
 sg13g2_fill_2 FILLER_64_97 ();
 sg13g2_fill_2 FILLER_64_117 ();
 sg13g2_fill_1 FILLER_64_119 ();
 sg13g2_fill_2 FILLER_64_151 ();
 sg13g2_fill_1 FILLER_64_158 ();
 sg13g2_decap_4 FILLER_64_178 ();
 sg13g2_decap_4 FILLER_64_191 ();
 sg13g2_fill_1 FILLER_64_223 ();
 sg13g2_fill_2 FILLER_64_232 ();
 sg13g2_fill_2 FILLER_64_243 ();
 sg13g2_fill_2 FILLER_64_253 ();
 sg13g2_decap_8 FILLER_64_270 ();
 sg13g2_decap_8 FILLER_64_277 ();
 sg13g2_fill_2 FILLER_64_284 ();
 sg13g2_fill_2 FILLER_64_295 ();
 sg13g2_decap_4 FILLER_64_306 ();
 sg13g2_fill_1 FILLER_64_310 ();
 sg13g2_decap_8 FILLER_64_341 ();
 sg13g2_decap_4 FILLER_64_348 ();
 sg13g2_fill_2 FILLER_64_352 ();
 sg13g2_fill_1 FILLER_64_381 ();
 sg13g2_decap_8 FILLER_64_410 ();
 sg13g2_decap_8 FILLER_64_417 ();
 sg13g2_decap_8 FILLER_64_424 ();
 sg13g2_decap_8 FILLER_64_431 ();
 sg13g2_fill_2 FILLER_64_438 ();
 sg13g2_fill_1 FILLER_64_440 ();
 sg13g2_fill_2 FILLER_64_486 ();
 sg13g2_decap_4 FILLER_64_597 ();
 sg13g2_fill_2 FILLER_64_649 ();
 sg13g2_fill_1 FILLER_64_651 ();
 sg13g2_decap_8 FILLER_64_657 ();
 sg13g2_fill_1 FILLER_64_664 ();
 sg13g2_decap_8 FILLER_64_674 ();
 sg13g2_decap_8 FILLER_64_681 ();
 sg13g2_decap_8 FILLER_64_688 ();
 sg13g2_decap_8 FILLER_64_695 ();
 sg13g2_decap_8 FILLER_64_702 ();
 sg13g2_fill_1 FILLER_64_709 ();
 sg13g2_decap_4 FILLER_64_715 ();
 sg13g2_fill_2 FILLER_64_719 ();
 sg13g2_fill_2 FILLER_64_739 ();
 sg13g2_fill_1 FILLER_64_746 ();
 sg13g2_fill_2 FILLER_64_752 ();
 sg13g2_decap_8 FILLER_64_774 ();
 sg13g2_decap_8 FILLER_64_781 ();
 sg13g2_decap_8 FILLER_64_788 ();
 sg13g2_decap_8 FILLER_64_795 ();
 sg13g2_decap_8 FILLER_64_802 ();
 sg13g2_decap_4 FILLER_64_809 ();
 sg13g2_fill_2 FILLER_64_813 ();
 sg13g2_fill_2 FILLER_64_842 ();
 sg13g2_fill_1 FILLER_64_844 ();
 sg13g2_decap_8 FILLER_64_861 ();
 sg13g2_decap_4 FILLER_64_868 ();
 sg13g2_fill_1 FILLER_64_934 ();
 sg13g2_decap_8 FILLER_64_963 ();
 sg13g2_fill_1 FILLER_64_970 ();
 sg13g2_fill_2 FILLER_64_1000 ();
 sg13g2_decap_4 FILLER_64_1029 ();
 sg13g2_decap_8 FILLER_64_1069 ();
 sg13g2_decap_8 FILLER_64_1076 ();
 sg13g2_decap_8 FILLER_64_1083 ();
 sg13g2_decap_4 FILLER_64_1090 ();
 sg13g2_fill_2 FILLER_64_1094 ();
 sg13g2_fill_2 FILLER_64_1113 ();
 sg13g2_fill_2 FILLER_64_1124 ();
 sg13g2_decap_8 FILLER_64_1154 ();
 sg13g2_decap_8 FILLER_64_1161 ();
 sg13g2_decap_8 FILLER_64_1168 ();
 sg13g2_fill_1 FILLER_64_1175 ();
 sg13g2_decap_4 FILLER_64_1193 ();
 sg13g2_decap_8 FILLER_64_1261 ();
 sg13g2_decap_8 FILLER_64_1268 ();
 sg13g2_fill_2 FILLER_64_1275 ();
 sg13g2_decap_4 FILLER_64_1281 ();
 sg13g2_fill_1 FILLER_64_1285 ();
 sg13g2_decap_8 FILLER_64_1308 ();
 sg13g2_decap_8 FILLER_64_1315 ();
 sg13g2_decap_8 FILLER_64_1322 ();
 sg13g2_decap_8 FILLER_64_1329 ();
 sg13g2_decap_4 FILLER_64_1336 ();
 sg13g2_fill_1 FILLER_64_1340 ();
 sg13g2_decap_8 FILLER_64_1350 ();
 sg13g2_decap_4 FILLER_64_1357 ();
 sg13g2_fill_2 FILLER_64_1392 ();
 sg13g2_fill_2 FILLER_64_1418 ();
 sg13g2_fill_1 FILLER_64_1420 ();
 sg13g2_decap_8 FILLER_64_1431 ();
 sg13g2_decap_8 FILLER_64_1460 ();
 sg13g2_decap_4 FILLER_64_1467 ();
 sg13g2_decap_8 FILLER_64_1498 ();
 sg13g2_decap_4 FILLER_64_1505 ();
 sg13g2_decap_8 FILLER_64_1518 ();
 sg13g2_decap_8 FILLER_64_1525 ();
 sg13g2_decap_8 FILLER_64_1571 ();
 sg13g2_decap_8 FILLER_64_1578 ();
 sg13g2_decap_8 FILLER_64_1585 ();
 sg13g2_fill_1 FILLER_64_1647 ();
 sg13g2_decap_4 FILLER_64_1686 ();
 sg13g2_decap_4 FILLER_64_1699 ();
 sg13g2_fill_2 FILLER_64_1703 ();
 sg13g2_decap_8 FILLER_64_1710 ();
 sg13g2_decap_8 FILLER_64_1745 ();
 sg13g2_decap_8 FILLER_64_1752 ();
 sg13g2_decap_8 FILLER_64_1759 ();
 sg13g2_decap_8 FILLER_64_1770 ();
 sg13g2_decap_4 FILLER_64_1777 ();
 sg13g2_decap_8 FILLER_64_1806 ();
 sg13g2_fill_1 FILLER_64_1813 ();
 sg13g2_decap_4 FILLER_64_1822 ();
 sg13g2_fill_1 FILLER_64_1826 ();
 sg13g2_fill_1 FILLER_64_1837 ();
 sg13g2_decap_8 FILLER_64_1851 ();
 sg13g2_decap_8 FILLER_64_1858 ();
 sg13g2_fill_2 FILLER_64_1891 ();
 sg13g2_decap_4 FILLER_64_1907 ();
 sg13g2_fill_1 FILLER_64_1927 ();
 sg13g2_fill_1 FILLER_64_1933 ();
 sg13g2_decap_8 FILLER_64_1949 ();
 sg13g2_fill_2 FILLER_64_1956 ();
 sg13g2_decap_4 FILLER_64_2013 ();
 sg13g2_decap_8 FILLER_64_2030 ();
 sg13g2_fill_2 FILLER_64_2042 ();
 sg13g2_fill_1 FILLER_64_2053 ();
 sg13g2_fill_2 FILLER_64_2072 ();
 sg13g2_fill_1 FILLER_64_2074 ();
 sg13g2_fill_1 FILLER_64_2089 ();
 sg13g2_decap_4 FILLER_64_2111 ();
 sg13g2_decap_8 FILLER_64_2127 ();
 sg13g2_decap_4 FILLER_64_2134 ();
 sg13g2_fill_2 FILLER_64_2138 ();
 sg13g2_decap_8 FILLER_64_2146 ();
 sg13g2_decap_8 FILLER_64_2153 ();
 sg13g2_decap_8 FILLER_64_2160 ();
 sg13g2_fill_1 FILLER_64_2167 ();
 sg13g2_fill_1 FILLER_64_2196 ();
 sg13g2_decap_8 FILLER_64_2223 ();
 sg13g2_decap_8 FILLER_64_2230 ();
 sg13g2_decap_8 FILLER_64_2237 ();
 sg13g2_decap_8 FILLER_64_2244 ();
 sg13g2_fill_1 FILLER_64_2251 ();
 sg13g2_decap_4 FILLER_64_2256 ();
 sg13g2_fill_1 FILLER_64_2260 ();
 sg13g2_decap_8 FILLER_64_2275 ();
 sg13g2_decap_4 FILLER_64_2282 ();
 sg13g2_fill_1 FILLER_64_2290 ();
 sg13g2_decap_4 FILLER_64_2304 ();
 sg13g2_decap_4 FILLER_64_2322 ();
 sg13g2_fill_1 FILLER_64_2326 ();
 sg13g2_decap_4 FILLER_64_2358 ();
 sg13g2_decap_8 FILLER_64_2417 ();
 sg13g2_decap_8 FILLER_64_2424 ();
 sg13g2_decap_8 FILLER_64_2431 ();
 sg13g2_decap_8 FILLER_64_2438 ();
 sg13g2_fill_1 FILLER_64_2445 ();
 sg13g2_fill_2 FILLER_64_2456 ();
 sg13g2_decap_8 FILLER_64_2479 ();
 sg13g2_decap_8 FILLER_64_2486 ();
 sg13g2_fill_1 FILLER_64_2493 ();
 sg13g2_fill_2 FILLER_64_2498 ();
 sg13g2_fill_2 FILLER_64_2504 ();
 sg13g2_fill_1 FILLER_64_2506 ();
 sg13g2_fill_2 FILLER_64_2526 ();
 sg13g2_fill_2 FILLER_64_2567 ();
 sg13g2_decap_8 FILLER_64_2596 ();
 sg13g2_decap_8 FILLER_64_2643 ();
 sg13g2_decap_8 FILLER_64_2650 ();
 sg13g2_fill_1 FILLER_64_2657 ();
 sg13g2_fill_2 FILLER_64_2668 ();
 sg13g2_decap_8 FILLER_64_2683 ();
 sg13g2_fill_2 FILLER_64_2690 ();
 sg13g2_decap_8 FILLER_64_2747 ();
 sg13g2_decap_8 FILLER_64_2754 ();
 sg13g2_fill_1 FILLER_64_2761 ();
 sg13g2_fill_2 FILLER_64_2766 ();
 sg13g2_fill_1 FILLER_64_2768 ();
 sg13g2_decap_4 FILLER_64_2804 ();
 sg13g2_decap_8 FILLER_64_2835 ();
 sg13g2_decap_8 FILLER_64_2842 ();
 sg13g2_fill_1 FILLER_64_2849 ();
 sg13g2_decap_8 FILLER_64_2907 ();
 sg13g2_decap_4 FILLER_64_2914 ();
 sg13g2_decap_8 FILLER_64_2980 ();
 sg13g2_fill_2 FILLER_64_2987 ();
 sg13g2_fill_1 FILLER_64_2989 ();
 sg13g2_fill_1 FILLER_64_3004 ();
 sg13g2_fill_2 FILLER_64_3014 ();
 sg13g2_fill_1 FILLER_64_3016 ();
 sg13g2_fill_2 FILLER_64_3021 ();
 sg13g2_fill_1 FILLER_64_3023 ();
 sg13g2_fill_1 FILLER_64_3034 ();
 sg13g2_decap_4 FILLER_64_3070 ();
 sg13g2_fill_2 FILLER_64_3074 ();
 sg13g2_decap_8 FILLER_64_3124 ();
 sg13g2_fill_2 FILLER_64_3131 ();
 sg13g2_decap_8 FILLER_64_3227 ();
 sg13g2_fill_2 FILLER_64_3234 ();
 sg13g2_fill_1 FILLER_64_3236 ();
 sg13g2_fill_2 FILLER_64_3241 ();
 sg13g2_fill_1 FILLER_64_3243 ();
 sg13g2_fill_1 FILLER_64_3248 ();
 sg13g2_decap_8 FILLER_64_3263 ();
 sg13g2_decap_8 FILLER_64_3270 ();
 sg13g2_decap_8 FILLER_64_3277 ();
 sg13g2_decap_8 FILLER_64_3284 ();
 sg13g2_decap_8 FILLER_64_3291 ();
 sg13g2_decap_4 FILLER_64_3298 ();
 sg13g2_fill_2 FILLER_64_3302 ();
 sg13g2_decap_8 FILLER_64_3350 ();
 sg13g2_decap_8 FILLER_64_3357 ();
 sg13g2_decap_4 FILLER_64_3364 ();
 sg13g2_fill_2 FILLER_64_3368 ();
 sg13g2_decap_8 FILLER_64_3400 ();
 sg13g2_decap_8 FILLER_64_3407 ();
 sg13g2_decap_8 FILLER_64_3414 ();
 sg13g2_decap_8 FILLER_64_3421 ();
 sg13g2_fill_1 FILLER_64_3428 ();
 sg13g2_fill_2 FILLER_64_3452 ();
 sg13g2_fill_1 FILLER_64_3454 ();
 sg13g2_decap_8 FILLER_64_3512 ();
 sg13g2_decap_8 FILLER_64_3519 ();
 sg13g2_decap_8 FILLER_64_3526 ();
 sg13g2_decap_4 FILLER_64_3533 ();
 sg13g2_decap_8 FILLER_64_3560 ();
 sg13g2_decap_8 FILLER_64_3567 ();
 sg13g2_decap_4 FILLER_64_3574 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_decap_4 FILLER_65_66 ();
 sg13g2_decap_8 FILLER_65_115 ();
 sg13g2_fill_2 FILLER_65_122 ();
 sg13g2_decap_4 FILLER_65_129 ();
 sg13g2_fill_2 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_179 ();
 sg13g2_decap_8 FILLER_65_186 ();
 sg13g2_decap_8 FILLER_65_193 ();
 sg13g2_decap_8 FILLER_65_200 ();
 sg13g2_fill_1 FILLER_65_207 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_4 FILLER_65_280 ();
 sg13g2_fill_1 FILLER_65_284 ();
 sg13g2_decap_8 FILLER_65_326 ();
 sg13g2_decap_8 FILLER_65_333 ();
 sg13g2_decap_8 FILLER_65_340 ();
 sg13g2_decap_8 FILLER_65_347 ();
 sg13g2_decap_8 FILLER_65_354 ();
 sg13g2_decap_8 FILLER_65_361 ();
 sg13g2_decap_4 FILLER_65_368 ();
 sg13g2_fill_2 FILLER_65_387 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_fill_2 FILLER_65_401 ();
 sg13g2_decap_8 FILLER_65_412 ();
 sg13g2_decap_8 FILLER_65_419 ();
 sg13g2_decap_8 FILLER_65_426 ();
 sg13g2_decap_8 FILLER_65_433 ();
 sg13g2_decap_8 FILLER_65_440 ();
 sg13g2_fill_1 FILLER_65_447 ();
 sg13g2_decap_4 FILLER_65_483 ();
 sg13g2_fill_2 FILLER_65_559 ();
 sg13g2_fill_1 FILLER_65_561 ();
 sg13g2_decap_8 FILLER_65_590 ();
 sg13g2_decap_8 FILLER_65_597 ();
 sg13g2_decap_4 FILLER_65_604 ();
 sg13g2_fill_2 FILLER_65_621 ();
 sg13g2_decap_8 FILLER_65_649 ();
 sg13g2_decap_8 FILLER_65_656 ();
 sg13g2_decap_8 FILLER_65_663 ();
 sg13g2_decap_8 FILLER_65_670 ();
 sg13g2_decap_8 FILLER_65_677 ();
 sg13g2_decap_4 FILLER_65_684 ();
 sg13g2_fill_1 FILLER_65_688 ();
 sg13g2_fill_2 FILLER_65_716 ();
 sg13g2_fill_2 FILLER_65_723 ();
 sg13g2_fill_1 FILLER_65_725 ();
 sg13g2_decap_4 FILLER_65_812 ();
 sg13g2_fill_1 FILLER_65_842 ();
 sg13g2_decap_8 FILLER_65_852 ();
 sg13g2_decap_8 FILLER_65_859 ();
 sg13g2_decap_8 FILLER_65_866 ();
 sg13g2_fill_1 FILLER_65_873 ();
 sg13g2_fill_1 FILLER_65_901 ();
 sg13g2_fill_1 FILLER_65_916 ();
 sg13g2_decap_8 FILLER_65_925 ();
 sg13g2_decap_8 FILLER_65_932 ();
 sg13g2_decap_8 FILLER_65_939 ();
 sg13g2_decap_8 FILLER_65_946 ();
 sg13g2_decap_8 FILLER_65_953 ();
 sg13g2_decap_8 FILLER_65_960 ();
 sg13g2_decap_4 FILLER_65_967 ();
 sg13g2_fill_1 FILLER_65_971 ();
 sg13g2_fill_1 FILLER_65_1005 ();
 sg13g2_decap_4 FILLER_65_1034 ();
 sg13g2_fill_2 FILLER_65_1038 ();
 sg13g2_fill_2 FILLER_65_1056 ();
 sg13g2_fill_1 FILLER_65_1058 ();
 sg13g2_decap_8 FILLER_65_1068 ();
 sg13g2_fill_2 FILLER_65_1075 ();
 sg13g2_decap_8 FILLER_65_1086 ();
 sg13g2_fill_1 FILLER_65_1093 ();
 sg13g2_fill_2 FILLER_65_1126 ();
 sg13g2_fill_1 FILLER_65_1128 ();
 sg13g2_fill_1 FILLER_65_1143 ();
 sg13g2_decap_8 FILLER_65_1153 ();
 sg13g2_decap_8 FILLER_65_1160 ();
 sg13g2_decap_4 FILLER_65_1167 ();
 sg13g2_fill_2 FILLER_65_1171 ();
 sg13g2_fill_2 FILLER_65_1182 ();
 sg13g2_decap_8 FILLER_65_1202 ();
 sg13g2_fill_2 FILLER_65_1222 ();
 sg13g2_fill_1 FILLER_65_1224 ();
 sg13g2_decap_8 FILLER_65_1242 ();
 sg13g2_decap_4 FILLER_65_1249 ();
 sg13g2_fill_2 FILLER_65_1273 ();
 sg13g2_fill_1 FILLER_65_1275 ();
 sg13g2_fill_1 FILLER_65_1334 ();
 sg13g2_fill_2 FILLER_65_1362 ();
 sg13g2_fill_1 FILLER_65_1364 ();
 sg13g2_fill_2 FILLER_65_1378 ();
 sg13g2_fill_2 FILLER_65_1405 ();
 sg13g2_fill_2 FILLER_65_1418 ();
 sg13g2_fill_2 FILLER_65_1428 ();
 sg13g2_fill_1 FILLER_65_1430 ();
 sg13g2_decap_8 FILLER_65_1471 ();
 sg13g2_fill_1 FILLER_65_1478 ();
 sg13g2_decap_8 FILLER_65_1525 ();
 sg13g2_decap_4 FILLER_65_1532 ();
 sg13g2_fill_1 FILLER_65_1536 ();
 sg13g2_decap_8 FILLER_65_1582 ();
 sg13g2_decap_4 FILLER_65_1589 ();
 sg13g2_fill_1 FILLER_65_1598 ();
 sg13g2_decap_8 FILLER_65_1636 ();
 sg13g2_decap_8 FILLER_65_1643 ();
 sg13g2_fill_2 FILLER_65_1650 ();
 sg13g2_decap_4 FILLER_65_1678 ();
 sg13g2_fill_2 FILLER_65_1715 ();
 sg13g2_fill_1 FILLER_65_1717 ();
 sg13g2_fill_2 FILLER_65_1725 ();
 sg13g2_decap_8 FILLER_65_1748 ();
 sg13g2_fill_2 FILLER_65_1755 ();
 sg13g2_fill_1 FILLER_65_1757 ();
 sg13g2_fill_2 FILLER_65_1785 ();
 sg13g2_fill_1 FILLER_65_1799 ();
 sg13g2_decap_8 FILLER_65_1809 ();
 sg13g2_fill_1 FILLER_65_1816 ();
 sg13g2_fill_2 FILLER_65_1831 ();
 sg13g2_decap_8 FILLER_65_1839 ();
 sg13g2_decap_8 FILLER_65_1846 ();
 sg13g2_decap_8 FILLER_65_1853 ();
 sg13g2_decap_4 FILLER_65_1860 ();
 sg13g2_fill_2 FILLER_65_1864 ();
 sg13g2_decap_4 FILLER_65_1879 ();
 sg13g2_fill_2 FILLER_65_1907 ();
 sg13g2_fill_2 FILLER_65_1935 ();
 sg13g2_decap_8 FILLER_65_1944 ();
 sg13g2_decap_8 FILLER_65_1951 ();
 sg13g2_decap_8 FILLER_65_1958 ();
 sg13g2_decap_8 FILLER_65_1965 ();
 sg13g2_decap_8 FILLER_65_1972 ();
 sg13g2_decap_8 FILLER_65_1984 ();
 sg13g2_fill_2 FILLER_65_1991 ();
 sg13g2_fill_1 FILLER_65_1993 ();
 sg13g2_decap_8 FILLER_65_1999 ();
 sg13g2_decap_8 FILLER_65_2006 ();
 sg13g2_decap_8 FILLER_65_2013 ();
 sg13g2_fill_1 FILLER_65_2020 ();
 sg13g2_fill_2 FILLER_65_2034 ();
 sg13g2_fill_1 FILLER_65_2036 ();
 sg13g2_fill_1 FILLER_65_2050 ();
 sg13g2_decap_8 FILLER_65_2056 ();
 sg13g2_decap_8 FILLER_65_2063 ();
 sg13g2_decap_4 FILLER_65_2070 ();
 sg13g2_fill_2 FILLER_65_2074 ();
 sg13g2_fill_2 FILLER_65_2094 ();
 sg13g2_fill_1 FILLER_65_2096 ();
 sg13g2_fill_1 FILLER_65_2107 ();
 sg13g2_decap_8 FILLER_65_2117 ();
 sg13g2_decap_4 FILLER_65_2124 ();
 sg13g2_fill_1 FILLER_65_2128 ();
 sg13g2_decap_8 FILLER_65_2137 ();
 sg13g2_fill_1 FILLER_65_2144 ();
 sg13g2_fill_2 FILLER_65_2163 ();
 sg13g2_decap_8 FILLER_65_2171 ();
 sg13g2_fill_2 FILLER_65_2189 ();
 sg13g2_decap_8 FILLER_65_2213 ();
 sg13g2_decap_8 FILLER_65_2220 ();
 sg13g2_decap_8 FILLER_65_2227 ();
 sg13g2_decap_8 FILLER_65_2234 ();
 sg13g2_decap_8 FILLER_65_2241 ();
 sg13g2_fill_2 FILLER_65_2288 ();
 sg13g2_fill_2 FILLER_65_2304 ();
 sg13g2_fill_1 FILLER_65_2306 ();
 sg13g2_fill_2 FILLER_65_2320 ();
 sg13g2_decap_8 FILLER_65_2342 ();
 sg13g2_decap_4 FILLER_65_2362 ();
 sg13g2_decap_8 FILLER_65_2400 ();
 sg13g2_decap_8 FILLER_65_2407 ();
 sg13g2_decap_8 FILLER_65_2414 ();
 sg13g2_decap_8 FILLER_65_2421 ();
 sg13g2_decap_8 FILLER_65_2428 ();
 sg13g2_fill_2 FILLER_65_2435 ();
 sg13g2_fill_2 FILLER_65_2468 ();
 sg13g2_decap_8 FILLER_65_2479 ();
 sg13g2_decap_8 FILLER_65_2486 ();
 sg13g2_decap_8 FILLER_65_2493 ();
 sg13g2_decap_8 FILLER_65_2500 ();
 sg13g2_decap_4 FILLER_65_2507 ();
 sg13g2_fill_1 FILLER_65_2511 ();
 sg13g2_decap_8 FILLER_65_2593 ();
 sg13g2_decap_8 FILLER_65_2600 ();
 sg13g2_fill_2 FILLER_65_2607 ();
 sg13g2_fill_2 FILLER_65_2613 ();
 sg13g2_decap_4 FILLER_65_2624 ();
 sg13g2_decap_8 FILLER_65_2637 ();
 sg13g2_fill_2 FILLER_65_2644 ();
 sg13g2_fill_2 FILLER_65_2656 ();
 sg13g2_decap_8 FILLER_65_2672 ();
 sg13g2_decap_8 FILLER_65_2679 ();
 sg13g2_decap_8 FILLER_65_2686 ();
 sg13g2_fill_1 FILLER_65_2693 ();
 sg13g2_fill_2 FILLER_65_2704 ();
 sg13g2_fill_1 FILLER_65_2706 ();
 sg13g2_decap_8 FILLER_65_2747 ();
 sg13g2_fill_2 FILLER_65_2754 ();
 sg13g2_fill_1 FILLER_65_2756 ();
 sg13g2_decap_4 FILLER_65_2770 ();
 sg13g2_fill_1 FILLER_65_2774 ();
 sg13g2_decap_4 FILLER_65_2790 ();
 sg13g2_fill_1 FILLER_65_2803 ();
 sg13g2_decap_8 FILLER_65_2836 ();
 sg13g2_decap_8 FILLER_65_2843 ();
 sg13g2_decap_8 FILLER_65_2850 ();
 sg13g2_fill_2 FILLER_65_2857 ();
 sg13g2_fill_1 FILLER_65_2859 ();
 sg13g2_fill_2 FILLER_65_2873 ();
 sg13g2_decap_4 FILLER_65_2917 ();
 sg13g2_decap_8 FILLER_65_2980 ();
 sg13g2_decap_8 FILLER_65_2987 ();
 sg13g2_fill_1 FILLER_65_2994 ();
 sg13g2_decap_8 FILLER_65_3008 ();
 sg13g2_decap_8 FILLER_65_3015 ();
 sg13g2_decap_8 FILLER_65_3022 ();
 sg13g2_fill_1 FILLER_65_3029 ();
 sg13g2_decap_8 FILLER_65_3065 ();
 sg13g2_decap_8 FILLER_65_3072 ();
 sg13g2_decap_8 FILLER_65_3079 ();
 sg13g2_fill_1 FILLER_65_3086 ();
 sg13g2_fill_2 FILLER_65_3144 ();
 sg13g2_fill_1 FILLER_65_3146 ();
 sg13g2_fill_2 FILLER_65_3174 ();
 sg13g2_fill_1 FILLER_65_3180 ();
 sg13g2_decap_8 FILLER_65_3236 ();
 sg13g2_decap_8 FILLER_65_3243 ();
 sg13g2_decap_8 FILLER_65_3250 ();
 sg13g2_fill_1 FILLER_65_3257 ();
 sg13g2_fill_2 FILLER_65_3268 ();
 sg13g2_decap_8 FILLER_65_3279 ();
 sg13g2_decap_4 FILLER_65_3286 ();
 sg13g2_fill_1 FILLER_65_3290 ();
 sg13g2_fill_2 FILLER_65_3294 ();
 sg13g2_fill_1 FILLER_65_3296 ();
 sg13g2_decap_8 FILLER_65_3345 ();
 sg13g2_decap_4 FILLER_65_3352 ();
 sg13g2_fill_2 FILLER_65_3356 ();
 sg13g2_fill_1 FILLER_65_3405 ();
 sg13g2_decap_8 FILLER_65_3410 ();
 sg13g2_fill_1 FILLER_65_3417 ();
 sg13g2_decap_8 FILLER_65_3431 ();
 sg13g2_decap_8 FILLER_65_3438 ();
 sg13g2_decap_8 FILLER_65_3445 ();
 sg13g2_decap_4 FILLER_65_3455 ();
 sg13g2_fill_1 FILLER_65_3459 ();
 sg13g2_fill_2 FILLER_65_3464 ();
 sg13g2_fill_1 FILLER_65_3466 ();
 sg13g2_fill_2 FILLER_65_3502 ();
 sg13g2_fill_1 FILLER_65_3504 ();
 sg13g2_decap_8 FILLER_65_3515 ();
 sg13g2_decap_8 FILLER_65_3568 ();
 sg13g2_fill_2 FILLER_65_3575 ();
 sg13g2_fill_1 FILLER_65_3577 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_fill_1 FILLER_66_45 ();
 sg13g2_fill_1 FILLER_66_61 ();
 sg13g2_decap_4 FILLER_66_71 ();
 sg13g2_fill_1 FILLER_66_111 ();
 sg13g2_decap_8 FILLER_66_117 ();
 sg13g2_fill_2 FILLER_66_124 ();
 sg13g2_decap_8 FILLER_66_131 ();
 sg13g2_decap_8 FILLER_66_138 ();
 sg13g2_fill_2 FILLER_66_159 ();
 sg13g2_fill_2 FILLER_66_197 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_decap_8 FILLER_66_204 ();
 sg13g2_decap_4 FILLER_66_211 ();
 sg13g2_decap_4 FILLER_66_251 ();
 sg13g2_fill_1 FILLER_66_255 ();
 sg13g2_decap_8 FILLER_66_284 ();
 sg13g2_decap_8 FILLER_66_291 ();
 sg13g2_fill_2 FILLER_66_298 ();
 sg13g2_decap_8 FILLER_66_304 ();
 sg13g2_decap_4 FILLER_66_311 ();
 sg13g2_fill_2 FILLER_66_315 ();
 sg13g2_decap_8 FILLER_66_330 ();
 sg13g2_fill_2 FILLER_66_337 ();
 sg13g2_fill_1 FILLER_66_339 ();
 sg13g2_fill_2 FILLER_66_344 ();
 sg13g2_decap_8 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_393 ();
 sg13g2_decap_8 FILLER_66_400 ();
 sg13g2_decap_8 FILLER_66_411 ();
 sg13g2_decap_8 FILLER_66_418 ();
 sg13g2_decap_8 FILLER_66_425 ();
 sg13g2_decap_8 FILLER_66_432 ();
 sg13g2_decap_8 FILLER_66_439 ();
 sg13g2_decap_4 FILLER_66_446 ();
 sg13g2_fill_2 FILLER_66_450 ();
 sg13g2_fill_2 FILLER_66_461 ();
 sg13g2_fill_1 FILLER_66_463 ();
 sg13g2_fill_2 FILLER_66_510 ();
 sg13g2_fill_1 FILLER_66_512 ();
 sg13g2_fill_2 FILLER_66_520 ();
 sg13g2_fill_1 FILLER_66_522 ();
 sg13g2_fill_1 FILLER_66_550 ();
 sg13g2_decap_8 FILLER_66_569 ();
 sg13g2_decap_4 FILLER_66_576 ();
 sg13g2_fill_1 FILLER_66_580 ();
 sg13g2_decap_8 FILLER_66_590 ();
 sg13g2_decap_8 FILLER_66_597 ();
 sg13g2_decap_8 FILLER_66_604 ();
 sg13g2_fill_2 FILLER_66_611 ();
 sg13g2_decap_8 FILLER_66_640 ();
 sg13g2_decap_8 FILLER_66_647 ();
 sg13g2_decap_8 FILLER_66_654 ();
 sg13g2_fill_2 FILLER_66_661 ();
 sg13g2_decap_8 FILLER_66_726 ();
 sg13g2_decap_4 FILLER_66_733 ();
 sg13g2_decap_8 FILLER_66_773 ();
 sg13g2_decap_8 FILLER_66_780 ();
 sg13g2_fill_2 FILLER_66_787 ();
 sg13g2_fill_1 FILLER_66_789 ();
 sg13g2_fill_1 FILLER_66_836 ();
 sg13g2_decap_8 FILLER_66_850 ();
 sg13g2_decap_8 FILLER_66_857 ();
 sg13g2_decap_4 FILLER_66_864 ();
 sg13g2_fill_2 FILLER_66_868 ();
 sg13g2_fill_1 FILLER_66_883 ();
 sg13g2_fill_2 FILLER_66_903 ();
 sg13g2_decap_8 FILLER_66_927 ();
 sg13g2_decap_8 FILLER_66_934 ();
 sg13g2_decap_8 FILLER_66_941 ();
 sg13g2_decap_8 FILLER_66_948 ();
 sg13g2_decap_8 FILLER_66_955 ();
 sg13g2_decap_8 FILLER_66_962 ();
 sg13g2_decap_8 FILLER_66_969 ();
 sg13g2_fill_2 FILLER_66_976 ();
 sg13g2_decap_4 FILLER_66_991 ();
 sg13g2_fill_1 FILLER_66_995 ();
 sg13g2_decap_8 FILLER_66_1018 ();
 sg13g2_decap_8 FILLER_66_1025 ();
 sg13g2_decap_8 FILLER_66_1032 ();
 sg13g2_decap_8 FILLER_66_1039 ();
 sg13g2_decap_8 FILLER_66_1046 ();
 sg13g2_fill_2 FILLER_66_1053 ();
 sg13g2_decap_8 FILLER_66_1086 ();
 sg13g2_fill_2 FILLER_66_1093 ();
 sg13g2_fill_1 FILLER_66_1095 ();
 sg13g2_decap_8 FILLER_66_1160 ();
 sg13g2_fill_2 FILLER_66_1194 ();
 sg13g2_fill_2 FILLER_66_1261 ();
 sg13g2_fill_1 FILLER_66_1263 ();
 sg13g2_fill_2 FILLER_66_1277 ();
 sg13g2_fill_1 FILLER_66_1279 ();
 sg13g2_fill_1 FILLER_66_1298 ();
 sg13g2_fill_1 FILLER_66_1308 ();
 sg13g2_decap_4 FILLER_66_1318 ();
 sg13g2_decap_4 FILLER_66_1356 ();
 sg13g2_fill_2 FILLER_66_1412 ();
 sg13g2_fill_1 FILLER_66_1429 ();
 sg13g2_fill_1 FILLER_66_1435 ();
 sg13g2_fill_2 FILLER_66_1455 ();
 sg13g2_decap_8 FILLER_66_1475 ();
 sg13g2_fill_1 FILLER_66_1482 ();
 sg13g2_decap_8 FILLER_66_1519 ();
 sg13g2_decap_8 FILLER_66_1526 ();
 sg13g2_fill_2 FILLER_66_1533 ();
 sg13g2_fill_1 FILLER_66_1552 ();
 sg13g2_decap_8 FILLER_66_1584 ();
 sg13g2_decap_8 FILLER_66_1628 ();
 sg13g2_decap_8 FILLER_66_1635 ();
 sg13g2_decap_8 FILLER_66_1642 ();
 sg13g2_decap_8 FILLER_66_1649 ();
 sg13g2_decap_4 FILLER_66_1662 ();
 sg13g2_fill_2 FILLER_66_1666 ();
 sg13g2_fill_1 FILLER_66_1694 ();
 sg13g2_fill_1 FILLER_66_1709 ();
 sg13g2_decap_8 FILLER_66_1742 ();
 sg13g2_decap_8 FILLER_66_1749 ();
 sg13g2_decap_4 FILLER_66_1756 ();
 sg13g2_fill_1 FILLER_66_1760 ();
 sg13g2_fill_2 FILLER_66_1788 ();
 sg13g2_fill_1 FILLER_66_1790 ();
 sg13g2_decap_8 FILLER_66_1797 ();
 sg13g2_fill_1 FILLER_66_1804 ();
 sg13g2_decap_4 FILLER_66_1811 ();
 sg13g2_fill_2 FILLER_66_1815 ();
 sg13g2_decap_4 FILLER_66_1822 ();
 sg13g2_decap_8 FILLER_66_1832 ();
 sg13g2_decap_8 FILLER_66_1839 ();
 sg13g2_decap_4 FILLER_66_1846 ();
 sg13g2_fill_2 FILLER_66_1850 ();
 sg13g2_fill_2 FILLER_66_1891 ();
 sg13g2_fill_1 FILLER_66_1893 ();
 sg13g2_fill_2 FILLER_66_1931 ();
 sg13g2_fill_1 FILLER_66_1933 ();
 sg13g2_decap_8 FILLER_66_1944 ();
 sg13g2_decap_8 FILLER_66_1951 ();
 sg13g2_decap_8 FILLER_66_1958 ();
 sg13g2_decap_8 FILLER_66_1973 ();
 sg13g2_fill_1 FILLER_66_1980 ();
 sg13g2_fill_2 FILLER_66_1986 ();
 sg13g2_fill_1 FILLER_66_1988 ();
 sg13g2_fill_2 FILLER_66_1997 ();
 sg13g2_fill_2 FILLER_66_2008 ();
 sg13g2_fill_2 FILLER_66_2015 ();
 sg13g2_fill_1 FILLER_66_2017 ();
 sg13g2_fill_2 FILLER_66_2031 ();
 sg13g2_fill_1 FILLER_66_2033 ();
 sg13g2_fill_1 FILLER_66_2053 ();
 sg13g2_decap_8 FILLER_66_2067 ();
 sg13g2_fill_2 FILLER_66_2074 ();
 sg13g2_fill_1 FILLER_66_2076 ();
 sg13g2_fill_1 FILLER_66_2082 ();
 sg13g2_decap_8 FILLER_66_2101 ();
 sg13g2_decap_4 FILLER_66_2121 ();
 sg13g2_decap_8 FILLER_66_2142 ();
 sg13g2_fill_2 FILLER_66_2149 ();
 sg13g2_fill_1 FILLER_66_2151 ();
 sg13g2_decap_8 FILLER_66_2161 ();
 sg13g2_decap_4 FILLER_66_2168 ();
 sg13g2_fill_2 FILLER_66_2185 ();
 sg13g2_fill_1 FILLER_66_2192 ();
 sg13g2_decap_8 FILLER_66_2198 ();
 sg13g2_fill_2 FILLER_66_2205 ();
 sg13g2_decap_8 FILLER_66_2215 ();
 sg13g2_decap_8 FILLER_66_2222 ();
 sg13g2_decap_8 FILLER_66_2229 ();
 sg13g2_decap_4 FILLER_66_2236 ();
 sg13g2_fill_2 FILLER_66_2240 ();
 sg13g2_decap_8 FILLER_66_2247 ();
 sg13g2_decap_4 FILLER_66_2254 ();
 sg13g2_decap_4 FILLER_66_2283 ();
 sg13g2_decap_8 FILLER_66_2300 ();
 sg13g2_decap_8 FILLER_66_2307 ();
 sg13g2_decap_8 FILLER_66_2314 ();
 sg13g2_decap_8 FILLER_66_2321 ();
 sg13g2_decap_4 FILLER_66_2328 ();
 sg13g2_fill_1 FILLER_66_2332 ();
 sg13g2_decap_8 FILLER_66_2343 ();
 sg13g2_decap_4 FILLER_66_2350 ();
 sg13g2_decap_8 FILLER_66_2359 ();
 sg13g2_decap_4 FILLER_66_2366 ();
 sg13g2_decap_8 FILLER_66_2404 ();
 sg13g2_decap_8 FILLER_66_2411 ();
 sg13g2_decap_8 FILLER_66_2418 ();
 sg13g2_decap_4 FILLER_66_2425 ();
 sg13g2_decap_8 FILLER_66_2487 ();
 sg13g2_decap_8 FILLER_66_2494 ();
 sg13g2_decap_8 FILLER_66_2501 ();
 sg13g2_decap_8 FILLER_66_2545 ();
 sg13g2_decap_4 FILLER_66_2552 ();
 sg13g2_decap_8 FILLER_66_2591 ();
 sg13g2_decap_8 FILLER_66_2598 ();
 sg13g2_decap_8 FILLER_66_2605 ();
 sg13g2_decap_4 FILLER_66_2612 ();
 sg13g2_fill_1 FILLER_66_2616 ();
 sg13g2_decap_8 FILLER_66_2675 ();
 sg13g2_decap_4 FILLER_66_2682 ();
 sg13g2_fill_2 FILLER_66_2686 ();
 sg13g2_decap_8 FILLER_66_2715 ();
 sg13g2_decap_4 FILLER_66_2722 ();
 sg13g2_decap_8 FILLER_66_2730 ();
 sg13g2_decap_8 FILLER_66_2737 ();
 sg13g2_decap_8 FILLER_66_2744 ();
 sg13g2_fill_1 FILLER_66_2751 ();
 sg13g2_fill_2 FILLER_66_2766 ();
 sg13g2_decap_8 FILLER_66_2781 ();
 sg13g2_decap_8 FILLER_66_2788 ();
 sg13g2_decap_8 FILLER_66_2795 ();
 sg13g2_fill_2 FILLER_66_2802 ();
 sg13g2_fill_1 FILLER_66_2818 ();
 sg13g2_fill_1 FILLER_66_2829 ();
 sg13g2_decap_8 FILLER_66_2839 ();
 sg13g2_decap_4 FILLER_66_2846 ();
 sg13g2_decap_8 FILLER_66_2863 ();
 sg13g2_fill_2 FILLER_66_2870 ();
 sg13g2_fill_1 FILLER_66_2872 ();
 sg13g2_decap_8 FILLER_66_2910 ();
 sg13g2_decap_4 FILLER_66_2917 ();
 sg13g2_decap_8 FILLER_66_2940 ();
 sg13g2_fill_1 FILLER_66_2947 ();
 sg13g2_decap_4 FILLER_66_2969 ();
 sg13g2_fill_1 FILLER_66_2973 ();
 sg13g2_decap_8 FILLER_66_2987 ();
 sg13g2_fill_2 FILLER_66_2994 ();
 sg13g2_fill_1 FILLER_66_2996 ();
 sg13g2_decap_8 FILLER_66_3010 ();
 sg13g2_decap_8 FILLER_66_3017 ();
 sg13g2_decap_4 FILLER_66_3024 ();
 sg13g2_fill_1 FILLER_66_3038 ();
 sg13g2_decap_8 FILLER_66_3061 ();
 sg13g2_decap_8 FILLER_66_3068 ();
 sg13g2_fill_2 FILLER_66_3075 ();
 sg13g2_fill_1 FILLER_66_3077 ();
 sg13g2_decap_8 FILLER_66_3115 ();
 sg13g2_decap_8 FILLER_66_3122 ();
 sg13g2_decap_4 FILLER_66_3129 ();
 sg13g2_fill_1 FILLER_66_3133 ();
 sg13g2_decap_8 FILLER_66_3173 ();
 sg13g2_decap_8 FILLER_66_3180 ();
 sg13g2_decap_4 FILLER_66_3187 ();
 sg13g2_fill_1 FILLER_66_3191 ();
 sg13g2_decap_8 FILLER_66_3242 ();
 sg13g2_fill_2 FILLER_66_3249 ();
 sg13g2_decap_8 FILLER_66_3278 ();
 sg13g2_decap_8 FILLER_66_3285 ();
 sg13g2_decap_8 FILLER_66_3292 ();
 sg13g2_fill_2 FILLER_66_3299 ();
 sg13g2_fill_1 FILLER_66_3301 ();
 sg13g2_fill_2 FILLER_66_3306 ();
 sg13g2_fill_1 FILLER_66_3339 ();
 sg13g2_decap_4 FILLER_66_3353 ();
 sg13g2_fill_2 FILLER_66_3357 ();
 sg13g2_fill_2 FILLER_66_3432 ();
 sg13g2_decap_8 FILLER_66_3460 ();
 sg13g2_fill_1 FILLER_66_3467 ();
 sg13g2_fill_2 FILLER_66_3481 ();
 sg13g2_fill_1 FILLER_66_3492 ();
 sg13g2_decap_4 FILLER_66_3503 ();
 sg13g2_fill_1 FILLER_66_3534 ();
 sg13g2_fill_2 FILLER_66_3575 ();
 sg13g2_fill_1 FILLER_66_3577 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_2 FILLER_67_14 ();
 sg13g2_fill_1 FILLER_67_16 ();
 sg13g2_fill_2 FILLER_67_74 ();
 sg13g2_fill_1 FILLER_67_76 ();
 sg13g2_fill_2 FILLER_67_109 ();
 sg13g2_fill_2 FILLER_67_121 ();
 sg13g2_fill_1 FILLER_67_123 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_fill_2 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_216 ();
 sg13g2_decap_8 FILLER_67_223 ();
 sg13g2_decap_8 FILLER_67_230 ();
 sg13g2_decap_4 FILLER_67_237 ();
 sg13g2_fill_1 FILLER_67_241 ();
 sg13g2_fill_1 FILLER_67_269 ();
 sg13g2_fill_1 FILLER_67_292 ();
 sg13g2_decap_8 FILLER_67_324 ();
 sg13g2_decap_4 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_384 ();
 sg13g2_decap_8 FILLER_67_391 ();
 sg13g2_decap_4 FILLER_67_398 ();
 sg13g2_fill_1 FILLER_67_402 ();
 sg13g2_decap_8 FILLER_67_439 ();
 sg13g2_decap_8 FILLER_67_446 ();
 sg13g2_decap_4 FILLER_67_453 ();
 sg13g2_fill_1 FILLER_67_457 ();
 sg13g2_fill_1 FILLER_67_485 ();
 sg13g2_decap_8 FILLER_67_499 ();
 sg13g2_decap_4 FILLER_67_506 ();
 sg13g2_decap_8 FILLER_67_542 ();
 sg13g2_fill_2 FILLER_67_549 ();
 sg13g2_fill_1 FILLER_67_551 ();
 sg13g2_fill_1 FILLER_67_611 ();
 sg13g2_decap_8 FILLER_67_639 ();
 sg13g2_decap_8 FILLER_67_646 ();
 sg13g2_decap_8 FILLER_67_653 ();
 sg13g2_decap_8 FILLER_67_660 ();
 sg13g2_fill_2 FILLER_67_667 ();
 sg13g2_decap_8 FILLER_67_696 ();
 sg13g2_fill_2 FILLER_67_703 ();
 sg13g2_decap_8 FILLER_67_714 ();
 sg13g2_decap_8 FILLER_67_721 ();
 sg13g2_decap_8 FILLER_67_728 ();
 sg13g2_decap_4 FILLER_67_735 ();
 sg13g2_fill_1 FILLER_67_739 ();
 sg13g2_fill_1 FILLER_67_753 ();
 sg13g2_fill_1 FILLER_67_763 ();
 sg13g2_decap_8 FILLER_67_768 ();
 sg13g2_decap_8 FILLER_67_775 ();
 sg13g2_decap_8 FILLER_67_782 ();
 sg13g2_decap_8 FILLER_67_817 ();
 sg13g2_decap_8 FILLER_67_850 ();
 sg13g2_fill_2 FILLER_67_857 ();
 sg13g2_fill_1 FILLER_67_859 ();
 sg13g2_fill_1 FILLER_67_887 ();
 sg13g2_fill_1 FILLER_67_910 ();
 sg13g2_decap_8 FILLER_67_929 ();
 sg13g2_decap_8 FILLER_67_936 ();
 sg13g2_decap_8 FILLER_67_943 ();
 sg13g2_fill_2 FILLER_67_950 ();
 sg13g2_fill_1 FILLER_67_952 ();
 sg13g2_decap_8 FILLER_67_980 ();
 sg13g2_decap_4 FILLER_67_987 ();
 sg13g2_decap_8 FILLER_67_1000 ();
 sg13g2_fill_2 FILLER_67_1007 ();
 sg13g2_decap_8 FILLER_67_1013 ();
 sg13g2_decap_4 FILLER_67_1020 ();
 sg13g2_fill_2 FILLER_67_1024 ();
 sg13g2_fill_2 FILLER_67_1054 ();
 sg13g2_fill_1 FILLER_67_1056 ();
 sg13g2_decap_8 FILLER_67_1084 ();
 sg13g2_decap_8 FILLER_67_1091 ();
 sg13g2_decap_8 FILLER_67_1098 ();
 sg13g2_decap_4 FILLER_67_1105 ();
 sg13g2_fill_2 FILLER_67_1137 ();
 sg13g2_decap_8 FILLER_67_1152 ();
 sg13g2_fill_2 FILLER_67_1159 ();
 sg13g2_fill_1 FILLER_67_1161 ();
 sg13g2_fill_1 FILLER_67_1205 ();
 sg13g2_decap_8 FILLER_67_1227 ();
 sg13g2_decap_8 FILLER_67_1234 ();
 sg13g2_fill_1 FILLER_67_1241 ();
 sg13g2_decap_4 FILLER_67_1251 ();
 sg13g2_fill_1 FILLER_67_1255 ();
 sg13g2_fill_1 FILLER_67_1295 ();
 sg13g2_decap_8 FILLER_67_1309 ();
 sg13g2_decap_8 FILLER_67_1316 ();
 sg13g2_decap_4 FILLER_67_1323 ();
 sg13g2_fill_1 FILLER_67_1327 ();
 sg13g2_fill_1 FILLER_67_1345 ();
 sg13g2_decap_8 FILLER_67_1352 ();
 sg13g2_decap_8 FILLER_67_1359 ();
 sg13g2_decap_8 FILLER_67_1366 ();
 sg13g2_fill_2 FILLER_67_1373 ();
 sg13g2_fill_1 FILLER_67_1375 ();
 sg13g2_decap_4 FILLER_67_1408 ();
 sg13g2_fill_1 FILLER_67_1422 ();
 sg13g2_fill_2 FILLER_67_1432 ();
 sg13g2_fill_1 FILLER_67_1434 ();
 sg13g2_fill_2 FILLER_67_1487 ();
 sg13g2_fill_1 FILLER_67_1498 ();
 sg13g2_fill_2 FILLER_67_1508 ();
 sg13g2_decap_4 FILLER_67_1514 ();
 sg13g2_decap_8 FILLER_67_1522 ();
 sg13g2_fill_2 FILLER_67_1529 ();
 sg13g2_decap_4 FILLER_67_1572 ();
 sg13g2_fill_1 FILLER_67_1576 ();
 sg13g2_decap_8 FILLER_67_1627 ();
 sg13g2_decap_8 FILLER_67_1634 ();
 sg13g2_decap_4 FILLER_67_1641 ();
 sg13g2_decap_8 FILLER_67_1673 ();
 sg13g2_decap_4 FILLER_67_1680 ();
 sg13g2_fill_1 FILLER_67_1684 ();
 sg13g2_fill_2 FILLER_67_1713 ();
 sg13g2_fill_1 FILLER_67_1715 ();
 sg13g2_decap_4 FILLER_67_1753 ();
 sg13g2_fill_1 FILLER_67_1778 ();
 sg13g2_decap_8 FILLER_67_1801 ();
 sg13g2_fill_2 FILLER_67_1825 ();
 sg13g2_fill_1 FILLER_67_1827 ();
 sg13g2_decap_4 FILLER_67_1832 ();
 sg13g2_decap_8 FILLER_67_1862 ();
 sg13g2_fill_1 FILLER_67_1869 ();
 sg13g2_fill_2 FILLER_67_1882 ();
 sg13g2_fill_1 FILLER_67_1884 ();
 sg13g2_decap_8 FILLER_67_1898 ();
 sg13g2_fill_1 FILLER_67_1905 ();
 sg13g2_decap_8 FILLER_67_1910 ();
 sg13g2_decap_8 FILLER_67_1917 ();
 sg13g2_fill_1 FILLER_67_1924 ();
 sg13g2_decap_8 FILLER_67_1951 ();
 sg13g2_decap_4 FILLER_67_1958 ();
 sg13g2_fill_1 FILLER_67_1962 ();
 sg13g2_decap_4 FILLER_67_1971 ();
 sg13g2_fill_1 FILLER_67_1975 ();
 sg13g2_fill_2 FILLER_67_1995 ();
 sg13g2_fill_2 FILLER_67_2005 ();
 sg13g2_decap_8 FILLER_67_2013 ();
 sg13g2_decap_4 FILLER_67_2020 ();
 sg13g2_fill_2 FILLER_67_2024 ();
 sg13g2_fill_2 FILLER_67_2041 ();
 sg13g2_fill_1 FILLER_67_2043 ();
 sg13g2_decap_8 FILLER_67_2057 ();
 sg13g2_decap_8 FILLER_67_2064 ();
 sg13g2_fill_2 FILLER_67_2071 ();
 sg13g2_fill_1 FILLER_67_2073 ();
 sg13g2_decap_8 FILLER_67_2092 ();
 sg13g2_decap_8 FILLER_67_2099 ();
 sg13g2_decap_8 FILLER_67_2106 ();
 sg13g2_decap_8 FILLER_67_2113 ();
 sg13g2_decap_8 FILLER_67_2120 ();
 sg13g2_decap_8 FILLER_67_2127 ();
 sg13g2_decap_8 FILLER_67_2134 ();
 sg13g2_fill_2 FILLER_67_2141 ();
 sg13g2_fill_1 FILLER_67_2143 ();
 sg13g2_fill_1 FILLER_67_2157 ();
 sg13g2_decap_8 FILLER_67_2168 ();
 sg13g2_decap_8 FILLER_67_2175 ();
 sg13g2_decap_8 FILLER_67_2182 ();
 sg13g2_decap_4 FILLER_67_2189 ();
 sg13g2_fill_2 FILLER_67_2193 ();
 sg13g2_decap_4 FILLER_67_2200 ();
 sg13g2_fill_1 FILLER_67_2204 ();
 sg13g2_fill_1 FILLER_67_2210 ();
 sg13g2_decap_8 FILLER_67_2217 ();
 sg13g2_decap_8 FILLER_67_2224 ();
 sg13g2_decap_8 FILLER_67_2238 ();
 sg13g2_fill_1 FILLER_67_2245 ();
 sg13g2_decap_8 FILLER_67_2275 ();
 sg13g2_decap_8 FILLER_67_2282 ();
 sg13g2_fill_2 FILLER_67_2289 ();
 sg13g2_fill_1 FILLER_67_2291 ();
 sg13g2_fill_2 FILLER_67_2307 ();
 sg13g2_fill_1 FILLER_67_2309 ();
 sg13g2_decap_8 FILLER_67_2320 ();
 sg13g2_decap_8 FILLER_67_2327 ();
 sg13g2_decap_8 FILLER_67_2334 ();
 sg13g2_decap_4 FILLER_67_2341 ();
 sg13g2_fill_1 FILLER_67_2345 ();
 sg13g2_decap_8 FILLER_67_2361 ();
 sg13g2_decap_4 FILLER_67_2368 ();
 sg13g2_fill_1 FILLER_67_2372 ();
 sg13g2_decap_8 FILLER_67_2406 ();
 sg13g2_decap_8 FILLER_67_2413 ();
 sg13g2_decap_8 FILLER_67_2420 ();
 sg13g2_decap_8 FILLER_67_2427 ();
 sg13g2_fill_2 FILLER_67_2434 ();
 sg13g2_fill_2 FILLER_67_2446 ();
 sg13g2_fill_1 FILLER_67_2448 ();
 sg13g2_decap_8 FILLER_67_2485 ();
 sg13g2_fill_2 FILLER_67_2492 ();
 sg13g2_decap_8 FILLER_67_2541 ();
 sg13g2_decap_8 FILLER_67_2548 ();
 sg13g2_decap_8 FILLER_67_2555 ();
 sg13g2_decap_4 FILLER_67_2562 ();
 sg13g2_fill_2 FILLER_67_2566 ();
 sg13g2_decap_8 FILLER_67_2595 ();
 sg13g2_fill_2 FILLER_67_2602 ();
 sg13g2_fill_1 FILLER_67_2604 ();
 sg13g2_fill_2 FILLER_67_2642 ();
 sg13g2_fill_1 FILLER_67_2644 ();
 sg13g2_decap_8 FILLER_67_2666 ();
 sg13g2_fill_1 FILLER_67_2673 ();
 sg13g2_decap_8 FILLER_67_2732 ();
 sg13g2_decap_8 FILLER_67_2739 ();
 sg13g2_fill_1 FILLER_67_2746 ();
 sg13g2_decap_8 FILLER_67_2784 ();
 sg13g2_decap_8 FILLER_67_2791 ();
 sg13g2_decap_8 FILLER_67_2798 ();
 sg13g2_decap_8 FILLER_67_2805 ();
 sg13g2_decap_8 FILLER_67_2839 ();
 sg13g2_decap_8 FILLER_67_2846 ();
 sg13g2_decap_8 FILLER_67_2853 ();
 sg13g2_decap_8 FILLER_67_2906 ();
 sg13g2_decap_8 FILLER_67_2913 ();
 sg13g2_decap_8 FILLER_67_2920 ();
 sg13g2_decap_4 FILLER_67_2927 ();
 sg13g2_fill_1 FILLER_67_2931 ();
 sg13g2_decap_8 FILLER_67_2973 ();
 sg13g2_decap_4 FILLER_67_2980 ();
 sg13g2_fill_2 FILLER_67_2984 ();
 sg13g2_fill_2 FILLER_67_2999 ();
 sg13g2_fill_1 FILLER_67_3001 ();
 sg13g2_fill_2 FILLER_67_3006 ();
 sg13g2_decap_8 FILLER_67_3055 ();
 sg13g2_fill_2 FILLER_67_3120 ();
 sg13g2_fill_1 FILLER_67_3122 ();
 sg13g2_decap_4 FILLER_67_3136 ();
 sg13g2_decap_8 FILLER_67_3178 ();
 sg13g2_decap_8 FILLER_67_3185 ();
 sg13g2_fill_1 FILLER_67_3192 ();
 sg13g2_decap_8 FILLER_67_3233 ();
 sg13g2_decap_8 FILLER_67_3240 ();
 sg13g2_fill_1 FILLER_67_3247 ();
 sg13g2_decap_8 FILLER_67_3283 ();
 sg13g2_decap_8 FILLER_67_3290 ();
 sg13g2_decap_8 FILLER_67_3297 ();
 sg13g2_decap_4 FILLER_67_3304 ();
 sg13g2_fill_2 FILLER_67_3308 ();
 sg13g2_decap_8 FILLER_67_3351 ();
 sg13g2_decap_4 FILLER_67_3358 ();
 sg13g2_fill_2 FILLER_67_3362 ();
 sg13g2_fill_1 FILLER_67_3368 ();
 sg13g2_decap_4 FILLER_67_3409 ();
 sg13g2_fill_2 FILLER_67_3413 ();
 sg13g2_decap_8 FILLER_67_3424 ();
 sg13g2_fill_2 FILLER_67_3431 ();
 sg13g2_decap_8 FILLER_67_3481 ();
 sg13g2_decap_8 FILLER_67_3488 ();
 sg13g2_fill_2 FILLER_67_3495 ();
 sg13g2_fill_1 FILLER_67_3497 ();
 sg13g2_fill_2 FILLER_67_3516 ();
 sg13g2_decap_8 FILLER_67_3522 ();
 sg13g2_decap_4 FILLER_67_3529 ();
 sg13g2_decap_8 FILLER_67_3570 ();
 sg13g2_fill_1 FILLER_67_3577 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_47 ();
 sg13g2_fill_1 FILLER_68_67 ();
 sg13g2_fill_1 FILLER_68_81 ();
 sg13g2_fill_2 FILLER_68_133 ();
 sg13g2_fill_1 FILLER_68_135 ();
 sg13g2_fill_2 FILLER_68_146 ();
 sg13g2_fill_1 FILLER_68_148 ();
 sg13g2_decap_4 FILLER_68_168 ();
 sg13g2_fill_1 FILLER_68_172 ();
 sg13g2_fill_1 FILLER_68_209 ();
 sg13g2_decap_4 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_236 ();
 sg13g2_decap_4 FILLER_68_243 ();
 sg13g2_fill_2 FILLER_68_295 ();
 sg13g2_fill_2 FILLER_68_333 ();
 sg13g2_decap_8 FILLER_68_387 ();
 sg13g2_fill_2 FILLER_68_394 ();
 sg13g2_fill_1 FILLER_68_396 ();
 sg13g2_decap_8 FILLER_68_447 ();
 sg13g2_decap_4 FILLER_68_454 ();
 sg13g2_decap_8 FILLER_68_485 ();
 sg13g2_decap_8 FILLER_68_492 ();
 sg13g2_decap_8 FILLER_68_499 ();
 sg13g2_decap_8 FILLER_68_506 ();
 sg13g2_decap_8 FILLER_68_513 ();
 sg13g2_decap_4 FILLER_68_520 ();
 sg13g2_fill_1 FILLER_68_524 ();
 sg13g2_decap_8 FILLER_68_530 ();
 sg13g2_decap_8 FILLER_68_537 ();
 sg13g2_decap_8 FILLER_68_544 ();
 sg13g2_decap_8 FILLER_68_551 ();
 sg13g2_decap_8 FILLER_68_558 ();
 sg13g2_fill_2 FILLER_68_565 ();
 sg13g2_decap_8 FILLER_68_573 ();
 sg13g2_decap_8 FILLER_68_580 ();
 sg13g2_decap_8 FILLER_68_587 ();
 sg13g2_decap_8 FILLER_68_643 ();
 sg13g2_decap_8 FILLER_68_650 ();
 sg13g2_decap_4 FILLER_68_657 ();
 sg13g2_fill_1 FILLER_68_661 ();
 sg13g2_decap_8 FILLER_68_689 ();
 sg13g2_decap_8 FILLER_68_696 ();
 sg13g2_decap_8 FILLER_68_703 ();
 sg13g2_fill_2 FILLER_68_710 ();
 sg13g2_fill_1 FILLER_68_712 ();
 sg13g2_decap_8 FILLER_68_717 ();
 sg13g2_decap_8 FILLER_68_724 ();
 sg13g2_decap_4 FILLER_68_731 ();
 sg13g2_fill_1 FILLER_68_735 ();
 sg13g2_fill_2 FILLER_68_749 ();
 sg13g2_fill_1 FILLER_68_751 ();
 sg13g2_decap_8 FILLER_68_756 ();
 sg13g2_decap_8 FILLER_68_763 ();
 sg13g2_decap_4 FILLER_68_770 ();
 sg13g2_fill_1 FILLER_68_774 ();
 sg13g2_fill_2 FILLER_68_830 ();
 sg13g2_fill_1 FILLER_68_943 ();
 sg13g2_fill_1 FILLER_68_972 ();
 sg13g2_fill_2 FILLER_68_1001 ();
 sg13g2_fill_1 FILLER_68_1003 ();
 sg13g2_decap_8 FILLER_68_1017 ();
 sg13g2_fill_2 FILLER_68_1052 ();
 sg13g2_decap_8 FILLER_68_1063 ();
 sg13g2_decap_4 FILLER_68_1070 ();
 sg13g2_decap_8 FILLER_68_1087 ();
 sg13g2_decap_8 FILLER_68_1094 ();
 sg13g2_decap_4 FILLER_68_1101 ();
 sg13g2_fill_2 FILLER_68_1105 ();
 sg13g2_fill_1 FILLER_68_1123 ();
 sg13g2_decap_8 FILLER_68_1137 ();
 sg13g2_decap_8 FILLER_68_1144 ();
 sg13g2_fill_2 FILLER_68_1151 ();
 sg13g2_decap_4 FILLER_68_1166 ();
 sg13g2_fill_1 FILLER_68_1170 ();
 sg13g2_decap_8 FILLER_68_1206 ();
 sg13g2_decap_8 FILLER_68_1213 ();
 sg13g2_decap_8 FILLER_68_1220 ();
 sg13g2_fill_2 FILLER_68_1227 ();
 sg13g2_decap_4 FILLER_68_1232 ();
 sg13g2_fill_2 FILLER_68_1236 ();
 sg13g2_fill_1 FILLER_68_1247 ();
 sg13g2_fill_1 FILLER_68_1255 ();
 sg13g2_decap_4 FILLER_68_1270 ();
 sg13g2_decap_8 FILLER_68_1314 ();
 sg13g2_fill_2 FILLER_68_1327 ();
 sg13g2_decap_8 FILLER_68_1342 ();
 sg13g2_decap_4 FILLER_68_1349 ();
 sg13g2_fill_1 FILLER_68_1353 ();
 sg13g2_fill_1 FILLER_68_1426 ();
 sg13g2_decap_8 FILLER_68_1482 ();
 sg13g2_fill_2 FILLER_68_1536 ();
 sg13g2_fill_1 FILLER_68_1538 ();
 sg13g2_decap_8 FILLER_68_1574 ();
 sg13g2_decap_8 FILLER_68_1581 ();
 sg13g2_fill_1 FILLER_68_1588 ();
 sg13g2_fill_2 FILLER_68_1635 ();
 sg13g2_fill_1 FILLER_68_1637 ();
 sg13g2_fill_2 FILLER_68_1642 ();
 sg13g2_fill_1 FILLER_68_1644 ();
 sg13g2_decap_8 FILLER_68_1673 ();
 sg13g2_decap_8 FILLER_68_1680 ();
 sg13g2_decap_8 FILLER_68_1687 ();
 sg13g2_decap_8 FILLER_68_1694 ();
 sg13g2_decap_8 FILLER_68_1710 ();
 sg13g2_decap_8 FILLER_68_1717 ();
 sg13g2_decap_4 FILLER_68_1724 ();
 sg13g2_fill_1 FILLER_68_1728 ();
 sg13g2_decap_8 FILLER_68_1739 ();
 sg13g2_decap_4 FILLER_68_1746 ();
 sg13g2_decap_8 FILLER_68_1802 ();
 sg13g2_fill_2 FILLER_68_1809 ();
 sg13g2_fill_1 FILLER_68_1811 ();
 sg13g2_decap_8 FILLER_68_1816 ();
 sg13g2_decap_4 FILLER_68_1823 ();
 sg13g2_fill_1 FILLER_68_1837 ();
 sg13g2_decap_8 FILLER_68_1844 ();
 sg13g2_decap_8 FILLER_68_1855 ();
 sg13g2_decap_8 FILLER_68_1862 ();
 sg13g2_decap_8 FILLER_68_1869 ();
 sg13g2_fill_2 FILLER_68_1876 ();
 sg13g2_fill_1 FILLER_68_1878 ();
 sg13g2_decap_8 FILLER_68_1890 ();
 sg13g2_decap_4 FILLER_68_1897 ();
 sg13g2_fill_1 FILLER_68_1901 ();
 sg13g2_decap_8 FILLER_68_1915 ();
 sg13g2_decap_4 FILLER_68_1926 ();
 sg13g2_fill_2 FILLER_68_1930 ();
 sg13g2_decap_4 FILLER_68_1936 ();
 sg13g2_fill_2 FILLER_68_1940 ();
 sg13g2_decap_8 FILLER_68_1950 ();
 sg13g2_fill_2 FILLER_68_1981 ();
 sg13g2_fill_1 FILLER_68_1983 ();
 sg13g2_fill_2 FILLER_68_1998 ();
 sg13g2_fill_1 FILLER_68_2000 ();
 sg13g2_fill_2 FILLER_68_2006 ();
 sg13g2_fill_1 FILLER_68_2008 ();
 sg13g2_decap_8 FILLER_68_2014 ();
 sg13g2_decap_4 FILLER_68_2021 ();
 sg13g2_decap_4 FILLER_68_2031 ();
 sg13g2_decap_8 FILLER_68_2048 ();
 sg13g2_decap_8 FILLER_68_2055 ();
 sg13g2_fill_1 FILLER_68_2062 ();
 sg13g2_decap_8 FILLER_68_2075 ();
 sg13g2_fill_2 FILLER_68_2082 ();
 sg13g2_fill_1 FILLER_68_2084 ();
 sg13g2_decap_8 FILLER_68_2103 ();
 sg13g2_fill_1 FILLER_68_2110 ();
 sg13g2_fill_2 FILLER_68_2123 ();
 sg13g2_decap_4 FILLER_68_2130 ();
 sg13g2_decap_8 FILLER_68_2139 ();
 sg13g2_decap_4 FILLER_68_2146 ();
 sg13g2_fill_1 FILLER_68_2150 ();
 sg13g2_decap_4 FILLER_68_2171 ();
 sg13g2_fill_1 FILLER_68_2175 ();
 sg13g2_decap_4 FILLER_68_2180 ();
 sg13g2_fill_1 FILLER_68_2184 ();
 sg13g2_decap_8 FILLER_68_2190 ();
 sg13g2_fill_2 FILLER_68_2197 ();
 sg13g2_fill_1 FILLER_68_2199 ();
 sg13g2_fill_1 FILLER_68_2223 ();
 sg13g2_fill_2 FILLER_68_2248 ();
 sg13g2_decap_8 FILLER_68_2265 ();
 sg13g2_decap_8 FILLER_68_2272 ();
 sg13g2_fill_1 FILLER_68_2279 ();
 sg13g2_fill_1 FILLER_68_2311 ();
 sg13g2_decap_8 FILLER_68_2317 ();
 sg13g2_decap_8 FILLER_68_2324 ();
 sg13g2_decap_8 FILLER_68_2331 ();
 sg13g2_fill_1 FILLER_68_2338 ();
 sg13g2_fill_1 FILLER_68_2353 ();
 sg13g2_decap_4 FILLER_68_2367 ();
 sg13g2_fill_1 FILLER_68_2371 ();
 sg13g2_fill_2 FILLER_68_2395 ();
 sg13g2_decap_8 FILLER_68_2415 ();
 sg13g2_decap_8 FILLER_68_2422 ();
 sg13g2_decap_8 FILLER_68_2429 ();
 sg13g2_decap_4 FILLER_68_2436 ();
 sg13g2_fill_2 FILLER_68_2440 ();
 sg13g2_decap_8 FILLER_68_2482 ();
 sg13g2_decap_8 FILLER_68_2489 ();
 sg13g2_decap_8 FILLER_68_2496 ();
 sg13g2_decap_8 FILLER_68_2547 ();
 sg13g2_decap_8 FILLER_68_2554 ();
 sg13g2_decap_8 FILLER_68_2561 ();
 sg13g2_fill_2 FILLER_68_2568 ();
 sg13g2_decap_8 FILLER_68_2578 ();
 sg13g2_decap_8 FILLER_68_2585 ();
 sg13g2_fill_2 FILLER_68_2592 ();
 sg13g2_fill_1 FILLER_68_2594 ();
 sg13g2_decap_8 FILLER_68_2608 ();
 sg13g2_fill_2 FILLER_68_2625 ();
 sg13g2_fill_1 FILLER_68_2627 ();
 sg13g2_decap_8 FILLER_68_2659 ();
 sg13g2_decap_8 FILLER_68_2666 ();
 sg13g2_decap_8 FILLER_68_2673 ();
 sg13g2_fill_2 FILLER_68_2680 ();
 sg13g2_fill_2 FILLER_68_2727 ();
 sg13g2_fill_1 FILLER_68_2738 ();
 sg13g2_decap_8 FILLER_68_2797 ();
 sg13g2_decap_4 FILLER_68_2804 ();
 sg13g2_fill_2 FILLER_68_2808 ();
 sg13g2_decap_8 FILLER_68_2837 ();
 sg13g2_decap_8 FILLER_68_2844 ();
 sg13g2_fill_2 FILLER_68_2851 ();
 sg13g2_fill_2 FILLER_68_2905 ();
 sg13g2_decap_8 FILLER_68_2920 ();
 sg13g2_fill_2 FILLER_68_2927 ();
 sg13g2_fill_1 FILLER_68_2929 ();
 sg13g2_decap_8 FILLER_68_2978 ();
 sg13g2_decap_8 FILLER_68_2985 ();
 sg13g2_decap_4 FILLER_68_2992 ();
 sg13g2_fill_1 FILLER_68_2996 ();
 sg13g2_decap_8 FILLER_68_3115 ();
 sg13g2_decap_8 FILLER_68_3122 ();
 sg13g2_decap_4 FILLER_68_3129 ();
 sg13g2_fill_1 FILLER_68_3133 ();
 sg13g2_decap_8 FILLER_68_3174 ();
 sg13g2_decap_8 FILLER_68_3181 ();
 sg13g2_decap_4 FILLER_68_3188 ();
 sg13g2_fill_2 FILLER_68_3192 ();
 sg13g2_decap_8 FILLER_68_3231 ();
 sg13g2_decap_4 FILLER_68_3238 ();
 sg13g2_fill_2 FILLER_68_3265 ();
 sg13g2_decap_4 FILLER_68_3301 ();
 sg13g2_decap_8 FILLER_68_3308 ();
 sg13g2_decap_8 FILLER_68_3315 ();
 sg13g2_fill_2 FILLER_68_3322 ();
 sg13g2_decap_4 FILLER_68_3338 ();
 sg13g2_decap_8 FILLER_68_3351 ();
 sg13g2_decap_8 FILLER_68_3358 ();
 sg13g2_decap_8 FILLER_68_3365 ();
 sg13g2_decap_4 FILLER_68_3372 ();
 sg13g2_fill_2 FILLER_68_3376 ();
 sg13g2_decap_8 FILLER_68_3406 ();
 sg13g2_decap_8 FILLER_68_3413 ();
 sg13g2_decap_8 FILLER_68_3420 ();
 sg13g2_fill_1 FILLER_68_3427 ();
 sg13g2_decap_8 FILLER_68_3465 ();
 sg13g2_decap_8 FILLER_68_3472 ();
 sg13g2_decap_8 FILLER_68_3479 ();
 sg13g2_decap_8 FILLER_68_3486 ();
 sg13g2_decap_8 FILLER_68_3493 ();
 sg13g2_decap_4 FILLER_68_3500 ();
 sg13g2_fill_1 FILLER_68_3504 ();
 sg13g2_decap_8 FILLER_68_3518 ();
 sg13g2_fill_2 FILLER_68_3525 ();
 sg13g2_fill_1 FILLER_68_3527 ();
 sg13g2_decap_8 FILLER_68_3565 ();
 sg13g2_decap_4 FILLER_68_3572 ();
 sg13g2_fill_2 FILLER_68_3576 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_58 ();
 sg13g2_decap_4 FILLER_69_65 ();
 sg13g2_fill_2 FILLER_69_69 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_118 ();
 sg13g2_fill_2 FILLER_69_125 ();
 sg13g2_decap_8 FILLER_69_162 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_210 ();
 sg13g2_decap_8 FILLER_69_229 ();
 sg13g2_fill_2 FILLER_69_268 ();
 sg13g2_fill_2 FILLER_69_293 ();
 sg13g2_fill_1 FILLER_69_333 ();
 sg13g2_fill_2 FILLER_69_428 ();
 sg13g2_fill_2 FILLER_69_445 ();
 sg13g2_fill_2 FILLER_69_474 ();
 sg13g2_fill_1 FILLER_69_476 ();
 sg13g2_decap_8 FILLER_69_495 ();
 sg13g2_decap_8 FILLER_69_506 ();
 sg13g2_decap_8 FILLER_69_513 ();
 sg13g2_fill_2 FILLER_69_533 ();
 sg13g2_decap_8 FILLER_69_539 ();
 sg13g2_decap_4 FILLER_69_546 ();
 sg13g2_decap_8 FILLER_69_554 ();
 sg13g2_decap_8 FILLER_69_561 ();
 sg13g2_decap_8 FILLER_69_568 ();
 sg13g2_fill_1 FILLER_69_602 ();
 sg13g2_decap_4 FILLER_69_648 ();
 sg13g2_fill_1 FILLER_69_652 ();
 sg13g2_fill_2 FILLER_69_690 ();
 sg13g2_fill_1 FILLER_69_697 ();
 sg13g2_fill_2 FILLER_69_735 ();
 sg13g2_fill_1 FILLER_69_737 ();
 sg13g2_decap_8 FILLER_69_766 ();
 sg13g2_decap_8 FILLER_69_773 ();
 sg13g2_fill_2 FILLER_69_780 ();
 sg13g2_fill_2 FILLER_69_809 ();
 sg13g2_fill_1 FILLER_69_811 ();
 sg13g2_fill_2 FILLER_69_821 ();
 sg13g2_fill_1 FILLER_69_823 ();
 sg13g2_decap_4 FILLER_69_850 ();
 sg13g2_fill_1 FILLER_69_854 ();
 sg13g2_decap_8 FILLER_69_868 ();
 sg13g2_fill_2 FILLER_69_894 ();
 sg13g2_fill_2 FILLER_69_961 ();
 sg13g2_fill_1 FILLER_69_963 ();
 sg13g2_decap_4 FILLER_69_986 ();
 sg13g2_decap_8 FILLER_69_999 ();
 sg13g2_decap_8 FILLER_69_1006 ();
 sg13g2_fill_1 FILLER_69_1013 ();
 sg13g2_fill_1 FILLER_69_1041 ();
 sg13g2_fill_2 FILLER_69_1056 ();
 sg13g2_fill_2 FILLER_69_1071 ();
 sg13g2_fill_1 FILLER_69_1073 ();
 sg13g2_decap_8 FILLER_69_1087 ();
 sg13g2_decap_8 FILLER_69_1094 ();
 sg13g2_decap_8 FILLER_69_1101 ();
 sg13g2_decap_8 FILLER_69_1108 ();
 sg13g2_decap_8 FILLER_69_1130 ();
 sg13g2_decap_8 FILLER_69_1137 ();
 sg13g2_decap_4 FILLER_69_1144 ();
 sg13g2_fill_2 FILLER_69_1148 ();
 sg13g2_decap_8 FILLER_69_1195 ();
 sg13g2_decap_8 FILLER_69_1202 ();
 sg13g2_decap_8 FILLER_69_1209 ();
 sg13g2_decap_4 FILLER_69_1216 ();
 sg13g2_fill_1 FILLER_69_1220 ();
 sg13g2_fill_1 FILLER_69_1240 ();
 sg13g2_fill_2 FILLER_69_1266 ();
 sg13g2_fill_1 FILLER_69_1268 ();
 sg13g2_fill_1 FILLER_69_1274 ();
 sg13g2_decap_8 FILLER_69_1339 ();
 sg13g2_decap_4 FILLER_69_1346 ();
 sg13g2_fill_2 FILLER_69_1350 ();
 sg13g2_decap_8 FILLER_69_1365 ();
 sg13g2_decap_8 FILLER_69_1372 ();
 sg13g2_fill_1 FILLER_69_1379 ();
 sg13g2_fill_1 FILLER_69_1407 ();
 sg13g2_decap_8 FILLER_69_1417 ();
 sg13g2_decap_4 FILLER_69_1424 ();
 sg13g2_decap_8 FILLER_69_1449 ();
 sg13g2_decap_8 FILLER_69_1469 ();
 sg13g2_decap_8 FILLER_69_1476 ();
 sg13g2_decap_8 FILLER_69_1483 ();
 sg13g2_decap_4 FILLER_69_1490 ();
 sg13g2_fill_1 FILLER_69_1494 ();
 sg13g2_fill_2 FILLER_69_1551 ();
 sg13g2_fill_1 FILLER_69_1553 ();
 sg13g2_fill_2 FILLER_69_1559 ();
 sg13g2_decap_8 FILLER_69_1574 ();
 sg13g2_fill_1 FILLER_69_1594 ();
 sg13g2_fill_2 FILLER_69_1600 ();
 sg13g2_fill_1 FILLER_69_1602 ();
 sg13g2_fill_1 FILLER_69_1612 ();
 sg13g2_fill_2 FILLER_69_1626 ();
 sg13g2_fill_1 FILLER_69_1628 ();
 sg13g2_decap_8 FILLER_69_1689 ();
 sg13g2_decap_4 FILLER_69_1696 ();
 sg13g2_fill_2 FILLER_69_1700 ();
 sg13g2_fill_2 FILLER_69_1716 ();
 sg13g2_fill_1 FILLER_69_1718 ();
 sg13g2_decap_8 FILLER_69_1745 ();
 sg13g2_decap_4 FILLER_69_1752 ();
 sg13g2_fill_1 FILLER_69_1756 ();
 sg13g2_fill_1 FILLER_69_1786 ();
 sg13g2_decap_8 FILLER_69_1792 ();
 sg13g2_decap_8 FILLER_69_1799 ();
 sg13g2_decap_8 FILLER_69_1806 ();
 sg13g2_decap_8 FILLER_69_1813 ();
 sg13g2_decap_4 FILLER_69_1820 ();
 sg13g2_fill_1 FILLER_69_1824 ();
 sg13g2_decap_4 FILLER_69_1830 ();
 sg13g2_decap_8 FILLER_69_1849 ();
 sg13g2_decap_8 FILLER_69_1856 ();
 sg13g2_decap_8 FILLER_69_1863 ();
 sg13g2_decap_8 FILLER_69_1870 ();
 sg13g2_fill_1 FILLER_69_1887 ();
 sg13g2_decap_4 FILLER_69_1898 ();
 sg13g2_fill_2 FILLER_69_1902 ();
 sg13g2_decap_4 FILLER_69_1909 ();
 sg13g2_fill_2 FILLER_69_1930 ();
 sg13g2_fill_1 FILLER_69_1947 ();
 sg13g2_fill_2 FILLER_69_1953 ();
 sg13g2_fill_2 FILLER_69_1964 ();
 sg13g2_decap_4 FILLER_69_1974 ();
 sg13g2_fill_1 FILLER_69_1978 ();
 sg13g2_fill_2 FILLER_69_1984 ();
 sg13g2_fill_1 FILLER_69_1998 ();
 sg13g2_fill_1 FILLER_69_2018 ();
 sg13g2_fill_2 FILLER_69_2045 ();
 sg13g2_decap_8 FILLER_69_2055 ();
 sg13g2_decap_8 FILLER_69_2062 ();
 sg13g2_decap_8 FILLER_69_2069 ();
 sg13g2_fill_1 FILLER_69_2076 ();
 sg13g2_fill_1 FILLER_69_2082 ();
 sg13g2_fill_1 FILLER_69_2091 ();
 sg13g2_decap_8 FILLER_69_2102 ();
 sg13g2_decap_8 FILLER_69_2109 ();
 sg13g2_fill_2 FILLER_69_2116 ();
 sg13g2_fill_1 FILLER_69_2123 ();
 sg13g2_decap_8 FILLER_69_2128 ();
 sg13g2_decap_8 FILLER_69_2135 ();
 sg13g2_decap_4 FILLER_69_2142 ();
 sg13g2_fill_1 FILLER_69_2180 ();
 sg13g2_fill_1 FILLER_69_2196 ();
 sg13g2_fill_1 FILLER_69_2202 ();
 sg13g2_fill_2 FILLER_69_2216 ();
 sg13g2_decap_8 FILLER_69_2233 ();
 sg13g2_fill_2 FILLER_69_2240 ();
 sg13g2_decap_8 FILLER_69_2260 ();
 sg13g2_decap_8 FILLER_69_2267 ();
 sg13g2_decap_8 FILLER_69_2274 ();
 sg13g2_decap_8 FILLER_69_2281 ();
 sg13g2_decap_8 FILLER_69_2288 ();
 sg13g2_fill_2 FILLER_69_2305 ();
 sg13g2_decap_8 FILLER_69_2312 ();
 sg13g2_fill_1 FILLER_69_2319 ();
 sg13g2_fill_1 FILLER_69_2328 ();
 sg13g2_fill_2 FILLER_69_2333 ();
 sg13g2_fill_1 FILLER_69_2335 ();
 sg13g2_fill_2 FILLER_69_2390 ();
 sg13g2_fill_1 FILLER_69_2392 ();
 sg13g2_decap_8 FILLER_69_2423 ();
 sg13g2_decap_8 FILLER_69_2430 ();
 sg13g2_decap_8 FILLER_69_2437 ();
 sg13g2_decap_8 FILLER_69_2444 ();
 sg13g2_decap_4 FILLER_69_2451 ();
 sg13g2_fill_2 FILLER_69_2455 ();
 sg13g2_decap_8 FILLER_69_2466 ();
 sg13g2_decap_8 FILLER_69_2473 ();
 sg13g2_fill_2 FILLER_69_2480 ();
 sg13g2_fill_1 FILLER_69_2482 ();
 sg13g2_decap_8 FILLER_69_2492 ();
 sg13g2_decap_8 FILLER_69_2499 ();
 sg13g2_fill_1 FILLER_69_2506 ();
 sg13g2_decap_8 FILLER_69_2538 ();
 sg13g2_decap_8 FILLER_69_2545 ();
 sg13g2_fill_2 FILLER_69_2552 ();
 sg13g2_fill_1 FILLER_69_2554 ();
 sg13g2_decap_4 FILLER_69_2564 ();
 sg13g2_decap_8 FILLER_69_2581 ();
 sg13g2_decap_8 FILLER_69_2602 ();
 sg13g2_fill_1 FILLER_69_2609 ();
 sg13g2_decap_8 FILLER_69_2652 ();
 sg13g2_decap_8 FILLER_69_2659 ();
 sg13g2_decap_8 FILLER_69_2666 ();
 sg13g2_decap_8 FILLER_69_2673 ();
 sg13g2_decap_8 FILLER_69_2680 ();
 sg13g2_fill_2 FILLER_69_2687 ();
 sg13g2_decap_8 FILLER_69_2703 ();
 sg13g2_decap_8 FILLER_69_2737 ();
 sg13g2_fill_1 FILLER_69_2744 ();
 sg13g2_decap_8 FILLER_69_2795 ();
 sg13g2_fill_1 FILLER_69_2802 ();
 sg13g2_fill_2 FILLER_69_2851 ();
 sg13g2_fill_1 FILLER_69_2889 ();
 sg13g2_decap_8 FILLER_69_2907 ();
 sg13g2_decap_8 FILLER_69_2914 ();
 sg13g2_fill_1 FILLER_69_2921 ();
 sg13g2_fill_1 FILLER_69_3001 ();
 sg13g2_fill_2 FILLER_69_3015 ();
 sg13g2_fill_1 FILLER_69_3017 ();
 sg13g2_decap_4 FILLER_69_3056 ();
 sg13g2_fill_2 FILLER_69_3060 ();
 sg13g2_decap_8 FILLER_69_3071 ();
 sg13g2_decap_8 FILLER_69_3078 ();
 sg13g2_decap_4 FILLER_69_3085 ();
 sg13g2_fill_2 FILLER_69_3099 ();
 sg13g2_fill_1 FILLER_69_3101 ();
 sg13g2_decap_8 FILLER_69_3112 ();
 sg13g2_decap_8 FILLER_69_3119 ();
 sg13g2_decap_8 FILLER_69_3126 ();
 sg13g2_decap_4 FILLER_69_3133 ();
 sg13g2_decap_8 FILLER_69_3195 ();
 sg13g2_fill_1 FILLER_69_3202 ();
 sg13g2_fill_2 FILLER_69_3213 ();
 sg13g2_decap_8 FILLER_69_3233 ();
 sg13g2_decap_8 FILLER_69_3240 ();
 sg13g2_fill_2 FILLER_69_3302 ();
 sg13g2_decap_8 FILLER_69_3313 ();
 sg13g2_decap_8 FILLER_69_3320 ();
 sg13g2_fill_2 FILLER_69_3327 ();
 sg13g2_decap_8 FILLER_69_3338 ();
 sg13g2_decap_8 FILLER_69_3345 ();
 sg13g2_decap_8 FILLER_69_3352 ();
 sg13g2_decap_8 FILLER_69_3359 ();
 sg13g2_fill_2 FILLER_69_3366 ();
 sg13g2_decap_8 FILLER_69_3400 ();
 sg13g2_decap_8 FILLER_69_3407 ();
 sg13g2_decap_8 FILLER_69_3414 ();
 sg13g2_fill_1 FILLER_69_3465 ();
 sg13g2_decap_8 FILLER_69_3475 ();
 sg13g2_fill_2 FILLER_69_3482 ();
 sg13g2_decap_4 FILLER_69_3494 ();
 sg13g2_fill_2 FILLER_69_3498 ();
 sg13g2_decap_8 FILLER_69_3513 ();
 sg13g2_decap_8 FILLER_69_3520 ();
 sg13g2_decap_8 FILLER_69_3527 ();
 sg13g2_decap_4 FILLER_69_3534 ();
 sg13g2_fill_2 FILLER_69_3548 ();
 sg13g2_decap_8 FILLER_69_3567 ();
 sg13g2_decap_4 FILLER_69_3574 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_4 FILLER_70_14 ();
 sg13g2_decap_4 FILLER_70_65 ();
 sg13g2_decap_8 FILLER_70_113 ();
 sg13g2_decap_8 FILLER_70_120 ();
 sg13g2_decap_8 FILLER_70_127 ();
 sg13g2_fill_2 FILLER_70_134 ();
 sg13g2_decap_8 FILLER_70_146 ();
 sg13g2_decap_8 FILLER_70_158 ();
 sg13g2_decap_8 FILLER_70_165 ();
 sg13g2_decap_4 FILLER_70_172 ();
 sg13g2_fill_2 FILLER_70_176 ();
 sg13g2_fill_1 FILLER_70_198 ();
 sg13g2_decap_8 FILLER_70_236 ();
 sg13g2_fill_2 FILLER_70_243 ();
 sg13g2_fill_1 FILLER_70_245 ();
 sg13g2_decap_4 FILLER_70_255 ();
 sg13g2_fill_1 FILLER_70_259 ();
 sg13g2_fill_2 FILLER_70_305 ();
 sg13g2_fill_1 FILLER_70_307 ();
 sg13g2_fill_1 FILLER_70_318 ();
 sg13g2_fill_2 FILLER_70_375 ();
 sg13g2_fill_1 FILLER_70_377 ();
 sg13g2_fill_2 FILLER_70_430 ();
 sg13g2_fill_1 FILLER_70_459 ();
 sg13g2_decap_4 FILLER_70_480 ();
 sg13g2_decap_4 FILLER_70_521 ();
 sg13g2_fill_1 FILLER_70_525 ();
 sg13g2_fill_2 FILLER_70_558 ();
 sg13g2_fill_2 FILLER_70_617 ();
 sg13g2_decap_8 FILLER_70_642 ();
 sg13g2_decap_4 FILLER_70_649 ();
 sg13g2_fill_1 FILLER_70_653 ();
 sg13g2_fill_2 FILLER_70_677 ();
 sg13g2_decap_4 FILLER_70_689 ();
 sg13g2_decap_8 FILLER_70_736 ();
 sg13g2_decap_8 FILLER_70_743 ();
 sg13g2_decap_4 FILLER_70_750 ();
 sg13g2_fill_1 FILLER_70_754 ();
 sg13g2_decap_8 FILLER_70_783 ();
 sg13g2_decap_8 FILLER_70_790 ();
 sg13g2_fill_2 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_829 ();
 sg13g2_decap_8 FILLER_70_836 ();
 sg13g2_decap_8 FILLER_70_843 ();
 sg13g2_fill_2 FILLER_70_850 ();
 sg13g2_fill_2 FILLER_70_861 ();
 sg13g2_decap_8 FILLER_70_876 ();
 sg13g2_fill_2 FILLER_70_886 ();
 sg13g2_decap_4 FILLER_70_920 ();
 sg13g2_decap_8 FILLER_70_930 ();
 sg13g2_decap_8 FILLER_70_937 ();
 sg13g2_decap_8 FILLER_70_944 ();
 sg13g2_decap_8 FILLER_70_951 ();
 sg13g2_fill_1 FILLER_70_958 ();
 sg13g2_decap_8 FILLER_70_972 ();
 sg13g2_decap_8 FILLER_70_979 ();
 sg13g2_decap_8 FILLER_70_986 ();
 sg13g2_decap_8 FILLER_70_993 ();
 sg13g2_decap_4 FILLER_70_1000 ();
 sg13g2_decap_8 FILLER_70_1019 ();
 sg13g2_decap_8 FILLER_70_1026 ();
 sg13g2_fill_1 FILLER_70_1033 ();
 sg13g2_decap_4 FILLER_70_1098 ();
 sg13g2_fill_2 FILLER_70_1102 ();
 sg13g2_decap_8 FILLER_70_1110 ();
 sg13g2_decap_4 FILLER_70_1121 ();
 sg13g2_fill_2 FILLER_70_1125 ();
 sg13g2_decap_4 FILLER_70_1136 ();
 sg13g2_fill_2 FILLER_70_1140 ();
 sg13g2_fill_2 FILLER_70_1152 ();
 sg13g2_fill_1 FILLER_70_1154 ();
 sg13g2_fill_1 FILLER_70_1164 ();
 sg13g2_fill_2 FILLER_70_1181 ();
 sg13g2_fill_2 FILLER_70_1192 ();
 sg13g2_decap_4 FILLER_70_1203 ();
 sg13g2_decap_4 FILLER_70_1262 ();
 sg13g2_decap_8 FILLER_70_1273 ();
 sg13g2_fill_2 FILLER_70_1294 ();
 sg13g2_fill_1 FILLER_70_1318 ();
 sg13g2_fill_1 FILLER_70_1334 ();
 sg13g2_decap_8 FILLER_70_1340 ();
 sg13g2_decap_8 FILLER_70_1347 ();
 sg13g2_decap_4 FILLER_70_1354 ();
 sg13g2_fill_1 FILLER_70_1358 ();
 sg13g2_fill_1 FILLER_70_1390 ();
 sg13g2_decap_8 FILLER_70_1415 ();
 sg13g2_decap_8 FILLER_70_1422 ();
 sg13g2_fill_1 FILLER_70_1429 ();
 sg13g2_fill_2 FILLER_70_1443 ();
 sg13g2_fill_1 FILLER_70_1445 ();
 sg13g2_fill_2 FILLER_70_1451 ();
 sg13g2_fill_1 FILLER_70_1453 ();
 sg13g2_fill_1 FILLER_70_1471 ();
 sg13g2_fill_2 FILLER_70_1485 ();
 sg13g2_fill_2 FILLER_70_1497 ();
 sg13g2_decap_8 FILLER_70_1531 ();
 sg13g2_fill_2 FILLER_70_1538 ();
 sg13g2_fill_1 FILLER_70_1540 ();
 sg13g2_fill_2 FILLER_70_1564 ();
 sg13g2_decap_4 FILLER_70_1579 ();
 sg13g2_fill_2 FILLER_70_1583 ();
 sg13g2_decap_4 FILLER_70_1639 ();
 sg13g2_fill_1 FILLER_70_1643 ();
 sg13g2_fill_2 FILLER_70_1654 ();
 sg13g2_fill_1 FILLER_70_1665 ();
 sg13g2_fill_1 FILLER_70_1679 ();
 sg13g2_decap_8 FILLER_70_1685 ();
 sg13g2_decap_4 FILLER_70_1692 ();
 sg13g2_fill_2 FILLER_70_1724 ();
 sg13g2_fill_1 FILLER_70_1726 ();
 sg13g2_decap_8 FILLER_70_1749 ();
 sg13g2_decap_4 FILLER_70_1756 ();
 sg13g2_fill_1 FILLER_70_1760 ();
 sg13g2_decap_8 FILLER_70_1788 ();
 sg13g2_decap_4 FILLER_70_1795 ();
 sg13g2_fill_2 FILLER_70_1799 ();
 sg13g2_decap_8 FILLER_70_1818 ();
 sg13g2_decap_4 FILLER_70_1825 ();
 sg13g2_fill_1 FILLER_70_1829 ();
 sg13g2_decap_8 FILLER_70_1846 ();
 sg13g2_decap_8 FILLER_70_1853 ();
 sg13g2_decap_4 FILLER_70_1860 ();
 sg13g2_fill_2 FILLER_70_1903 ();
 sg13g2_fill_1 FILLER_70_1905 ();
 sg13g2_fill_2 FILLER_70_1926 ();
 sg13g2_fill_1 FILLER_70_1928 ();
 sg13g2_fill_2 FILLER_70_1944 ();
 sg13g2_decap_8 FILLER_70_1981 ();
 sg13g2_fill_1 FILLER_70_2018 ();
 sg13g2_fill_2 FILLER_70_2032 ();
 sg13g2_fill_1 FILLER_70_2034 ();
 sg13g2_decap_4 FILLER_70_2041 ();
 sg13g2_decap_4 FILLER_70_2076 ();
 sg13g2_decap_8 FILLER_70_2095 ();
 sg13g2_decap_4 FILLER_70_2102 ();
 sg13g2_fill_1 FILLER_70_2106 ();
 sg13g2_fill_2 FILLER_70_2139 ();
 sg13g2_fill_1 FILLER_70_2141 ();
 sg13g2_fill_1 FILLER_70_2156 ();
 sg13g2_decap_8 FILLER_70_2167 ();
 sg13g2_decap_4 FILLER_70_2174 ();
 sg13g2_fill_2 FILLER_70_2193 ();
 sg13g2_decap_8 FILLER_70_2200 ();
 sg13g2_fill_2 FILLER_70_2207 ();
 sg13g2_fill_1 FILLER_70_2209 ();
 sg13g2_decap_8 FILLER_70_2228 ();
 sg13g2_decap_8 FILLER_70_2235 ();
 sg13g2_fill_1 FILLER_70_2242 ();
 sg13g2_decap_8 FILLER_70_2256 ();
 sg13g2_fill_2 FILLER_70_2263 ();
 sg13g2_decap_8 FILLER_70_2275 ();
 sg13g2_fill_2 FILLER_70_2282 ();
 sg13g2_fill_1 FILLER_70_2284 ();
 sg13g2_fill_2 FILLER_70_2295 ();
 sg13g2_fill_1 FILLER_70_2297 ();
 sg13g2_decap_8 FILLER_70_2334 ();
 sg13g2_fill_2 FILLER_70_2341 ();
 sg13g2_fill_1 FILLER_70_2343 ();
 sg13g2_fill_1 FILLER_70_2370 ();
 sg13g2_fill_1 FILLER_70_2375 ();
 sg13g2_fill_1 FILLER_70_2397 ();
 sg13g2_fill_2 FILLER_70_2413 ();
 sg13g2_decap_8 FILLER_70_2443 ();
 sg13g2_decap_4 FILLER_70_2450 ();
 sg13g2_decap_4 FILLER_70_2502 ();
 sg13g2_decap_8 FILLER_70_2528 ();
 sg13g2_decap_8 FILLER_70_2535 ();
 sg13g2_fill_2 FILLER_70_2542 ();
 sg13g2_fill_1 FILLER_70_2544 ();
 sg13g2_decap_8 FILLER_70_2568 ();
 sg13g2_decap_8 FILLER_70_2575 ();
 sg13g2_fill_1 FILLER_70_2582 ();
 sg13g2_fill_2 FILLER_70_2631 ();
 sg13g2_fill_1 FILLER_70_2633 ();
 sg13g2_decap_8 FILLER_70_2638 ();
 sg13g2_decap_4 FILLER_70_2645 ();
 sg13g2_fill_2 FILLER_70_2649 ();
 sg13g2_decap_4 FILLER_70_2672 ();
 sg13g2_fill_1 FILLER_70_2676 ();
 sg13g2_decap_8 FILLER_70_2687 ();
 sg13g2_fill_2 FILLER_70_2694 ();
 sg13g2_fill_1 FILLER_70_2696 ();
 sg13g2_decap_4 FILLER_70_2719 ();
 sg13g2_fill_2 FILLER_70_2723 ();
 sg13g2_decap_8 FILLER_70_2738 ();
 sg13g2_decap_4 FILLER_70_2745 ();
 sg13g2_fill_1 FILLER_70_2749 ();
 sg13g2_decap_8 FILLER_70_2790 ();
 sg13g2_fill_2 FILLER_70_2797 ();
 sg13g2_decap_4 FILLER_70_2845 ();
 sg13g2_fill_2 FILLER_70_2849 ();
 sg13g2_decap_8 FILLER_70_2900 ();
 sg13g2_decap_8 FILLER_70_2907 ();
 sg13g2_decap_8 FILLER_70_2914 ();
 sg13g2_fill_1 FILLER_70_2921 ();
 sg13g2_fill_2 FILLER_70_2945 ();
 sg13g2_decap_8 FILLER_70_2978 ();
 sg13g2_decap_8 FILLER_70_2985 ();
 sg13g2_decap_8 FILLER_70_2992 ();
 sg13g2_decap_4 FILLER_70_2999 ();
 sg13g2_fill_2 FILLER_70_3003 ();
 sg13g2_fill_2 FILLER_70_3032 ();
 sg13g2_decap_8 FILLER_70_3053 ();
 sg13g2_decap_8 FILLER_70_3060 ();
 sg13g2_decap_8 FILLER_70_3067 ();
 sg13g2_decap_4 FILLER_70_3074 ();
 sg13g2_fill_1 FILLER_70_3078 ();
 sg13g2_decap_8 FILLER_70_3125 ();
 sg13g2_decap_8 FILLER_70_3132 ();
 sg13g2_decap_4 FILLER_70_3139 ();
 sg13g2_fill_2 FILLER_70_3143 ();
 sg13g2_decap_8 FILLER_70_3190 ();
 sg13g2_decap_8 FILLER_70_3197 ();
 sg13g2_decap_8 FILLER_70_3204 ();
 sg13g2_fill_2 FILLER_70_3211 ();
 sg13g2_decap_8 FILLER_70_3221 ();
 sg13g2_decap_4 FILLER_70_3228 ();
 sg13g2_fill_2 FILLER_70_3232 ();
 sg13g2_fill_2 FILLER_70_3247 ();
 sg13g2_decap_4 FILLER_70_3290 ();
 sg13g2_fill_2 FILLER_70_3294 ();
 sg13g2_fill_2 FILLER_70_3333 ();
 sg13g2_fill_1 FILLER_70_3335 ();
 sg13g2_decap_4 FILLER_70_3349 ();
 sg13g2_fill_1 FILLER_70_3353 ();
 sg13g2_decap_8 FILLER_70_3407 ();
 sg13g2_decap_8 FILLER_70_3414 ();
 sg13g2_decap_8 FILLER_70_3466 ();
 sg13g2_decap_8 FILLER_70_3473 ();
 sg13g2_fill_2 FILLER_70_3480 ();
 sg13g2_fill_1 FILLER_70_3482 ();
 sg13g2_decap_4 FILLER_70_3510 ();
 sg13g2_decap_4 FILLER_70_3524 ();
 sg13g2_fill_2 FILLER_70_3528 ();
 sg13g2_decap_8 FILLER_70_3567 ();
 sg13g2_decap_4 FILLER_70_3574 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_37 ();
 sg13g2_decap_4 FILLER_71_56 ();
 sg13g2_fill_2 FILLER_71_65 ();
 sg13g2_fill_1 FILLER_71_67 ();
 sg13g2_fill_1 FILLER_71_73 ();
 sg13g2_decap_4 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_93 ();
 sg13g2_decap_8 FILLER_71_100 ();
 sg13g2_decap_8 FILLER_71_107 ();
 sg13g2_decap_8 FILLER_71_114 ();
 sg13g2_decap_8 FILLER_71_121 ();
 sg13g2_decap_4 FILLER_71_175 ();
 sg13g2_fill_1 FILLER_71_179 ();
 sg13g2_fill_2 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_246 ();
 sg13g2_decap_4 FILLER_71_253 ();
 sg13g2_fill_1 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_285 ();
 sg13g2_fill_2 FILLER_71_310 ();
 sg13g2_fill_1 FILLER_71_312 ();
 sg13g2_fill_2 FILLER_71_323 ();
 sg13g2_decap_4 FILLER_71_384 ();
 sg13g2_fill_1 FILLER_71_428 ();
 sg13g2_fill_1 FILLER_71_443 ();
 sg13g2_fill_2 FILLER_71_458 ();
 sg13g2_decap_4 FILLER_71_476 ();
 sg13g2_fill_1 FILLER_71_480 ();
 sg13g2_fill_1 FILLER_71_559 ();
 sg13g2_fill_1 FILLER_71_586 ();
 sg13g2_decap_8 FILLER_71_641 ();
 sg13g2_decap_8 FILLER_71_648 ();
 sg13g2_decap_4 FILLER_71_655 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_decap_4 FILLER_71_691 ();
 sg13g2_decap_4 FILLER_71_714 ();
 sg13g2_decap_4 FILLER_71_727 ();
 sg13g2_decap_8 FILLER_71_773 ();
 sg13g2_decap_8 FILLER_71_780 ();
 sg13g2_fill_2 FILLER_71_787 ();
 sg13g2_fill_1 FILLER_71_789 ();
 sg13g2_fill_1 FILLER_71_820 ();
 sg13g2_fill_2 FILLER_71_830 ();
 sg13g2_decap_4 FILLER_71_836 ();
 sg13g2_fill_2 FILLER_71_840 ();
 sg13g2_decap_4 FILLER_71_880 ();
 sg13g2_fill_1 FILLER_71_884 ();
 sg13g2_decap_8 FILLER_71_894 ();
 sg13g2_decap_4 FILLER_71_920 ();
 sg13g2_fill_2 FILLER_71_924 ();
 sg13g2_decap_8 FILLER_71_967 ();
 sg13g2_decap_8 FILLER_71_974 ();
 sg13g2_fill_1 FILLER_71_981 ();
 sg13g2_decap_8 FILLER_71_1028 ();
 sg13g2_decap_4 FILLER_71_1035 ();
 sg13g2_fill_1 FILLER_71_1039 ();
 sg13g2_decap_8 FILLER_71_1050 ();
 sg13g2_decap_8 FILLER_71_1057 ();
 sg13g2_decap_4 FILLER_71_1064 ();
 sg13g2_fill_1 FILLER_71_1068 ();
 sg13g2_fill_2 FILLER_71_1091 ();
 sg13g2_fill_1 FILLER_71_1106 ();
 sg13g2_fill_1 FILLER_71_1116 ();
 sg13g2_fill_2 FILLER_71_1131 ();
 sg13g2_fill_2 FILLER_71_1139 ();
 sg13g2_fill_1 FILLER_71_1141 ();
 sg13g2_decap_8 FILLER_71_1153 ();
 sg13g2_decap_8 FILLER_71_1160 ();
 sg13g2_decap_8 FILLER_71_1167 ();
 sg13g2_fill_2 FILLER_71_1174 ();
 sg13g2_fill_1 FILLER_71_1176 ();
 sg13g2_fill_2 FILLER_71_1207 ();
 sg13g2_fill_1 FILLER_71_1222 ();
 sg13g2_fill_1 FILLER_71_1266 ();
 sg13g2_fill_2 FILLER_71_1281 ();
 sg13g2_fill_1 FILLER_71_1283 ();
 sg13g2_decap_4 FILLER_71_1320 ();
 sg13g2_fill_2 FILLER_71_1324 ();
 sg13g2_decap_8 FILLER_71_1329 ();
 sg13g2_decap_8 FILLER_71_1336 ();
 sg13g2_fill_1 FILLER_71_1390 ();
 sg13g2_decap_8 FILLER_71_1397 ();
 sg13g2_decap_4 FILLER_71_1404 ();
 sg13g2_fill_1 FILLER_71_1408 ();
 sg13g2_decap_4 FILLER_71_1414 ();
 sg13g2_decap_8 FILLER_71_1486 ();
 sg13g2_fill_1 FILLER_71_1493 ();
 sg13g2_decap_8 FILLER_71_1522 ();
 sg13g2_decap_4 FILLER_71_1529 ();
 sg13g2_fill_2 FILLER_71_1533 ();
 sg13g2_decap_8 FILLER_71_1589 ();
 sg13g2_fill_1 FILLER_71_1596 ();
 sg13g2_fill_1 FILLER_71_1647 ();
 sg13g2_decap_8 FILLER_71_1657 ();
 sg13g2_fill_2 FILLER_71_1664 ();
 sg13g2_fill_2 FILLER_71_1688 ();
 sg13g2_fill_1 FILLER_71_1690 ();
 sg13g2_fill_2 FILLER_71_1719 ();
 sg13g2_fill_2 FILLER_71_1734 ();
 sg13g2_fill_1 FILLER_71_1736 ();
 sg13g2_decap_8 FILLER_71_1741 ();
 sg13g2_decap_8 FILLER_71_1748 ();
 sg13g2_decap_8 FILLER_71_1755 ();
 sg13g2_decap_8 FILLER_71_1798 ();
 sg13g2_fill_2 FILLER_71_1805 ();
 sg13g2_fill_2 FILLER_71_1813 ();
 sg13g2_fill_1 FILLER_71_1815 ();
 sg13g2_fill_2 FILLER_71_1821 ();
 sg13g2_fill_1 FILLER_71_1823 ();
 sg13g2_decap_8 FILLER_71_1857 ();
 sg13g2_fill_1 FILLER_71_1864 ();
 sg13g2_fill_2 FILLER_71_1870 ();
 sg13g2_decap_8 FILLER_71_1907 ();
 sg13g2_fill_2 FILLER_71_1914 ();
 sg13g2_fill_1 FILLER_71_1920 ();
 sg13g2_fill_1 FILLER_71_1931 ();
 sg13g2_decap_8 FILLER_71_1943 ();
 sg13g2_fill_2 FILLER_71_1950 ();
 sg13g2_fill_1 FILLER_71_1952 ();
 sg13g2_decap_4 FILLER_71_1967 ();
 sg13g2_fill_2 FILLER_71_1971 ();
 sg13g2_decap_8 FILLER_71_1986 ();
 sg13g2_decap_4 FILLER_71_1993 ();
 sg13g2_fill_1 FILLER_71_1997 ();
 sg13g2_fill_1 FILLER_71_2008 ();
 sg13g2_decap_8 FILLER_71_2015 ();
 sg13g2_decap_4 FILLER_71_2022 ();
 sg13g2_fill_2 FILLER_71_2026 ();
 sg13g2_fill_1 FILLER_71_2034 ();
 sg13g2_fill_1 FILLER_71_2045 ();
 sg13g2_decap_8 FILLER_71_2064 ();
 sg13g2_decap_8 FILLER_71_2071 ();
 sg13g2_decap_8 FILLER_71_2105 ();
 sg13g2_decap_4 FILLER_71_2112 ();
 sg13g2_fill_1 FILLER_71_2116 ();
 sg13g2_fill_2 FILLER_71_2127 ();
 sg13g2_fill_1 FILLER_71_2139 ();
 sg13g2_decap_8 FILLER_71_2144 ();
 sg13g2_decap_8 FILLER_71_2151 ();
 sg13g2_decap_8 FILLER_71_2158 ();
 sg13g2_decap_4 FILLER_71_2165 ();
 sg13g2_fill_1 FILLER_71_2169 ();
 sg13g2_decap_8 FILLER_71_2174 ();
 sg13g2_decap_4 FILLER_71_2181 ();
 sg13g2_fill_2 FILLER_71_2185 ();
 sg13g2_decap_4 FILLER_71_2191 ();
 sg13g2_fill_2 FILLER_71_2195 ();
 sg13g2_decap_4 FILLER_71_2208 ();
 sg13g2_decap_8 FILLER_71_2222 ();
 sg13g2_decap_8 FILLER_71_2229 ();
 sg13g2_decap_8 FILLER_71_2236 ();
 sg13g2_decap_8 FILLER_71_2243 ();
 sg13g2_fill_1 FILLER_71_2263 ();
 sg13g2_decap_4 FILLER_71_2269 ();
 sg13g2_fill_2 FILLER_71_2273 ();
 sg13g2_fill_2 FILLER_71_2298 ();
 sg13g2_decap_8 FILLER_71_2331 ();
 sg13g2_fill_2 FILLER_71_2346 ();
 sg13g2_fill_1 FILLER_71_2348 ();
 sg13g2_decap_8 FILLER_71_2362 ();
 sg13g2_decap_8 FILLER_71_2369 ();
 sg13g2_decap_8 FILLER_71_2376 ();
 sg13g2_decap_8 FILLER_71_2428 ();
 sg13g2_decap_8 FILLER_71_2435 ();
 sg13g2_decap_8 FILLER_71_2442 ();
 sg13g2_decap_4 FILLER_71_2449 ();
 sg13g2_fill_1 FILLER_71_2453 ();
 sg13g2_fill_1 FILLER_71_2495 ();
 sg13g2_decap_8 FILLER_71_2523 ();
 sg13g2_decap_8 FILLER_71_2530 ();
 sg13g2_decap_4 FILLER_71_2537 ();
 sg13g2_decap_8 FILLER_71_2578 ();
 sg13g2_decap_4 FILLER_71_2585 ();
 sg13g2_fill_2 FILLER_71_2589 ();
 sg13g2_decap_8 FILLER_71_2636 ();
 sg13g2_decap_8 FILLER_71_2643 ();
 sg13g2_decap_8 FILLER_71_2650 ();
 sg13g2_decap_4 FILLER_71_2657 ();
 sg13g2_fill_1 FILLER_71_2661 ();
 sg13g2_fill_2 FILLER_71_2694 ();
 sg13g2_decap_8 FILLER_71_2717 ();
 sg13g2_decap_8 FILLER_71_2724 ();
 sg13g2_decap_8 FILLER_71_2731 ();
 sg13g2_decap_8 FILLER_71_2738 ();
 sg13g2_decap_8 FILLER_71_2745 ();
 sg13g2_fill_1 FILLER_71_2752 ();
 sg13g2_fill_1 FILLER_71_2766 ();
 sg13g2_decap_8 FILLER_71_2780 ();
 sg13g2_decap_4 FILLER_71_2787 ();
 sg13g2_fill_1 FILLER_71_2791 ();
 sg13g2_decap_8 FILLER_71_2829 ();
 sg13g2_decap_8 FILLER_71_2836 ();
 sg13g2_decap_8 FILLER_71_2843 ();
 sg13g2_decap_8 FILLER_71_2850 ();
 sg13g2_decap_8 FILLER_71_2857 ();
 sg13g2_decap_4 FILLER_71_2864 ();
 sg13g2_fill_1 FILLER_71_2868 ();
 sg13g2_decap_8 FILLER_71_2912 ();
 sg13g2_decap_8 FILLER_71_2919 ();
 sg13g2_fill_1 FILLER_71_2926 ();
 sg13g2_decap_8 FILLER_71_2982 ();
 sg13g2_decap_8 FILLER_71_2989 ();
 sg13g2_decap_4 FILLER_71_2996 ();
 sg13g2_fill_1 FILLER_71_3000 ();
 sg13g2_fill_2 FILLER_71_3028 ();
 sg13g2_fill_2 FILLER_71_3040 ();
 sg13g2_fill_1 FILLER_71_3042 ();
 sg13g2_decap_8 FILLER_71_3056 ();
 sg13g2_decap_8 FILLER_71_3063 ();
 sg13g2_fill_2 FILLER_71_3070 ();
 sg13g2_fill_1 FILLER_71_3072 ();
 sg13g2_decap_8 FILLER_71_3130 ();
 sg13g2_decap_8 FILLER_71_3137 ();
 sg13g2_decap_4 FILLER_71_3144 ();
 sg13g2_fill_1 FILLER_71_3148 ();
 sg13g2_decap_8 FILLER_71_3186 ();
 sg13g2_fill_2 FILLER_71_3193 ();
 sg13g2_fill_1 FILLER_71_3195 ();
 sg13g2_decap_4 FILLER_71_3206 ();
 sg13g2_fill_2 FILLER_71_3214 ();
 sg13g2_decap_8 FILLER_71_3225 ();
 sg13g2_decap_4 FILLER_71_3232 ();
 sg13g2_decap_4 FILLER_71_3249 ();
 sg13g2_fill_1 FILLER_71_3253 ();
 sg13g2_fill_1 FILLER_71_3268 ();
 sg13g2_fill_2 FILLER_71_3296 ();
 sg13g2_decap_8 FILLER_71_3399 ();
 sg13g2_decap_8 FILLER_71_3406 ();
 sg13g2_decap_8 FILLER_71_3413 ();
 sg13g2_decap_4 FILLER_71_3420 ();
 sg13g2_fill_2 FILLER_71_3434 ();
 sg13g2_fill_1 FILLER_71_3455 ();
 sg13g2_decap_8 FILLER_71_3469 ();
 sg13g2_fill_1 FILLER_71_3476 ();
 sg13g2_decap_8 FILLER_71_3571 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_53 ();
 sg13g2_decap_4 FILLER_72_63 ();
 sg13g2_decap_4 FILLER_72_80 ();
 sg13g2_fill_1 FILLER_72_116 ();
 sg13g2_fill_2 FILLER_72_154 ();
 sg13g2_fill_1 FILLER_72_156 ();
 sg13g2_fill_2 FILLER_72_170 ();
 sg13g2_fill_2 FILLER_72_217 ();
 sg13g2_fill_1 FILLER_72_219 ();
 sg13g2_decap_8 FILLER_72_229 ();
 sg13g2_decap_8 FILLER_72_236 ();
 sg13g2_decap_8 FILLER_72_243 ();
 sg13g2_fill_1 FILLER_72_296 ();
 sg13g2_fill_2 FILLER_72_333 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_fill_2 FILLER_72_367 ();
 sg13g2_fill_1 FILLER_72_369 ();
 sg13g2_decap_8 FILLER_72_375 ();
 sg13g2_fill_2 FILLER_72_382 ();
 sg13g2_fill_1 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_431 ();
 sg13g2_fill_1 FILLER_72_438 ();
 sg13g2_decap_8 FILLER_72_453 ();
 sg13g2_fill_1 FILLER_72_460 ();
 sg13g2_fill_2 FILLER_72_521 ();
 sg13g2_fill_1 FILLER_72_523 ();
 sg13g2_fill_1 FILLER_72_533 ();
 sg13g2_fill_2 FILLER_72_543 ();
 sg13g2_fill_1 FILLER_72_555 ();
 sg13g2_decap_8 FILLER_72_560 ();
 sg13g2_decap_8 FILLER_72_567 ();
 sg13g2_decap_4 FILLER_72_574 ();
 sg13g2_fill_1 FILLER_72_578 ();
 sg13g2_fill_2 FILLER_72_584 ();
 sg13g2_fill_1 FILLER_72_586 ();
 sg13g2_fill_1 FILLER_72_600 ();
 sg13g2_decap_4 FILLER_72_656 ();
 sg13g2_fill_2 FILLER_72_691 ();
 sg13g2_fill_1 FILLER_72_693 ();
 sg13g2_fill_2 FILLER_72_713 ();
 sg13g2_decap_4 FILLER_72_728 ();
 sg13g2_decap_8 FILLER_72_785 ();
 sg13g2_decap_8 FILLER_72_792 ();
 sg13g2_decap_4 FILLER_72_799 ();
 sg13g2_fill_1 FILLER_72_803 ();
 sg13g2_fill_2 FILLER_72_844 ();
 sg13g2_fill_1 FILLER_72_846 ();
 sg13g2_decap_4 FILLER_72_894 ();
 sg13g2_decap_4 FILLER_72_907 ();
 sg13g2_fill_2 FILLER_72_911 ();
 sg13g2_fill_2 FILLER_72_917 ();
 sg13g2_fill_1 FILLER_72_919 ();
 sg13g2_fill_1 FILLER_72_965 ();
 sg13g2_decap_4 FILLER_72_970 ();
 sg13g2_fill_2 FILLER_72_974 ();
 sg13g2_fill_2 FILLER_72_995 ();
 sg13g2_fill_1 FILLER_72_997 ();
 sg13g2_fill_2 FILLER_72_1017 ();
 sg13g2_fill_1 FILLER_72_1019 ();
 sg13g2_decap_8 FILLER_72_1033 ();
 sg13g2_decap_8 FILLER_72_1040 ();
 sg13g2_decap_4 FILLER_72_1047 ();
 sg13g2_fill_2 FILLER_72_1051 ();
 sg13g2_decap_4 FILLER_72_1060 ();
 sg13g2_fill_2 FILLER_72_1104 ();
 sg13g2_fill_2 FILLER_72_1117 ();
 sg13g2_fill_1 FILLER_72_1119 ();
 sg13g2_decap_8 FILLER_72_1157 ();
 sg13g2_decap_8 FILLER_72_1164 ();
 sg13g2_decap_4 FILLER_72_1171 ();
 sg13g2_fill_1 FILLER_72_1198 ();
 sg13g2_fill_2 FILLER_72_1208 ();
 sg13g2_fill_1 FILLER_72_1210 ();
 sg13g2_fill_2 FILLER_72_1232 ();
 sg13g2_fill_1 FILLER_72_1339 ();
 sg13g2_fill_2 FILLER_72_1345 ();
 sg13g2_decap_8 FILLER_72_1351 ();
 sg13g2_decap_8 FILLER_72_1358 ();
 sg13g2_decap_8 FILLER_72_1365 ();
 sg13g2_fill_2 FILLER_72_1372 ();
 sg13g2_fill_2 FILLER_72_1401 ();
 sg13g2_fill_1 FILLER_72_1403 ();
 sg13g2_decap_8 FILLER_72_1409 ();
 sg13g2_decap_8 FILLER_72_1416 ();
 sg13g2_decap_8 FILLER_72_1423 ();
 sg13g2_fill_1 FILLER_72_1443 ();
 sg13g2_fill_2 FILLER_72_1448 ();
 sg13g2_decap_4 FILLER_72_1469 ();
 sg13g2_fill_1 FILLER_72_1473 ();
 sg13g2_decap_8 FILLER_72_1492 ();
 sg13g2_fill_1 FILLER_72_1499 ();
 sg13g2_fill_1 FILLER_72_1505 ();
 sg13g2_decap_4 FILLER_72_1525 ();
 sg13g2_fill_2 FILLER_72_1529 ();
 sg13g2_fill_2 FILLER_72_1597 ();
 sg13g2_fill_2 FILLER_72_1614 ();
 sg13g2_fill_1 FILLER_72_1616 ();
 sg13g2_fill_1 FILLER_72_1623 ();
 sg13g2_fill_2 FILLER_72_1641 ();
 sg13g2_fill_1 FILLER_72_1643 ();
 sg13g2_decap_4 FILLER_72_1677 ();
 sg13g2_fill_2 FILLER_72_1681 ();
 sg13g2_fill_1 FILLER_72_1702 ();
 sg13g2_decap_8 FILLER_72_1753 ();
 sg13g2_decap_8 FILLER_72_1760 ();
 sg13g2_fill_2 FILLER_72_1767 ();
 sg13g2_fill_1 FILLER_72_1789 ();
 sg13g2_fill_1 FILLER_72_1802 ();
 sg13g2_decap_4 FILLER_72_1825 ();
 sg13g2_fill_2 FILLER_72_1834 ();
 sg13g2_fill_2 FILLER_72_1851 ();
 sg13g2_fill_1 FILLER_72_1853 ();
 sg13g2_decap_8 FILLER_72_1865 ();
 sg13g2_decap_4 FILLER_72_1872 ();
 sg13g2_fill_2 FILLER_72_1876 ();
 sg13g2_decap_8 FILLER_72_1905 ();
 sg13g2_decap_4 FILLER_72_1912 ();
 sg13g2_fill_2 FILLER_72_1916 ();
 sg13g2_fill_1 FILLER_72_1926 ();
 sg13g2_decap_8 FILLER_72_1937 ();
 sg13g2_decap_8 FILLER_72_1944 ();
 sg13g2_decap_8 FILLER_72_1951 ();
 sg13g2_decap_8 FILLER_72_1958 ();
 sg13g2_decap_8 FILLER_72_1965 ();
 sg13g2_decap_4 FILLER_72_1972 ();
 sg13g2_fill_1 FILLER_72_1976 ();
 sg13g2_decap_8 FILLER_72_1982 ();
 sg13g2_decap_8 FILLER_72_1989 ();
 sg13g2_decap_8 FILLER_72_1996 ();
 sg13g2_decap_8 FILLER_72_2003 ();
 sg13g2_decap_8 FILLER_72_2010 ();
 sg13g2_decap_8 FILLER_72_2017 ();
 sg13g2_fill_2 FILLER_72_2024 ();
 sg13g2_decap_8 FILLER_72_2039 ();
 sg13g2_decap_8 FILLER_72_2051 ();
 sg13g2_fill_1 FILLER_72_2058 ();
 sg13g2_fill_1 FILLER_72_2067 ();
 sg13g2_fill_2 FILLER_72_2081 ();
 sg13g2_decap_8 FILLER_72_2104 ();
 sg13g2_decap_8 FILLER_72_2111 ();
 sg13g2_fill_2 FILLER_72_2118 ();
 sg13g2_fill_1 FILLER_72_2120 ();
 sg13g2_decap_4 FILLER_72_2125 ();
 sg13g2_decap_8 FILLER_72_2139 ();
 sg13g2_decap_8 FILLER_72_2146 ();
 sg13g2_decap_8 FILLER_72_2153 ();
 sg13g2_fill_2 FILLER_72_2160 ();
 sg13g2_fill_2 FILLER_72_2166 ();
 sg13g2_fill_2 FILLER_72_2206 ();
 sg13g2_fill_1 FILLER_72_2208 ();
 sg13g2_decap_8 FILLER_72_2214 ();
 sg13g2_decap_8 FILLER_72_2221 ();
 sg13g2_decap_8 FILLER_72_2233 ();
 sg13g2_decap_8 FILLER_72_2240 ();
 sg13g2_decap_8 FILLER_72_2247 ();
 sg13g2_decap_8 FILLER_72_2293 ();
 sg13g2_decap_8 FILLER_72_2300 ();
 sg13g2_fill_2 FILLER_72_2307 ();
 sg13g2_decap_8 FILLER_72_2327 ();
 sg13g2_decap_8 FILLER_72_2334 ();
 sg13g2_fill_2 FILLER_72_2346 ();
 sg13g2_decap_4 FILLER_72_2359 ();
 sg13g2_fill_2 FILLER_72_2363 ();
 sg13g2_fill_2 FILLER_72_2370 ();
 sg13g2_fill_1 FILLER_72_2372 ();
 sg13g2_decap_8 FILLER_72_2414 ();
 sg13g2_decap_8 FILLER_72_2421 ();
 sg13g2_decap_8 FILLER_72_2428 ();
 sg13g2_decap_8 FILLER_72_2435 ();
 sg13g2_decap_8 FILLER_72_2442 ();
 sg13g2_decap_4 FILLER_72_2449 ();
 sg13g2_fill_1 FILLER_72_2453 ();
 sg13g2_fill_2 FILLER_72_2499 ();
 sg13g2_fill_1 FILLER_72_2535 ();
 sg13g2_decap_8 FILLER_72_2584 ();
 sg13g2_fill_2 FILLER_72_2591 ();
 sg13g2_fill_1 FILLER_72_2593 ();
 sg13g2_decap_8 FILLER_72_2648 ();
 sg13g2_decap_4 FILLER_72_2655 ();
 sg13g2_fill_2 FILLER_72_2707 ();
 sg13g2_fill_1 FILLER_72_2709 ();
 sg13g2_decap_8 FILLER_72_2737 ();
 sg13g2_decap_8 FILLER_72_2744 ();
 sg13g2_decap_8 FILLER_72_2751 ();
 sg13g2_decap_4 FILLER_72_2758 ();
 sg13g2_decap_8 FILLER_72_2771 ();
 sg13g2_decap_8 FILLER_72_2778 ();
 sg13g2_decap_8 FILLER_72_2785 ();
 sg13g2_decap_4 FILLER_72_2792 ();
 sg13g2_fill_1 FILLER_72_2796 ();
 sg13g2_fill_2 FILLER_72_2801 ();
 sg13g2_fill_1 FILLER_72_2803 ();
 sg13g2_decap_8 FILLER_72_2808 ();
 sg13g2_decap_4 FILLER_72_2815 ();
 sg13g2_decap_8 FILLER_72_2838 ();
 sg13g2_decap_4 FILLER_72_2845 ();
 sg13g2_fill_2 FILLER_72_2849 ();
 sg13g2_fill_2 FILLER_72_2861 ();
 sg13g2_fill_1 FILLER_72_2863 ();
 sg13g2_decap_8 FILLER_72_2922 ();
 sg13g2_fill_2 FILLER_72_2929 ();
 sg13g2_decap_4 FILLER_72_3002 ();
 sg13g2_decap_8 FILLER_72_3010 ();
 sg13g2_decap_4 FILLER_72_3017 ();
 sg13g2_fill_1 FILLER_72_3021 ();
 sg13g2_decap_4 FILLER_72_3073 ();
 sg13g2_fill_1 FILLER_72_3077 ();
 sg13g2_fill_2 FILLER_72_3082 ();
 sg13g2_fill_1 FILLER_72_3084 ();
 sg13g2_fill_1 FILLER_72_3138 ();
 sg13g2_fill_2 FILLER_72_3149 ();
 sg13g2_fill_1 FILLER_72_3151 ();
 sg13g2_decap_4 FILLER_72_3177 ();
 sg13g2_fill_1 FILLER_72_3181 ();
 sg13g2_fill_2 FILLER_72_3202 ();
 sg13g2_fill_1 FILLER_72_3204 ();
 sg13g2_decap_8 FILLER_72_3232 ();
 sg13g2_decap_8 FILLER_72_3239 ();
 sg13g2_fill_2 FILLER_72_3246 ();
 sg13g2_fill_1 FILLER_72_3248 ();
 sg13g2_fill_2 FILLER_72_3286 ();
 sg13g2_fill_1 FILLER_72_3288 ();
 sg13g2_decap_4 FILLER_72_3328 ();
 sg13g2_fill_2 FILLER_72_3332 ();
 sg13g2_fill_2 FILLER_72_3348 ();
 sg13g2_fill_1 FILLER_72_3350 ();
 sg13g2_fill_2 FILLER_72_3370 ();
 sg13g2_fill_1 FILLER_72_3372 ();
 sg13g2_decap_8 FILLER_72_3400 ();
 sg13g2_decap_8 FILLER_72_3407 ();
 sg13g2_decap_4 FILLER_72_3414 ();
 sg13g2_fill_2 FILLER_72_3418 ();
 sg13g2_decap_8 FILLER_72_3460 ();
 sg13g2_decap_8 FILLER_72_3467 ();
 sg13g2_decap_4 FILLER_72_3474 ();
 sg13g2_decap_8 FILLER_72_3509 ();
 sg13g2_fill_2 FILLER_72_3516 ();
 sg13g2_fill_1 FILLER_72_3518 ();
 sg13g2_fill_2 FILLER_72_3542 ();
 sg13g2_fill_1 FILLER_72_3544 ();
 sg13g2_decap_4 FILLER_72_3572 ();
 sg13g2_fill_2 FILLER_72_3576 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_7 ();
 sg13g2_fill_2 FILLER_73_11 ();
 sg13g2_fill_1 FILLER_73_60 ();
 sg13g2_fill_2 FILLER_73_98 ();
 sg13g2_fill_1 FILLER_73_100 ();
 sg13g2_fill_1 FILLER_73_161 ();
 sg13g2_fill_2 FILLER_73_176 ();
 sg13g2_fill_1 FILLER_73_178 ();
 sg13g2_decap_8 FILLER_73_228 ();
 sg13g2_fill_2 FILLER_73_299 ();
 sg13g2_decap_8 FILLER_73_342 ();
 sg13g2_decap_8 FILLER_73_349 ();
 sg13g2_decap_8 FILLER_73_356 ();
 sg13g2_decap_4 FILLER_73_363 ();
 sg13g2_fill_2 FILLER_73_391 ();
 sg13g2_decap_8 FILLER_73_440 ();
 sg13g2_decap_4 FILLER_73_447 ();
 sg13g2_fill_1 FILLER_73_451 ();
 sg13g2_decap_8 FILLER_73_465 ();
 sg13g2_fill_2 FILLER_73_472 ();
 sg13g2_fill_2 FILLER_73_500 ();
 sg13g2_fill_1 FILLER_73_502 ();
 sg13g2_fill_2 FILLER_73_515 ();
 sg13g2_fill_1 FILLER_73_586 ();
 sg13g2_fill_1 FILLER_73_624 ();
 sg13g2_fill_2 FILLER_73_652 ();
 sg13g2_decap_4 FILLER_73_701 ();
 sg13g2_fill_1 FILLER_73_724 ();
 sg13g2_decap_4 FILLER_73_750 ();
 sg13g2_fill_1 FILLER_73_754 ();
 sg13g2_decap_8 FILLER_73_783 ();
 sg13g2_decap_8 FILLER_73_790 ();
 sg13g2_decap_8 FILLER_73_797 ();
 sg13g2_decap_4 FILLER_73_804 ();
 sg13g2_fill_1 FILLER_73_808 ();
 sg13g2_fill_1 FILLER_73_819 ();
 sg13g2_decap_8 FILLER_73_855 ();
 sg13g2_fill_1 FILLER_73_862 ();
 sg13g2_decap_4 FILLER_73_890 ();
 sg13g2_fill_1 FILLER_73_894 ();
 sg13g2_fill_1 FILLER_73_923 ();
 sg13g2_fill_2 FILLER_73_987 ();
 sg13g2_fill_1 FILLER_73_999 ();
 sg13g2_decap_8 FILLER_73_1035 ();
 sg13g2_decap_8 FILLER_73_1042 ();
 sg13g2_decap_8 FILLER_73_1049 ();
 sg13g2_decap_8 FILLER_73_1056 ();
 sg13g2_fill_2 FILLER_73_1063 ();
 sg13g2_fill_1 FILLER_73_1065 ();
 sg13g2_fill_2 FILLER_73_1107 ();
 sg13g2_decap_8 FILLER_73_1161 ();
 sg13g2_decap_8 FILLER_73_1168 ();
 sg13g2_decap_4 FILLER_73_1175 ();
 sg13g2_fill_1 FILLER_73_1189 ();
 sg13g2_decap_8 FILLER_73_1204 ();
 sg13g2_decap_8 FILLER_73_1211 ();
 sg13g2_fill_2 FILLER_73_1218 ();
 sg13g2_fill_1 FILLER_73_1220 ();
 sg13g2_decap_4 FILLER_73_1249 ();
 sg13g2_fill_2 FILLER_73_1258 ();
 sg13g2_fill_1 FILLER_73_1260 ();
 sg13g2_decap_8 FILLER_73_1275 ();
 sg13g2_decap_4 FILLER_73_1282 ();
 sg13g2_fill_2 FILLER_73_1295 ();
 sg13g2_fill_1 FILLER_73_1297 ();
 sg13g2_fill_2 FILLER_73_1302 ();
 sg13g2_fill_2 FILLER_73_1331 ();
 sg13g2_fill_2 FILLER_73_1350 ();
 sg13g2_fill_2 FILLER_73_1370 ();
 sg13g2_fill_2 FILLER_73_1390 ();
 sg13g2_fill_1 FILLER_73_1392 ();
 sg13g2_decap_8 FILLER_73_1412 ();
 sg13g2_decap_8 FILLER_73_1419 ();
 sg13g2_decap_8 FILLER_73_1426 ();
 sg13g2_decap_4 FILLER_73_1438 ();
 sg13g2_fill_2 FILLER_73_1442 ();
 sg13g2_fill_2 FILLER_73_1452 ();
 sg13g2_decap_4 FILLER_73_1468 ();
 sg13g2_decap_8 FILLER_73_1498 ();
 sg13g2_decap_8 FILLER_73_1505 ();
 sg13g2_decap_8 FILLER_73_1512 ();
 sg13g2_decap_8 FILLER_73_1519 ();
 sg13g2_decap_8 FILLER_73_1526 ();
 sg13g2_fill_2 FILLER_73_1533 ();
 sg13g2_fill_1 FILLER_73_1535 ();
 sg13g2_decap_8 FILLER_73_1592 ();
 sg13g2_fill_2 FILLER_73_1599 ();
 sg13g2_fill_2 FILLER_73_1642 ();
 sg13g2_fill_1 FILLER_73_1644 ();
 sg13g2_fill_1 FILLER_73_1650 ();
 sg13g2_fill_1 FILLER_73_1683 ();
 sg13g2_fill_2 FILLER_73_1738 ();
 sg13g2_decap_4 FILLER_73_1745 ();
 sg13g2_fill_2 FILLER_73_1749 ();
 sg13g2_fill_2 FILLER_73_1755 ();
 sg13g2_fill_2 FILLER_73_1774 ();
 sg13g2_decap_4 FILLER_73_1789 ();
 sg13g2_fill_1 FILLER_73_1793 ();
 sg13g2_decap_8 FILLER_73_1799 ();
 sg13g2_decap_8 FILLER_73_1806 ();
 sg13g2_decap_8 FILLER_73_1852 ();
 sg13g2_decap_8 FILLER_73_1859 ();
 sg13g2_decap_8 FILLER_73_1866 ();
 sg13g2_decap_8 FILLER_73_1873 ();
 sg13g2_decap_4 FILLER_73_1880 ();
 sg13g2_decap_4 FILLER_73_1888 ();
 sg13g2_fill_2 FILLER_73_1892 ();
 sg13g2_fill_2 FILLER_73_1899 ();
 sg13g2_fill_1 FILLER_73_1901 ();
 sg13g2_fill_2 FILLER_73_1913 ();
 sg13g2_fill_1 FILLER_73_1915 ();
 sg13g2_decap_8 FILLER_73_1921 ();
 sg13g2_decap_8 FILLER_73_1928 ();
 sg13g2_decap_8 FILLER_73_1935 ();
 sg13g2_decap_8 FILLER_73_1942 ();
 sg13g2_decap_8 FILLER_73_1949 ();
 sg13g2_decap_4 FILLER_73_1956 ();
 sg13g2_fill_1 FILLER_73_1960 ();
 sg13g2_fill_2 FILLER_73_1980 ();
 sg13g2_fill_1 FILLER_73_1982 ();
 sg13g2_decap_8 FILLER_73_1996 ();
 sg13g2_decap_8 FILLER_73_2003 ();
 sg13g2_fill_2 FILLER_73_2010 ();
 sg13g2_fill_1 FILLER_73_2012 ();
 sg13g2_decap_8 FILLER_73_2018 ();
 sg13g2_fill_2 FILLER_73_2025 ();
 sg13g2_fill_2 FILLER_73_2036 ();
 sg13g2_fill_1 FILLER_73_2038 ();
 sg13g2_fill_2 FILLER_73_2053 ();
 sg13g2_decap_8 FILLER_73_2060 ();
 sg13g2_fill_2 FILLER_73_2067 ();
 sg13g2_decap_4 FILLER_73_2073 ();
 sg13g2_decap_8 FILLER_73_2102 ();
 sg13g2_decap_8 FILLER_73_2109 ();
 sg13g2_decap_8 FILLER_73_2116 ();
 sg13g2_decap_8 FILLER_73_2123 ();
 sg13g2_decap_4 FILLER_73_2130 ();
 sg13g2_fill_2 FILLER_73_2134 ();
 sg13g2_fill_2 FILLER_73_2156 ();
 sg13g2_fill_1 FILLER_73_2158 ();
 sg13g2_fill_2 FILLER_73_2171 ();
 sg13g2_fill_2 FILLER_73_2178 ();
 sg13g2_fill_1 FILLER_73_2188 ();
 sg13g2_decap_4 FILLER_73_2193 ();
 sg13g2_fill_2 FILLER_73_2197 ();
 sg13g2_decap_4 FILLER_73_2226 ();
 sg13g2_fill_1 FILLER_73_2230 ();
 sg13g2_decap_8 FILLER_73_2253 ();
 sg13g2_fill_2 FILLER_73_2260 ();
 sg13g2_fill_1 FILLER_73_2262 ();
 sg13g2_decap_8 FILLER_73_2268 ();
 sg13g2_fill_2 FILLER_73_2275 ();
 sg13g2_fill_1 FILLER_73_2277 ();
 sg13g2_decap_8 FILLER_73_2291 ();
 sg13g2_fill_2 FILLER_73_2298 ();
 sg13g2_decap_4 FILLER_73_2305 ();
 sg13g2_fill_1 FILLER_73_2309 ();
 sg13g2_decap_8 FILLER_73_2333 ();
 sg13g2_decap_4 FILLER_73_2340 ();
 sg13g2_fill_2 FILLER_73_2400 ();
 sg13g2_decap_8 FILLER_73_2415 ();
 sg13g2_decap_8 FILLER_73_2422 ();
 sg13g2_decap_8 FILLER_73_2429 ();
 sg13g2_decap_8 FILLER_73_2436 ();
 sg13g2_decap_8 FILLER_73_2443 ();
 sg13g2_decap_8 FILLER_73_2450 ();
 sg13g2_decap_4 FILLER_73_2461 ();
 sg13g2_fill_2 FILLER_73_2465 ();
 sg13g2_decap_4 FILLER_73_2486 ();
 sg13g2_fill_1 FILLER_73_2490 ();
 sg13g2_decap_8 FILLER_73_2519 ();
 sg13g2_decap_8 FILLER_73_2526 ();
 sg13g2_decap_8 FILLER_73_2533 ();
 sg13g2_fill_1 FILLER_73_2540 ();
 sg13g2_fill_1 FILLER_73_2545 ();
 sg13g2_fill_2 FILLER_73_2573 ();
 sg13g2_decap_8 FILLER_73_2588 ();
 sg13g2_decap_4 FILLER_73_2595 ();
 sg13g2_fill_2 FILLER_73_2599 ();
 sg13g2_decap_8 FILLER_73_2636 ();
 sg13g2_decap_8 FILLER_73_2643 ();
 sg13g2_fill_1 FILLER_73_2691 ();
 sg13g2_decap_4 FILLER_73_2701 ();
 sg13g2_decap_4 FILLER_73_2719 ();
 sg13g2_decap_8 FILLER_73_2753 ();
 sg13g2_fill_2 FILLER_73_2760 ();
 sg13g2_decap_8 FILLER_73_2775 ();
 sg13g2_decap_8 FILLER_73_2782 ();
 sg13g2_decap_8 FILLER_73_2789 ();
 sg13g2_decap_4 FILLER_73_2848 ();
 sg13g2_fill_2 FILLER_73_2879 ();
 sg13g2_decap_8 FILLER_73_2921 ();
 sg13g2_decap_4 FILLER_73_2955 ();
 sg13g2_fill_1 FILLER_73_2959 ();
 sg13g2_decap_8 FILLER_73_2997 ();
 sg13g2_decap_8 FILLER_73_3004 ();
 sg13g2_fill_2 FILLER_73_3011 ();
 sg13g2_fill_1 FILLER_73_3013 ();
 sg13g2_decap_8 FILLER_73_3078 ();
 sg13g2_decap_4 FILLER_73_3085 ();
 sg13g2_fill_2 FILLER_73_3103 ();
 sg13g2_fill_1 FILLER_73_3105 ();
 sg13g2_fill_2 FILLER_73_3146 ();
 sg13g2_fill_1 FILLER_73_3148 ();
 sg13g2_decap_4 FILLER_73_3176 ();
 sg13g2_decap_8 FILLER_73_3229 ();
 sg13g2_decap_8 FILLER_73_3236 ();
 sg13g2_decap_8 FILLER_73_3243 ();
 sg13g2_decap_4 FILLER_73_3250 ();
 sg13g2_decap_8 FILLER_73_3258 ();
 sg13g2_decap_4 FILLER_73_3265 ();
 sg13g2_decap_4 FILLER_73_3291 ();
 sg13g2_fill_1 FILLER_73_3295 ();
 sg13g2_decap_4 FILLER_73_3309 ();
 sg13g2_decap_8 FILLER_73_3321 ();
 sg13g2_decap_8 FILLER_73_3328 ();
 sg13g2_decap_8 FILLER_73_3335 ();
 sg13g2_decap_8 FILLER_73_3342 ();
 sg13g2_decap_8 FILLER_73_3349 ();
 sg13g2_decap_4 FILLER_73_3360 ();
 sg13g2_fill_2 FILLER_73_3364 ();
 sg13g2_fill_1 FILLER_73_3376 ();
 sg13g2_decap_8 FILLER_73_3399 ();
 sg13g2_decap_8 FILLER_73_3406 ();
 sg13g2_fill_2 FILLER_73_3413 ();
 sg13g2_fill_2 FILLER_73_3430 ();
 sg13g2_decap_8 FILLER_73_3468 ();
 sg13g2_decap_4 FILLER_73_3475 ();
 sg13g2_fill_1 FILLER_73_3479 ();
 sg13g2_decap_8 FILLER_73_3513 ();
 sg13g2_decap_8 FILLER_73_3520 ();
 sg13g2_decap_4 FILLER_73_3527 ();
 sg13g2_fill_2 FILLER_73_3531 ();
 sg13g2_fill_2 FILLER_73_3554 ();
 sg13g2_fill_1 FILLER_73_3556 ();
 sg13g2_decap_8 FILLER_73_3566 ();
 sg13g2_decap_4 FILLER_73_3573 ();
 sg13g2_fill_1 FILLER_73_3577 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_11 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_102 ();
 sg13g2_fill_1 FILLER_74_109 ();
 sg13g2_decap_4 FILLER_74_124 ();
 sg13g2_fill_1 FILLER_74_218 ();
 sg13g2_fill_2 FILLER_74_247 ();
 sg13g2_fill_1 FILLER_74_249 ();
 sg13g2_fill_1 FILLER_74_296 ();
 sg13g2_decap_8 FILLER_74_339 ();
 sg13g2_decap_8 FILLER_74_346 ();
 sg13g2_decap_8 FILLER_74_353 ();
 sg13g2_fill_2 FILLER_74_372 ();
 sg13g2_fill_1 FILLER_74_374 ();
 sg13g2_fill_1 FILLER_74_388 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_4 FILLER_74_418 ();
 sg13g2_fill_1 FILLER_74_422 ();
 sg13g2_decap_8 FILLER_74_436 ();
 sg13g2_decap_8 FILLER_74_443 ();
 sg13g2_decap_8 FILLER_74_450 ();
 sg13g2_fill_2 FILLER_74_457 ();
 sg13g2_decap_8 FILLER_74_463 ();
 sg13g2_fill_1 FILLER_74_470 ();
 sg13g2_fill_2 FILLER_74_475 ();
 sg13g2_decap_8 FILLER_74_490 ();
 sg13g2_fill_2 FILLER_74_523 ();
 sg13g2_fill_1 FILLER_74_525 ();
 sg13g2_fill_1 FILLER_74_530 ();
 sg13g2_fill_2 FILLER_74_558 ();
 sg13g2_decap_8 FILLER_74_564 ();
 sg13g2_fill_2 FILLER_74_571 ();
 sg13g2_fill_1 FILLER_74_573 ();
 sg13g2_decap_4 FILLER_74_578 ();
 sg13g2_fill_2 FILLER_74_582 ();
 sg13g2_fill_1 FILLER_74_606 ();
 sg13g2_fill_2 FILLER_74_653 ();
 sg13g2_fill_1 FILLER_74_678 ();
 sg13g2_fill_2 FILLER_74_692 ();
 sg13g2_fill_2 FILLER_74_699 ();
 sg13g2_fill_1 FILLER_74_701 ();
 sg13g2_fill_2 FILLER_74_707 ();
 sg13g2_fill_1 FILLER_74_748 ();
 sg13g2_decap_8 FILLER_74_777 ();
 sg13g2_decap_8 FILLER_74_784 ();
 sg13g2_decap_4 FILLER_74_791 ();
 sg13g2_fill_2 FILLER_74_846 ();
 sg13g2_fill_1 FILLER_74_848 ();
 sg13g2_decap_4 FILLER_74_881 ();
 sg13g2_fill_2 FILLER_74_913 ();
 sg13g2_fill_1 FILLER_74_915 ();
 sg13g2_decap_4 FILLER_74_957 ();
 sg13g2_fill_2 FILLER_74_961 ();
 sg13g2_fill_2 FILLER_74_968 ();
 sg13g2_fill_1 FILLER_74_970 ();
 sg13g2_fill_2 FILLER_74_990 ();
 sg13g2_fill_1 FILLER_74_1017 ();
 sg13g2_fill_1 FILLER_74_1024 ();
 sg13g2_fill_1 FILLER_74_1040 ();
 sg13g2_decap_4 FILLER_74_1046 ();
 sg13g2_fill_1 FILLER_74_1050 ();
 sg13g2_decap_8 FILLER_74_1055 ();
 sg13g2_decap_8 FILLER_74_1065 ();
 sg13g2_decap_8 FILLER_74_1072 ();
 sg13g2_fill_1 FILLER_74_1104 ();
 sg13g2_fill_1 FILLER_74_1109 ();
 sg13g2_decap_8 FILLER_74_1153 ();
 sg13g2_decap_8 FILLER_74_1160 ();
 sg13g2_decap_8 FILLER_74_1167 ();
 sg13g2_decap_8 FILLER_74_1174 ();
 sg13g2_fill_2 FILLER_74_1181 ();
 sg13g2_fill_2 FILLER_74_1189 ();
 sg13g2_decap_8 FILLER_74_1195 ();
 sg13g2_fill_1 FILLER_74_1202 ();
 sg13g2_fill_1 FILLER_74_1209 ();
 sg13g2_decap_4 FILLER_74_1226 ();
 sg13g2_decap_8 FILLER_74_1241 ();
 sg13g2_decap_8 FILLER_74_1248 ();
 sg13g2_fill_1 FILLER_74_1255 ();
 sg13g2_fill_1 FILLER_74_1292 ();
 sg13g2_fill_2 FILLER_74_1375 ();
 sg13g2_fill_2 FILLER_74_1394 ();
 sg13g2_fill_1 FILLER_74_1396 ();
 sg13g2_fill_2 FILLER_74_1437 ();
 sg13g2_fill_1 FILLER_74_1439 ();
 sg13g2_decap_8 FILLER_74_1444 ();
 sg13g2_decap_8 FILLER_74_1451 ();
 sg13g2_fill_2 FILLER_74_1472 ();
 sg13g2_fill_1 FILLER_74_1474 ();
 sg13g2_fill_1 FILLER_74_1495 ();
 sg13g2_fill_2 FILLER_74_1502 ();
 sg13g2_fill_1 FILLER_74_1504 ();
 sg13g2_fill_2 FILLER_74_1523 ();
 sg13g2_decap_8 FILLER_74_1533 ();
 sg13g2_decap_8 FILLER_74_1591 ();
 sg13g2_decap_4 FILLER_74_1598 ();
 sg13g2_fill_1 FILLER_74_1602 ();
 sg13g2_decap_4 FILLER_74_1641 ();
 sg13g2_fill_1 FILLER_74_1712 ();
 sg13g2_fill_1 FILLER_74_1719 ();
 sg13g2_fill_1 FILLER_74_1729 ();
 sg13g2_fill_2 FILLER_74_1735 ();
 sg13g2_fill_1 FILLER_74_1737 ();
 sg13g2_fill_2 FILLER_74_1765 ();
 sg13g2_decap_8 FILLER_74_1786 ();
 sg13g2_decap_8 FILLER_74_1793 ();
 sg13g2_decap_8 FILLER_74_1800 ();
 sg13g2_decap_8 FILLER_74_1807 ();
 sg13g2_fill_2 FILLER_74_1814 ();
 sg13g2_fill_1 FILLER_74_1816 ();
 sg13g2_fill_1 FILLER_74_1838 ();
 sg13g2_decap_8 FILLER_74_1849 ();
 sg13g2_decap_8 FILLER_74_1856 ();
 sg13g2_decap_8 FILLER_74_1863 ();
 sg13g2_decap_8 FILLER_74_1870 ();
 sg13g2_decap_4 FILLER_74_1877 ();
 sg13g2_fill_1 FILLER_74_1894 ();
 sg13g2_decap_8 FILLER_74_1916 ();
 sg13g2_decap_8 FILLER_74_1923 ();
 sg13g2_decap_8 FILLER_74_1930 ();
 sg13g2_decap_4 FILLER_74_1937 ();
 sg13g2_fill_1 FILLER_74_1941 ();
 sg13g2_fill_1 FILLER_74_1945 ();
 sg13g2_decap_4 FILLER_74_1966 ();
 sg13g2_fill_2 FILLER_74_1970 ();
 sg13g2_decap_8 FILLER_74_1977 ();
 sg13g2_fill_2 FILLER_74_1984 ();
 sg13g2_fill_1 FILLER_74_1986 ();
 sg13g2_decap_8 FILLER_74_1995 ();
 sg13g2_fill_2 FILLER_74_2002 ();
 sg13g2_decap_8 FILLER_74_2019 ();
 sg13g2_decap_8 FILLER_74_2026 ();
 sg13g2_decap_8 FILLER_74_2033 ();
 sg13g2_decap_8 FILLER_74_2040 ();
 sg13g2_fill_1 FILLER_74_2047 ();
 sg13g2_decap_4 FILLER_74_2052 ();
 sg13g2_fill_1 FILLER_74_2056 ();
 sg13g2_decap_8 FILLER_74_2061 ();
 sg13g2_decap_4 FILLER_74_2083 ();
 sg13g2_fill_1 FILLER_74_2087 ();
 sg13g2_decap_8 FILLER_74_2098 ();
 sg13g2_decap_4 FILLER_74_2105 ();
 sg13g2_decap_4 FILLER_74_2119 ();
 sg13g2_fill_2 FILLER_74_2123 ();
 sg13g2_decap_4 FILLER_74_2155 ();
 sg13g2_decap_8 FILLER_74_2188 ();
 sg13g2_decap_8 FILLER_74_2195 ();
 sg13g2_decap_8 FILLER_74_2202 ();
 sg13g2_decap_8 FILLER_74_2209 ();
 sg13g2_fill_2 FILLER_74_2216 ();
 sg13g2_fill_1 FILLER_74_2218 ();
 sg13g2_decap_4 FILLER_74_2224 ();
 sg13g2_decap_8 FILLER_74_2233 ();
 sg13g2_decap_8 FILLER_74_2240 ();
 sg13g2_decap_8 FILLER_74_2267 ();
 sg13g2_fill_1 FILLER_74_2285 ();
 sg13g2_decap_8 FILLER_74_2302 ();
 sg13g2_fill_2 FILLER_74_2309 ();
 sg13g2_fill_1 FILLER_74_2311 ();
 sg13g2_decap_4 FILLER_74_2345 ();
 sg13g2_fill_1 FILLER_74_2349 ();
 sg13g2_fill_2 FILLER_74_2355 ();
 sg13g2_fill_1 FILLER_74_2375 ();
 sg13g2_fill_2 FILLER_74_2386 ();
 sg13g2_fill_1 FILLER_74_2398 ();
 sg13g2_decap_8 FILLER_74_2416 ();
 sg13g2_decap_8 FILLER_74_2423 ();
 sg13g2_decap_8 FILLER_74_2430 ();
 sg13g2_decap_8 FILLER_74_2437 ();
 sg13g2_fill_2 FILLER_74_2444 ();
 sg13g2_fill_2 FILLER_74_2456 ();
 sg13g2_decap_8 FILLER_74_2467 ();
 sg13g2_decap_8 FILLER_74_2474 ();
 sg13g2_decap_4 FILLER_74_2481 ();
 sg13g2_fill_2 FILLER_74_2485 ();
 sg13g2_decap_8 FILLER_74_2510 ();
 sg13g2_decap_8 FILLER_74_2517 ();
 sg13g2_decap_8 FILLER_74_2524 ();
 sg13g2_decap_8 FILLER_74_2531 ();
 sg13g2_decap_8 FILLER_74_2538 ();
 sg13g2_fill_2 FILLER_74_2545 ();
 sg13g2_decap_8 FILLER_74_2580 ();
 sg13g2_decap_8 FILLER_74_2587 ();
 sg13g2_decap_8 FILLER_74_2594 ();
 sg13g2_decap_8 FILLER_74_2601 ();
 sg13g2_fill_1 FILLER_74_2608 ();
 sg13g2_decap_8 FILLER_74_2641 ();
 sg13g2_decap_8 FILLER_74_2648 ();
 sg13g2_fill_2 FILLER_74_2672 ();
 sg13g2_fill_1 FILLER_74_2674 ();
 sg13g2_decap_8 FILLER_74_2702 ();
 sg13g2_fill_1 FILLER_74_2709 ();
 sg13g2_decap_8 FILLER_74_2737 ();
 sg13g2_fill_2 FILLER_74_2744 ();
 sg13g2_decap_8 FILLER_74_2773 ();
 sg13g2_decap_8 FILLER_74_2780 ();
 sg13g2_decap_4 FILLER_74_2787 ();
 sg13g2_decap_8 FILLER_74_2923 ();
 sg13g2_fill_2 FILLER_74_2930 ();
 sg13g2_fill_1 FILLER_74_2932 ();
 sg13g2_fill_2 FILLER_74_2968 ();
 sg13g2_decap_8 FILLER_74_2997 ();
 sg13g2_decap_8 FILLER_74_3004 ();
 sg13g2_fill_2 FILLER_74_3011 ();
 sg13g2_fill_2 FILLER_74_3053 ();
 sg13g2_decap_8 FILLER_74_3064 ();
 sg13g2_decap_8 FILLER_74_3071 ();
 sg13g2_decap_8 FILLER_74_3078 ();
 sg13g2_decap_8 FILLER_74_3085 ();
 sg13g2_decap_8 FILLER_74_3092 ();
 sg13g2_decap_8 FILLER_74_3099 ();
 sg13g2_decap_8 FILLER_74_3106 ();
 sg13g2_fill_1 FILLER_74_3113 ();
 sg13g2_decap_4 FILLER_74_3128 ();
 sg13g2_decap_8 FILLER_74_3141 ();
 sg13g2_decap_4 FILLER_74_3148 ();
 sg13g2_decap_8 FILLER_74_3190 ();
 sg13g2_fill_1 FILLER_74_3197 ();
 sg13g2_decap_8 FILLER_74_3229 ();
 sg13g2_decap_8 FILLER_74_3236 ();
 sg13g2_fill_2 FILLER_74_3243 ();
 sg13g2_fill_1 FILLER_74_3245 ();
 sg13g2_fill_2 FILLER_74_3256 ();
 sg13g2_decap_4 FILLER_74_3289 ();
 sg13g2_fill_2 FILLER_74_3293 ();
 sg13g2_decap_8 FILLER_74_3322 ();
 sg13g2_decap_8 FILLER_74_3329 ();
 sg13g2_fill_2 FILLER_74_3346 ();
 sg13g2_fill_1 FILLER_74_3348 ();
 sg13g2_fill_1 FILLER_74_3383 ();
 sg13g2_decap_8 FILLER_74_3393 ();
 sg13g2_decap_8 FILLER_74_3400 ();
 sg13g2_decap_4 FILLER_74_3407 ();
 sg13g2_fill_2 FILLER_74_3411 ();
 sg13g2_fill_1 FILLER_74_3440 ();
 sg13g2_decap_4 FILLER_74_3481 ();
 sg13g2_fill_1 FILLER_74_3485 ();
 sg13g2_decap_8 FILLER_74_3517 ();
 sg13g2_decap_8 FILLER_74_3524 ();
 sg13g2_decap_8 FILLER_74_3531 ();
 sg13g2_decap_8 FILLER_74_3538 ();
 sg13g2_decap_4 FILLER_74_3549 ();
 sg13g2_decap_8 FILLER_74_3562 ();
 sg13g2_decap_8 FILLER_74_3569 ();
 sg13g2_fill_2 FILLER_74_3576 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_fill_2 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_16 ();
 sg13g2_decap_8 FILLER_75_57 ();
 sg13g2_decap_8 FILLER_75_64 ();
 sg13g2_decap_4 FILLER_75_71 ();
 sg13g2_fill_2 FILLER_75_75 ();
 sg13g2_decap_8 FILLER_75_90 ();
 sg13g2_decap_8 FILLER_75_97 ();
 sg13g2_decap_4 FILLER_75_104 ();
 sg13g2_fill_2 FILLER_75_135 ();
 sg13g2_fill_1 FILLER_75_137 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_fill_2 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_235 ();
 sg13g2_decap_8 FILLER_75_242 ();
 sg13g2_decap_8 FILLER_75_249 ();
 sg13g2_fill_2 FILLER_75_256 ();
 sg13g2_fill_1 FILLER_75_267 ();
 sg13g2_fill_1 FILLER_75_277 ();
 sg13g2_fill_1 FILLER_75_290 ();
 sg13g2_decap_4 FILLER_75_324 ();
 sg13g2_fill_2 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_decap_8 FILLER_75_342 ();
 sg13g2_fill_2 FILLER_75_349 ();
 sg13g2_fill_1 FILLER_75_351 ();
 sg13g2_decap_8 FILLER_75_445 ();
 sg13g2_decap_8 FILLER_75_452 ();
 sg13g2_decap_8 FILLER_75_459 ();
 sg13g2_fill_2 FILLER_75_502 ();
 sg13g2_fill_1 FILLER_75_504 ();
 sg13g2_decap_4 FILLER_75_509 ();
 sg13g2_decap_4 FILLER_75_563 ();
 sg13g2_fill_2 FILLER_75_567 ();
 sg13g2_fill_2 FILLER_75_609 ();
 sg13g2_fill_2 FILLER_75_615 ();
 sg13g2_fill_1 FILLER_75_617 ();
 sg13g2_decap_8 FILLER_75_622 ();
 sg13g2_fill_2 FILLER_75_629 ();
 sg13g2_fill_2 FILLER_75_662 ();
 sg13g2_fill_1 FILLER_75_673 ();
 sg13g2_decap_4 FILLER_75_706 ();
 sg13g2_decap_4 FILLER_75_720 ();
 sg13g2_fill_2 FILLER_75_724 ();
 sg13g2_decap_8 FILLER_75_753 ();
 sg13g2_decap_8 FILLER_75_760 ();
 sg13g2_decap_8 FILLER_75_767 ();
 sg13g2_decap_8 FILLER_75_774 ();
 sg13g2_decap_8 FILLER_75_781 ();
 sg13g2_fill_2 FILLER_75_788 ();
 sg13g2_fill_1 FILLER_75_790 ();
 sg13g2_decap_8 FILLER_75_888 ();
 sg13g2_decap_8 FILLER_75_913 ();
 sg13g2_fill_1 FILLER_75_920 ();
 sg13g2_decap_8 FILLER_75_939 ();
 sg13g2_fill_2 FILLER_75_946 ();
 sg13g2_fill_1 FILLER_75_948 ();
 sg13g2_decap_8 FILLER_75_954 ();
 sg13g2_decap_8 FILLER_75_961 ();
 sg13g2_decap_8 FILLER_75_968 ();
 sg13g2_fill_2 FILLER_75_975 ();
 sg13g2_fill_2 FILLER_75_992 ();
 sg13g2_fill_1 FILLER_75_994 ();
 sg13g2_decap_8 FILLER_75_1039 ();
 sg13g2_decap_4 FILLER_75_1046 ();
 sg13g2_fill_1 FILLER_75_1050 ();
 sg13g2_fill_2 FILLER_75_1058 ();
 sg13g2_decap_4 FILLER_75_1084 ();
 sg13g2_fill_2 FILLER_75_1092 ();
 sg13g2_fill_1 FILLER_75_1110 ();
 sg13g2_decap_8 FILLER_75_1153 ();
 sg13g2_decap_8 FILLER_75_1160 ();
 sg13g2_decap_4 FILLER_75_1167 ();
 sg13g2_fill_2 FILLER_75_1192 ();
 sg13g2_fill_2 FILLER_75_1230 ();
 sg13g2_decap_8 FILLER_75_1241 ();
 sg13g2_decap_8 FILLER_75_1248 ();
 sg13g2_fill_2 FILLER_75_1255 ();
 sg13g2_decap_4 FILLER_75_1266 ();
 sg13g2_decap_8 FILLER_75_1283 ();
 sg13g2_decap_4 FILLER_75_1290 ();
 sg13g2_fill_1 FILLER_75_1294 ();
 sg13g2_fill_2 FILLER_75_1340 ();
 sg13g2_fill_1 FILLER_75_1342 ();
 sg13g2_fill_1 FILLER_75_1403 ();
 sg13g2_decap_8 FILLER_75_1497 ();
 sg13g2_fill_2 FILLER_75_1504 ();
 sg13g2_decap_8 FILLER_75_1515 ();
 sg13g2_decap_8 FILLER_75_1522 ();
 sg13g2_decap_8 FILLER_75_1529 ();
 sg13g2_decap_4 FILLER_75_1536 ();
 sg13g2_fill_2 FILLER_75_1540 ();
 sg13g2_decap_8 FILLER_75_1554 ();
 sg13g2_fill_1 FILLER_75_1561 ();
 sg13g2_decap_8 FILLER_75_1579 ();
 sg13g2_decap_8 FILLER_75_1586 ();
 sg13g2_decap_8 FILLER_75_1593 ();
 sg13g2_decap_8 FILLER_75_1600 ();
 sg13g2_decap_8 FILLER_75_1607 ();
 sg13g2_decap_4 FILLER_75_1614 ();
 sg13g2_decap_8 FILLER_75_1631 ();
 sg13g2_decap_8 FILLER_75_1638 ();
 sg13g2_fill_1 FILLER_75_1645 ();
 sg13g2_fill_2 FILLER_75_1751 ();
 sg13g2_fill_2 FILLER_75_1774 ();
 sg13g2_decap_8 FILLER_75_1789 ();
 sg13g2_decap_4 FILLER_75_1796 ();
 sg13g2_decap_4 FILLER_75_1816 ();
 sg13g2_fill_1 FILLER_75_1820 ();
 sg13g2_decap_4 FILLER_75_1831 ();
 sg13g2_fill_1 FILLER_75_1835 ();
 sg13g2_decap_8 FILLER_75_1853 ();
 sg13g2_decap_8 FILLER_75_1860 ();
 sg13g2_decap_8 FILLER_75_1867 ();
 sg13g2_fill_2 FILLER_75_1874 ();
 sg13g2_fill_1 FILLER_75_1876 ();
 sg13g2_decap_8 FILLER_75_1917 ();
 sg13g2_decap_8 FILLER_75_1924 ();
 sg13g2_fill_1 FILLER_75_1931 ();
 sg13g2_fill_2 FILLER_75_1963 ();
 sg13g2_decap_8 FILLER_75_1973 ();
 sg13g2_fill_2 FILLER_75_1980 ();
 sg13g2_fill_1 FILLER_75_1982 ();
 sg13g2_fill_1 FILLER_75_2034 ();
 sg13g2_decap_4 FILLER_75_2048 ();
 sg13g2_fill_1 FILLER_75_2057 ();
 sg13g2_fill_1 FILLER_75_2073 ();
 sg13g2_decap_8 FILLER_75_2094 ();
 sg13g2_decap_8 FILLER_75_2101 ();
 sg13g2_decap_8 FILLER_75_2108 ();
 sg13g2_decap_8 FILLER_75_2115 ();
 sg13g2_fill_2 FILLER_75_2122 ();
 sg13g2_decap_8 FILLER_75_2154 ();
 sg13g2_decap_4 FILLER_75_2161 ();
 sg13g2_fill_1 FILLER_75_2170 ();
 sg13g2_decap_8 FILLER_75_2184 ();
 sg13g2_decap_8 FILLER_75_2191 ();
 sg13g2_fill_2 FILLER_75_2198 ();
 sg13g2_fill_1 FILLER_75_2200 ();
 sg13g2_decap_4 FILLER_75_2206 ();
 sg13g2_decap_8 FILLER_75_2220 ();
 sg13g2_fill_2 FILLER_75_2227 ();
 sg13g2_fill_1 FILLER_75_2229 ();
 sg13g2_decap_8 FILLER_75_2235 ();
 sg13g2_decap_8 FILLER_75_2242 ();
 sg13g2_decap_8 FILLER_75_2254 ();
 sg13g2_decap_8 FILLER_75_2261 ();
 sg13g2_decap_4 FILLER_75_2268 ();
 sg13g2_decap_8 FILLER_75_2278 ();
 sg13g2_decap_8 FILLER_75_2285 ();
 sg13g2_decap_4 FILLER_75_2292 ();
 sg13g2_decap_8 FILLER_75_2304 ();
 sg13g2_decap_8 FILLER_75_2311 ();
 sg13g2_decap_8 FILLER_75_2318 ();
 sg13g2_decap_4 FILLER_75_2325 ();
 sg13g2_decap_8 FILLER_75_2341 ();
 sg13g2_decap_8 FILLER_75_2348 ();
 sg13g2_decap_8 FILLER_75_2355 ();
 sg13g2_fill_2 FILLER_75_2362 ();
 sg13g2_fill_1 FILLER_75_2373 ();
 sg13g2_fill_2 FILLER_75_2388 ();
 sg13g2_decap_8 FILLER_75_2411 ();
 sg13g2_decap_4 FILLER_75_2418 ();
 sg13g2_fill_1 FILLER_75_2422 ();
 sg13g2_fill_2 FILLER_75_2432 ();
 sg13g2_fill_1 FILLER_75_2434 ();
 sg13g2_fill_2 FILLER_75_2479 ();
 sg13g2_fill_1 FILLER_75_2481 ();
 sg13g2_decap_8 FILLER_75_2513 ();
 sg13g2_decap_8 FILLER_75_2520 ();
 sg13g2_decap_8 FILLER_75_2527 ();
 sg13g2_fill_1 FILLER_75_2534 ();
 sg13g2_fill_2 FILLER_75_2576 ();
 sg13g2_fill_2 FILLER_75_2591 ();
 sg13g2_fill_1 FILLER_75_2593 ();
 sg13g2_decap_8 FILLER_75_2625 ();
 sg13g2_decap_8 FILLER_75_2632 ();
 sg13g2_decap_8 FILLER_75_2639 ();
 sg13g2_fill_1 FILLER_75_2646 ();
 sg13g2_fill_1 FILLER_75_2651 ();
 sg13g2_fill_2 FILLER_75_2662 ();
 sg13g2_fill_1 FILLER_75_2664 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_decap_8 FILLER_75_2679 ();
 sg13g2_decap_8 FILLER_75_2686 ();
 sg13g2_decap_4 FILLER_75_2693 ();
 sg13g2_decap_4 FILLER_75_2734 ();
 sg13g2_fill_1 FILLER_75_2738 ();
 sg13g2_fill_2 FILLER_75_2749 ();
 sg13g2_fill_1 FILLER_75_2751 ();
 sg13g2_decap_8 FILLER_75_2779 ();
 sg13g2_decap_4 FILLER_75_2786 ();
 sg13g2_fill_2 FILLER_75_2837 ();
 sg13g2_fill_2 FILLER_75_2849 ();
 sg13g2_fill_2 FILLER_75_2860 ();
 sg13g2_fill_1 FILLER_75_2862 ();
 sg13g2_fill_1 FILLER_75_2886 ();
 sg13g2_decap_4 FILLER_75_2891 ();
 sg13g2_decap_8 FILLER_75_2916 ();
 sg13g2_decap_8 FILLER_75_2923 ();
 sg13g2_decap_8 FILLER_75_2930 ();
 sg13g2_decap_8 FILLER_75_2937 ();
 sg13g2_fill_1 FILLER_75_2944 ();
 sg13g2_decap_8 FILLER_75_2973 ();
 sg13g2_decap_8 FILLER_75_2989 ();
 sg13g2_decap_8 FILLER_75_2996 ();
 sg13g2_decap_8 FILLER_75_3003 ();
 sg13g2_fill_2 FILLER_75_3010 ();
 sg13g2_fill_1 FILLER_75_3012 ();
 sg13g2_fill_2 FILLER_75_3043 ();
 sg13g2_decap_8 FILLER_75_3064 ();
 sg13g2_decap_8 FILLER_75_3071 ();
 sg13g2_fill_1 FILLER_75_3078 ();
 sg13g2_decap_8 FILLER_75_3088 ();
 sg13g2_decap_4 FILLER_75_3095 ();
 sg13g2_fill_1 FILLER_75_3099 ();
 sg13g2_decap_4 FILLER_75_3114 ();
 sg13g2_fill_1 FILLER_75_3118 ();
 sg13g2_decap_8 FILLER_75_3146 ();
 sg13g2_decap_4 FILLER_75_3153 ();
 sg13g2_fill_1 FILLER_75_3157 ();
 sg13g2_decap_8 FILLER_75_3180 ();
 sg13g2_decap_8 FILLER_75_3187 ();
 sg13g2_decap_4 FILLER_75_3194 ();
 sg13g2_fill_1 FILLER_75_3198 ();
 sg13g2_decap_8 FILLER_75_3221 ();
 sg13g2_decap_8 FILLER_75_3228 ();
 sg13g2_decap_8 FILLER_75_3235 ();
 sg13g2_fill_1 FILLER_75_3242 ();
 sg13g2_decap_4 FILLER_75_3270 ();
 sg13g2_fill_2 FILLER_75_3274 ();
 sg13g2_decap_4 FILLER_75_3303 ();
 sg13g2_fill_2 FILLER_75_3307 ();
 sg13g2_decap_8 FILLER_75_3318 ();
 sg13g2_fill_1 FILLER_75_3325 ();
 sg13g2_decap_4 FILLER_75_3357 ();
 sg13g2_fill_2 FILLER_75_3371 ();
 sg13g2_decap_8 FILLER_75_3400 ();
 sg13g2_decap_8 FILLER_75_3457 ();
 sg13g2_decap_8 FILLER_75_3464 ();
 sg13g2_decap_8 FILLER_75_3471 ();
 sg13g2_fill_2 FILLER_75_3478 ();
 sg13g2_fill_1 FILLER_75_3480 ();
 sg13g2_decap_8 FILLER_75_3517 ();
 sg13g2_decap_8 FILLER_75_3524 ();
 sg13g2_decap_8 FILLER_75_3531 ();
 sg13g2_decap_8 FILLER_75_3538 ();
 sg13g2_decap_8 FILLER_75_3545 ();
 sg13g2_decap_8 FILLER_75_3552 ();
 sg13g2_decap_8 FILLER_75_3559 ();
 sg13g2_decap_8 FILLER_75_3566 ();
 sg13g2_decap_4 FILLER_75_3573 ();
 sg13g2_fill_1 FILLER_75_3577 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_fill_1 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_48 ();
 sg13g2_decap_8 FILLER_76_55 ();
 sg13g2_decap_8 FILLER_76_62 ();
 sg13g2_decap_8 FILLER_76_69 ();
 sg13g2_decap_8 FILLER_76_76 ();
 sg13g2_decap_8 FILLER_76_83 ();
 sg13g2_decap_8 FILLER_76_90 ();
 sg13g2_decap_8 FILLER_76_97 ();
 sg13g2_decap_8 FILLER_76_104 ();
 sg13g2_fill_2 FILLER_76_111 ();
 sg13g2_decap_4 FILLER_76_117 ();
 sg13g2_fill_2 FILLER_76_121 ();
 sg13g2_decap_4 FILLER_76_153 ();
 sg13g2_fill_1 FILLER_76_157 ();
 sg13g2_decap_4 FILLER_76_166 ();
 sg13g2_fill_2 FILLER_76_170 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_2 FILLER_76_186 ();
 sg13g2_fill_1 FILLER_76_188 ();
 sg13g2_decap_8 FILLER_76_202 ();
 sg13g2_decap_8 FILLER_76_209 ();
 sg13g2_decap_8 FILLER_76_216 ();
 sg13g2_decap_8 FILLER_76_223 ();
 sg13g2_fill_2 FILLER_76_230 ();
 sg13g2_fill_1 FILLER_76_249 ();
 sg13g2_decap_4 FILLER_76_259 ();
 sg13g2_fill_1 FILLER_76_263 ();
 sg13g2_decap_8 FILLER_76_332 ();
 sg13g2_decap_8 FILLER_76_339 ();
 sg13g2_decap_8 FILLER_76_346 ();
 sg13g2_decap_4 FILLER_76_375 ();
 sg13g2_fill_2 FILLER_76_401 ();
 sg13g2_fill_1 FILLER_76_403 ();
 sg13g2_fill_2 FILLER_76_453 ();
 sg13g2_decap_4 FILLER_76_513 ();
 sg13g2_decap_4 FILLER_76_547 ();
 sg13g2_fill_1 FILLER_76_551 ();
 sg13g2_fill_2 FILLER_76_561 ();
 sg13g2_decap_4 FILLER_76_576 ();
 sg13g2_fill_1 FILLER_76_580 ();
 sg13g2_fill_2 FILLER_76_591 ();
 sg13g2_decap_8 FILLER_76_614 ();
 sg13g2_decap_4 FILLER_76_621 ();
 sg13g2_fill_1 FILLER_76_625 ();
 sg13g2_fill_2 FILLER_76_691 ();
 sg13g2_decap_8 FILLER_76_698 ();
 sg13g2_decap_8 FILLER_76_705 ();
 sg13g2_decap_8 FILLER_76_712 ();
 sg13g2_decap_4 FILLER_76_719 ();
 sg13g2_fill_1 FILLER_76_732 ();
 sg13g2_decap_8 FILLER_76_746 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_decap_8 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_767 ();
 sg13g2_decap_4 FILLER_76_774 ();
 sg13g2_fill_2 FILLER_76_778 ();
 sg13g2_fill_2 FILLER_76_789 ();
 sg13g2_fill_1 FILLER_76_791 ();
 sg13g2_fill_2 FILLER_76_834 ();
 sg13g2_fill_1 FILLER_76_836 ();
 sg13g2_fill_1 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_856 ();
 sg13g2_decap_8 FILLER_76_863 ();
 sg13g2_fill_2 FILLER_76_870 ();
 sg13g2_fill_1 FILLER_76_872 ();
 sg13g2_decap_8 FILLER_76_878 ();
 sg13g2_fill_2 FILLER_76_885 ();
 sg13g2_decap_8 FILLER_76_896 ();
 sg13g2_fill_1 FILLER_76_907 ();
 sg13g2_decap_8 FILLER_76_912 ();
 sg13g2_fill_1 FILLER_76_919 ();
 sg13g2_fill_2 FILLER_76_925 ();
 sg13g2_decap_8 FILLER_76_931 ();
 sg13g2_decap_8 FILLER_76_938 ();
 sg13g2_decap_8 FILLER_76_945 ();
 sg13g2_decap_8 FILLER_76_952 ();
 sg13g2_decap_4 FILLER_76_959 ();
 sg13g2_decap_8 FILLER_76_989 ();
 sg13g2_decap_8 FILLER_76_996 ();
 sg13g2_fill_1 FILLER_76_1003 ();
 sg13g2_fill_1 FILLER_76_1022 ();
 sg13g2_decap_8 FILLER_76_1028 ();
 sg13g2_decap_8 FILLER_76_1035 ();
 sg13g2_decap_8 FILLER_76_1042 ();
 sg13g2_decap_8 FILLER_76_1049 ();
 sg13g2_decap_8 FILLER_76_1056 ();
 sg13g2_decap_8 FILLER_76_1063 ();
 sg13g2_decap_8 FILLER_76_1070 ();
 sg13g2_decap_8 FILLER_76_1077 ();
 sg13g2_decap_8 FILLER_76_1084 ();
 sg13g2_decap_4 FILLER_76_1091 ();
 sg13g2_fill_2 FILLER_76_1095 ();
 sg13g2_decap_4 FILLER_76_1119 ();
 sg13g2_decap_8 FILLER_76_1148 ();
 sg13g2_decap_8 FILLER_76_1155 ();
 sg13g2_fill_1 FILLER_76_1162 ();
 sg13g2_decap_8 FILLER_76_1180 ();
 sg13g2_fill_1 FILLER_76_1187 ();
 sg13g2_decap_8 FILLER_76_1197 ();
 sg13g2_fill_2 FILLER_76_1204 ();
 sg13g2_fill_1 FILLER_76_1206 ();
 sg13g2_fill_2 FILLER_76_1210 ();
 sg13g2_decap_4 FILLER_76_1263 ();
 sg13g2_decap_8 FILLER_76_1280 ();
 sg13g2_decap_8 FILLER_76_1287 ();
 sg13g2_decap_4 FILLER_76_1294 ();
 sg13g2_fill_1 FILLER_76_1349 ();
 sg13g2_fill_2 FILLER_76_1397 ();
 sg13g2_fill_1 FILLER_76_1399 ();
 sg13g2_fill_2 FILLER_76_1440 ();
 sg13g2_fill_1 FILLER_76_1447 ();
 sg13g2_fill_2 FILLER_76_1480 ();
 sg13g2_fill_1 FILLER_76_1482 ();
 sg13g2_decap_8 FILLER_76_1524 ();
 sg13g2_decap_4 FILLER_76_1531 ();
 sg13g2_fill_2 FILLER_76_1535 ();
 sg13g2_fill_1 FILLER_76_1546 ();
 sg13g2_fill_2 FILLER_76_1564 ();
 sg13g2_fill_1 FILLER_76_1566 ();
 sg13g2_decap_8 FILLER_76_1590 ();
 sg13g2_decap_8 FILLER_76_1597 ();
 sg13g2_decap_4 FILLER_76_1604 ();
 sg13g2_fill_2 FILLER_76_1608 ();
 sg13g2_decap_8 FILLER_76_1615 ();
 sg13g2_fill_2 FILLER_76_1622 ();
 sg13g2_decap_4 FILLER_76_1637 ();
 sg13g2_fill_2 FILLER_76_1641 ();
 sg13g2_fill_1 FILLER_76_1674 ();
 sg13g2_fill_1 FILLER_76_1729 ();
 sg13g2_fill_2 FILLER_76_1757 ();
 sg13g2_decap_8 FILLER_76_1785 ();
 sg13g2_decap_8 FILLER_76_1792 ();
 sg13g2_decap_4 FILLER_76_1799 ();
 sg13g2_fill_2 FILLER_76_1803 ();
 sg13g2_fill_2 FILLER_76_1813 ();
 sg13g2_fill_2 FILLER_76_1823 ();
 sg13g2_decap_8 FILLER_76_1846 ();
 sg13g2_decap_4 FILLER_76_1853 ();
 sg13g2_fill_1 FILLER_76_1857 ();
 sg13g2_decap_8 FILLER_76_1871 ();
 sg13g2_decap_4 FILLER_76_1878 ();
 sg13g2_fill_2 FILLER_76_1882 ();
 sg13g2_fill_2 FILLER_76_1894 ();
 sg13g2_decap_8 FILLER_76_1907 ();
 sg13g2_fill_2 FILLER_76_1914 ();
 sg13g2_fill_2 FILLER_76_1921 ();
 sg13g2_fill_1 FILLER_76_1923 ();
 sg13g2_fill_1 FILLER_76_1938 ();
 sg13g2_fill_2 FILLER_76_1957 ();
 sg13g2_fill_1 FILLER_76_1959 ();
 sg13g2_fill_2 FILLER_76_1972 ();
 sg13g2_fill_2 FILLER_76_1983 ();
 sg13g2_fill_1 FILLER_76_1991 ();
 sg13g2_decap_4 FILLER_76_2007 ();
 sg13g2_fill_1 FILLER_76_2023 ();
 sg13g2_decap_8 FILLER_76_2035 ();
 sg13g2_decap_8 FILLER_76_2042 ();
 sg13g2_decap_8 FILLER_76_2049 ();
 sg13g2_fill_1 FILLER_76_2067 ();
 sg13g2_fill_2 FILLER_76_2093 ();
 sg13g2_fill_2 FILLER_76_2105 ();
 sg13g2_fill_1 FILLER_76_2107 ();
 sg13g2_decap_8 FILLER_76_2113 ();
 sg13g2_fill_1 FILLER_76_2120 ();
 sg13g2_decap_8 FILLER_76_2131 ();
 sg13g2_decap_8 FILLER_76_2138 ();
 sg13g2_decap_4 FILLER_76_2145 ();
 sg13g2_fill_2 FILLER_76_2149 ();
 sg13g2_decap_8 FILLER_76_2170 ();
 sg13g2_decap_8 FILLER_76_2177 ();
 sg13g2_decap_8 FILLER_76_2184 ();
 sg13g2_decap_8 FILLER_76_2191 ();
 sg13g2_fill_1 FILLER_76_2198 ();
 sg13g2_fill_2 FILLER_76_2254 ();
 sg13g2_fill_1 FILLER_76_2265 ();
 sg13g2_fill_1 FILLER_76_2281 ();
 sg13g2_decap_8 FILLER_76_2291 ();
 sg13g2_decap_8 FILLER_76_2298 ();
 sg13g2_decap_8 FILLER_76_2305 ();
 sg13g2_decap_4 FILLER_76_2312 ();
 sg13g2_fill_1 FILLER_76_2316 ();
 sg13g2_fill_1 FILLER_76_2322 ();
 sg13g2_decap_8 FILLER_76_2357 ();
 sg13g2_fill_1 FILLER_76_2376 ();
 sg13g2_decap_8 FILLER_76_2410 ();
 sg13g2_decap_8 FILLER_76_2417 ();
 sg13g2_decap_8 FILLER_76_2424 ();
 sg13g2_decap_4 FILLER_76_2431 ();
 sg13g2_decap_4 FILLER_76_2472 ();
 sg13g2_fill_2 FILLER_76_2476 ();
 sg13g2_decap_8 FILLER_76_2518 ();
 sg13g2_fill_2 FILLER_76_2525 ();
 sg13g2_decap_4 FILLER_76_2584 ();
 sg13g2_fill_1 FILLER_76_2588 ();
 sg13g2_decap_8 FILLER_76_2629 ();
 sg13g2_decap_8 FILLER_76_2636 ();
 sg13g2_fill_2 FILLER_76_2653 ();
 sg13g2_decap_8 FILLER_76_2691 ();
 sg13g2_decap_4 FILLER_76_2698 ();
 sg13g2_fill_2 FILLER_76_2702 ();
 sg13g2_fill_1 FILLER_76_2718 ();
 sg13g2_fill_2 FILLER_76_2741 ();
 sg13g2_fill_1 FILLER_76_2757 ();
 sg13g2_decap_8 FILLER_76_2776 ();
 sg13g2_decap_8 FILLER_76_2783 ();
 sg13g2_decap_4 FILLER_76_2790 ();
 sg13g2_fill_1 FILLER_76_2794 ();
 sg13g2_fill_1 FILLER_76_2799 ();
 sg13g2_decap_8 FILLER_76_2804 ();
 sg13g2_decap_8 FILLER_76_2850 ();
 sg13g2_fill_2 FILLER_76_2857 ();
 sg13g2_decap_8 FILLER_76_2863 ();
 sg13g2_decap_8 FILLER_76_2870 ();
 sg13g2_fill_1 FILLER_76_2877 ();
 sg13g2_decap_8 FILLER_76_2887 ();
 sg13g2_decap_8 FILLER_76_2894 ();
 sg13g2_decap_4 FILLER_76_2901 ();
 sg13g2_fill_1 FILLER_76_2905 ();
 sg13g2_decap_8 FILLER_76_2916 ();
 sg13g2_decap_8 FILLER_76_2923 ();
 sg13g2_decap_8 FILLER_76_2930 ();
 sg13g2_decap_8 FILLER_76_2937 ();
 sg13g2_decap_8 FILLER_76_2944 ();
 sg13g2_decap_4 FILLER_76_2951 ();
 sg13g2_fill_2 FILLER_76_2955 ();
 sg13g2_decap_8 FILLER_76_2978 ();
 sg13g2_decap_8 FILLER_76_2985 ();
 sg13g2_decap_8 FILLER_76_2992 ();
 sg13g2_decap_8 FILLER_76_2999 ();
 sg13g2_decap_8 FILLER_76_3006 ();
 sg13g2_fill_2 FILLER_76_3013 ();
 sg13g2_decap_8 FILLER_76_3046 ();
 sg13g2_decap_4 FILLER_76_3053 ();
 sg13g2_fill_2 FILLER_76_3057 ();
 sg13g2_decap_8 FILLER_76_3096 ();
 sg13g2_fill_2 FILLER_76_3103 ();
 sg13g2_fill_2 FILLER_76_3153 ();
 sg13g2_fill_1 FILLER_76_3155 ();
 sg13g2_decap_8 FILLER_76_3166 ();
 sg13g2_decap_8 FILLER_76_3182 ();
 sg13g2_decap_4 FILLER_76_3189 ();
 sg13g2_fill_2 FILLER_76_3203 ();
 sg13g2_fill_1 FILLER_76_3205 ();
 sg13g2_fill_2 FILLER_76_3246 ();
 sg13g2_fill_1 FILLER_76_3248 ();
 sg13g2_fill_2 FILLER_76_3253 ();
 sg13g2_decap_8 FILLER_76_3305 ();
 sg13g2_decap_8 FILLER_76_3312 ();
 sg13g2_decap_8 FILLER_76_3319 ();
 sg13g2_decap_8 FILLER_76_3326 ();
 sg13g2_decap_8 FILLER_76_3343 ();
 sg13g2_decap_8 FILLER_76_3350 ();
 sg13g2_fill_2 FILLER_76_3357 ();
 sg13g2_decap_8 FILLER_76_3390 ();
 sg13g2_decap_8 FILLER_76_3397 ();
 sg13g2_decap_8 FILLER_76_3404 ();
 sg13g2_decap_4 FILLER_76_3411 ();
 sg13g2_fill_2 FILLER_76_3429 ();
 sg13g2_fill_1 FILLER_76_3431 ();
 sg13g2_fill_2 FILLER_76_3445 ();
 sg13g2_fill_1 FILLER_76_3447 ();
 sg13g2_decap_8 FILLER_76_3452 ();
 sg13g2_decap_8 FILLER_76_3459 ();
 sg13g2_decap_8 FILLER_76_3466 ();
 sg13g2_decap_8 FILLER_76_3473 ();
 sg13g2_decap_4 FILLER_76_3480 ();
 sg13g2_fill_2 FILLER_76_3484 ();
 sg13g2_decap_4 FILLER_76_3490 ();
 sg13g2_fill_2 FILLER_76_3494 ();
 sg13g2_decap_8 FILLER_76_3505 ();
 sg13g2_decap_8 FILLER_76_3512 ();
 sg13g2_decap_8 FILLER_76_3519 ();
 sg13g2_decap_8 FILLER_76_3526 ();
 sg13g2_decap_8 FILLER_76_3533 ();
 sg13g2_decap_8 FILLER_76_3540 ();
 sg13g2_decap_8 FILLER_76_3547 ();
 sg13g2_decap_8 FILLER_76_3554 ();
 sg13g2_decap_8 FILLER_76_3561 ();
 sg13g2_decap_8 FILLER_76_3568 ();
 sg13g2_fill_2 FILLER_76_3575 ();
 sg13g2_fill_1 FILLER_76_3577 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_fill_2 FILLER_77_112 ();
 sg13g2_fill_1 FILLER_77_114 ();
 sg13g2_decap_4 FILLER_77_119 ();
 sg13g2_fill_2 FILLER_77_156 ();
 sg13g2_decap_8 FILLER_77_167 ();
 sg13g2_decap_8 FILLER_77_218 ();
 sg13g2_decap_4 FILLER_77_225 ();
 sg13g2_fill_1 FILLER_77_229 ();
 sg13g2_decap_8 FILLER_77_339 ();
 sg13g2_decap_4 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_379 ();
 sg13g2_fill_1 FILLER_77_395 ();
 sg13g2_fill_1 FILLER_77_456 ();
 sg13g2_fill_2 FILLER_77_512 ();
 sg13g2_fill_1 FILLER_77_514 ();
 sg13g2_decap_8 FILLER_77_564 ();
 sg13g2_fill_2 FILLER_77_581 ();
 sg13g2_fill_1 FILLER_77_583 ();
 sg13g2_decap_4 FILLER_77_615 ();
 sg13g2_fill_2 FILLER_77_619 ();
 sg13g2_fill_2 FILLER_77_680 ();
 sg13g2_decap_8 FILLER_77_766 ();
 sg13g2_decap_4 FILLER_77_773 ();
 sg13g2_fill_2 FILLER_77_777 ();
 sg13g2_fill_1 FILLER_77_848 ();
 sg13g2_fill_2 FILLER_77_859 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_fill_1 FILLER_77_902 ();
 sg13g2_fill_1 FILLER_77_939 ();
 sg13g2_fill_2 FILLER_77_945 ();
 sg13g2_decap_8 FILLER_77_1001 ();
 sg13g2_fill_2 FILLER_77_1008 ();
 sg13g2_fill_1 FILLER_77_1020 ();
 sg13g2_decap_8 FILLER_77_1049 ();
 sg13g2_decap_8 FILLER_77_1056 ();
 sg13g2_decap_8 FILLER_77_1063 ();
 sg13g2_decap_8 FILLER_77_1070 ();
 sg13g2_fill_1 FILLER_77_1077 ();
 sg13g2_decap_8 FILLER_77_1087 ();
 sg13g2_fill_2 FILLER_77_1094 ();
 sg13g2_fill_1 FILLER_77_1119 ();
 sg13g2_decap_8 FILLER_77_1146 ();
 sg13g2_fill_1 FILLER_77_1153 ();
 sg13g2_decap_8 FILLER_77_1191 ();
 sg13g2_decap_8 FILLER_77_1198 ();
 sg13g2_fill_2 FILLER_77_1205 ();
 sg13g2_fill_1 FILLER_77_1249 ();
 sg13g2_decap_8 FILLER_77_1277 ();
 sg13g2_decap_8 FILLER_77_1284 ();
 sg13g2_decap_4 FILLER_77_1291 ();
 sg13g2_fill_1 FILLER_77_1295 ();
 sg13g2_fill_2 FILLER_77_1337 ();
 sg13g2_fill_2 FILLER_77_1348 ();
 sg13g2_fill_1 FILLER_77_1350 ();
 sg13g2_fill_2 FILLER_77_1418 ();
 sg13g2_fill_2 FILLER_77_1424 ();
 sg13g2_fill_2 FILLER_77_1435 ();
 sg13g2_fill_1 FILLER_77_1437 ();
 sg13g2_fill_1 FILLER_77_1496 ();
 sg13g2_fill_2 FILLER_77_1544 ();
 sg13g2_fill_1 FILLER_77_1546 ();
 sg13g2_fill_2 FILLER_77_1588 ();
 sg13g2_fill_1 FILLER_77_1590 ();
 sg13g2_decap_4 FILLER_77_1622 ();
 sg13g2_decap_4 FILLER_77_1665 ();
 sg13g2_fill_1 FILLER_77_1684 ();
 sg13g2_fill_2 FILLER_77_1731 ();
 sg13g2_fill_1 FILLER_77_1733 ();
 sg13g2_decap_8 FILLER_77_1789 ();
 sg13g2_decap_4 FILLER_77_1796 ();
 sg13g2_fill_1 FILLER_77_1800 ();
 sg13g2_fill_2 FILLER_77_1809 ();
 sg13g2_fill_1 FILLER_77_1811 ();
 sg13g2_fill_1 FILLER_77_1857 ();
 sg13g2_fill_2 FILLER_77_1892 ();
 sg13g2_fill_1 FILLER_77_1894 ();
 sg13g2_decap_4 FILLER_77_1913 ();
 sg13g2_decap_8 FILLER_77_1921 ();
 sg13g2_decap_4 FILLER_77_1928 ();
 sg13g2_fill_2 FILLER_77_1932 ();
 sg13g2_fill_2 FILLER_77_1972 ();
 sg13g2_fill_1 FILLER_77_1974 ();
 sg13g2_fill_1 FILLER_77_1983 ();
 sg13g2_decap_4 FILLER_77_1999 ();
 sg13g2_decap_4 FILLER_77_2008 ();
 sg13g2_decap_8 FILLER_77_2046 ();
 sg13g2_decap_8 FILLER_77_2053 ();
 sg13g2_fill_1 FILLER_77_2060 ();
 sg13g2_fill_1 FILLER_77_2088 ();
 sg13g2_decap_4 FILLER_77_2097 ();
 sg13g2_fill_1 FILLER_77_2101 ();
 sg13g2_fill_2 FILLER_77_2130 ();
 sg13g2_fill_1 FILLER_77_2162 ();
 sg13g2_fill_1 FILLER_77_2184 ();
 sg13g2_fill_2 FILLER_77_2194 ();
 sg13g2_fill_1 FILLER_77_2196 ();
 sg13g2_fill_1 FILLER_77_2215 ();
 sg13g2_fill_1 FILLER_77_2254 ();
 sg13g2_decap_8 FILLER_77_2294 ();
 sg13g2_fill_1 FILLER_77_2314 ();
 sg13g2_fill_2 FILLER_77_2367 ();
 sg13g2_fill_2 FILLER_77_2374 ();
 sg13g2_fill_1 FILLER_77_2391 ();
 sg13g2_decap_8 FILLER_77_2405 ();
 sg13g2_decap_8 FILLER_77_2412 ();
 sg13g2_decap_8 FILLER_77_2419 ();
 sg13g2_decap_4 FILLER_77_2426 ();
 sg13g2_fill_1 FILLER_77_2430 ();
 sg13g2_decap_4 FILLER_77_2475 ();
 sg13g2_fill_2 FILLER_77_2479 ();
 sg13g2_fill_1 FILLER_77_2491 ();
 sg13g2_decap_8 FILLER_77_2513 ();
 sg13g2_decap_8 FILLER_77_2520 ();
 sg13g2_fill_2 FILLER_77_2581 ();
 sg13g2_fill_1 FILLER_77_2583 ();
 sg13g2_decap_8 FILLER_77_2693 ();
 sg13g2_decap_8 FILLER_77_2700 ();
 sg13g2_fill_2 FILLER_77_2707 ();
 sg13g2_fill_2 FILLER_77_2719 ();
 sg13g2_fill_1 FILLER_77_2721 ();
 sg13g2_fill_2 FILLER_77_2753 ();
 sg13g2_decap_8 FILLER_77_2781 ();
 sg13g2_decap_8 FILLER_77_2788 ();
 sg13g2_decap_4 FILLER_77_2795 ();
 sg13g2_fill_2 FILLER_77_2799 ();
 sg13g2_fill_1 FILLER_77_2833 ();
 sg13g2_decap_8 FILLER_77_2847 ();
 sg13g2_decap_8 FILLER_77_2854 ();
 sg13g2_decap_8 FILLER_77_2861 ();
 sg13g2_decap_8 FILLER_77_2868 ();
 sg13g2_decap_4 FILLER_77_2875 ();
 sg13g2_decap_4 FILLER_77_2963 ();
 sg13g2_fill_2 FILLER_77_2967 ();
 sg13g2_decap_8 FILLER_77_2996 ();
 sg13g2_fill_2 FILLER_77_3003 ();
 sg13g2_fill_2 FILLER_77_3009 ();
 sg13g2_fill_1 FILLER_77_3011 ();
 sg13g2_decap_8 FILLER_77_3052 ();
 sg13g2_decap_8 FILLER_77_3059 ();
 sg13g2_decap_8 FILLER_77_3066 ();
 sg13g2_fill_1 FILLER_77_3073 ();
 sg13g2_fill_1 FILLER_77_3078 ();
 sg13g2_fill_1 FILLER_77_3110 ();
 sg13g2_decap_4 FILLER_77_3140 ();
 sg13g2_fill_2 FILLER_77_3144 ();
 sg13g2_decap_4 FILLER_77_3155 ();
 sg13g2_fill_1 FILLER_77_3159 ();
 sg13g2_fill_1 FILLER_77_3187 ();
 sg13g2_fill_2 FILLER_77_3201 ();
 sg13g2_fill_1 FILLER_77_3203 ();
 sg13g2_decap_4 FILLER_77_3217 ();
 sg13g2_fill_2 FILLER_77_3221 ();
 sg13g2_decap_8 FILLER_77_3250 ();
 sg13g2_decap_8 FILLER_77_3257 ();
 sg13g2_decap_4 FILLER_77_3264 ();
 sg13g2_fill_1 FILLER_77_3268 ();
 sg13g2_decap_8 FILLER_77_3301 ();
 sg13g2_decap_8 FILLER_77_3308 ();
 sg13g2_decap_8 FILLER_77_3315 ();
 sg13g2_fill_2 FILLER_77_3322 ();
 sg13g2_fill_1 FILLER_77_3324 ();
 sg13g2_decap_8 FILLER_77_3361 ();
 sg13g2_fill_1 FILLER_77_3368 ();
 sg13g2_decap_8 FILLER_77_3397 ();
 sg13g2_decap_8 FILLER_77_3404 ();
 sg13g2_decap_8 FILLER_77_3411 ();
 sg13g2_decap_8 FILLER_77_3418 ();
 sg13g2_decap_4 FILLER_77_3425 ();
 sg13g2_fill_2 FILLER_77_3429 ();
 sg13g2_decap_8 FILLER_77_3440 ();
 sg13g2_decap_8 FILLER_77_3447 ();
 sg13g2_decap_8 FILLER_77_3454 ();
 sg13g2_decap_8 FILLER_77_3461 ();
 sg13g2_decap_8 FILLER_77_3468 ();
 sg13g2_decap_8 FILLER_77_3475 ();
 sg13g2_decap_8 FILLER_77_3482 ();
 sg13g2_decap_8 FILLER_77_3489 ();
 sg13g2_decap_8 FILLER_77_3496 ();
 sg13g2_decap_8 FILLER_77_3503 ();
 sg13g2_decap_8 FILLER_77_3510 ();
 sg13g2_decap_8 FILLER_77_3517 ();
 sg13g2_decap_8 FILLER_77_3524 ();
 sg13g2_decap_8 FILLER_77_3531 ();
 sg13g2_decap_8 FILLER_77_3538 ();
 sg13g2_decap_8 FILLER_77_3545 ();
 sg13g2_decap_8 FILLER_77_3552 ();
 sg13g2_decap_8 FILLER_77_3559 ();
 sg13g2_decap_8 FILLER_77_3566 ();
 sg13g2_decap_4 FILLER_77_3573 ();
 sg13g2_fill_1 FILLER_77_3577 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_fill_1 FILLER_78_105 ();
 sg13g2_fill_2 FILLER_78_173 ();
 sg13g2_fill_1 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_243 ();
 sg13g2_fill_1 FILLER_78_296 ();
 sg13g2_fill_2 FILLER_78_355 ();
 sg13g2_fill_1 FILLER_78_396 ();
 sg13g2_fill_2 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_445 ();
 sg13g2_fill_1 FILLER_78_452 ();
 sg13g2_fill_2 FILLER_78_512 ();
 sg13g2_fill_1 FILLER_78_514 ();
 sg13g2_decap_8 FILLER_78_561 ();
 sg13g2_decap_8 FILLER_78_614 ();
 sg13g2_fill_2 FILLER_78_621 ();
 sg13g2_fill_1 FILLER_78_623 ();
 sg13g2_fill_2 FILLER_78_681 ();
 sg13g2_fill_1 FILLER_78_683 ();
 sg13g2_fill_2 FILLER_78_752 ();
 sg13g2_fill_2 FILLER_78_781 ();
 sg13g2_fill_1 FILLER_78_783 ();
 sg13g2_fill_1 FILLER_78_820 ();
 sg13g2_fill_1 FILLER_78_831 ();
 sg13g2_decap_8 FILLER_78_860 ();
 sg13g2_decap_4 FILLER_78_867 ();
 sg13g2_fill_2 FILLER_78_898 ();
 sg13g2_fill_2 FILLER_78_940 ();
 sg13g2_fill_2 FILLER_78_978 ();
 sg13g2_fill_1 FILLER_78_980 ();
 sg13g2_decap_8 FILLER_78_1014 ();
 sg13g2_fill_1 FILLER_78_1021 ();
 sg13g2_decap_4 FILLER_78_1073 ();
 sg13g2_fill_2 FILLER_78_1077 ();
 sg13g2_decap_4 FILLER_78_1107 ();
 sg13g2_fill_2 FILLER_78_1138 ();
 sg13g2_decap_8 FILLER_78_1167 ();
 sg13g2_fill_1 FILLER_78_1184 ();
 sg13g2_fill_2 FILLER_78_1221 ();
 sg13g2_fill_2 FILLER_78_1232 ();
 sg13g2_decap_8 FILLER_78_1276 ();
 sg13g2_decap_8 FILLER_78_1283 ();
 sg13g2_decap_8 FILLER_78_1290 ();
 sg13g2_decap_4 FILLER_78_1297 ();
 sg13g2_fill_2 FILLER_78_1331 ();
 sg13g2_fill_2 FILLER_78_1366 ();
 sg13g2_decap_4 FILLER_78_1423 ();
 sg13g2_fill_2 FILLER_78_1489 ();
 sg13g2_fill_1 FILLER_78_1491 ();
 sg13g2_fill_1 FILLER_78_1586 ();
 sg13g2_fill_2 FILLER_78_1615 ();
 sg13g2_fill_1 FILLER_78_1617 ();
 sg13g2_decap_8 FILLER_78_1646 ();
 sg13g2_fill_1 FILLER_78_1653 ();
 sg13g2_decap_4 FILLER_78_1720 ();
 sg13g2_fill_2 FILLER_78_1729 ();
 sg13g2_fill_1 FILLER_78_1731 ();
 sg13g2_decap_8 FILLER_78_1781 ();
 sg13g2_decap_8 FILLER_78_1788 ();
 sg13g2_fill_2 FILLER_78_1858 ();
 sg13g2_fill_1 FILLER_78_1860 ();
 sg13g2_fill_1 FILLER_78_1874 ();
 sg13g2_decap_8 FILLER_78_1913 ();
 sg13g2_fill_1 FILLER_78_1920 ();
 sg13g2_decap_8 FILLER_78_1936 ();
 sg13g2_fill_1 FILLER_78_1943 ();
 sg13g2_fill_2 FILLER_78_1976 ();
 sg13g2_decap_8 FILLER_78_1991 ();
 sg13g2_fill_1 FILLER_78_1998 ();
 sg13g2_fill_2 FILLER_78_2004 ();
 sg13g2_fill_2 FILLER_78_2024 ();
 sg13g2_decap_4 FILLER_78_2047 ();
 sg13g2_fill_1 FILLER_78_2051 ();
 sg13g2_decap_4 FILLER_78_2073 ();
 sg13g2_fill_2 FILLER_78_2077 ();
 sg13g2_decap_8 FILLER_78_2100 ();
 sg13g2_fill_1 FILLER_78_2154 ();
 sg13g2_fill_1 FILLER_78_2202 ();
 sg13g2_fill_1 FILLER_78_2213 ();
 sg13g2_decap_8 FILLER_78_2255 ();
 sg13g2_fill_1 FILLER_78_2262 ();
 sg13g2_decap_8 FILLER_78_2280 ();
 sg13g2_fill_1 FILLER_78_2287 ();
 sg13g2_decap_4 FILLER_78_2396 ();
 sg13g2_decap_8 FILLER_78_2413 ();
 sg13g2_decap_8 FILLER_78_2420 ();
 sg13g2_decap_8 FILLER_78_2427 ();
 sg13g2_decap_8 FILLER_78_2434 ();
 sg13g2_fill_1 FILLER_78_2441 ();
 sg13g2_decap_8 FILLER_78_2469 ();
 sg13g2_decap_8 FILLER_78_2516 ();
 sg13g2_decap_8 FILLER_78_2523 ();
 sg13g2_decap_4 FILLER_78_2567 ();
 sg13g2_fill_2 FILLER_78_2571 ();
 sg13g2_decap_8 FILLER_78_2582 ();
 sg13g2_fill_2 FILLER_78_2589 ();
 sg13g2_fill_1 FILLER_78_2591 ();
 sg13g2_decap_8 FILLER_78_2619 ();
 sg13g2_fill_1 FILLER_78_2626 ();
 sg13g2_fill_1 FILLER_78_2640 ();
 sg13g2_fill_1 FILLER_78_2645 ();
 sg13g2_decap_8 FILLER_78_2682 ();
 sg13g2_decap_8 FILLER_78_2689 ();
 sg13g2_fill_2 FILLER_78_2743 ();
 sg13g2_decap_8 FILLER_78_2776 ();
 sg13g2_fill_2 FILLER_78_2783 ();
 sg13g2_fill_1 FILLER_78_2785 ();
 sg13g2_decap_4 FILLER_78_2867 ();
 sg13g2_fill_1 FILLER_78_2871 ();
 sg13g2_fill_2 FILLER_78_2909 ();
 sg13g2_decap_8 FILLER_78_2992 ();
 sg13g2_fill_1 FILLER_78_2999 ();
 sg13g2_decap_4 FILLER_78_3027 ();
 sg13g2_fill_1 FILLER_78_3031 ();
 sg13g2_decap_8 FILLER_78_3059 ();
 sg13g2_decap_4 FILLER_78_3066 ();
 sg13g2_decap_4 FILLER_78_3080 ();
 sg13g2_decap_8 FILLER_78_3120 ();
 sg13g2_fill_1 FILLER_78_3127 ();
 sg13g2_decap_4 FILLER_78_3159 ();
 sg13g2_fill_2 FILLER_78_3163 ();
 sg13g2_decap_8 FILLER_78_3169 ();
 sg13g2_decap_8 FILLER_78_3176 ();
 sg13g2_decap_8 FILLER_78_3183 ();
 sg13g2_decap_4 FILLER_78_3190 ();
 sg13g2_fill_2 FILLER_78_3194 ();
 sg13g2_decap_8 FILLER_78_3250 ();
 sg13g2_decap_8 FILLER_78_3257 ();
 sg13g2_decap_8 FILLER_78_3264 ();
 sg13g2_decap_8 FILLER_78_3271 ();
 sg13g2_decap_4 FILLER_78_3278 ();
 sg13g2_fill_1 FILLER_78_3282 ();
 sg13g2_decap_8 FILLER_78_3287 ();
 sg13g2_decap_4 FILLER_78_3294 ();
 sg13g2_decap_8 FILLER_78_3311 ();
 sg13g2_decap_8 FILLER_78_3318 ();
 sg13g2_decap_4 FILLER_78_3325 ();
 sg13g2_fill_1 FILLER_78_3329 ();
 sg13g2_decap_8 FILLER_78_3334 ();
 sg13g2_decap_8 FILLER_78_3341 ();
 sg13g2_decap_8 FILLER_78_3348 ();
 sg13g2_decap_8 FILLER_78_3355 ();
 sg13g2_decap_8 FILLER_78_3362 ();
 sg13g2_decap_8 FILLER_78_3369 ();
 sg13g2_fill_2 FILLER_78_3376 ();
 sg13g2_fill_1 FILLER_78_3378 ();
 sg13g2_decap_8 FILLER_78_3383 ();
 sg13g2_decap_8 FILLER_78_3390 ();
 sg13g2_decap_8 FILLER_78_3397 ();
 sg13g2_decap_8 FILLER_78_3404 ();
 sg13g2_decap_8 FILLER_78_3411 ();
 sg13g2_decap_8 FILLER_78_3418 ();
 sg13g2_decap_8 FILLER_78_3425 ();
 sg13g2_decap_8 FILLER_78_3432 ();
 sg13g2_decap_8 FILLER_78_3439 ();
 sg13g2_decap_8 FILLER_78_3446 ();
 sg13g2_decap_8 FILLER_78_3453 ();
 sg13g2_decap_8 FILLER_78_3460 ();
 sg13g2_decap_8 FILLER_78_3467 ();
 sg13g2_decap_8 FILLER_78_3474 ();
 sg13g2_decap_8 FILLER_78_3481 ();
 sg13g2_decap_8 FILLER_78_3488 ();
 sg13g2_decap_8 FILLER_78_3495 ();
 sg13g2_decap_8 FILLER_78_3502 ();
 sg13g2_decap_8 FILLER_78_3509 ();
 sg13g2_decap_8 FILLER_78_3516 ();
 sg13g2_decap_8 FILLER_78_3523 ();
 sg13g2_decap_8 FILLER_78_3530 ();
 sg13g2_decap_8 FILLER_78_3537 ();
 sg13g2_decap_8 FILLER_78_3544 ();
 sg13g2_decap_8 FILLER_78_3551 ();
 sg13g2_decap_8 FILLER_78_3558 ();
 sg13g2_decap_8 FILLER_78_3565 ();
 sg13g2_decap_4 FILLER_78_3572 ();
 sg13g2_fill_2 FILLER_78_3576 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_4 FILLER_79_98 ();
 sg13g2_fill_1 FILLER_79_102 ();
 sg13g2_fill_1 FILLER_79_149 ();
 sg13g2_decap_8 FILLER_79_167 ();
 sg13g2_decap_8 FILLER_79_174 ();
 sg13g2_fill_2 FILLER_79_181 ();
 sg13g2_decap_8 FILLER_79_191 ();
 sg13g2_fill_2 FILLER_79_198 ();
 sg13g2_fill_1 FILLER_79_240 ();
 sg13g2_fill_2 FILLER_79_286 ();
 sg13g2_fill_2 FILLER_79_297 ();
 sg13g2_decap_8 FILLER_79_358 ();
 sg13g2_fill_2 FILLER_79_397 ();
 sg13g2_fill_1 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_436 ();
 sg13g2_fill_1 FILLER_79_443 ();
 sg13g2_decap_4 FILLER_79_573 ();
 sg13g2_fill_2 FILLER_79_618 ();
 sg13g2_fill_2 FILLER_79_691 ();
 sg13g2_fill_2 FILLER_79_713 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_fill_2 FILLER_79_753 ();
 sg13g2_fill_2 FILLER_79_818 ();
 sg13g2_fill_1 FILLER_79_825 ();
 sg13g2_fill_1 FILLER_79_881 ();
 sg13g2_decap_8 FILLER_79_972 ();
 sg13g2_fill_2 FILLER_79_979 ();
 sg13g2_fill_1 FILLER_79_981 ();
 sg13g2_decap_4 FILLER_79_1001 ();
 sg13g2_fill_2 FILLER_79_1005 ();
 sg13g2_fill_1 FILLER_79_1016 ();
 sg13g2_fill_2 FILLER_79_1030 ();
 sg13g2_decap_4 FILLER_79_1072 ();
 sg13g2_fill_2 FILLER_79_1126 ();
 sg13g2_fill_1 FILLER_79_1128 ();
 sg13g2_decap_8 FILLER_79_1132 ();
 sg13g2_decap_4 FILLER_79_1139 ();
 sg13g2_fill_1 FILLER_79_1179 ();
 sg13g2_fill_1 FILLER_79_1226 ();
 sg13g2_fill_2 FILLER_79_1240 ();
 sg13g2_decap_8 FILLER_79_1274 ();
 sg13g2_decap_8 FILLER_79_1281 ();
 sg13g2_decap_8 FILLER_79_1288 ();
 sg13g2_decap_4 FILLER_79_1295 ();
 sg13g2_fill_1 FILLER_79_1299 ();
 sg13g2_fill_1 FILLER_79_1331 ();
 sg13g2_decap_4 FILLER_79_1396 ();
 sg13g2_fill_1 FILLER_79_1400 ();
 sg13g2_decap_4 FILLER_79_1438 ();
 sg13g2_decap_4 FILLER_79_1475 ();
 sg13g2_fill_1 FILLER_79_1479 ();
 sg13g2_decap_4 FILLER_79_1484 ();
 sg13g2_fill_2 FILLER_79_1488 ();
 sg13g2_fill_1 FILLER_79_1536 ();
 sg13g2_fill_1 FILLER_79_1541 ();
 sg13g2_fill_2 FILLER_79_1546 ();
 sg13g2_fill_2 FILLER_79_1598 ();
 sg13g2_fill_1 FILLER_79_1600 ();
 sg13g2_decap_8 FILLER_79_1610 ();
 sg13g2_fill_2 FILLER_79_1617 ();
 sg13g2_fill_1 FILLER_79_1619 ();
 sg13g2_fill_2 FILLER_79_1660 ();
 sg13g2_decap_4 FILLER_79_1726 ();
 sg13g2_fill_1 FILLER_79_1730 ();
 sg13g2_decap_8 FILLER_79_1776 ();
 sg13g2_decap_8 FILLER_79_1783 ();
 sg13g2_decap_8 FILLER_79_1790 ();
 sg13g2_decap_8 FILLER_79_1797 ();
 sg13g2_fill_2 FILLER_79_1804 ();
 sg13g2_fill_1 FILLER_79_1806 ();
 sg13g2_fill_2 FILLER_79_1845 ();
 sg13g2_fill_1 FILLER_79_1847 ();
 sg13g2_fill_2 FILLER_79_1861 ();
 sg13g2_decap_8 FILLER_79_1871 ();
 sg13g2_decap_8 FILLER_79_1878 ();
 sg13g2_fill_1 FILLER_79_1885 ();
 sg13g2_decap_8 FILLER_79_1907 ();
 sg13g2_decap_4 FILLER_79_1940 ();
 sg13g2_fill_2 FILLER_79_1944 ();
 sg13g2_fill_2 FILLER_79_1972 ();
 sg13g2_decap_4 FILLER_79_1978 ();
 sg13g2_decap_8 FILLER_79_1989 ();
 sg13g2_decap_8 FILLER_79_1996 ();
 sg13g2_decap_8 FILLER_79_2003 ();
 sg13g2_fill_1 FILLER_79_2010 ();
 sg13g2_decap_8 FILLER_79_2050 ();
 sg13g2_fill_2 FILLER_79_2057 ();
 sg13g2_fill_1 FILLER_79_2059 ();
 sg13g2_decap_8 FILLER_79_2093 ();
 sg13g2_decap_8 FILLER_79_2100 ();
 sg13g2_decap_8 FILLER_79_2107 ();
 sg13g2_decap_4 FILLER_79_2114 ();
 sg13g2_fill_1 FILLER_79_2118 ();
 sg13g2_decap_8 FILLER_79_2163 ();
 sg13g2_fill_1 FILLER_79_2170 ();
 sg13g2_decap_8 FILLER_79_2176 ();
 sg13g2_decap_8 FILLER_79_2183 ();
 sg13g2_decap_8 FILLER_79_2190 ();
 sg13g2_decap_8 FILLER_79_2197 ();
 sg13g2_fill_2 FILLER_79_2204 ();
 sg13g2_fill_1 FILLER_79_2206 ();
 sg13g2_fill_2 FILLER_79_2224 ();
 sg13g2_fill_1 FILLER_79_2226 ();
 sg13g2_fill_1 FILLER_79_2240 ();
 sg13g2_decap_8 FILLER_79_2250 ();
 sg13g2_decap_8 FILLER_79_2257 ();
 sg13g2_fill_1 FILLER_79_2264 ();
 sg13g2_decap_4 FILLER_79_2285 ();
 sg13g2_fill_2 FILLER_79_2289 ();
 sg13g2_decap_8 FILLER_79_2314 ();
 sg13g2_decap_4 FILLER_79_2321 ();
 sg13g2_fill_2 FILLER_79_2325 ();
 sg13g2_decap_4 FILLER_79_2341 ();
 sg13g2_decap_8 FILLER_79_2349 ();
 sg13g2_fill_2 FILLER_79_2356 ();
 sg13g2_fill_1 FILLER_79_2358 ();
 sg13g2_decap_8 FILLER_79_2385 ();
 sg13g2_fill_2 FILLER_79_2392 ();
 sg13g2_decap_8 FILLER_79_2407 ();
 sg13g2_decap_8 FILLER_79_2414 ();
 sg13g2_decap_8 FILLER_79_2421 ();
 sg13g2_decap_4 FILLER_79_2428 ();
 sg13g2_fill_1 FILLER_79_2432 ();
 sg13g2_decap_4 FILLER_79_2464 ();
 sg13g2_decap_8 FILLER_79_2523 ();
 sg13g2_fill_2 FILLER_79_2530 ();
 sg13g2_fill_1 FILLER_79_2532 ();
 sg13g2_decap_8 FILLER_79_2569 ();
 sg13g2_decap_4 FILLER_79_2576 ();
 sg13g2_fill_2 FILLER_79_2580 ();
 sg13g2_decap_4 FILLER_79_2622 ();
 sg13g2_fill_1 FILLER_79_2626 ();
 sg13g2_decap_4 FILLER_79_2636 ();
 sg13g2_fill_1 FILLER_79_2640 ();
 sg13g2_fill_1 FILLER_79_2672 ();
 sg13g2_decap_8 FILLER_79_2677 ();
 sg13g2_decap_8 FILLER_79_2684 ();
 sg13g2_decap_8 FILLER_79_2691 ();
 sg13g2_fill_1 FILLER_79_2698 ();
 sg13g2_decap_4 FILLER_79_2735 ();
 sg13g2_fill_1 FILLER_79_2739 ();
 sg13g2_decap_8 FILLER_79_2767 ();
 sg13g2_decap_8 FILLER_79_2774 ();
 sg13g2_decap_8 FILLER_79_2781 ();
 sg13g2_fill_2 FILLER_79_2788 ();
 sg13g2_fill_1 FILLER_79_2790 ();
 sg13g2_decap_4 FILLER_79_2795 ();
 sg13g2_fill_2 FILLER_79_2799 ();
 sg13g2_decap_4 FILLER_79_2834 ();
 sg13g2_fill_2 FILLER_79_2838 ();
 sg13g2_decap_8 FILLER_79_2862 ();
 sg13g2_fill_2 FILLER_79_2869 ();
 sg13g2_fill_1 FILLER_79_2871 ();
 sg13g2_decap_8 FILLER_79_2920 ();
 sg13g2_decap_4 FILLER_79_2927 ();
 sg13g2_fill_1 FILLER_79_2931 ();
 sg13g2_fill_2 FILLER_79_2950 ();
 sg13g2_fill_1 FILLER_79_2952 ();
 sg13g2_fill_2 FILLER_79_2991 ();
 sg13g2_decap_4 FILLER_79_3061 ();
 sg13g2_fill_1 FILLER_79_3065 ();
 sg13g2_decap_8 FILLER_79_3120 ();
 sg13g2_decap_4 FILLER_79_3127 ();
 sg13g2_decap_8 FILLER_79_3158 ();
 sg13g2_decap_8 FILLER_79_3165 ();
 sg13g2_decap_8 FILLER_79_3172 ();
 sg13g2_decap_8 FILLER_79_3179 ();
 sg13g2_decap_8 FILLER_79_3186 ();
 sg13g2_decap_8 FILLER_79_3193 ();
 sg13g2_fill_1 FILLER_79_3200 ();
 sg13g2_decap_8 FILLER_79_3205 ();
 sg13g2_fill_2 FILLER_79_3212 ();
 sg13g2_decap_8 FILLER_79_3251 ();
 sg13g2_decap_8 FILLER_79_3258 ();
 sg13g2_decap_8 FILLER_79_3265 ();
 sg13g2_decap_8 FILLER_79_3272 ();
 sg13g2_decap_8 FILLER_79_3279 ();
 sg13g2_decap_8 FILLER_79_3286 ();
 sg13g2_decap_8 FILLER_79_3293 ();
 sg13g2_decap_8 FILLER_79_3300 ();
 sg13g2_decap_8 FILLER_79_3307 ();
 sg13g2_decap_8 FILLER_79_3314 ();
 sg13g2_decap_8 FILLER_79_3321 ();
 sg13g2_decap_8 FILLER_79_3328 ();
 sg13g2_decap_8 FILLER_79_3335 ();
 sg13g2_decap_8 FILLER_79_3342 ();
 sg13g2_decap_8 FILLER_79_3349 ();
 sg13g2_decap_8 FILLER_79_3356 ();
 sg13g2_decap_8 FILLER_79_3363 ();
 sg13g2_decap_8 FILLER_79_3370 ();
 sg13g2_decap_8 FILLER_79_3377 ();
 sg13g2_decap_8 FILLER_79_3384 ();
 sg13g2_decap_8 FILLER_79_3391 ();
 sg13g2_decap_8 FILLER_79_3398 ();
 sg13g2_decap_8 FILLER_79_3405 ();
 sg13g2_decap_8 FILLER_79_3412 ();
 sg13g2_decap_8 FILLER_79_3419 ();
 sg13g2_decap_8 FILLER_79_3426 ();
 sg13g2_decap_8 FILLER_79_3433 ();
 sg13g2_decap_8 FILLER_79_3440 ();
 sg13g2_decap_8 FILLER_79_3447 ();
 sg13g2_decap_8 FILLER_79_3454 ();
 sg13g2_decap_8 FILLER_79_3461 ();
 sg13g2_decap_8 FILLER_79_3468 ();
 sg13g2_decap_8 FILLER_79_3475 ();
 sg13g2_decap_8 FILLER_79_3482 ();
 sg13g2_decap_8 FILLER_79_3489 ();
 sg13g2_decap_8 FILLER_79_3496 ();
 sg13g2_decap_8 FILLER_79_3503 ();
 sg13g2_decap_8 FILLER_79_3510 ();
 sg13g2_decap_8 FILLER_79_3517 ();
 sg13g2_decap_8 FILLER_79_3524 ();
 sg13g2_decap_8 FILLER_79_3531 ();
 sg13g2_decap_8 FILLER_79_3538 ();
 sg13g2_decap_8 FILLER_79_3545 ();
 sg13g2_decap_8 FILLER_79_3552 ();
 sg13g2_decap_8 FILLER_79_3559 ();
 sg13g2_decap_8 FILLER_79_3566 ();
 sg13g2_decap_4 FILLER_79_3573 ();
 sg13g2_fill_1 FILLER_79_3577 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_decap_8 FILLER_80_84 ();
 sg13g2_decap_8 FILLER_80_91 ();
 sg13g2_decap_8 FILLER_80_98 ();
 sg13g2_fill_2 FILLER_80_105 ();
 sg13g2_decap_8 FILLER_80_152 ();
 sg13g2_decap_8 FILLER_80_159 ();
 sg13g2_decap_8 FILLER_80_166 ();
 sg13g2_decap_8 FILLER_80_173 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_4 FILLER_80_194 ();
 sg13g2_fill_1 FILLER_80_198 ();
 sg13g2_decap_8 FILLER_80_212 ();
 sg13g2_decap_8 FILLER_80_219 ();
 sg13g2_decap_4 FILLER_80_226 ();
 sg13g2_fill_2 FILLER_80_230 ();
 sg13g2_fill_2 FILLER_80_320 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_fill_1 FILLER_80_396 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_425 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_decap_4 FILLER_80_451 ();
 sg13g2_fill_2 FILLER_80_504 ();
 sg13g2_fill_1 FILLER_80_506 ();
 sg13g2_decap_4 FILLER_80_622 ();
 sg13g2_fill_1 FILLER_80_626 ();
 sg13g2_fill_1 FILLER_80_653 ();
 sg13g2_decap_4 FILLER_80_672 ();
 sg13g2_fill_2 FILLER_80_690 ();
 sg13g2_fill_1 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_751 ();
 sg13g2_decap_8 FILLER_80_758 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_fill_2 FILLER_80_823 ();
 sg13g2_fill_1 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_865 ();
 sg13g2_decap_8 FILLER_80_872 ();
 sg13g2_decap_8 FILLER_80_879 ();
 sg13g2_decap_4 FILLER_80_886 ();
 sg13g2_fill_2 FILLER_80_890 ();
 sg13g2_fill_2 FILLER_80_913 ();
 sg13g2_fill_2 FILLER_80_943 ();
 sg13g2_fill_1 FILLER_80_945 ();
 sg13g2_fill_2 FILLER_80_950 ();
 sg13g2_fill_1 FILLER_80_952 ();
 sg13g2_decap_8 FILLER_80_962 ();
 sg13g2_decap_8 FILLER_80_969 ();
 sg13g2_decap_8 FILLER_80_976 ();
 sg13g2_decap_8 FILLER_80_983 ();
 sg13g2_decap_8 FILLER_80_990 ();
 sg13g2_decap_8 FILLER_80_997 ();
 sg13g2_decap_8 FILLER_80_1004 ();
 sg13g2_decap_8 FILLER_80_1011 ();
 sg13g2_fill_2 FILLER_80_1018 ();
 sg13g2_fill_1 FILLER_80_1020 ();
 sg13g2_decap_8 FILLER_80_1057 ();
 sg13g2_decap_8 FILLER_80_1064 ();
 sg13g2_decap_8 FILLER_80_1080 ();
 sg13g2_decap_4 FILLER_80_1087 ();
 sg13g2_fill_1 FILLER_80_1091 ();
 sg13g2_decap_8 FILLER_80_1119 ();
 sg13g2_decap_8 FILLER_80_1126 ();
 sg13g2_decap_8 FILLER_80_1133 ();
 sg13g2_decap_8 FILLER_80_1140 ();
 sg13g2_decap_8 FILLER_80_1147 ();
 sg13g2_decap_8 FILLER_80_1154 ();
 sg13g2_decap_8 FILLER_80_1161 ();
 sg13g2_decap_8 FILLER_80_1168 ();
 sg13g2_decap_8 FILLER_80_1175 ();
 sg13g2_decap_8 FILLER_80_1191 ();
 sg13g2_decap_8 FILLER_80_1198 ();
 sg13g2_fill_2 FILLER_80_1205 ();
 sg13g2_fill_1 FILLER_80_1207 ();
 sg13g2_fill_2 FILLER_80_1256 ();
 sg13g2_fill_1 FILLER_80_1258 ();
 sg13g2_decap_8 FILLER_80_1273 ();
 sg13g2_decap_8 FILLER_80_1280 ();
 sg13g2_decap_8 FILLER_80_1287 ();
 sg13g2_decap_8 FILLER_80_1294 ();
 sg13g2_decap_4 FILLER_80_1301 ();
 sg13g2_fill_1 FILLER_80_1305 ();
 sg13g2_fill_1 FILLER_80_1333 ();
 sg13g2_fill_2 FILLER_80_1338 ();
 sg13g2_fill_1 FILLER_80_1340 ();
 sg13g2_fill_2 FILLER_80_1358 ();
 sg13g2_decap_4 FILLER_80_1368 ();
 sg13g2_fill_1 FILLER_80_1372 ();
 sg13g2_decap_8 FILLER_80_1382 ();
 sg13g2_decap_8 FILLER_80_1389 ();
 sg13g2_decap_8 FILLER_80_1396 ();
 sg13g2_decap_8 FILLER_80_1403 ();
 sg13g2_decap_8 FILLER_80_1410 ();
 sg13g2_decap_8 FILLER_80_1417 ();
 sg13g2_decap_8 FILLER_80_1424 ();
 sg13g2_decap_8 FILLER_80_1431 ();
 sg13g2_decap_4 FILLER_80_1438 ();
 sg13g2_decap_8 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1480 ();
 sg13g2_decap_8 FILLER_80_1487 ();
 sg13g2_decap_4 FILLER_80_1494 ();
 sg13g2_decap_8 FILLER_80_1533 ();
 sg13g2_decap_4 FILLER_80_1540 ();
 sg13g2_fill_2 FILLER_80_1544 ();
 sg13g2_fill_2 FILLER_80_1550 ();
 sg13g2_fill_2 FILLER_80_1557 ();
 sg13g2_fill_1 FILLER_80_1559 ();
 sg13g2_decap_8 FILLER_80_1582 ();
 sg13g2_decap_8 FILLER_80_1589 ();
 sg13g2_decap_4 FILLER_80_1596 ();
 sg13g2_decap_8 FILLER_80_1609 ();
 sg13g2_decap_8 FILLER_80_1616 ();
 sg13g2_decap_8 FILLER_80_1623 ();
 sg13g2_decap_8 FILLER_80_1630 ();
 sg13g2_fill_2 FILLER_80_1637 ();
 sg13g2_decap_8 FILLER_80_1648 ();
 sg13g2_decap_8 FILLER_80_1655 ();
 sg13g2_decap_8 FILLER_80_1662 ();
 sg13g2_decap_8 FILLER_80_1669 ();
 sg13g2_decap_8 FILLER_80_1676 ();
 sg13g2_decap_8 FILLER_80_1683 ();
 sg13g2_fill_2 FILLER_80_1690 ();
 sg13g2_fill_1 FILLER_80_1706 ();
 sg13g2_decap_8 FILLER_80_1716 ();
 sg13g2_decap_8 FILLER_80_1723 ();
 sg13g2_decap_8 FILLER_80_1730 ();
 sg13g2_decap_8 FILLER_80_1737 ();
 sg13g2_decap_8 FILLER_80_1744 ();
 sg13g2_decap_8 FILLER_80_1751 ();
 sg13g2_decap_8 FILLER_80_1758 ();
 sg13g2_decap_8 FILLER_80_1765 ();
 sg13g2_decap_8 FILLER_80_1772 ();
 sg13g2_decap_8 FILLER_80_1779 ();
 sg13g2_decap_8 FILLER_80_1786 ();
 sg13g2_decap_8 FILLER_80_1793 ();
 sg13g2_decap_8 FILLER_80_1800 ();
 sg13g2_decap_8 FILLER_80_1807 ();
 sg13g2_decap_4 FILLER_80_1814 ();
 sg13g2_fill_2 FILLER_80_1818 ();
 sg13g2_fill_2 FILLER_80_1834 ();
 sg13g2_decap_8 FILLER_80_1844 ();
 sg13g2_fill_2 FILLER_80_1851 ();
 sg13g2_decap_8 FILLER_80_1857 ();
 sg13g2_decap_8 FILLER_80_1864 ();
 sg13g2_decap_8 FILLER_80_1871 ();
 sg13g2_decap_8 FILLER_80_1878 ();
 sg13g2_decap_8 FILLER_80_1885 ();
 sg13g2_fill_1 FILLER_80_1892 ();
 sg13g2_decap_8 FILLER_80_1901 ();
 sg13g2_decap_8 FILLER_80_1908 ();
 sg13g2_decap_8 FILLER_80_1915 ();
 sg13g2_decap_8 FILLER_80_1922 ();
 sg13g2_decap_8 FILLER_80_1929 ();
 sg13g2_decap_8 FILLER_80_1936 ();
 sg13g2_decap_8 FILLER_80_1943 ();
 sg13g2_decap_8 FILLER_80_1950 ();
 sg13g2_decap_8 FILLER_80_1957 ();
 sg13g2_decap_8 FILLER_80_1964 ();
 sg13g2_decap_8 FILLER_80_1971 ();
 sg13g2_decap_8 FILLER_80_1978 ();
 sg13g2_decap_8 FILLER_80_1985 ();
 sg13g2_decap_8 FILLER_80_1992 ();
 sg13g2_decap_8 FILLER_80_1999 ();
 sg13g2_decap_8 FILLER_80_2006 ();
 sg13g2_fill_2 FILLER_80_2013 ();
 sg13g2_decap_8 FILLER_80_2020 ();
 sg13g2_decap_8 FILLER_80_2027 ();
 sg13g2_decap_8 FILLER_80_2034 ();
 sg13g2_decap_8 FILLER_80_2041 ();
 sg13g2_decap_8 FILLER_80_2048 ();
 sg13g2_decap_8 FILLER_80_2055 ();
 sg13g2_fill_1 FILLER_80_2062 ();
 sg13g2_decap_8 FILLER_80_2073 ();
 sg13g2_decap_8 FILLER_80_2080 ();
 sg13g2_decap_8 FILLER_80_2087 ();
 sg13g2_decap_8 FILLER_80_2094 ();
 sg13g2_decap_8 FILLER_80_2101 ();
 sg13g2_decap_8 FILLER_80_2108 ();
 sg13g2_decap_8 FILLER_80_2115 ();
 sg13g2_decap_8 FILLER_80_2122 ();
 sg13g2_decap_8 FILLER_80_2129 ();
 sg13g2_decap_8 FILLER_80_2136 ();
 sg13g2_decap_4 FILLER_80_2147 ();
 sg13g2_fill_2 FILLER_80_2151 ();
 sg13g2_decap_8 FILLER_80_2166 ();
 sg13g2_decap_8 FILLER_80_2173 ();
 sg13g2_decap_8 FILLER_80_2180 ();
 sg13g2_decap_8 FILLER_80_2187 ();
 sg13g2_decap_8 FILLER_80_2194 ();
 sg13g2_decap_8 FILLER_80_2201 ();
 sg13g2_decap_8 FILLER_80_2208 ();
 sg13g2_decap_8 FILLER_80_2215 ();
 sg13g2_decap_4 FILLER_80_2222 ();
 sg13g2_fill_2 FILLER_80_2226 ();
 sg13g2_fill_2 FILLER_80_2233 ();
 sg13g2_fill_1 FILLER_80_2235 ();
 sg13g2_decap_8 FILLER_80_2239 ();
 sg13g2_decap_8 FILLER_80_2246 ();
 sg13g2_decap_8 FILLER_80_2253 ();
 sg13g2_decap_8 FILLER_80_2260 ();
 sg13g2_decap_8 FILLER_80_2267 ();
 sg13g2_decap_8 FILLER_80_2274 ();
 sg13g2_decap_8 FILLER_80_2281 ();
 sg13g2_decap_8 FILLER_80_2288 ();
 sg13g2_decap_8 FILLER_80_2305 ();
 sg13g2_decap_8 FILLER_80_2312 ();
 sg13g2_decap_8 FILLER_80_2319 ();
 sg13g2_decap_8 FILLER_80_2326 ();
 sg13g2_decap_8 FILLER_80_2333 ();
 sg13g2_decap_8 FILLER_80_2340 ();
 sg13g2_decap_8 FILLER_80_2347 ();
 sg13g2_decap_4 FILLER_80_2354 ();
 sg13g2_fill_2 FILLER_80_2358 ();
 sg13g2_decap_8 FILLER_80_2373 ();
 sg13g2_decap_8 FILLER_80_2380 ();
 sg13g2_decap_8 FILLER_80_2387 ();
 sg13g2_decap_8 FILLER_80_2394 ();
 sg13g2_decap_8 FILLER_80_2401 ();
 sg13g2_decap_8 FILLER_80_2408 ();
 sg13g2_decap_8 FILLER_80_2415 ();
 sg13g2_decap_8 FILLER_80_2422 ();
 sg13g2_decap_8 FILLER_80_2429 ();
 sg13g2_decap_8 FILLER_80_2436 ();
 sg13g2_fill_1 FILLER_80_2447 ();
 sg13g2_decap_8 FILLER_80_2467 ();
 sg13g2_decap_8 FILLER_80_2474 ();
 sg13g2_fill_2 FILLER_80_2481 ();
 sg13g2_fill_2 FILLER_80_2487 ();
 sg13g2_fill_1 FILLER_80_2489 ();
 sg13g2_decap_8 FILLER_80_2513 ();
 sg13g2_decap_8 FILLER_80_2520 ();
 sg13g2_decap_8 FILLER_80_2527 ();
 sg13g2_decap_4 FILLER_80_2534 ();
 sg13g2_fill_2 FILLER_80_2542 ();
 sg13g2_fill_1 FILLER_80_2544 ();
 sg13g2_fill_1 FILLER_80_2559 ();
 sg13g2_decap_8 FILLER_80_2569 ();
 sg13g2_decap_8 FILLER_80_2576 ();
 sg13g2_decap_8 FILLER_80_2583 ();
 sg13g2_fill_1 FILLER_80_2590 ();
 sg13g2_fill_2 FILLER_80_2595 ();
 sg13g2_fill_1 FILLER_80_2597 ();
 sg13g2_fill_2 FILLER_80_2608 ();
 sg13g2_fill_1 FILLER_80_2610 ();
 sg13g2_decap_8 FILLER_80_2620 ();
 sg13g2_decap_8 FILLER_80_2627 ();
 sg13g2_decap_4 FILLER_80_2634 ();
 sg13g2_fill_2 FILLER_80_2638 ();
 sg13g2_fill_1 FILLER_80_2654 ();
 sg13g2_decap_8 FILLER_80_2673 ();
 sg13g2_decap_8 FILLER_80_2680 ();
 sg13g2_decap_8 FILLER_80_2687 ();
 sg13g2_decap_8 FILLER_80_2694 ();
 sg13g2_fill_2 FILLER_80_2701 ();
 sg13g2_fill_1 FILLER_80_2703 ();
 sg13g2_fill_1 FILLER_80_2708 ();
 sg13g2_decap_8 FILLER_80_2722 ();
 sg13g2_decap_8 FILLER_80_2729 ();
 sg13g2_decap_8 FILLER_80_2736 ();
 sg13g2_decap_8 FILLER_80_2743 ();
 sg13g2_fill_2 FILLER_80_2750 ();
 sg13g2_decap_8 FILLER_80_2765 ();
 sg13g2_decap_8 FILLER_80_2772 ();
 sg13g2_decap_8 FILLER_80_2779 ();
 sg13g2_decap_8 FILLER_80_2786 ();
 sg13g2_decap_8 FILLER_80_2793 ();
 sg13g2_decap_8 FILLER_80_2800 ();
 sg13g2_fill_2 FILLER_80_2807 ();
 sg13g2_fill_1 FILLER_80_2809 ();
 sg13g2_decap_4 FILLER_80_2814 ();
 sg13g2_fill_1 FILLER_80_2818 ();
 sg13g2_fill_1 FILLER_80_2829 ();
 sg13g2_decap_8 FILLER_80_2862 ();
 sg13g2_decap_8 FILLER_80_2869 ();
 sg13g2_fill_2 FILLER_80_2890 ();
 sg13g2_fill_1 FILLER_80_2892 ();
 sg13g2_fill_2 FILLER_80_2903 ();
 sg13g2_decap_8 FILLER_80_2923 ();
 sg13g2_decap_8 FILLER_80_2930 ();
 sg13g2_decap_4 FILLER_80_2937 ();
 sg13g2_fill_1 FILLER_80_2941 ();
 sg13g2_fill_2 FILLER_80_2952 ();
 sg13g2_fill_1 FILLER_80_2954 ();
 sg13g2_decap_4 FILLER_80_2964 ();
 sg13g2_fill_1 FILLER_80_2968 ();
 sg13g2_decap_8 FILLER_80_2986 ();
 sg13g2_decap_8 FILLER_80_2993 ();
 sg13g2_fill_2 FILLER_80_3000 ();
 sg13g2_fill_1 FILLER_80_3002 ();
 sg13g2_decap_8 FILLER_80_3053 ();
 sg13g2_decap_8 FILLER_80_3060 ();
 sg13g2_decap_4 FILLER_80_3067 ();
 sg13g2_fill_1 FILLER_80_3075 ();
 sg13g2_fill_1 FILLER_80_3103 ();
 sg13g2_decap_8 FILLER_80_3113 ();
 sg13g2_decap_8 FILLER_80_3120 ();
 sg13g2_decap_8 FILLER_80_3127 ();
 sg13g2_fill_2 FILLER_80_3134 ();
 sg13g2_fill_1 FILLER_80_3140 ();
 sg13g2_decap_8 FILLER_80_3150 ();
 sg13g2_decap_8 FILLER_80_3157 ();
 sg13g2_decap_8 FILLER_80_3164 ();
 sg13g2_decap_8 FILLER_80_3171 ();
 sg13g2_decap_8 FILLER_80_3178 ();
 sg13g2_decap_8 FILLER_80_3185 ();
 sg13g2_decap_8 FILLER_80_3192 ();
 sg13g2_decap_8 FILLER_80_3199 ();
 sg13g2_decap_4 FILLER_80_3206 ();
 sg13g2_fill_1 FILLER_80_3210 ();
 sg13g2_fill_2 FILLER_80_3225 ();
 sg13g2_fill_2 FILLER_80_3231 ();
 sg13g2_fill_1 FILLER_80_3233 ();
 sg13g2_decap_8 FILLER_80_3256 ();
 sg13g2_decap_8 FILLER_80_3263 ();
 sg13g2_decap_8 FILLER_80_3270 ();
 sg13g2_decap_8 FILLER_80_3277 ();
 sg13g2_decap_8 FILLER_80_3284 ();
 sg13g2_decap_8 FILLER_80_3291 ();
 sg13g2_decap_8 FILLER_80_3298 ();
 sg13g2_decap_8 FILLER_80_3305 ();
 sg13g2_decap_8 FILLER_80_3312 ();
 sg13g2_decap_8 FILLER_80_3319 ();
 sg13g2_decap_8 FILLER_80_3326 ();
 sg13g2_decap_8 FILLER_80_3333 ();
 sg13g2_decap_8 FILLER_80_3340 ();
 sg13g2_decap_8 FILLER_80_3347 ();
 sg13g2_decap_8 FILLER_80_3354 ();
 sg13g2_decap_8 FILLER_80_3361 ();
 sg13g2_decap_8 FILLER_80_3368 ();
 sg13g2_decap_8 FILLER_80_3375 ();
 sg13g2_decap_8 FILLER_80_3382 ();
 sg13g2_decap_8 FILLER_80_3389 ();
 sg13g2_decap_8 FILLER_80_3396 ();
 sg13g2_decap_8 FILLER_80_3403 ();
 sg13g2_decap_8 FILLER_80_3410 ();
 sg13g2_decap_8 FILLER_80_3417 ();
 sg13g2_decap_8 FILLER_80_3424 ();
 sg13g2_decap_8 FILLER_80_3431 ();
 sg13g2_decap_8 FILLER_80_3438 ();
 sg13g2_decap_8 FILLER_80_3445 ();
 sg13g2_decap_8 FILLER_80_3452 ();
 sg13g2_decap_8 FILLER_80_3459 ();
 sg13g2_decap_8 FILLER_80_3466 ();
 sg13g2_decap_8 FILLER_80_3473 ();
 sg13g2_decap_8 FILLER_80_3480 ();
 sg13g2_decap_8 FILLER_80_3487 ();
 sg13g2_decap_8 FILLER_80_3494 ();
 sg13g2_decap_8 FILLER_80_3501 ();
 sg13g2_decap_8 FILLER_80_3508 ();
 sg13g2_decap_8 FILLER_80_3515 ();
 sg13g2_decap_8 FILLER_80_3522 ();
 sg13g2_decap_8 FILLER_80_3529 ();
 sg13g2_decap_8 FILLER_80_3536 ();
 sg13g2_decap_8 FILLER_80_3543 ();
 sg13g2_decap_8 FILLER_80_3550 ();
 sg13g2_decap_8 FILLER_80_3557 ();
 sg13g2_decap_8 FILLER_80_3564 ();
 sg13g2_decap_8 FILLER_80_3571 ();
endmodule
