module tt_um_flummer_ltc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire \ltc.bit_clk ;
 wire \ltc.bit_counter[0] ;
 wire \ltc.bit_counter[10] ;
 wire \ltc.bit_counter[11] ;
 wire \ltc.bit_counter[1] ;
 wire \ltc.bit_counter[2] ;
 wire \ltc.bit_counter[3] ;
 wire \ltc.bit_counter[4] ;
 wire \ltc.bit_counter[5] ;
 wire \ltc.bit_counter[6] ;
 wire \ltc.bit_counter[7] ;
 wire \ltc.bit_counter[8] ;
 wire \ltc.bit_counter[9] ;
 wire \ltc.frm_counter[0] ;
 wire \ltc.frm_counter[10] ;
 wire \ltc.frm_counter[11] ;
 wire \ltc.frm_counter[12] ;
 wire \ltc.frm_counter[13] ;
 wire \ltc.frm_counter[14] ;
 wire \ltc.frm_counter[15] ;
 wire \ltc.frm_counter[16] ;
 wire \ltc.frm_counter[17] ;
 wire \ltc.frm_counter[18] ;
 wire \ltc.frm_counter[19] ;
 wire \ltc.frm_counter[1] ;
 wire \ltc.frm_counter[20] ;
 wire \ltc.frm_counter[21] ;
 wire \ltc.frm_counter[22] ;
 wire \ltc.frm_counter[23] ;
 wire \ltc.frm_counter[2] ;
 wire \ltc.frm_counter[3] ;
 wire \ltc.frm_counter[4] ;
 wire \ltc.frm_counter[5] ;
 wire \ltc.frm_counter[6] ;
 wire \ltc.frm_counter[7] ;
 wire \ltc.frm_counter[8] ;
 wire \ltc.frm_counter[9] ;
 wire \ltc.frm_d[0] ;
 wire \ltc.frm_d[1] ;
 wire \ltc.frm_u[0] ;
 wire \ltc.frm_u[1] ;
 wire \ltc.frm_u[2] ;
 wire \ltc.frm_u[3] ;
 wire \ltc.hrs_d[0] ;
 wire \ltc.hrs_d[1] ;
 wire \ltc.hrs_u[0] ;
 wire \ltc.hrs_u[1] ;
 wire \ltc.hrs_u[2] ;
 wire \ltc.hrs_u[3] ;
 wire \ltc.min_d[0] ;
 wire \ltc.min_d[1] ;
 wire \ltc.min_d[2] ;
 wire \ltc.min_u[0] ;
 wire \ltc.min_u[1] ;
 wire \ltc.min_u[2] ;
 wire \ltc.min_u[3] ;
 wire \ltc.output_buffer[0] ;
 wire \ltc.output_buffer[10] ;
 wire \ltc.output_buffer[11] ;
 wire \ltc.output_buffer[12] ;
 wire \ltc.output_buffer[13] ;
 wire \ltc.output_buffer[14] ;
 wire \ltc.output_buffer[15] ;
 wire \ltc.output_buffer[16] ;
 wire \ltc.output_buffer[17] ;
 wire \ltc.output_buffer[18] ;
 wire \ltc.output_buffer[19] ;
 wire \ltc.output_buffer[1] ;
 wire \ltc.output_buffer[20] ;
 wire \ltc.output_buffer[21] ;
 wire \ltc.output_buffer[22] ;
 wire \ltc.output_buffer[23] ;
 wire \ltc.output_buffer[24] ;
 wire \ltc.output_buffer[25] ;
 wire \ltc.output_buffer[26] ;
 wire \ltc.output_buffer[27] ;
 wire \ltc.output_buffer[28] ;
 wire \ltc.output_buffer[29] ;
 wire \ltc.output_buffer[2] ;
 wire \ltc.output_buffer[30] ;
 wire \ltc.output_buffer[31] ;
 wire \ltc.output_buffer[32] ;
 wire \ltc.output_buffer[33] ;
 wire \ltc.output_buffer[34] ;
 wire \ltc.output_buffer[35] ;
 wire \ltc.output_buffer[36] ;
 wire \ltc.output_buffer[37] ;
 wire \ltc.output_buffer[38] ;
 wire \ltc.output_buffer[39] ;
 wire \ltc.output_buffer[3] ;
 wire \ltc.output_buffer[40] ;
 wire \ltc.output_buffer[41] ;
 wire \ltc.output_buffer[42] ;
 wire \ltc.output_buffer[43] ;
 wire \ltc.output_buffer[44] ;
 wire \ltc.output_buffer[45] ;
 wire \ltc.output_buffer[46] ;
 wire \ltc.output_buffer[47] ;
 wire \ltc.output_buffer[48] ;
 wire \ltc.output_buffer[49] ;
 wire \ltc.output_buffer[4] ;
 wire \ltc.output_buffer[50] ;
 wire \ltc.output_buffer[51] ;
 wire \ltc.output_buffer[52] ;
 wire \ltc.output_buffer[53] ;
 wire \ltc.output_buffer[54] ;
 wire \ltc.output_buffer[55] ;
 wire \ltc.output_buffer[56] ;
 wire \ltc.output_buffer[57] ;
 wire \ltc.output_buffer[58] ;
 wire \ltc.output_buffer[59] ;
 wire \ltc.output_buffer[5] ;
 wire \ltc.output_buffer[60] ;
 wire \ltc.output_buffer[61] ;
 wire \ltc.output_buffer[62] ;
 wire \ltc.output_buffer[63] ;
 wire \ltc.output_buffer[64] ;
 wire \ltc.output_buffer[65] ;
 wire \ltc.output_buffer[66] ;
 wire \ltc.output_buffer[67] ;
 wire \ltc.output_buffer[68] ;
 wire \ltc.output_buffer[69] ;
 wire \ltc.output_buffer[6] ;
 wire \ltc.output_buffer[70] ;
 wire \ltc.output_buffer[71] ;
 wire \ltc.output_buffer[72] ;
 wire \ltc.output_buffer[73] ;
 wire \ltc.output_buffer[74] ;
 wire \ltc.output_buffer[75] ;
 wire \ltc.output_buffer[76] ;
 wire \ltc.output_buffer[77] ;
 wire \ltc.output_buffer[78] ;
 wire \ltc.output_buffer[79] ;
 wire \ltc.output_buffer[7] ;
 wire \ltc.output_buffer[8] ;
 wire \ltc.output_buffer[9] ;
 wire \ltc.sec_d[0] ;
 wire \ltc.sec_d[1] ;
 wire \ltc.sec_d[2] ;
 wire \ltc.sec_u[0] ;
 wire \ltc.sec_u[1] ;
 wire \ltc.sec_u[2] ;
 wire \ltc.sec_u[3] ;
 wire \ltc.timecode ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;

 sg13g2_inv_1 _0714_ (.Y(_0144_),
    .A(net444));
 sg13g2_inv_1 _0715_ (.Y(_0145_),
    .A(net390));
 sg13g2_inv_1 _0716_ (.Y(_0146_),
    .A(net294));
 sg13g2_inv_1 _0717_ (.Y(_0147_),
    .A(net467));
 sg13g2_inv_1 _0718_ (.Y(_0148_),
    .A(net463));
 sg13g2_inv_1 _0719_ (.Y(_0149_),
    .A(net424));
 sg13g2_inv_1 _0720_ (.Y(_0150_),
    .A(net330));
 sg13g2_inv_1 _0721_ (.Y(_0151_),
    .A(net439));
 sg13g2_inv_1 _0722_ (.Y(_0152_),
    .A(\ltc.frm_counter[12] ));
 sg13g2_inv_1 _0723_ (.Y(_0153_),
    .A(net473));
 sg13g2_inv_1 _0724_ (.Y(_0154_),
    .A(\ltc.bit_counter[6] ));
 sg13g2_inv_1 _0725_ (.Y(_0155_),
    .A(net175));
 sg13g2_inv_1 _0726_ (.Y(_0156_),
    .A(net238));
 sg13g2_inv_1 _0727_ (.Y(_0157_),
    .A(net253));
 sg13g2_inv_1 _0728_ (.Y(_0158_),
    .A(\ltc.output_buffer[3] ));
 sg13g2_inv_1 _0729_ (.Y(_0159_),
    .A(net256));
 sg13g2_inv_1 _0730_ (.Y(_0160_),
    .A(net240));
 sg13g2_inv_1 _0731_ (.Y(_0161_),
    .A(net233));
 sg13g2_inv_1 _0732_ (.Y(_0162_),
    .A(net251));
 sg13g2_inv_1 _0733_ (.Y(_0163_),
    .A(net249));
 sg13g2_inv_1 _0734_ (.Y(_0164_),
    .A(net247));
 sg13g2_inv_1 _0735_ (.Y(_0165_),
    .A(net252));
 sg13g2_inv_1 _0736_ (.Y(_0166_),
    .A(net243));
 sg13g2_inv_1 _0737_ (.Y(_0167_),
    .A(net259));
 sg13g2_inv_1 _0738_ (.Y(_0168_),
    .A(net245));
 sg13g2_nand2_1 _0739_ (.Y(_0169_),
    .A(net7),
    .B(net8));
 sg13g2_nand4_1 _0740_ (.B(net5),
    .C(net2),
    .A(net6),
    .Y(_0170_),
    .D(net1));
 sg13g2_nor2_1 _0741_ (.A(_0169_),
    .B(_0170_),
    .Y(uo_out[0]));
 sg13g2_nor2_1 _0742_ (.A(net383),
    .B(net227),
    .Y(_0171_));
 sg13g2_nor3_1 _0743_ (.A(\ltc.bit_counter[2] ),
    .B(\ltc.bit_counter[10] ),
    .C(\ltc.bit_counter[11] ),
    .Y(_0172_));
 sg13g2_nor2_1 _0744_ (.A(\ltc.bit_counter[5] ),
    .B(\ltc.bit_counter[4] ),
    .Y(_0173_));
 sg13g2_nor2_1 _0745_ (.A(\ltc.bit_counter[8] ),
    .B(\ltc.bit_counter[9] ),
    .Y(_0174_));
 sg13g2_nor4_1 _0746_ (.A(\ltc.bit_counter[1] ),
    .B(net227),
    .C(\ltc.bit_counter[6] ),
    .D(\ltc.bit_counter[7] ),
    .Y(_0175_));
 sg13g2_nor3_1 _0747_ (.A(\ltc.bit_counter[5] ),
    .B(\ltc.bit_counter[4] ),
    .C(\ltc.bit_counter[3] ),
    .Y(_0176_));
 sg13g2_nand4_1 _0748_ (.B(_0174_),
    .C(_0175_),
    .A(_0172_),
    .Y(_0177_),
    .D(_0176_));
 sg13g2_nor2_2 _0749_ (.A(net231),
    .B(_0177_),
    .Y(_0178_));
 sg13g2_nor2_2 _0750_ (.A(net163),
    .B(net152),
    .Y(_0179_));
 sg13g2_nor3_1 _0751_ (.A(\ltc.frm_counter[16] ),
    .B(\ltc.frm_counter[17] ),
    .C(\ltc.frm_counter[18] ),
    .Y(_0180_));
 sg13g2_nor4_1 _0752_ (.A(\ltc.frm_counter[10] ),
    .B(\ltc.frm_counter[11] ),
    .C(\ltc.frm_counter[12] ),
    .D(\ltc.frm_counter[13] ),
    .Y(_0181_));
 sg13g2_nor4_1 _0753_ (.A(\ltc.frm_counter[3] ),
    .B(\ltc.frm_counter[2] ),
    .C(\ltc.frm_counter[6] ),
    .D(\ltc.frm_counter[7] ),
    .Y(_0182_));
 sg13g2_nand3_1 _0754_ (.B(_0181_),
    .C(_0182_),
    .A(_0180_),
    .Y(_0183_));
 sg13g2_nor2_1 _0755_ (.A(\ltc.frm_counter[19] ),
    .B(\ltc.frm_counter[20] ),
    .Y(_0184_));
 sg13g2_nor3_1 _0756_ (.A(\ltc.frm_counter[21] ),
    .B(\ltc.frm_counter[22] ),
    .C(\ltc.frm_counter[23] ),
    .Y(_0185_));
 sg13g2_nand2_1 _0757_ (.Y(_0186_),
    .A(_0184_),
    .B(_0185_));
 sg13g2_nor2_1 _0758_ (.A(\ltc.frm_counter[14] ),
    .B(\ltc.frm_counter[15] ),
    .Y(_0187_));
 sg13g2_nor2_1 _0759_ (.A(net469),
    .B(net466),
    .Y(_0188_));
 sg13g2_nor2_1 _0760_ (.A(\ltc.frm_counter[5] ),
    .B(\ltc.frm_counter[4] ),
    .Y(_0189_));
 sg13g2_nand3_1 _0761_ (.B(_0188_),
    .C(_0189_),
    .A(_0187_),
    .Y(_0190_));
 sg13g2_nor3_1 _0762_ (.A(_0183_),
    .B(_0186_),
    .C(_0190_),
    .Y(_0191_));
 sg13g2_nor2b_1 _0763_ (.A(net428),
    .B_N(net228),
    .Y(_0192_));
 sg13g2_and2_1 _0764_ (.A(_0191_),
    .B(_0192_),
    .X(_0193_));
 sg13g2_nand2_1 _0765_ (.Y(_0194_),
    .A(_0191_),
    .B(_0192_));
 sg13g2_o21ai_1 _0766_ (.B1(net146),
    .Y(_0195_),
    .A1(net242),
    .A2(net141));
 sg13g2_inv_1 _0767_ (.Y(_0000_),
    .A(_0195_));
 sg13g2_nor2_1 _0768_ (.A(net151),
    .B(net138),
    .Y(_0196_));
 sg13g2_a22oi_1 _0769_ (.Y(_0197_),
    .B1(net129),
    .B2(net238),
    .A2(net157),
    .A1(net242));
 sg13g2_nor2_1 _0770_ (.A(net164),
    .B(_0197_),
    .Y(_0001_));
 sg13g2_a221oi_1 _0771_ (.B2(_0157_),
    .C1(net164),
    .B1(net129),
    .A1(_0156_),
    .Y(_0002_),
    .A2(net157));
 sg13g2_a221oi_1 _0772_ (.B2(_0158_),
    .C1(net164),
    .B1(net129),
    .A1(_0157_),
    .Y(_0003_),
    .A2(net155));
 sg13g2_a221oi_1 _0773_ (.B2(_0159_),
    .C1(net165),
    .B1(net127),
    .A1(_0158_),
    .Y(_0004_),
    .A2(net155));
 sg13g2_a221oi_1 _0774_ (.B2(_0160_),
    .C1(net165),
    .B1(net127),
    .A1(_0159_),
    .Y(_0005_),
    .A2(net155));
 sg13g2_a221oi_1 _0775_ (.B2(_0161_),
    .C1(net165),
    .B1(net127),
    .A1(_0160_),
    .Y(_0006_),
    .A2(net155));
 sg13g2_a221oi_1 _0776_ (.B2(_0162_),
    .C1(net165),
    .B1(net127),
    .A1(_0161_),
    .Y(_0007_),
    .A2(net155));
 sg13g2_a221oi_1 _0777_ (.B2(_0163_),
    .C1(net165),
    .B1(net127),
    .A1(_0162_),
    .Y(_0008_),
    .A2(net155));
 sg13g2_a221oi_1 _0778_ (.B2(_0164_),
    .C1(net165),
    .B1(net127),
    .A1(_0163_),
    .Y(_0009_),
    .A2(net156));
 sg13g2_a221oi_1 _0779_ (.B2(_0165_),
    .C1(net166),
    .B1(net127),
    .A1(_0164_),
    .Y(_0010_),
    .A2(net156));
 sg13g2_a221oi_1 _0780_ (.B2(_0166_),
    .C1(net166),
    .B1(net128),
    .A1(_0165_),
    .Y(_0011_),
    .A2(net156));
 sg13g2_a221oi_1 _0781_ (.B2(_0167_),
    .C1(net166),
    .B1(net128),
    .A1(_0166_),
    .Y(_0012_),
    .A2(net156));
 sg13g2_a221oi_1 _0782_ (.B2(_0168_),
    .C1(net165),
    .B1(net128),
    .A1(_0167_),
    .Y(_0013_),
    .A2(net160));
 sg13g2_a22oi_1 _0783_ (.Y(_0198_),
    .B1(net128),
    .B2(net255),
    .A2(net155),
    .A1(net245));
 sg13g2_nor2_1 _0784_ (.A(net165),
    .B(_0198_),
    .Y(_0014_));
 sg13g2_a22oi_1 _0785_ (.Y(_0199_),
    .B1(net127),
    .B2(net258),
    .A2(net155),
    .A1(net255));
 sg13g2_nor2_1 _0786_ (.A(net164),
    .B(_0199_),
    .Y(_0015_));
 sg13g2_a22oi_1 _0787_ (.Y(_0200_),
    .B1(net129),
    .B2(net282),
    .A2(net157),
    .A1(net258));
 sg13g2_nor2_1 _0788_ (.A(net167),
    .B(_0200_),
    .Y(_0016_));
 sg13g2_a22oi_1 _0789_ (.Y(_0201_),
    .B1(net129),
    .B2(net387),
    .A2(net157),
    .A1(net282));
 sg13g2_nor2_1 _0790_ (.A(net167),
    .B(_0201_),
    .Y(_0017_));
 sg13g2_a22oi_1 _0791_ (.Y(_0202_),
    .B1(net129),
    .B2(net307),
    .A2(net157),
    .A1(\ltc.output_buffer[17] ));
 sg13g2_nor2_1 _0792_ (.A(net167),
    .B(net308),
    .Y(_0018_));
 sg13g2_a22oi_1 _0793_ (.Y(_0203_),
    .B1(net126),
    .B2(net328),
    .A2(net157),
    .A1(net307));
 sg13g2_nor2_1 _0794_ (.A(net161),
    .B(_0203_),
    .Y(_0019_));
 sg13g2_nand2_1 _0795_ (.Y(_0204_),
    .A(net328),
    .B(net149));
 sg13g2_nor2b_1 _0796_ (.A(net228),
    .B_N(net428),
    .Y(_0205_));
 sg13g2_and2_1 _0797_ (.A(_0191_),
    .B(_0205_),
    .X(_0206_));
 sg13g2_nor2b_2 _0798_ (.A(net4),
    .B_N(net3),
    .Y(_0207_));
 sg13g2_nand2_1 _0799_ (.Y(_0208_),
    .A(_0206_),
    .B(_0207_));
 sg13g2_xor2_1 _0800_ (.B(\ltc.output_buffer[66] ),
    .A(\ltc.output_buffer[67] ),
    .X(_0209_));
 sg13g2_xor2_1 _0801_ (.B(\ltc.output_buffer[64] ),
    .A(\ltc.output_buffer[65] ),
    .X(_0210_));
 sg13g2_xnor2_1 _0802_ (.Y(_0211_),
    .A(_0209_),
    .B(_0210_));
 sg13g2_xnor2_1 _0803_ (.Y(_0212_),
    .A(\ltc.output_buffer[71] ),
    .B(\ltc.output_buffer[70] ));
 sg13g2_xor2_1 _0804_ (.B(\ltc.output_buffer[68] ),
    .A(\ltc.output_buffer[69] ),
    .X(_0213_));
 sg13g2_xnor2_1 _0805_ (.Y(_0214_),
    .A(_0212_),
    .B(_0213_));
 sg13g2_xnor2_1 _0806_ (.Y(_0215_),
    .A(_0211_),
    .B(_0214_));
 sg13g2_xnor2_1 _0807_ (.Y(_0216_),
    .A(\ltc.output_buffer[51] ),
    .B(\ltc.output_buffer[50] ));
 sg13g2_xor2_1 _0808_ (.B(\ltc.output_buffer[48] ),
    .A(\ltc.output_buffer[49] ),
    .X(_0217_));
 sg13g2_xnor2_1 _0809_ (.Y(_0218_),
    .A(_0216_),
    .B(_0217_));
 sg13g2_xnor2_1 _0810_ (.Y(_0219_),
    .A(\ltc.output_buffer[55] ),
    .B(\ltc.output_buffer[54] ));
 sg13g2_xor2_1 _0811_ (.B(\ltc.output_buffer[53] ),
    .A(\ltc.output_buffer[52] ),
    .X(_0220_));
 sg13g2_xnor2_1 _0812_ (.Y(_0221_),
    .A(_0219_),
    .B(_0220_));
 sg13g2_xnor2_1 _0813_ (.Y(_0222_),
    .A(_0218_),
    .B(_0221_));
 sg13g2_xnor2_1 _0814_ (.Y(_0223_),
    .A(_0215_),
    .B(_0222_));
 sg13g2_xnor2_1 _0815_ (.Y(_0224_),
    .A(\ltc.output_buffer[63] ),
    .B(\ltc.output_buffer[62] ));
 sg13g2_xor2_1 _0816_ (.B(\ltc.output_buffer[60] ),
    .A(\ltc.output_buffer[61] ),
    .X(_0225_));
 sg13g2_xnor2_1 _0817_ (.Y(_0226_),
    .A(_0224_),
    .B(_0225_));
 sg13g2_xnor2_1 _0818_ (.Y(_0227_),
    .A(\ltc.output_buffer[76] ),
    .B(\ltc.output_buffer[78] ));
 sg13g2_xor2_1 _0819_ (.B(\ltc.output_buffer[77] ),
    .A(\ltc.output_buffer[79] ),
    .X(_0228_));
 sg13g2_xnor2_1 _0820_ (.Y(_0229_),
    .A(_0227_),
    .B(_0228_));
 sg13g2_xnor2_1 _0821_ (.Y(_0230_),
    .A(_0226_),
    .B(_0229_));
 sg13g2_xnor2_1 _0822_ (.Y(_0231_),
    .A(\ltc.output_buffer[59] ),
    .B(\ltc.output_buffer[58] ));
 sg13g2_xnor2_1 _0823_ (.Y(_0232_),
    .A(\ltc.output_buffer[73] ),
    .B(\ltc.output_buffer[72] ));
 sg13g2_xnor2_1 _0824_ (.Y(_0233_),
    .A(_0231_),
    .B(_0232_));
 sg13g2_xor2_1 _0825_ (.B(\ltc.output_buffer[56] ),
    .A(\ltc.output_buffer[57] ),
    .X(_0234_));
 sg13g2_xnor2_1 _0826_ (.Y(_0235_),
    .A(\ltc.output_buffer[75] ),
    .B(\ltc.output_buffer[74] ));
 sg13g2_xnor2_1 _0827_ (.Y(_0236_),
    .A(_0234_),
    .B(_0235_));
 sg13g2_xnor2_1 _0828_ (.Y(_0237_),
    .A(_0233_),
    .B(_0236_));
 sg13g2_xnor2_1 _0829_ (.Y(_0238_),
    .A(_0230_),
    .B(_0237_));
 sg13g2_xnor2_1 _0830_ (.Y(_0239_),
    .A(_0223_),
    .B(_0238_));
 sg13g2_xnor2_1 _0831_ (.Y(_0240_),
    .A(\ltc.output_buffer[19] ),
    .B(\ltc.output_buffer[18] ));
 sg13g2_xor2_1 _0832_ (.B(\ltc.output_buffer[16] ),
    .A(\ltc.output_buffer[17] ),
    .X(_0241_));
 sg13g2_xnor2_1 _0833_ (.Y(_0242_),
    .A(_0240_),
    .B(_0241_));
 sg13g2_xnor2_1 _0834_ (.Y(_0243_),
    .A(\ltc.output_buffer[23] ),
    .B(\ltc.output_buffer[22] ));
 sg13g2_xor2_1 _0835_ (.B(\ltc.output_buffer[20] ),
    .A(\ltc.output_buffer[21] ),
    .X(_0244_));
 sg13g2_xnor2_1 _0836_ (.Y(_0245_),
    .A(_0243_),
    .B(_0244_));
 sg13g2_xnor2_1 _0837_ (.Y(_0246_),
    .A(_0242_),
    .B(_0245_));
 sg13g2_xor2_1 _0838_ (.B(\ltc.output_buffer[34] ),
    .A(\ltc.output_buffer[35] ),
    .X(_0247_));
 sg13g2_xnor2_1 _0839_ (.Y(_0248_),
    .A(\ltc.output_buffer[37] ),
    .B(\ltc.output_buffer[36] ));
 sg13g2_xnor2_1 _0840_ (.Y(_0249_),
    .A(_0247_),
    .B(_0248_));
 sg13g2_xor2_1 _0841_ (.B(\ltc.output_buffer[32] ),
    .A(\ltc.output_buffer[33] ),
    .X(_0250_));
 sg13g2_xnor2_1 _0842_ (.Y(_0251_),
    .A(\ltc.output_buffer[39] ),
    .B(\ltc.output_buffer[38] ));
 sg13g2_xnor2_1 _0843_ (.Y(_0252_),
    .A(_0250_),
    .B(_0251_));
 sg13g2_xnor2_1 _0844_ (.Y(_0253_),
    .A(_0249_),
    .B(_0252_));
 sg13g2_xnor2_1 _0845_ (.Y(_0254_),
    .A(_0246_),
    .B(_0253_));
 sg13g2_xor2_1 _0846_ (.B(\ltc.output_buffer[30] ),
    .A(\ltc.output_buffer[31] ),
    .X(_0255_));
 sg13g2_xor2_1 _0847_ (.B(\ltc.output_buffer[28] ),
    .A(\ltc.output_buffer[29] ),
    .X(_0256_));
 sg13g2_xnor2_1 _0848_ (.Y(_0257_),
    .A(_0255_),
    .B(_0256_));
 sg13g2_xnor2_1 _0849_ (.Y(_0258_),
    .A(\ltc.output_buffer[47] ),
    .B(\ltc.output_buffer[46] ));
 sg13g2_xor2_1 _0850_ (.B(\ltc.output_buffer[44] ),
    .A(\ltc.output_buffer[45] ),
    .X(_0259_));
 sg13g2_xnor2_1 _0851_ (.Y(_0260_),
    .A(_0258_),
    .B(_0259_));
 sg13g2_xnor2_1 _0852_ (.Y(_0261_),
    .A(_0257_),
    .B(_0260_));
 sg13g2_xnor2_1 _0853_ (.Y(_0262_),
    .A(\ltc.output_buffer[27] ),
    .B(\ltc.output_buffer[26] ));
 sg13g2_xnor2_1 _0854_ (.Y(_0263_),
    .A(\ltc.output_buffer[41] ),
    .B(\ltc.output_buffer[40] ));
 sg13g2_xnor2_1 _0855_ (.Y(_0264_),
    .A(_0262_),
    .B(_0263_));
 sg13g2_xor2_1 _0856_ (.B(\ltc.output_buffer[24] ),
    .A(\ltc.output_buffer[25] ),
    .X(_0265_));
 sg13g2_xnor2_1 _0857_ (.Y(_0266_),
    .A(\ltc.output_buffer[43] ),
    .B(\ltc.output_buffer[42] ));
 sg13g2_xnor2_1 _0858_ (.Y(_0267_),
    .A(_0265_),
    .B(_0266_));
 sg13g2_xnor2_1 _0859_ (.Y(_0268_),
    .A(_0264_),
    .B(_0267_));
 sg13g2_xnor2_1 _0860_ (.Y(_0269_),
    .A(_0261_),
    .B(_0268_));
 sg13g2_xnor2_1 _0861_ (.Y(_0270_),
    .A(_0254_),
    .B(_0269_));
 sg13g2_xnor2_1 _0862_ (.Y(_0271_),
    .A(_0239_),
    .B(_0270_));
 sg13g2_nand2_1 _0863_ (.Y(_0272_),
    .A(\ltc.output_buffer[20] ),
    .B(net136));
 sg13g2_a21oi_1 _0864_ (.A1(_0208_),
    .A2(_0272_),
    .Y(_0273_),
    .B1(net153));
 sg13g2_o21ai_1 _0865_ (.B1(_0273_),
    .Y(_0274_),
    .A1(_0208_),
    .A2(_0271_));
 sg13g2_a21oi_1 _0866_ (.A1(_0204_),
    .A2(_0274_),
    .Y(_0020_),
    .B1(net161));
 sg13g2_a22oi_1 _0867_ (.Y(_0275_),
    .B1(net132),
    .B2(net319),
    .A2(net150),
    .A1(\ltc.output_buffer[20] ));
 sg13g2_nor2_1 _0868_ (.A(net163),
    .B(net320),
    .Y(_0021_));
 sg13g2_nand3_1 _0869_ (.B(net319),
    .C(net150),
    .A(net172),
    .Y(_0276_));
 sg13g2_nor2_1 _0870_ (.A(net330),
    .B(net134),
    .Y(_0277_));
 sg13g2_o21ai_1 _0871_ (.B1(net143),
    .Y(_0278_),
    .A1(net276),
    .A2(net139));
 sg13g2_o21ai_1 _0872_ (.B1(_0276_),
    .Y(_0022_),
    .A1(_0277_),
    .A2(_0278_));
 sg13g2_nor2_1 _0873_ (.A(\ltc.hrs_d[0] ),
    .B(net134),
    .Y(_0279_));
 sg13g2_o21ai_1 _0874_ (.B1(net144),
    .Y(_0280_),
    .A1(\ltc.output_buffer[23] ),
    .A2(net139));
 sg13g2_nand3_1 _0875_ (.B(net276),
    .C(net150),
    .A(net172),
    .Y(_0281_));
 sg13g2_o21ai_1 _0876_ (.B1(_0281_),
    .Y(_0023_),
    .A1(_0279_),
    .A2(_0280_));
 sg13g2_a22oi_1 _0877_ (.Y(_0282_),
    .B1(net125),
    .B2(net358),
    .A2(net149),
    .A1(\ltc.output_buffer[23] ));
 sg13g2_nor2_1 _0878_ (.A(net161),
    .B(net359),
    .Y(_0024_));
 sg13g2_a22oi_1 _0879_ (.Y(_0283_),
    .B1(net125),
    .B2(net384),
    .A2(net149),
    .A1(net358));
 sg13g2_nor2_1 _0880_ (.A(net161),
    .B(_0283_),
    .Y(_0025_));
 sg13g2_a22oi_1 _0881_ (.Y(_0284_),
    .B1(net124),
    .B2(net380),
    .A2(net149),
    .A1(\ltc.output_buffer[25] ));
 sg13g2_nor2_1 _0882_ (.A(net161),
    .B(net381),
    .Y(_0026_));
 sg13g2_a22oi_1 _0883_ (.Y(_0285_),
    .B1(net125),
    .B2(net366),
    .A2(net149),
    .A1(\ltc.output_buffer[26] ));
 sg13g2_nor2_1 _0884_ (.A(net161),
    .B(net367),
    .Y(_0027_));
 sg13g2_nand3_1 _0885_ (.B(net366),
    .C(net149),
    .A(net172),
    .Y(_0286_));
 sg13g2_nor2_1 _0886_ (.A(net374),
    .B(net133),
    .Y(_0287_));
 sg13g2_o21ai_1 _0887_ (.B1(net143),
    .Y(_0288_),
    .A1(net315),
    .A2(net138));
 sg13g2_o21ai_1 _0888_ (.B1(_0286_),
    .Y(_0028_),
    .A1(_0287_),
    .A2(_0288_));
 sg13g2_nor2_1 _0889_ (.A(\ltc.hrs_u[2] ),
    .B(net133),
    .Y(_0289_));
 sg13g2_o21ai_1 _0890_ (.B1(net143),
    .Y(_0290_),
    .A1(net288),
    .A2(net138));
 sg13g2_nand3_1 _0891_ (.B(net315),
    .C(net148),
    .A(net170),
    .Y(_0291_));
 sg13g2_o21ai_1 _0892_ (.B1(_0291_),
    .Y(_0029_),
    .A1(_0289_),
    .A2(_0290_));
 sg13g2_nor2_1 _0893_ (.A(\ltc.hrs_u[1] ),
    .B(net133),
    .Y(_0292_));
 sg13g2_o21ai_1 _0894_ (.B1(net143),
    .Y(_0293_),
    .A1(\ltc.output_buffer[30] ),
    .A2(net138));
 sg13g2_nand3_1 _0895_ (.B(net288),
    .C(net148),
    .A(net170),
    .Y(_0294_));
 sg13g2_o21ai_1 _0896_ (.B1(_0294_),
    .Y(_0030_),
    .A1(_0292_),
    .A2(_0293_));
 sg13g2_nor2_1 _0897_ (.A(\ltc.output_buffer[31] ),
    .B(net138),
    .Y(_0295_));
 sg13g2_o21ai_1 _0898_ (.B1(net143),
    .Y(_0296_),
    .A1(\ltc.hrs_u[0] ),
    .A2(net133));
 sg13g2_nand3_1 _0899_ (.B(net290),
    .C(net148),
    .A(net170),
    .Y(_0297_));
 sg13g2_o21ai_1 _0900_ (.B1(_0297_),
    .Y(_0031_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_a22oi_1 _0901_ (.Y(_0298_),
    .B1(net124),
    .B2(net360),
    .A2(net147),
    .A1(\ltc.output_buffer[31] ));
 sg13g2_nor2_1 _0902_ (.A(net162),
    .B(net361),
    .Y(_0032_));
 sg13g2_a22oi_1 _0903_ (.Y(_0299_),
    .B1(net124),
    .B2(net313),
    .A2(net148),
    .A1(\ltc.output_buffer[32] ));
 sg13g2_nor2_1 _0904_ (.A(net162),
    .B(net314),
    .Y(_0033_));
 sg13g2_a22oi_1 _0905_ (.Y(_0300_),
    .B1(net124),
    .B2(net368),
    .A2(net147),
    .A1(net313));
 sg13g2_nor2_1 _0906_ (.A(net162),
    .B(_0300_),
    .Y(_0034_));
 sg13g2_a22oi_1 _0907_ (.Y(_0301_),
    .B1(net124),
    .B2(net333),
    .A2(net147),
    .A1(\ltc.output_buffer[34] ));
 sg13g2_nor2_1 _0908_ (.A(net162),
    .B(net334),
    .Y(_0035_));
 sg13g2_a22oi_1 _0909_ (.Y(_0302_),
    .B1(net124),
    .B2(net292),
    .A2(net147),
    .A1(net333));
 sg13g2_nor2_1 _0910_ (.A(net162),
    .B(_0302_),
    .Y(_0036_));
 sg13g2_nand3_1 _0911_ (.B(net292),
    .C(net147),
    .A(net170),
    .Y(_0303_));
 sg13g2_nor2_1 _0912_ (.A(\ltc.output_buffer[37] ),
    .B(net138),
    .Y(_0304_));
 sg13g2_o21ai_1 _0913_ (.B1(net143),
    .Y(_0305_),
    .A1(\ltc.min_d[2] ),
    .A2(net133));
 sg13g2_o21ai_1 _0914_ (.B1(_0303_),
    .Y(_0037_),
    .A1(_0304_),
    .A2(_0305_));
 sg13g2_nor2_1 _0915_ (.A(\ltc.min_d[1] ),
    .B(net133),
    .Y(_0306_));
 sg13g2_o21ai_1 _0916_ (.B1(net143),
    .Y(_0307_),
    .A1(net305),
    .A2(net138));
 sg13g2_nand3_1 _0917_ (.B(net317),
    .C(net147),
    .A(net170),
    .Y(_0308_));
 sg13g2_o21ai_1 _0918_ (.B1(_0308_),
    .Y(_0038_),
    .A1(_0306_),
    .A2(_0307_));
 sg13g2_nor2_1 _0919_ (.A(\ltc.min_d[0] ),
    .B(net133),
    .Y(_0309_));
 sg13g2_o21ai_1 _0920_ (.B1(net143),
    .Y(_0310_),
    .A1(\ltc.output_buffer[39] ),
    .A2(net138));
 sg13g2_nand3_1 _0921_ (.B(net305),
    .C(net147),
    .A(net171),
    .Y(_0311_));
 sg13g2_o21ai_1 _0922_ (.B1(_0311_),
    .Y(_0039_),
    .A1(_0309_),
    .A2(_0310_));
 sg13g2_a22oi_1 _0923_ (.Y(_0312_),
    .B1(net124),
    .B2(net369),
    .A2(net147),
    .A1(\ltc.output_buffer[39] ));
 sg13g2_nor2_1 _0924_ (.A(net162),
    .B(net370),
    .Y(_0040_));
 sg13g2_a22oi_1 _0925_ (.Y(_0313_),
    .B1(net125),
    .B2(net386),
    .A2(net149),
    .A1(net369));
 sg13g2_nor2_1 _0926_ (.A(net161),
    .B(_0313_),
    .Y(_0041_));
 sg13g2_a22oi_1 _0927_ (.Y(_0314_),
    .B1(net125),
    .B2(net354),
    .A2(net149),
    .A1(\ltc.output_buffer[41] ));
 sg13g2_nor2_1 _0928_ (.A(net161),
    .B(net355),
    .Y(_0042_));
 sg13g2_a22oi_1 _0929_ (.Y(_0315_),
    .B1(net124),
    .B2(net350),
    .A2(net150),
    .A1(\ltc.output_buffer[42] ));
 sg13g2_nor2_1 _0930_ (.A(net162),
    .B(net351),
    .Y(_0043_));
 sg13g2_nand3_1 _0931_ (.B(net350),
    .C(net148),
    .A(net172),
    .Y(_0316_));
 sg13g2_nor2_1 _0932_ (.A(net392),
    .B(net133),
    .Y(_0317_));
 sg13g2_o21ai_1 _0933_ (.B1(net144),
    .Y(_0318_),
    .A1(net324),
    .A2(net139));
 sg13g2_o21ai_1 _0934_ (.B1(_0316_),
    .Y(_0044_),
    .A1(_0317_),
    .A2(_0318_));
 sg13g2_nor2_1 _0935_ (.A(\ltc.min_u[2] ),
    .B(net134),
    .Y(_0319_));
 sg13g2_o21ai_1 _0936_ (.B1(net144),
    .Y(_0320_),
    .A1(net299),
    .A2(net139));
 sg13g2_nand3_1 _0937_ (.B(net324),
    .C(net151),
    .A(net171),
    .Y(_0321_));
 sg13g2_o21ai_1 _0938_ (.B1(_0321_),
    .Y(_0045_),
    .A1(_0319_),
    .A2(_0320_));
 sg13g2_nor2_1 _0939_ (.A(\ltc.min_u[1] ),
    .B(net137),
    .Y(_0322_));
 sg13g2_o21ai_1 _0940_ (.B1(net144),
    .Y(_0323_),
    .A1(\ltc.output_buffer[46] ),
    .A2(net139));
 sg13g2_nand3_1 _0941_ (.B(net299),
    .C(net151),
    .A(net171),
    .Y(_0324_));
 sg13g2_o21ai_1 _0942_ (.B1(_0324_),
    .Y(_0046_),
    .A1(_0322_),
    .A2(_0323_));
 sg13g2_nor2_1 _0943_ (.A(\ltc.min_u[0] ),
    .B(net137),
    .Y(_0325_));
 sg13g2_o21ai_1 _0944_ (.B1(net144),
    .Y(_0326_),
    .A1(\ltc.output_buffer[47] ),
    .A2(net139));
 sg13g2_nand3_1 _0945_ (.B(net301),
    .C(net151),
    .A(net173),
    .Y(_0327_));
 sg13g2_o21ai_1 _0946_ (.B1(_0327_),
    .Y(_0047_),
    .A1(_0325_),
    .A2(_0326_));
 sg13g2_a22oi_1 _0947_ (.Y(_0328_),
    .B1(net132),
    .B2(net348),
    .A2(net152),
    .A1(\ltc.output_buffer[47] ));
 sg13g2_nor2_1 _0948_ (.A(net169),
    .B(net349),
    .Y(_0048_));
 sg13g2_a22oi_1 _0949_ (.Y(_0329_),
    .B1(net126),
    .B2(net373),
    .A2(net151),
    .A1(net348));
 sg13g2_nor2_1 _0950_ (.A(net163),
    .B(_0329_),
    .Y(_0049_));
 sg13g2_a22oi_1 _0951_ (.Y(_0330_),
    .B1(net126),
    .B2(net371),
    .A2(net151),
    .A1(\ltc.output_buffer[49] ));
 sg13g2_nor2_1 _0952_ (.A(net163),
    .B(net372),
    .Y(_0050_));
 sg13g2_a22oi_1 _0953_ (.Y(_0331_),
    .B1(net126),
    .B2(net263),
    .A2(net151),
    .A1(net371));
 sg13g2_nor2_1 _0954_ (.A(net169),
    .B(_0331_),
    .Y(_0051_));
 sg13g2_nand2_1 _0955_ (.Y(_0332_),
    .A(net263),
    .B(net151));
 sg13g2_nor2_2 _0956_ (.A(net4),
    .B(net3),
    .Y(_0333_));
 sg13g2_and2_1 _0957_ (.A(net4),
    .B(net3),
    .X(_0334_));
 sg13g2_o21ai_1 _0958_ (.B1(_0206_),
    .Y(_0335_),
    .A1(_0333_),
    .A2(_0334_));
 sg13g2_nand2_1 _0959_ (.Y(_0336_),
    .A(\ltc.output_buffer[52] ),
    .B(net134));
 sg13g2_a21oi_1 _0960_ (.A1(_0335_),
    .A2(_0336_),
    .Y(_0337_),
    .B1(net153));
 sg13g2_o21ai_1 _0961_ (.B1(_0337_),
    .Y(_0338_),
    .A1(_0271_),
    .A2(_0335_));
 sg13g2_a21oi_1 _0962_ (.A1(_0332_),
    .A2(_0338_),
    .Y(_0052_),
    .B1(net163));
 sg13g2_nor2_1 _0963_ (.A(\ltc.sec_d[2] ),
    .B(net134),
    .Y(_0339_));
 sg13g2_o21ai_1 _0964_ (.B1(net144),
    .Y(_0340_),
    .A1(\ltc.output_buffer[53] ),
    .A2(net142));
 sg13g2_nand3_1 _0965_ (.B(net278),
    .C(net152),
    .A(net173),
    .Y(_0341_));
 sg13g2_o21ai_1 _0966_ (.B1(_0341_),
    .Y(_0053_),
    .A1(_0339_),
    .A2(_0340_));
 sg13g2_nor2_1 _0967_ (.A(\ltc.sec_d[1] ),
    .B(net134),
    .Y(_0342_));
 sg13g2_o21ai_1 _0968_ (.B1(_0179_),
    .Y(_0343_),
    .A1(\ltc.output_buffer[54] ),
    .A2(net142));
 sg13g2_nand3_1 _0969_ (.B(net342),
    .C(net152),
    .A(net173),
    .Y(_0344_));
 sg13g2_o21ai_1 _0970_ (.B1(_0344_),
    .Y(_0054_),
    .A1(_0342_),
    .A2(_0343_));
 sg13g2_nor2_1 _0971_ (.A(\ltc.sec_d[0] ),
    .B(net134),
    .Y(_0345_));
 sg13g2_o21ai_1 _0972_ (.B1(net144),
    .Y(_0346_),
    .A1(\ltc.output_buffer[55] ),
    .A2(net139));
 sg13g2_nand3_1 _0973_ (.B(net344),
    .C(net152),
    .A(net173),
    .Y(_0347_));
 sg13g2_o21ai_1 _0974_ (.B1(_0347_),
    .Y(_0055_),
    .A1(_0345_),
    .A2(_0346_));
 sg13g2_a22oi_1 _0975_ (.Y(_0348_),
    .B1(net126),
    .B2(net346),
    .A2(net153),
    .A1(\ltc.output_buffer[55] ));
 sg13g2_nor2_1 _0976_ (.A(net163),
    .B(net347),
    .Y(_0056_));
 sg13g2_a22oi_1 _0977_ (.Y(_0349_),
    .B1(net126),
    .B2(net303),
    .A2(net153),
    .A1(\ltc.output_buffer[56] ));
 sg13g2_nor2_1 _0978_ (.A(net163),
    .B(net304),
    .Y(_0057_));
 sg13g2_a22oi_1 _0979_ (.Y(_0350_),
    .B1(net130),
    .B2(net382),
    .A2(net158),
    .A1(net303));
 sg13g2_nor2_1 _0980_ (.A(net164),
    .B(_0350_),
    .Y(_0058_));
 sg13g2_a22oi_1 _0981_ (.Y(_0351_),
    .B1(net130),
    .B2(net364),
    .A2(net158),
    .A1(net382));
 sg13g2_nor2_1 _0982_ (.A(net164),
    .B(_0351_),
    .Y(_0059_));
 sg13g2_nand3_1 _0983_ (.B(net364),
    .C(net158),
    .A(net175),
    .Y(_0352_));
 sg13g2_nor2_1 _0984_ (.A(\ltc.sec_u[3] ),
    .B(net135),
    .Y(_0353_));
 sg13g2_o21ai_1 _0985_ (.B1(net145),
    .Y(_0354_),
    .A1(net356),
    .A2(net140));
 sg13g2_o21ai_1 _0986_ (.B1(_0352_),
    .Y(_0060_),
    .A1(_0353_),
    .A2(_0354_));
 sg13g2_nor2_1 _0987_ (.A(net335),
    .B(net140),
    .Y(_0355_));
 sg13g2_o21ai_1 _0988_ (.B1(net145),
    .Y(_0356_),
    .A1(\ltc.sec_u[2] ),
    .A2(net135));
 sg13g2_nand3_1 _0989_ (.B(net356),
    .C(net153),
    .A(net175),
    .Y(_0357_));
 sg13g2_o21ai_1 _0990_ (.B1(_0357_),
    .Y(_0061_),
    .A1(_0355_),
    .A2(_0356_));
 sg13g2_nor2_1 _0991_ (.A(\ltc.sec_u[1] ),
    .B(net135),
    .Y(_0358_));
 sg13g2_o21ai_1 _0992_ (.B1(net145),
    .Y(_0359_),
    .A1(net295),
    .A2(net140));
 sg13g2_nand3_1 _0993_ (.B(net335),
    .C(net158),
    .A(net175),
    .Y(_0360_));
 sg13g2_o21ai_1 _0994_ (.B1(_0360_),
    .Y(_0062_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_nor2_1 _0995_ (.A(\ltc.output_buffer[63] ),
    .B(net140),
    .Y(_0361_));
 sg13g2_o21ai_1 _0996_ (.B1(net145),
    .Y(_0362_),
    .A1(\ltc.sec_u[0] ),
    .A2(net135));
 sg13g2_nand3_1 _0997_ (.B(net295),
    .C(net158),
    .A(net175),
    .Y(_0363_));
 sg13g2_o21ai_1 _0998_ (.B1(_0363_),
    .Y(_0063_),
    .A1(_0361_),
    .A2(_0362_));
 sg13g2_a22oi_1 _0999_ (.Y(_0364_),
    .B1(net130),
    .B2(net362),
    .A2(net158),
    .A1(\ltc.output_buffer[63] ));
 sg13g2_nor2_1 _1000_ (.A(net164),
    .B(net363),
    .Y(_0064_));
 sg13g2_a22oi_1 _1001_ (.Y(_0365_),
    .B1(net130),
    .B2(net423),
    .A2(net157),
    .A1(net362));
 sg13g2_nor2_1 _1002_ (.A(net164),
    .B(_0365_),
    .Y(_0065_));
 sg13g2_a22oi_1 _1003_ (.Y(_0366_),
    .B1(net131),
    .B2(net331),
    .A2(net156),
    .A1(\ltc.output_buffer[65] ));
 sg13g2_nor2_1 _1004_ (.A(net166),
    .B(net332),
    .Y(_0066_));
 sg13g2_a22oi_1 _1005_ (.Y(_0367_),
    .B1(net131),
    .B2(net321),
    .A2(net156),
    .A1(\ltc.output_buffer[66] ));
 sg13g2_nor2_1 _1006_ (.A(net166),
    .B(net322),
    .Y(_0067_));
 sg13g2_a22oi_1 _1007_ (.Y(_0368_),
    .B1(net131),
    .B2(net311),
    .A2(net156),
    .A1(\ltc.output_buffer[67] ));
 sg13g2_nor2_1 _1008_ (.A(net166),
    .B(net312),
    .Y(_0068_));
 sg13g2_a22oi_1 _1009_ (.Y(_0369_),
    .B1(net130),
    .B2(net280),
    .A2(net159),
    .A1(net311));
 sg13g2_nor2_1 _1010_ (.A(net166),
    .B(_0369_),
    .Y(_0069_));
 sg13g2_nand3_1 _1011_ (.B(net280),
    .C(net159),
    .A(net175),
    .Y(_0370_));
 sg13g2_nor2_1 _1012_ (.A(\ltc.frm_d[1] ),
    .B(net135),
    .Y(_0371_));
 sg13g2_o21ai_1 _1013_ (.B1(net145),
    .Y(_0372_),
    .A1(\ltc.output_buffer[70] ),
    .A2(net140));
 sg13g2_o21ai_1 _1014_ (.B1(_0370_),
    .Y(_0070_),
    .A1(_0371_),
    .A2(_0372_));
 sg13g2_nor2_1 _1015_ (.A(\ltc.frm_d[0] ),
    .B(net135),
    .Y(_0373_));
 sg13g2_o21ai_1 _1016_ (.B1(net145),
    .Y(_0374_),
    .A1(\ltc.output_buffer[71] ),
    .A2(net140));
 sg13g2_nand3_1 _1017_ (.B(net297),
    .C(net160),
    .A(net175),
    .Y(_0375_));
 sg13g2_o21ai_1 _1018_ (.B1(_0375_),
    .Y(_0071_),
    .A1(_0373_),
    .A2(_0374_));
 sg13g2_a22oi_1 _1019_ (.Y(_0376_),
    .B1(net130),
    .B2(net340),
    .A2(net159),
    .A1(\ltc.output_buffer[71] ));
 sg13g2_nor2_1 _1020_ (.A(net168),
    .B(net341),
    .Y(_0072_));
 sg13g2_a22oi_1 _1021_ (.Y(_0377_),
    .B1(net130),
    .B2(net385),
    .A2(net159),
    .A1(net340));
 sg13g2_nor2_1 _1022_ (.A(net168),
    .B(_0377_),
    .Y(_0073_));
 sg13g2_a22oi_1 _1023_ (.Y(_0378_),
    .B1(net130),
    .B2(net326),
    .A2(net159),
    .A1(\ltc.output_buffer[73] ));
 sg13g2_nor2_1 _1024_ (.A(net168),
    .B(net327),
    .Y(_0074_));
 sg13g2_a22oi_1 _1025_ (.Y(_0379_),
    .B1(net131),
    .B2(net271),
    .A2(net159),
    .A1(net326));
 sg13g2_nor2_1 _1026_ (.A(net168),
    .B(_0379_),
    .Y(_0075_));
 sg13g2_nand3_1 _1027_ (.B(net271),
    .C(net160),
    .A(net174),
    .Y(_0380_));
 sg13g2_nor2_1 _1028_ (.A(\ltc.frm_u[3] ),
    .B(net135),
    .Y(_0381_));
 sg13g2_o21ai_1 _1029_ (.B1(net146),
    .Y(_0382_),
    .A1(\ltc.output_buffer[76] ),
    .A2(net141));
 sg13g2_o21ai_1 _1030_ (.B1(_0380_),
    .Y(_0076_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_nor2_1 _1031_ (.A(\ltc.output_buffer[77] ),
    .B(net141),
    .Y(_0383_));
 sg13g2_o21ai_1 _1032_ (.B1(net146),
    .Y(_0384_),
    .A1(\ltc.frm_u[2] ),
    .A2(net136));
 sg13g2_nand3_1 _1033_ (.B(net283),
    .C(net158),
    .A(net176),
    .Y(_0385_));
 sg13g2_o21ai_1 _1034_ (.B1(_0385_),
    .Y(_0077_),
    .A1(_0383_),
    .A2(_0384_));
 sg13g2_nor2_1 _1035_ (.A(\ltc.frm_u[1] ),
    .B(net136),
    .Y(_0386_));
 sg13g2_o21ai_1 _1036_ (.B1(net145),
    .Y(_0387_),
    .A1(net309),
    .A2(net140));
 sg13g2_nand3_1 _1037_ (.B(net352),
    .C(net158),
    .A(net174),
    .Y(_0388_));
 sg13g2_o21ai_1 _1038_ (.B1(_0388_),
    .Y(_0078_),
    .A1(_0386_),
    .A2(_0387_));
 sg13g2_nor2_1 _1039_ (.A(net294),
    .B(net135),
    .Y(_0389_));
 sg13g2_o21ai_1 _1040_ (.B1(net145),
    .Y(_0390_),
    .A1(\ltc.output_buffer[79] ),
    .A2(net140));
 sg13g2_nand3_1 _1041_ (.B(net309),
    .C(net159),
    .A(net174),
    .Y(_0391_));
 sg13g2_o21ai_1 _1042_ (.B1(_0391_),
    .Y(_0079_),
    .A1(_0389_),
    .A2(_0390_));
 sg13g2_nand3b_1 _1043_ (.B(net429),
    .C(net402),
    .Y(_0392_),
    .A_N(net407));
 sg13g2_nor2_1 _1044_ (.A(_0151_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_nor4_1 _1045_ (.A(net416),
    .B(_0150_),
    .C(net430),
    .D(net439),
    .Y(_0394_));
 sg13g2_nand3b_1 _1046_ (.B(net441),
    .C(_0394_),
    .Y(_0395_),
    .A_N(net374));
 sg13g2_nand2_1 _1047_ (.Y(_0396_),
    .A(net374),
    .B(net416));
 sg13g2_nor3_2 _1048_ (.A(net441),
    .B(net439),
    .C(_0396_),
    .Y(_0397_));
 sg13g2_nor2_1 _1049_ (.A(_0392_),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_a21oi_1 _1050_ (.A1(_0395_),
    .A2(_0398_),
    .Y(_0399_),
    .B1(net439));
 sg13g2_o21ai_1 _1051_ (.B1(net170),
    .Y(_0080_),
    .A1(_0393_),
    .A2(net440));
 sg13g2_and4_1 _1052_ (.A(\ltc.frm_counter[3] ),
    .B(net260),
    .C(net228),
    .D(net428),
    .X(_0400_));
 sg13g2_nand4_1 _1053_ (.B(net260),
    .C(net228),
    .A(net450),
    .Y(_0401_),
    .D(net428));
 sg13g2_nand2_1 _1054_ (.Y(_0402_),
    .A(\ltc.frm_counter[6] ),
    .B(\ltc.frm_counter[7] ));
 sg13g2_and4_1 _1055_ (.A(\ltc.frm_counter[5] ),
    .B(\ltc.frm_counter[4] ),
    .C(\ltc.frm_counter[6] ),
    .D(\ltc.frm_counter[7] ),
    .X(_0403_));
 sg13g2_nand4_1 _1056_ (.B(\ltc.frm_counter[4] ),
    .C(\ltc.frm_counter[6] ),
    .A(\ltc.frm_counter[5] ),
    .Y(_0404_),
    .D(\ltc.frm_counter[7] ));
 sg13g2_nor2_1 _1057_ (.A(_0401_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_nand2_1 _1058_ (.Y(_0406_),
    .A(_0400_),
    .B(_0403_));
 sg13g2_nand4_1 _1059_ (.B(\ltc.frm_counter[8] ),
    .C(\ltc.frm_counter[10] ),
    .A(\ltc.frm_counter[9] ),
    .Y(_0407_),
    .D(net399));
 sg13g2_nor3_1 _1060_ (.A(_0401_),
    .B(_0404_),
    .C(_0407_),
    .Y(_0408_));
 sg13g2_nor4_2 _1061_ (.A(_0152_),
    .B(_0401_),
    .C(_0404_),
    .Y(_0409_),
    .D(_0407_));
 sg13g2_nand2_1 _1062_ (.Y(_0410_),
    .A(net461),
    .B(_0409_));
 sg13g2_nand3_1 _1063_ (.B(net471),
    .C(_0409_),
    .A(net461),
    .Y(_0411_));
 sg13g2_and4_1 _1064_ (.A(net461),
    .B(\ltc.frm_counter[14] ),
    .C(net459),
    .D(_0409_),
    .X(_0412_));
 sg13g2_and2_1 _1065_ (.A(net464),
    .B(_0412_),
    .X(_0413_));
 sg13g2_nand3_1 _1066_ (.B(\ltc.frm_counter[17] ),
    .C(_0412_),
    .A(\ltc.frm_counter[16] ),
    .Y(_0414_));
 sg13g2_nand3_1 _1067_ (.B(\ltc.frm_counter[18] ),
    .C(_0413_),
    .A(\ltc.frm_counter[17] ),
    .Y(_0415_));
 sg13g2_xor2_1 _1068_ (.B(_0414_),
    .A(net454),
    .X(_0416_));
 sg13g2_or2_1 _1069_ (.X(_0417_),
    .B(_0416_),
    .A(_0186_));
 sg13g2_xnor2_1 _1070_ (.Y(_0418_),
    .A(_0153_),
    .B(_0413_));
 sg13g2_xnor2_1 _1071_ (.Y(_0419_),
    .A(net464),
    .B(_0412_));
 sg13g2_xnor2_1 _1072_ (.Y(_0420_),
    .A(net468),
    .B(_0408_));
 sg13g2_or2_1 _1073_ (.X(_0421_),
    .B(_0409_),
    .A(net461));
 sg13g2_nor2_1 _1074_ (.A(net474),
    .B(_0420_),
    .Y(_0422_));
 sg13g2_and3_1 _1075_ (.X(_0423_),
    .A(net425),
    .B(net436),
    .C(_0400_));
 sg13g2_and4_1 _1076_ (.A(net425),
    .B(net436),
    .C(net453),
    .D(_0400_),
    .X(_0424_));
 sg13g2_nor2b_1 _1077_ (.A(\ltc.frm_counter[8] ),
    .B_N(\ltc.frm_counter[9] ),
    .Y(_0425_));
 sg13g2_nand2_1 _1078_ (.Y(_0426_),
    .A(\ltc.frm_counter[11] ),
    .B(_0425_));
 sg13g2_nand3_1 _1079_ (.B(_0334_),
    .C(_0402_),
    .A(_0187_),
    .Y(_0427_));
 sg13g2_nor3_1 _1080_ (.A(\ltc.frm_counter[10] ),
    .B(_0426_),
    .C(_0427_),
    .Y(_0428_));
 sg13g2_and2_1 _1081_ (.A(_0424_),
    .B(_0428_),
    .X(_0429_));
 sg13g2_nand4_1 _1082_ (.B(_0419_),
    .C(_0422_),
    .A(_0418_),
    .Y(_0430_),
    .D(_0429_));
 sg13g2_and4_1 _1083_ (.A(\ltc.frm_counter[9] ),
    .B(\ltc.frm_counter[8] ),
    .C(_0400_),
    .D(_0403_),
    .X(_0431_));
 sg13g2_a21oi_1 _1084_ (.A1(\ltc.frm_counter[10] ),
    .A2(_0431_),
    .Y(_0432_),
    .B1(net399));
 sg13g2_xnor2_1 _1085_ (.Y(_0433_),
    .A(net457),
    .B(_0431_));
 sg13g2_o21ai_1 _1086_ (.B1(_0433_),
    .Y(_0434_),
    .A1(_0408_),
    .A2(_0432_));
 sg13g2_nor3_1 _1087_ (.A(_0153_),
    .B(_0419_),
    .C(_0434_),
    .Y(_0435_));
 sg13g2_xor2_1 _1088_ (.B(_0411_),
    .A(net459),
    .X(_0436_));
 sg13g2_a21oi_1 _1089_ (.A1(_0400_),
    .A2(_0403_),
    .Y(_0437_),
    .B1(net469));
 sg13g2_or3_1 _1090_ (.A(_0188_),
    .B(_0431_),
    .C(_0437_),
    .X(_0438_));
 sg13g2_o21ai_1 _1091_ (.B1(_0406_),
    .Y(_0439_),
    .A1(net470),
    .A2(_0424_));
 sg13g2_nand4_1 _1092_ (.B(_0421_),
    .C(_0438_),
    .A(_0420_),
    .Y(_0440_),
    .D(_0439_));
 sg13g2_xnor2_1 _1093_ (.Y(_0441_),
    .A(net453),
    .B(_0423_));
 sg13g2_and2_1 _1094_ (.A(net436),
    .B(_0400_),
    .X(_0442_));
 sg13g2_nor3_1 _1095_ (.A(\ltc.frm_counter[5] ),
    .B(net4),
    .C(net3),
    .Y(_0443_));
 sg13g2_xnor2_1 _1096_ (.Y(_0444_),
    .A(net466),
    .B(_0406_));
 sg13g2_nand4_1 _1097_ (.B(_0442_),
    .C(_0443_),
    .A(_0441_),
    .Y(_0445_),
    .D(_0444_));
 sg13g2_a21o_1 _1098_ (.A2(_0409_),
    .A1(net461),
    .B1(net471),
    .X(_0446_));
 sg13g2_nor4_1 _1099_ (.A(_0436_),
    .B(_0440_),
    .C(_0445_),
    .D(_0446_),
    .Y(_0447_));
 sg13g2_nand4_1 _1100_ (.B(_0405_),
    .C(_0425_),
    .A(_0207_),
    .Y(_0448_),
    .D(_0446_));
 sg13g2_nor4_1 _1101_ (.A(\ltc.frm_counter[13] ),
    .B(\ltc.frm_counter[15] ),
    .C(_0420_),
    .D(_0448_),
    .Y(_0449_));
 sg13g2_o21ai_1 _1102_ (.B1(_0435_),
    .Y(_0450_),
    .A1(_0447_),
    .A2(_0449_));
 sg13g2_a21oi_2 _1103_ (.B1(_0417_),
    .Y(_0451_),
    .A2(_0450_),
    .A1(_0430_));
 sg13g2_a21o_2 _1104_ (.A2(_0450_),
    .A1(_0430_),
    .B1(_0417_),
    .X(_0452_));
 sg13g2_nand2_1 _1105_ (.Y(_0453_),
    .A(net174),
    .B(net123));
 sg13g2_nor2_1 _1106_ (.A(net228),
    .B(net120),
    .Y(_0081_));
 sg13g2_nor2_1 _1107_ (.A(_0192_),
    .B(_0205_),
    .Y(_0454_));
 sg13g2_nor2_1 _1108_ (.A(net120),
    .B(_0454_),
    .Y(_0082_));
 sg13g2_and3_1 _1109_ (.X(_0455_),
    .A(net260),
    .B(net228),
    .C(net428));
 sg13g2_a21oi_1 _1110_ (.A1(net228),
    .A2(\ltc.frm_counter[1] ),
    .Y(_0456_),
    .B1(net260));
 sg13g2_nor3_1 _1111_ (.A(net120),
    .B(_0455_),
    .C(net261),
    .Y(_0083_));
 sg13g2_o21ai_1 _1112_ (.B1(_0401_),
    .Y(_0457_),
    .A1(net450),
    .A2(_0455_));
 sg13g2_nor2_1 _1113_ (.A(net120),
    .B(_0457_),
    .Y(_0084_));
 sg13g2_nor2_1 _1114_ (.A(net436),
    .B(_0400_),
    .Y(_0458_));
 sg13g2_nor3_1 _1115_ (.A(_0442_),
    .B(net121),
    .C(net437),
    .Y(_0085_));
 sg13g2_nor2_1 _1116_ (.A(net425),
    .B(_0442_),
    .Y(_0459_));
 sg13g2_nor3_1 _1117_ (.A(_0423_),
    .B(net121),
    .C(net426),
    .Y(_0086_));
 sg13g2_nor2_1 _1118_ (.A(_0441_),
    .B(net121),
    .Y(_0087_));
 sg13g2_nor2_1 _1119_ (.A(_0439_),
    .B(net122),
    .Y(_0088_));
 sg13g2_nor2b_1 _1120_ (.A(net120),
    .B_N(_0444_),
    .Y(_0089_));
 sg13g2_nor2_1 _1121_ (.A(_0438_),
    .B(net122),
    .Y(_0090_));
 sg13g2_nor2_1 _1122_ (.A(net458),
    .B(net120),
    .Y(_0091_));
 sg13g2_nor3_1 _1123_ (.A(_0408_),
    .B(net400),
    .C(net120),
    .Y(_0092_));
 sg13g2_nor2_1 _1124_ (.A(_0420_),
    .B(net120),
    .Y(_0093_));
 sg13g2_and4_1 _1125_ (.A(net174),
    .B(_0410_),
    .C(_0421_),
    .D(net123),
    .X(_0094_));
 sg13g2_and4_1 _1126_ (.A(net174),
    .B(_0411_),
    .C(net472),
    .D(_0452_),
    .X(_0095_));
 sg13g2_nor2_1 _1127_ (.A(net460),
    .B(net121),
    .Y(_0096_));
 sg13g2_nor2_1 _1128_ (.A(net465),
    .B(net121),
    .Y(_0097_));
 sg13g2_and3_1 _1129_ (.X(_0098_),
    .A(net176),
    .B(_0418_),
    .C(net123));
 sg13g2_nor2_1 _1130_ (.A(net455),
    .B(net121),
    .Y(_0099_));
 sg13g2_and4_1 _1131_ (.A(\ltc.frm_counter[17] ),
    .B(\ltc.frm_counter[18] ),
    .C(net265),
    .D(_0413_),
    .X(_0460_));
 sg13g2_nor2b_1 _1132_ (.A(net265),
    .B_N(_0415_),
    .Y(_0461_));
 sg13g2_nor3_1 _1133_ (.A(net121),
    .B(_0460_),
    .C(net266),
    .Y(_0100_));
 sg13g2_xnor2_1 _1134_ (.Y(_0462_),
    .A(net405),
    .B(_0460_));
 sg13g2_nor2_1 _1135_ (.A(net121),
    .B(net406),
    .Y(_0101_));
 sg13g2_and3_1 _1136_ (.X(_0463_),
    .A(\ltc.frm_counter[20] ),
    .B(net235),
    .C(_0460_));
 sg13g2_a21oi_1 _1137_ (.A1(\ltc.frm_counter[20] ),
    .A2(_0460_),
    .Y(_0464_),
    .B1(net235));
 sg13g2_nor3_1 _1138_ (.A(net122),
    .B(_0463_),
    .C(net236),
    .Y(_0102_));
 sg13g2_nor2_1 _1139_ (.A(net377),
    .B(_0463_),
    .Y(_0465_));
 sg13g2_and2_1 _1140_ (.A(net377),
    .B(_0463_),
    .X(_0466_));
 sg13g2_nor3_1 _1141_ (.A(net122),
    .B(net378),
    .C(_0466_),
    .Y(_0103_));
 sg13g2_nor2_1 _1142_ (.A(net337),
    .B(_0466_),
    .Y(_0467_));
 sg13g2_and2_1 _1143_ (.A(net337),
    .B(_0466_),
    .X(_0468_));
 sg13g2_nor3_1 _1144_ (.A(net122),
    .B(net338),
    .C(_0468_),
    .Y(_0104_));
 sg13g2_nand2_1 _1145_ (.Y(_0469_),
    .A(net170),
    .B(_0395_));
 sg13g2_nand2_1 _1146_ (.Y(_0470_),
    .A(net430),
    .B(_0397_));
 sg13g2_xnor2_1 _1147_ (.Y(_0471_),
    .A(net430),
    .B(_0397_));
 sg13g2_nor2_1 _1148_ (.A(_0469_),
    .B(net431),
    .Y(_0105_));
 sg13g2_xnor2_1 _1149_ (.Y(_0472_),
    .A(_0150_),
    .B(_0470_));
 sg13g2_nor2_1 _1150_ (.A(_0469_),
    .B(_0472_),
    .Y(_0106_));
 sg13g2_or2_1 _1151_ (.X(_0473_),
    .B(_0469_),
    .A(_0397_));
 sg13g2_and2_1 _1152_ (.A(net416),
    .B(_0393_),
    .X(_0474_));
 sg13g2_nor2_1 _1153_ (.A(net416),
    .B(_0393_),
    .Y(_0475_));
 sg13g2_nor3_1 _1154_ (.A(_0473_),
    .B(_0474_),
    .C(net417),
    .Y(_0107_));
 sg13g2_nand2_1 _1155_ (.Y(_0476_),
    .A(net441),
    .B(_0474_));
 sg13g2_xnor2_1 _1156_ (.Y(_0477_),
    .A(net441),
    .B(_0474_));
 sg13g2_nor2_1 _1157_ (.A(_0473_),
    .B(_0477_),
    .Y(_0108_));
 sg13g2_xor2_1 _1158_ (.B(_0476_),
    .A(net374),
    .X(_0478_));
 sg13g2_nor2_1 _1159_ (.A(_0473_),
    .B(_0478_),
    .Y(_0109_));
 sg13g2_nand2_1 _1160_ (.Y(_0479_),
    .A(net392),
    .B(net388));
 sg13g2_nor3_1 _1161_ (.A(net413),
    .B(net424),
    .C(_0479_),
    .Y(_0480_));
 sg13g2_and2_1 _1162_ (.A(net407),
    .B(_0480_),
    .X(_0481_));
 sg13g2_nand2_1 _1163_ (.Y(_0482_),
    .A(net170),
    .B(_0392_));
 sg13g2_nor2_1 _1164_ (.A(net407),
    .B(_0480_),
    .Y(_0483_));
 sg13g2_nor3_1 _1165_ (.A(_0481_),
    .B(_0482_),
    .C(net408),
    .Y(_0110_));
 sg13g2_nor2_1 _1166_ (.A(net429),
    .B(_0481_),
    .Y(_0484_));
 sg13g2_and2_1 _1167_ (.A(net429),
    .B(_0481_),
    .X(_0485_));
 sg13g2_nor3_1 _1168_ (.A(_0482_),
    .B(_0484_),
    .C(_0485_),
    .Y(_0111_));
 sg13g2_xnor2_1 _1169_ (.Y(_0486_),
    .A(net402),
    .B(_0485_));
 sg13g2_nor2_1 _1170_ (.A(_0482_),
    .B(net403),
    .Y(_0112_));
 sg13g2_nand3b_1 _1171_ (.B(net421),
    .C(net410),
    .Y(_0487_),
    .A_N(net393));
 sg13g2_nor2_1 _1172_ (.A(_0149_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_nand2b_2 _1173_ (.Y(_0489_),
    .B(net171),
    .A_N(_0480_));
 sg13g2_and2_1 _1174_ (.A(_0149_),
    .B(_0487_),
    .X(_0490_));
 sg13g2_nor3_1 _1175_ (.A(_0488_),
    .B(_0489_),
    .C(_0490_),
    .Y(_0113_));
 sg13g2_and2_1 _1176_ (.A(net388),
    .B(_0488_),
    .X(_0491_));
 sg13g2_nor2_1 _1177_ (.A(net388),
    .B(_0488_),
    .Y(_0492_));
 sg13g2_nor3_1 _1178_ (.A(_0489_),
    .B(_0491_),
    .C(net389),
    .Y(_0114_));
 sg13g2_nand2_1 _1179_ (.Y(_0493_),
    .A(net413),
    .B(_0491_));
 sg13g2_xnor2_1 _1180_ (.Y(_0494_),
    .A(net413),
    .B(_0491_));
 sg13g2_nor2_1 _1181_ (.A(_0489_),
    .B(net414),
    .Y(_0115_));
 sg13g2_xor2_1 _1182_ (.B(_0493_),
    .A(net392),
    .X(_0495_));
 sg13g2_nor2_1 _1183_ (.A(_0489_),
    .B(_0495_),
    .Y(_0116_));
 sg13g2_nand2_1 _1184_ (.Y(_0496_),
    .A(\ltc.sec_u[3] ),
    .B(net418));
 sg13g2_nor3_1 _1185_ (.A(net433),
    .B(\ltc.sec_u[0] ),
    .C(_0496_),
    .Y(_0497_));
 sg13g2_and2_1 _1186_ (.A(net393),
    .B(_0497_),
    .X(_0498_));
 sg13g2_nand2_1 _1187_ (.Y(_0499_),
    .A(net173),
    .B(_0487_));
 sg13g2_nor2_1 _1188_ (.A(net393),
    .B(_0497_),
    .Y(_0500_));
 sg13g2_nor3_1 _1189_ (.A(_0498_),
    .B(_0499_),
    .C(net394),
    .Y(_0117_));
 sg13g2_nor2_1 _1190_ (.A(net421),
    .B(_0498_),
    .Y(_0501_));
 sg13g2_and2_1 _1191_ (.A(net421),
    .B(_0498_),
    .X(_0502_));
 sg13g2_nor3_1 _1192_ (.A(_0499_),
    .B(net422),
    .C(_0502_),
    .Y(_0118_));
 sg13g2_xnor2_1 _1193_ (.Y(_0503_),
    .A(net410),
    .B(_0502_));
 sg13g2_nor2_1 _1194_ (.A(_0499_),
    .B(net411),
    .Y(_0119_));
 sg13g2_nor2_1 _1195_ (.A(net438),
    .B(net294),
    .Y(_0504_));
 sg13g2_nor2b_1 _1196_ (.A(\ltc.frm_u[1] ),
    .B_N(\ltc.frm_u[0] ),
    .Y(_0505_));
 sg13g2_a22oi_1 _1197_ (.Y(_0506_),
    .B1(_0505_),
    .B2(_0207_),
    .A2(_0504_),
    .A1(_0333_));
 sg13g2_nand2_1 _1198_ (.Y(_0507_),
    .A(\ltc.frm_u[2] ),
    .B(_0147_));
 sg13g2_nand4_1 _1199_ (.B(\ltc.frm_d[0] ),
    .C(_0334_),
    .A(_0145_),
    .Y(_0508_),
    .D(_0504_));
 sg13g2_o21ai_1 _1200_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0506_),
    .A2(_0507_));
 sg13g2_nand3_1 _1201_ (.B(net375),
    .C(_0509_),
    .A(_0144_),
    .Y(_0510_));
 sg13g2_nor2_1 _1202_ (.A(_0148_),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_nand2b_2 _1203_ (.Y(_0512_),
    .B(net173),
    .A_N(_0497_));
 sg13g2_a21oi_1 _1204_ (.A1(_0148_),
    .A2(_0510_),
    .Y(_0513_),
    .B1(_0512_));
 sg13g2_nor2b_1 _1205_ (.A(_0511_),
    .B_N(_0513_),
    .Y(_0120_));
 sg13g2_nor2_1 _1206_ (.A(net418),
    .B(_0511_),
    .Y(_0514_));
 sg13g2_and2_1 _1207_ (.A(net418),
    .B(_0511_),
    .X(_0515_));
 sg13g2_nor3_1 _1208_ (.A(_0512_),
    .B(net419),
    .C(_0515_),
    .Y(_0121_));
 sg13g2_nand2_1 _1209_ (.Y(_0516_),
    .A(net433),
    .B(_0515_));
 sg13g2_xnor2_1 _1210_ (.Y(_0517_),
    .A(net433),
    .B(_0515_));
 sg13g2_nor2_1 _1211_ (.A(_0512_),
    .B(net434),
    .Y(_0122_));
 sg13g2_xor2_1 _1212_ (.B(_0516_),
    .A(net448),
    .X(_0518_));
 sg13g2_nor2_1 _1213_ (.A(_0512_),
    .B(_0518_),
    .Y(_0123_));
 sg13g2_nand2_1 _1214_ (.Y(_0519_),
    .A(net174),
    .B(_0510_));
 sg13g2_nand4_1 _1215_ (.B(_0145_),
    .C(net438),
    .A(net444),
    .Y(_0520_),
    .D(_0146_));
 sg13g2_and2_1 _1216_ (.A(_0147_),
    .B(_0520_),
    .X(_0521_));
 sg13g2_nor2_1 _1217_ (.A(_0147_),
    .B(_0520_),
    .Y(_0522_));
 sg13g2_nor3_1 _1218_ (.A(_0519_),
    .B(_0521_),
    .C(_0522_),
    .Y(_0124_));
 sg13g2_xnor2_1 _1219_ (.Y(_0523_),
    .A(net375),
    .B(_0522_));
 sg13g2_nor2_1 _1220_ (.A(_0519_),
    .B(net376),
    .Y(_0125_));
 sg13g2_nand3_1 _1221_ (.B(_0510_),
    .C(_0520_),
    .A(net123),
    .Y(_0524_));
 sg13g2_o21ai_1 _1222_ (.B1(net174),
    .Y(_0525_),
    .A1(net294),
    .A2(_0451_));
 sg13g2_a21oi_1 _1223_ (.A1(net294),
    .A2(_0524_),
    .Y(_0126_),
    .B1(_0525_));
 sg13g2_nand4_1 _1224_ (.B(net123),
    .C(_0510_),
    .A(net438),
    .Y(_0526_),
    .D(_0520_));
 sg13g2_nand2_1 _1225_ (.Y(_0527_),
    .A(net438),
    .B(net294));
 sg13g2_nand3b_1 _1226_ (.B(_0527_),
    .C(_0451_),
    .Y(_0528_),
    .A_N(_0504_));
 sg13g2_a21oi_1 _1227_ (.A1(_0526_),
    .A2(_0528_),
    .Y(_0127_),
    .B1(net168));
 sg13g2_nand4_1 _1228_ (.B(net123),
    .C(_0510_),
    .A(net390),
    .Y(_0529_),
    .D(_0520_));
 sg13g2_nand2_1 _1229_ (.Y(_0530_),
    .A(_0145_),
    .B(_0527_));
 sg13g2_nand3_1 _1230_ (.B(net438),
    .C(net294),
    .A(net390),
    .Y(_0531_));
 sg13g2_nand2_1 _1231_ (.Y(_0532_),
    .A(_0451_),
    .B(_0531_));
 sg13g2_nand3_1 _1232_ (.B(_0530_),
    .C(_0531_),
    .A(_0451_),
    .Y(_0533_));
 sg13g2_a21oi_1 _1233_ (.A1(_0529_),
    .A2(_0533_),
    .Y(_0128_),
    .B1(net168));
 sg13g2_a21oi_1 _1234_ (.A1(net123),
    .A2(_0520_),
    .Y(_0534_),
    .B1(_0144_));
 sg13g2_or2_1 _1235_ (.X(_0535_),
    .B(_0531_),
    .A(net123));
 sg13g2_a221oi_1 _1236_ (.B2(_0144_),
    .C1(net168),
    .B1(_0535_),
    .A1(_0532_),
    .Y(_0129_),
    .A2(_0534_));
 sg13g2_nor2_1 _1237_ (.A(\ltc.bit_clk ),
    .B(\ltc.output_buffer[79] ),
    .Y(_0536_));
 sg13g2_nor2_1 _1238_ (.A(_0177_),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_o21ai_1 _1239_ (.B1(net173),
    .Y(_0538_),
    .A1(net229),
    .A2(_0537_));
 sg13g2_a21oi_1 _1240_ (.A1(net229),
    .A2(_0537_),
    .Y(_0130_),
    .B1(_0538_));
 sg13g2_and2_1 _1241_ (.A(net383),
    .B(net227),
    .X(_0539_));
 sg13g2_and4_1 _1242_ (.A(net273),
    .B(\ltc.bit_counter[2] ),
    .C(net383),
    .D(net227),
    .X(_0540_));
 sg13g2_nand2_1 _1243_ (.Y(_0541_),
    .A(\ltc.bit_counter[5] ),
    .B(\ltc.bit_counter[4] ));
 sg13g2_and3_2 _1244_ (.X(_0542_),
    .A(net268),
    .B(net442),
    .C(_0540_));
 sg13g2_and3_1 _1245_ (.X(_0543_),
    .A(\ltc.bit_counter[6] ),
    .B(net285),
    .C(_0542_));
 sg13g2_and4_1 _1246_ (.A(\ltc.bit_counter[6] ),
    .B(net285),
    .C(net396),
    .D(_0542_),
    .X(_0544_));
 sg13g2_nand3_1 _1247_ (.B(net452),
    .C(_0544_),
    .A(net446),
    .Y(_0545_));
 sg13g2_xor2_1 _1248_ (.B(_0545_),
    .A(net323),
    .X(_0546_));
 sg13g2_a21o_1 _1249_ (.A2(_0544_),
    .A1(net446),
    .B1(net452),
    .X(_0547_));
 sg13g2_nand2_1 _1250_ (.Y(_0548_),
    .A(_0545_),
    .B(_0547_));
 sg13g2_nand3_1 _1251_ (.B(\ltc.bit_counter[9] ),
    .C(_0207_),
    .A(\ltc.bit_counter[2] ),
    .Y(_0549_));
 sg13g2_nor3_1 _1252_ (.A(\ltc.bit_counter[6] ),
    .B(_0541_),
    .C(_0549_),
    .Y(_0550_));
 sg13g2_nor3_1 _1253_ (.A(\ltc.bit_counter[2] ),
    .B(_0154_),
    .C(\ltc.bit_counter[9] ),
    .Y(_0551_));
 sg13g2_and2_1 _1254_ (.A(_0173_),
    .B(_0334_),
    .X(_0552_));
 sg13g2_a21oi_1 _1255_ (.A1(_0551_),
    .A2(_0552_),
    .Y(_0553_),
    .B1(_0550_));
 sg13g2_nand3_1 _1256_ (.B(\ltc.bit_counter[8] ),
    .C(_0539_),
    .A(\ltc.bit_counter[7] ),
    .Y(_0554_));
 sg13g2_nor3_1 _1257_ (.A(\ltc.bit_counter[3] ),
    .B(_0553_),
    .C(_0554_),
    .Y(_0555_));
 sg13g2_xnor2_1 _1258_ (.Y(_0556_),
    .A(net456),
    .B(_0539_));
 sg13g2_nand3_1 _1259_ (.B(_0175_),
    .C(_0333_),
    .A(_0174_),
    .Y(_0557_));
 sg13g2_nor4_1 _1260_ (.A(\ltc.bit_counter[3] ),
    .B(_0541_),
    .C(_0556_),
    .D(_0557_),
    .Y(_0558_));
 sg13g2_mux2_1 _1261_ (.A0(_0558_),
    .A1(_0555_),
    .S(_0548_),
    .X(_0559_));
 sg13g2_nor2b_1 _1262_ (.A(_0546_),
    .B_N(_0559_),
    .Y(_0560_));
 sg13g2_nand2b_1 _1263_ (.Y(_0561_),
    .B(net173),
    .A_N(_0560_));
 sg13g2_nor2_1 _1264_ (.A(net227),
    .B(net119),
    .Y(_0131_));
 sg13g2_nor3_1 _1265_ (.A(_0171_),
    .B(_0539_),
    .C(net119),
    .Y(_0132_));
 sg13g2_nor2_1 _1266_ (.A(_0556_),
    .B(net118),
    .Y(_0133_));
 sg13g2_a21oi_1 _1267_ (.A1(\ltc.bit_counter[2] ),
    .A2(_0539_),
    .Y(_0562_),
    .B1(net273));
 sg13g2_nor3_1 _1268_ (.A(_0540_),
    .B(net119),
    .C(net274),
    .Y(_0134_));
 sg13g2_xnor2_1 _1269_ (.Y(_0563_),
    .A(net442),
    .B(_0540_));
 sg13g2_nor2_1 _1270_ (.A(net118),
    .B(net443),
    .Y(_0135_));
 sg13g2_a21oi_1 _1271_ (.A1(\ltc.bit_counter[4] ),
    .A2(_0540_),
    .Y(_0564_),
    .B1(net268));
 sg13g2_nor3_1 _1272_ (.A(_0542_),
    .B(net119),
    .C(net269),
    .Y(_0136_));
 sg13g2_xnor2_1 _1273_ (.Y(_0565_),
    .A(net451),
    .B(_0542_));
 sg13g2_nor2_1 _1274_ (.A(net118),
    .B(_0565_),
    .Y(_0137_));
 sg13g2_a21oi_1 _1275_ (.A1(\ltc.bit_counter[6] ),
    .A2(_0542_),
    .Y(_0566_),
    .B1(net285));
 sg13g2_nor3_1 _1276_ (.A(_0543_),
    .B(net118),
    .C(net286),
    .Y(_0138_));
 sg13g2_nor2_1 _1277_ (.A(net396),
    .B(_0543_),
    .Y(_0567_));
 sg13g2_nor3_1 _1278_ (.A(_0544_),
    .B(net118),
    .C(net397),
    .Y(_0139_));
 sg13g2_xnor2_1 _1279_ (.Y(_0568_),
    .A(net446),
    .B(_0544_));
 sg13g2_nor2_1 _1280_ (.A(net118),
    .B(net447),
    .Y(_0140_));
 sg13g2_nor2_1 _1281_ (.A(_0548_),
    .B(net118),
    .Y(_0141_));
 sg13g2_nor2_1 _1282_ (.A(_0546_),
    .B(net118),
    .Y(_0142_));
 sg13g2_o21ai_1 _1283_ (.B1(net176),
    .Y(_0569_),
    .A1(net231),
    .A2(_0560_));
 sg13g2_a21oi_1 _1284_ (.A1(net231),
    .A2(_0560_),
    .Y(_0143_),
    .B1(_0569_));
 sg13g2_dfrbpq_1 _1285_ (.RESET_B(net105),
    .D(_0000_),
    .Q(\ltc.output_buffer[0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1286_ (.RESET_B(net89),
    .D(_0001_),
    .Q(\ltc.output_buffer[1] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1287_ (.RESET_B(net88),
    .D(net239),
    .Q(\ltc.output_buffer[2] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1288_ (.RESET_B(net87),
    .D(net254),
    .Q(\ltc.output_buffer[3] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1289_ (.RESET_B(net86),
    .D(net257),
    .Q(\ltc.output_buffer[4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1290_ (.RESET_B(net85),
    .D(net241),
    .Q(\ltc.output_buffer[5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1291_ (.RESET_B(net84),
    .D(net234),
    .Q(\ltc.output_buffer[6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1292_ (.RESET_B(net83),
    .D(_0007_),
    .Q(\ltc.output_buffer[7] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1293_ (.RESET_B(net82),
    .D(net250),
    .Q(\ltc.output_buffer[8] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1294_ (.RESET_B(net81),
    .D(net248),
    .Q(\ltc.output_buffer[9] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1295_ (.RESET_B(net80),
    .D(_0010_),
    .Q(\ltc.output_buffer[10] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1296_ (.RESET_B(net79),
    .D(net244),
    .Q(\ltc.output_buffer[11] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1297_ (.RESET_B(net78),
    .D(_0012_),
    .Q(\ltc.output_buffer[12] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1298_ (.RESET_B(net77),
    .D(net246),
    .Q(\ltc.output_buffer[13] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1299_ (.RESET_B(net76),
    .D(_0014_),
    .Q(\ltc.output_buffer[14] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1300_ (.RESET_B(net75),
    .D(_0015_),
    .Q(\ltc.output_buffer[15] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1301_ (.RESET_B(net74),
    .D(_0016_),
    .Q(\ltc.output_buffer[16] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1302_ (.RESET_B(net73),
    .D(_0017_),
    .Q(\ltc.output_buffer[17] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1303_ (.RESET_B(net72),
    .D(_0018_),
    .Q(\ltc.output_buffer[18] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1304_ (.RESET_B(net71),
    .D(_0019_),
    .Q(\ltc.output_buffer[19] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1305_ (.RESET_B(net70),
    .D(net329),
    .Q(\ltc.output_buffer[20] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _1306_ (.RESET_B(net69),
    .D(_0021_),
    .Q(\ltc.output_buffer[21] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1307_ (.RESET_B(net68),
    .D(_0022_),
    .Q(\ltc.output_buffer[22] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1308_ (.RESET_B(net67),
    .D(net277),
    .Q(\ltc.output_buffer[23] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1309_ (.RESET_B(net66),
    .D(_0024_),
    .Q(\ltc.output_buffer[24] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1310_ (.RESET_B(net65),
    .D(_0025_),
    .Q(\ltc.output_buffer[25] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1311_ (.RESET_B(net64),
    .D(_0026_),
    .Q(\ltc.output_buffer[26] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1312_ (.RESET_B(net63),
    .D(_0027_),
    .Q(\ltc.output_buffer[27] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1313_ (.RESET_B(net62),
    .D(_0028_),
    .Q(\ltc.output_buffer[28] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1314_ (.RESET_B(net61),
    .D(net316),
    .Q(\ltc.output_buffer[29] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1315_ (.RESET_B(net60),
    .D(net289),
    .Q(\ltc.output_buffer[30] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1316_ (.RESET_B(net59),
    .D(net291),
    .Q(\ltc.output_buffer[31] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1317_ (.RESET_B(net58),
    .D(_0032_),
    .Q(\ltc.output_buffer[32] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1318_ (.RESET_B(net57),
    .D(_0033_),
    .Q(\ltc.output_buffer[33] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1319_ (.RESET_B(net56),
    .D(_0034_),
    .Q(\ltc.output_buffer[34] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1320_ (.RESET_B(net55),
    .D(_0035_),
    .Q(\ltc.output_buffer[35] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1321_ (.RESET_B(net54),
    .D(_0036_),
    .Q(\ltc.output_buffer[36] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1322_ (.RESET_B(net53),
    .D(net293),
    .Q(\ltc.output_buffer[37] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1323_ (.RESET_B(net52),
    .D(net318),
    .Q(\ltc.output_buffer[38] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1324_ (.RESET_B(net51),
    .D(net306),
    .Q(\ltc.output_buffer[39] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1325_ (.RESET_B(net50),
    .D(_0040_),
    .Q(\ltc.output_buffer[40] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1326_ (.RESET_B(net49),
    .D(_0041_),
    .Q(\ltc.output_buffer[41] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1327_ (.RESET_B(net48),
    .D(_0042_),
    .Q(\ltc.output_buffer[42] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _1328_ (.RESET_B(net47),
    .D(_0043_),
    .Q(\ltc.output_buffer[43] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1329_ (.RESET_B(net46),
    .D(_0044_),
    .Q(\ltc.output_buffer[44] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1330_ (.RESET_B(net45),
    .D(net325),
    .Q(\ltc.output_buffer[45] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1331_ (.RESET_B(net44),
    .D(net300),
    .Q(\ltc.output_buffer[46] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _1332_ (.RESET_B(net43),
    .D(net302),
    .Q(\ltc.output_buffer[47] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1333_ (.RESET_B(net42),
    .D(_0048_),
    .Q(\ltc.output_buffer[48] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1334_ (.RESET_B(net41),
    .D(_0049_),
    .Q(\ltc.output_buffer[49] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1335_ (.RESET_B(net40),
    .D(_0050_),
    .Q(\ltc.output_buffer[50] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1336_ (.RESET_B(net39),
    .D(_0051_),
    .Q(\ltc.output_buffer[51] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1337_ (.RESET_B(net38),
    .D(net264),
    .Q(\ltc.output_buffer[52] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1338_ (.RESET_B(net37),
    .D(net279),
    .Q(\ltc.output_buffer[53] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1339_ (.RESET_B(net36),
    .D(net343),
    .Q(\ltc.output_buffer[54] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1340_ (.RESET_B(net35),
    .D(net345),
    .Q(\ltc.output_buffer[55] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1341_ (.RESET_B(net34),
    .D(_0056_),
    .Q(\ltc.output_buffer[56] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _1342_ (.RESET_B(net33),
    .D(_0057_),
    .Q(\ltc.output_buffer[57] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1343_ (.RESET_B(net32),
    .D(_0058_),
    .Q(\ltc.output_buffer[58] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1344_ (.RESET_B(net31),
    .D(_0059_),
    .Q(\ltc.output_buffer[59] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1345_ (.RESET_B(net30),
    .D(net365),
    .Q(\ltc.output_buffer[60] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1346_ (.RESET_B(net29),
    .D(net357),
    .Q(\ltc.output_buffer[61] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1347_ (.RESET_B(net28),
    .D(net336),
    .Q(\ltc.output_buffer[62] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1348_ (.RESET_B(net27),
    .D(net296),
    .Q(\ltc.output_buffer[63] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1349_ (.RESET_B(net26),
    .D(_0064_),
    .Q(\ltc.output_buffer[64] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1350_ (.RESET_B(net25),
    .D(_0065_),
    .Q(\ltc.output_buffer[65] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1351_ (.RESET_B(net24),
    .D(_0066_),
    .Q(\ltc.output_buffer[66] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1352_ (.RESET_B(net23),
    .D(_0067_),
    .Q(\ltc.output_buffer[67] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1353_ (.RESET_B(net225),
    .D(_0068_),
    .Q(\ltc.output_buffer[68] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1354_ (.RESET_B(net224),
    .D(_0069_),
    .Q(\ltc.output_buffer[69] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1355_ (.RESET_B(net223),
    .D(net281),
    .Q(\ltc.output_buffer[70] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1356_ (.RESET_B(net222),
    .D(net298),
    .Q(\ltc.output_buffer[71] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1357_ (.RESET_B(net221),
    .D(_0072_),
    .Q(\ltc.output_buffer[72] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1358_ (.RESET_B(net220),
    .D(_0073_),
    .Q(\ltc.output_buffer[73] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1359_ (.RESET_B(net219),
    .D(_0074_),
    .Q(\ltc.output_buffer[74] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1360_ (.RESET_B(net218),
    .D(_0075_),
    .Q(\ltc.output_buffer[75] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _1361_ (.RESET_B(net217),
    .D(net272),
    .Q(\ltc.output_buffer[76] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1362_ (.RESET_B(net216),
    .D(net284),
    .Q(\ltc.output_buffer[77] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1363_ (.RESET_B(net215),
    .D(net353),
    .Q(\ltc.output_buffer[78] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1364_ (.RESET_B(net214),
    .D(net310),
    .Q(\ltc.output_buffer[79] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1365_ (.RESET_B(net213),
    .D(_0080_),
    .Q(\ltc.hrs_u[0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1366_ (.RESET_B(net211),
    .D(_0081_),
    .Q(\ltc.frm_counter[0] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1367_ (.RESET_B(net210),
    .D(_0082_),
    .Q(\ltc.frm_counter[1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1368_ (.RESET_B(net209),
    .D(net262),
    .Q(\ltc.frm_counter[2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1369_ (.RESET_B(net208),
    .D(_0084_),
    .Q(\ltc.frm_counter[3] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1370_ (.RESET_B(net207),
    .D(_0085_),
    .Q(\ltc.frm_counter[4] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1371_ (.RESET_B(net206),
    .D(net427),
    .Q(\ltc.frm_counter[5] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1372_ (.RESET_B(net205),
    .D(_0087_),
    .Q(\ltc.frm_counter[6] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1373_ (.RESET_B(net204),
    .D(_0088_),
    .Q(\ltc.frm_counter[7] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1374_ (.RESET_B(net203),
    .D(_0089_),
    .Q(\ltc.frm_counter[8] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1375_ (.RESET_B(net202),
    .D(_0090_),
    .Q(\ltc.frm_counter[9] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1376_ (.RESET_B(net201),
    .D(_0091_),
    .Q(\ltc.frm_counter[10] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1377_ (.RESET_B(net200),
    .D(net401),
    .Q(\ltc.frm_counter[11] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1378_ (.RESET_B(net199),
    .D(_0093_),
    .Q(\ltc.frm_counter[12] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1379_ (.RESET_B(net198),
    .D(net462),
    .Q(\ltc.frm_counter[13] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1380_ (.RESET_B(net197),
    .D(_0095_),
    .Q(\ltc.frm_counter[14] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1381_ (.RESET_B(net196),
    .D(_0096_),
    .Q(\ltc.frm_counter[15] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1382_ (.RESET_B(net195),
    .D(_0097_),
    .Q(\ltc.frm_counter[16] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1383_ (.RESET_B(net194),
    .D(_0098_),
    .Q(\ltc.frm_counter[17] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1384_ (.RESET_B(net193),
    .D(_0099_),
    .Q(\ltc.frm_counter[18] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1385_ (.RESET_B(net192),
    .D(net267),
    .Q(\ltc.frm_counter[19] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1386_ (.RESET_B(net191),
    .D(_0101_),
    .Q(\ltc.frm_counter[20] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net190),
    .D(net237),
    .Q(\ltc.frm_counter[21] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1388_ (.RESET_B(net189),
    .D(net379),
    .Q(\ltc.frm_counter[22] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1389_ (.RESET_B(net188),
    .D(net339),
    .Q(\ltc.frm_counter[23] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1390_ (.RESET_B(net187),
    .D(net432),
    .Q(\ltc.hrs_d[0] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net185),
    .D(_0106_),
    .Q(\ltc.hrs_d[1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1392_ (.RESET_B(net183),
    .D(_0107_),
    .Q(\ltc.hrs_u[1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1393_ (.RESET_B(net181),
    .D(_0108_),
    .Q(\ltc.hrs_u[2] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1394_ (.RESET_B(net179),
    .D(_0109_),
    .Q(\ltc.hrs_u[3] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1395_ (.RESET_B(net177),
    .D(net409),
    .Q(\ltc.min_d[0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1396_ (.RESET_B(net116),
    .D(_0111_),
    .Q(\ltc.min_d[1] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1397_ (.RESET_B(net114),
    .D(net404),
    .Q(\ltc.min_d[2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1398_ (.RESET_B(net112),
    .D(_0113_),
    .Q(\ltc.min_u[0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _1399_ (.RESET_B(net110),
    .D(_0114_),
    .Q(\ltc.min_u[1] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _1400_ (.RESET_B(net108),
    .D(net415),
    .Q(\ltc.min_u[2] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _1401_ (.RESET_B(net106),
    .D(_0116_),
    .Q(\ltc.min_u[3] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1402_ (.RESET_B(net104),
    .D(net395),
    .Q(\ltc.sec_d[0] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1403_ (.RESET_B(net102),
    .D(_0118_),
    .Q(\ltc.sec_d[1] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1404_ (.RESET_B(net100),
    .D(net412),
    .Q(\ltc.sec_d[2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1405_ (.RESET_B(net98),
    .D(_0120_),
    .Q(\ltc.sec_u[0] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1406_ (.RESET_B(net96),
    .D(net420),
    .Q(\ltc.sec_u[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1407_ (.RESET_B(net94),
    .D(net435),
    .Q(\ltc.sec_u[2] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1408_ (.RESET_B(net92),
    .D(net449),
    .Q(\ltc.sec_u[3] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1409_ (.RESET_B(net90),
    .D(_0124_),
    .Q(\ltc.frm_d[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1410_ (.RESET_B(net186),
    .D(_0125_),
    .Q(\ltc.frm_d[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1411_ (.RESET_B(net182),
    .D(_0126_),
    .Q(\ltc.frm_u[0] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1412_ (.RESET_B(net178),
    .D(_0127_),
    .Q(\ltc.frm_u[1] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1413_ (.RESET_B(net115),
    .D(net391),
    .Q(\ltc.frm_u[2] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1414_ (.RESET_B(net111),
    .D(net445),
    .Q(\ltc.frm_u[3] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1415_ (.RESET_B(net107),
    .D(net230),
    .Q(\ltc.timecode ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1416_ (.RESET_B(net103),
    .D(_0131_),
    .Q(\ltc.bit_counter[0] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net101),
    .D(_0132_),
    .Q(\ltc.bit_counter[1] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1418_ (.RESET_B(net99),
    .D(_0133_),
    .Q(\ltc.bit_counter[2] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1419_ (.RESET_B(net97),
    .D(net275),
    .Q(\ltc.bit_counter[3] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1420_ (.RESET_B(net95),
    .D(_0135_),
    .Q(\ltc.bit_counter[4] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1421_ (.RESET_B(net93),
    .D(net270),
    .Q(\ltc.bit_counter[5] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1422_ (.RESET_B(net91),
    .D(_0137_),
    .Q(\ltc.bit_counter[6] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1423_ (.RESET_B(net212),
    .D(net287),
    .Q(\ltc.bit_counter[7] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net184),
    .D(net398),
    .Q(\ltc.bit_counter[8] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1425_ (.RESET_B(net180),
    .D(_0140_),
    .Q(\ltc.bit_counter[9] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1426_ (.RESET_B(net117),
    .D(_0141_),
    .Q(\ltc.bit_counter[10] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net113),
    .D(_0142_),
    .Q(\ltc.bit_counter[11] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1428_ (.RESET_B(net109),
    .D(net232),
    .Q(\ltc.bit_clk ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_tiehi _1351__24 (.L_HI(net24));
 sg13g2_tiehi _1350__25 (.L_HI(net25));
 sg13g2_tiehi _1349__26 (.L_HI(net26));
 sg13g2_tiehi _1348__27 (.L_HI(net27));
 sg13g2_tiehi _1347__28 (.L_HI(net28));
 sg13g2_tiehi _1346__29 (.L_HI(net29));
 sg13g2_tiehi _1345__30 (.L_HI(net30));
 sg13g2_tiehi _1344__31 (.L_HI(net31));
 sg13g2_tiehi _1343__32 (.L_HI(net32));
 sg13g2_tiehi _1342__33 (.L_HI(net33));
 sg13g2_tiehi _1341__34 (.L_HI(net34));
 sg13g2_tiehi _1340__35 (.L_HI(net35));
 sg13g2_tiehi _1339__36 (.L_HI(net36));
 sg13g2_tiehi _1338__37 (.L_HI(net37));
 sg13g2_tiehi _1337__38 (.L_HI(net38));
 sg13g2_tiehi _1336__39 (.L_HI(net39));
 sg13g2_tiehi _1335__40 (.L_HI(net40));
 sg13g2_tiehi _1334__41 (.L_HI(net41));
 sg13g2_tiehi _1333__42 (.L_HI(net42));
 sg13g2_tiehi _1332__43 (.L_HI(net43));
 sg13g2_tiehi _1331__44 (.L_HI(net44));
 sg13g2_tiehi _1330__45 (.L_HI(net45));
 sg13g2_tiehi _1329__46 (.L_HI(net46));
 sg13g2_tiehi _1328__47 (.L_HI(net47));
 sg13g2_tiehi _1327__48 (.L_HI(net48));
 sg13g2_tiehi _1326__49 (.L_HI(net49));
 sg13g2_tiehi _1325__50 (.L_HI(net50));
 sg13g2_tiehi _1324__51 (.L_HI(net51));
 sg13g2_tiehi _1323__52 (.L_HI(net52));
 sg13g2_tiehi _1322__53 (.L_HI(net53));
 sg13g2_tiehi _1321__54 (.L_HI(net54));
 sg13g2_tiehi _1320__55 (.L_HI(net55));
 sg13g2_tiehi _1319__56 (.L_HI(net56));
 sg13g2_tiehi _1318__57 (.L_HI(net57));
 sg13g2_tiehi _1317__58 (.L_HI(net58));
 sg13g2_tiehi _1316__59 (.L_HI(net59));
 sg13g2_tiehi _1315__60 (.L_HI(net60));
 sg13g2_tiehi _1314__61 (.L_HI(net61));
 sg13g2_tiehi _1313__62 (.L_HI(net62));
 sg13g2_tiehi _1312__63 (.L_HI(net63));
 sg13g2_tiehi _1311__64 (.L_HI(net64));
 sg13g2_tiehi _1310__65 (.L_HI(net65));
 sg13g2_tiehi _1309__66 (.L_HI(net66));
 sg13g2_tiehi _1308__67 (.L_HI(net67));
 sg13g2_tiehi _1307__68 (.L_HI(net68));
 sg13g2_tiehi _1306__69 (.L_HI(net69));
 sg13g2_tiehi _1305__70 (.L_HI(net70));
 sg13g2_tiehi _1304__71 (.L_HI(net71));
 sg13g2_tiehi _1303__72 (.L_HI(net72));
 sg13g2_tiehi _1302__73 (.L_HI(net73));
 sg13g2_tiehi _1301__74 (.L_HI(net74));
 sg13g2_tiehi _1300__75 (.L_HI(net75));
 sg13g2_tiehi _1299__76 (.L_HI(net76));
 sg13g2_tiehi _1298__77 (.L_HI(net77));
 sg13g2_tiehi _1297__78 (.L_HI(net78));
 sg13g2_tiehi _1296__79 (.L_HI(net79));
 sg13g2_tiehi _1295__80 (.L_HI(net80));
 sg13g2_tiehi _1294__81 (.L_HI(net81));
 sg13g2_tiehi _1293__82 (.L_HI(net82));
 sg13g2_tiehi _1292__83 (.L_HI(net83));
 sg13g2_tiehi _1291__84 (.L_HI(net84));
 sg13g2_tiehi _1290__85 (.L_HI(net85));
 sg13g2_tiehi _1289__86 (.L_HI(net86));
 sg13g2_tiehi _1288__87 (.L_HI(net87));
 sg13g2_tiehi _1287__88 (.L_HI(net88));
 sg13g2_tiehi _1286__89 (.L_HI(net89));
 sg13g2_tiehi _1409__90 (.L_HI(net90));
 sg13g2_tiehi _1422__91 (.L_HI(net91));
 sg13g2_tiehi _1408__92 (.L_HI(net92));
 sg13g2_tiehi _1421__93 (.L_HI(net93));
 sg13g2_tiehi _1407__94 (.L_HI(net94));
 sg13g2_tiehi _1420__95 (.L_HI(net95));
 sg13g2_tiehi _1406__96 (.L_HI(net96));
 sg13g2_tiehi _1419__97 (.L_HI(net97));
 sg13g2_tiehi _1405__98 (.L_HI(net98));
 sg13g2_tiehi _1418__99 (.L_HI(net99));
 sg13g2_tiehi _1404__100 (.L_HI(net100));
 sg13g2_tiehi _1417__101 (.L_HI(net101));
 sg13g2_tiehi _1403__102 (.L_HI(net102));
 sg13g2_tiehi _1416__103 (.L_HI(net103));
 sg13g2_tiehi _1402__104 (.L_HI(net104));
 sg13g2_tiehi _1285__105 (.L_HI(net105));
 sg13g2_tiehi _1401__106 (.L_HI(net106));
 sg13g2_tiehi _1415__107 (.L_HI(net107));
 sg13g2_tiehi _1400__108 (.L_HI(net108));
 sg13g2_tiehi _1428__109 (.L_HI(net109));
 sg13g2_tiehi _1399__110 (.L_HI(net110));
 sg13g2_tiehi _1414__111 (.L_HI(net111));
 sg13g2_tiehi _1398__112 (.L_HI(net112));
 sg13g2_tiehi _1427__113 (.L_HI(net113));
 sg13g2_tiehi _1397__114 (.L_HI(net114));
 sg13g2_tiehi _1413__115 (.L_HI(net115));
 sg13g2_tiehi _1396__116 (.L_HI(net116));
 sg13g2_tiehi _1426__117 (.L_HI(net117));
 sg13g2_tiehi _1395__118 (.L_HI(net177));
 sg13g2_tiehi _1412__119 (.L_HI(net178));
 sg13g2_tiehi _1394__120 (.L_HI(net179));
 sg13g2_tiehi _1425__121 (.L_HI(net180));
 sg13g2_tiehi _1393__122 (.L_HI(net181));
 sg13g2_tiehi _1411__123 (.L_HI(net182));
 sg13g2_tiehi _1392__124 (.L_HI(net183));
 sg13g2_tiehi _1424__125 (.L_HI(net184));
 sg13g2_tiehi _1391__126 (.L_HI(net185));
 sg13g2_tiehi _1410__127 (.L_HI(net186));
 sg13g2_tiehi _1390__128 (.L_HI(net187));
 sg13g2_tiehi _1389__129 (.L_HI(net188));
 sg13g2_tiehi _1388__130 (.L_HI(net189));
 sg13g2_tiehi _1387__131 (.L_HI(net190));
 sg13g2_tiehi _1386__132 (.L_HI(net191));
 sg13g2_tiehi _1385__133 (.L_HI(net192));
 sg13g2_tiehi _1384__134 (.L_HI(net193));
 sg13g2_tiehi _1383__135 (.L_HI(net194));
 sg13g2_tiehi _1382__136 (.L_HI(net195));
 sg13g2_tiehi _1381__137 (.L_HI(net196));
 sg13g2_tiehi _1380__138 (.L_HI(net197));
 sg13g2_tiehi _1379__139 (.L_HI(net198));
 sg13g2_tiehi _1378__140 (.L_HI(net199));
 sg13g2_tiehi _1377__141 (.L_HI(net200));
 sg13g2_tiehi _1376__142 (.L_HI(net201));
 sg13g2_tiehi _1375__143 (.L_HI(net202));
 sg13g2_tiehi _1374__144 (.L_HI(net203));
 sg13g2_tiehi _1373__145 (.L_HI(net204));
 sg13g2_tiehi _1372__146 (.L_HI(net205));
 sg13g2_tiehi _1371__147 (.L_HI(net206));
 sg13g2_tiehi _1370__148 (.L_HI(net207));
 sg13g2_tiehi _1369__149 (.L_HI(net208));
 sg13g2_tiehi _1368__150 (.L_HI(net209));
 sg13g2_tiehi _1367__151 (.L_HI(net210));
 sg13g2_tiehi _1366__152 (.L_HI(net211));
 sg13g2_tiehi _1423__153 (.L_HI(net212));
 sg13g2_tiehi _1365__154 (.L_HI(net213));
 sg13g2_tiehi _1364__155 (.L_HI(net214));
 sg13g2_tiehi _1363__156 (.L_HI(net215));
 sg13g2_tiehi _1362__157 (.L_HI(net216));
 sg13g2_tiehi _1361__158 (.L_HI(net217));
 sg13g2_tiehi _1360__159 (.L_HI(net218));
 sg13g2_tiehi _1359__160 (.L_HI(net219));
 sg13g2_tiehi _1358__161 (.L_HI(net220));
 sg13g2_tiehi _1357__162 (.L_HI(net221));
 sg13g2_tiehi _1356__163 (.L_HI(net222));
 sg13g2_tiehi _1355__164 (.L_HI(net223));
 sg13g2_tiehi _1354__165 (.L_HI(net224));
 sg13g2_tiehi _1353__166 (.L_HI(net225));
 sg13g2_tiehi tt_um_flummer_ltc_167 (.L_HI(net226));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_flummer_ltc_10 (.L_LO(net10));
 sg13g2_tielo tt_um_flummer_ltc_11 (.L_LO(net11));
 sg13g2_tielo tt_um_flummer_ltc_12 (.L_LO(net12));
 sg13g2_tielo tt_um_flummer_ltc_13 (.L_LO(net13));
 sg13g2_tielo tt_um_flummer_ltc_14 (.L_LO(net14));
 sg13g2_tielo tt_um_flummer_ltc_15 (.L_LO(net15));
 sg13g2_tielo tt_um_flummer_ltc_16 (.L_LO(net16));
 sg13g2_tielo tt_um_flummer_ltc_17 (.L_LO(net17));
 sg13g2_tielo tt_um_flummer_ltc_18 (.L_LO(net18));
 sg13g2_tielo tt_um_flummer_ltc_19 (.L_LO(net19));
 sg13g2_tielo tt_um_flummer_ltc_20 (.L_LO(net20));
 sg13g2_tielo tt_um_flummer_ltc_21 (.L_LO(net21));
 sg13g2_tielo tt_um_flummer_ltc_22 (.L_LO(net22));
 sg13g2_tiehi _1352__23 (.L_HI(net23));
 sg13g2_buf_1 _1588_ (.A(\ltc.timecode ),
    .X(uio_out[7]));
 sg13g2_buf_1 _1589_ (.A(uio_in[0]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1590_ (.A(uio_in[1]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1591_ (.A(uio_in[2]),
    .X(uo_out[3]));
 sg13g2_buf_1 _1592_ (.A(uio_in[3]),
    .X(uo_out[4]));
 sg13g2_buf_1 _1593_ (.A(uio_in[4]),
    .X(uo_out[5]));
 sg13g2_buf_1 _1594_ (.A(uio_in[5]),
    .X(uo_out[6]));
 sg13g2_buf_1 _1595_ (.A(uio_in[6]),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout118 (.A(_0561_),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(_0561_),
    .X(net119));
 sg13g2_buf_8 fanout120 (.A(net122),
    .X(net120));
 sg13g2_buf_8 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_8 fanout122 (.A(_0453_),
    .X(net122));
 sg13g2_buf_8 fanout123 (.A(_0452_),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(net126),
    .X(net124));
 sg13g2_buf_1 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(net132),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(net129),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(net129),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(net132),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(net132),
    .X(net130));
 sg13g2_buf_1 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(_0196_),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(net137),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(_0194_),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(net142),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_1 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(_0193_),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0179_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_0179_),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(net154),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net154),
    .X(net149));
 sg13g2_buf_1 fanout150 (.A(net154),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net153),
    .X(net151));
 sg13g2_buf_1 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_0178_),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net160),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(net159),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(_0178_),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net169),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(net167),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(net167),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(_0155_),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_1 fanout172 (.A(net176),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net176),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(rst_n),
    .X(net176));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_flummer_ltc_9 (.L_LO(net9));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ltc.bit_counter[0] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ltc.frm_counter[0] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ltc.timecode ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0130_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ltc.bit_clk ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0143_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold7 (.A(\ltc.output_buffer[6] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0006_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ltc.frm_counter[21] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0464_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0102_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold12 (.A(\ltc.output_buffer[1] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0002_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ltc.output_buffer[5] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0005_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ltc.output_buffer[0] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ltc.output_buffer[11] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0011_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ltc.output_buffer[13] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0013_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold21 (.A(\ltc.output_buffer[9] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0009_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ltc.output_buffer[8] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0008_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold25 (.A(\ltc.output_buffer[7] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ltc.output_buffer[10] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold27 (.A(\ltc.output_buffer[2] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0003_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ltc.output_buffer[14] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ltc.output_buffer[4] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0004_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ltc.output_buffer[15] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold33 (.A(\ltc.output_buffer[12] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ltc.frm_counter[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0456_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0083_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold37 (.A(\ltc.output_buffer[51] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0052_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold39 (.A(\ltc.frm_counter[19] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0461_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0100_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold42 (.A(\ltc.bit_counter[5] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0564_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0136_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold45 (.A(\ltc.output_buffer[75] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0076_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold47 (.A(\ltc.bit_counter[3] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0562_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0134_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ltc.output_buffer[22] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0023_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ltc.output_buffer[52] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0053_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ltc.output_buffer[69] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0070_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold56 (.A(\ltc.output_buffer[16] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ltc.output_buffer[76] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0077_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold59 (.A(\ltc.bit_counter[7] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0566_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0138_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ltc.output_buffer[29] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0030_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ltc.output_buffer[30] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0031_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold66 (.A(\ltc.output_buffer[36] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0037_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold68 (.A(\ltc.frm_u[0] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ltc.output_buffer[62] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0063_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ltc.output_buffer[70] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0071_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ltc.output_buffer[45] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0046_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold75 (.A(\ltc.output_buffer[46] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0047_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ltc.output_buffer[57] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0349_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ltc.output_buffer[38] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0039_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold81 (.A(\ltc.output_buffer[18] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0202_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold83 (.A(\ltc.output_buffer[78] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0079_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold85 (.A(\ltc.output_buffer[68] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0368_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold87 (.A(\ltc.output_buffer[33] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0299_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold89 (.A(\ltc.output_buffer[28] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0029_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ltc.output_buffer[37] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0038_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold93 (.A(\ltc.output_buffer[21] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0275_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold95 (.A(\ltc.output_buffer[67] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0367_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold97 (.A(\ltc.bit_counter[11] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ltc.output_buffer[44] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0045_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold100 (.A(\ltc.output_buffer[74] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0378_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold102 (.A(\ltc.output_buffer[19] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0020_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold104 (.A(\ltc.hrs_d[1] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold105 (.A(\ltc.output_buffer[66] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0366_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold107 (.A(\ltc.output_buffer[35] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0301_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ltc.output_buffer[61] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0062_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ltc.frm_counter[23] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0467_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0104_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold114 (.A(\ltc.output_buffer[72] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0376_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold116 (.A(\ltc.output_buffer[53] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0054_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold118 (.A(\ltc.output_buffer[54] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0055_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ltc.output_buffer[56] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0348_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold122 (.A(\ltc.output_buffer[48] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0328_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold124 (.A(\ltc.output_buffer[43] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0315_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold126 (.A(\ltc.output_buffer[77] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0078_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold128 (.A(\ltc.output_buffer[42] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0314_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold130 (.A(\ltc.output_buffer[60] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0061_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold132 (.A(\ltc.output_buffer[24] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0282_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold134 (.A(\ltc.output_buffer[32] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0298_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ltc.output_buffer[64] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0364_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold138 (.A(\ltc.output_buffer[59] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0060_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold140 (.A(\ltc.output_buffer[27] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0285_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold142 (.A(\ltc.output_buffer[34] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold143 (.A(\ltc.output_buffer[40] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0312_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold145 (.A(\ltc.output_buffer[50] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0330_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold147 (.A(\ltc.output_buffer[49] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ltc.hrs_u[3] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold149 (.A(\ltc.frm_d[1] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0523_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold151 (.A(\ltc.frm_counter[22] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0465_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0103_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold154 (.A(\ltc.output_buffer[26] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0284_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold156 (.A(\ltc.output_buffer[58] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold157 (.A(\ltc.bit_counter[1] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold158 (.A(\ltc.output_buffer[25] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ltc.output_buffer[73] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold160 (.A(\ltc.output_buffer[41] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold161 (.A(\ltc.output_buffer[17] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold162 (.A(\ltc.min_u[1] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0492_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold164 (.A(\ltc.frm_u[2] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0128_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold166 (.A(\ltc.min_u[3] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold167 (.A(\ltc.sec_d[0] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0500_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0117_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold170 (.A(\ltc.bit_counter[8] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0567_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0139_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold173 (.A(\ltc.frm_counter[11] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0432_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0092_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold176 (.A(\ltc.min_d[2] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0486_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0112_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ltc.frm_counter[20] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0462_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold181 (.A(\ltc.min_d[0] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0483_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0110_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold184 (.A(\ltc.sec_d[2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0503_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0119_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold187 (.A(\ltc.min_u[2] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0494_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0115_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ltc.hrs_u[1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0475_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold192 (.A(\ltc.sec_u[1] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0514_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0121_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold195 (.A(\ltc.sec_d[1] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0501_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold197 (.A(\ltc.output_buffer[65] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold198 (.A(\ltc.min_u[0] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold199 (.A(\ltc.frm_counter[5] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0459_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0086_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold202 (.A(\ltc.frm_counter[1] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold203 (.A(\ltc.min_d[1] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold204 (.A(\ltc.hrs_d[0] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0471_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0105_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold207 (.A(\ltc.sec_u[2] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0517_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0122_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold210 (.A(\ltc.frm_counter[4] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0458_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold212 (.A(\ltc.frm_u[1] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold213 (.A(\ltc.hrs_u[0] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0399_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold215 (.A(\ltc.hrs_u[2] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold216 (.A(\ltc.bit_counter[4] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0563_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold218 (.A(\ltc.frm_u[3] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0129_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold220 (.A(\ltc.bit_counter[9] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0568_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold222 (.A(\ltc.sec_u[3] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0123_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold224 (.A(\ltc.frm_counter[3] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold225 (.A(\ltc.bit_counter[6] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold226 (.A(\ltc.bit_counter[10] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold227 (.A(\ltc.frm_counter[6] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold228 (.A(\ltc.frm_counter[18] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0416_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold230 (.A(\ltc.bit_counter[2] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold231 (.A(\ltc.frm_counter[10] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0433_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold233 (.A(\ltc.frm_counter[15] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0436_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold235 (.A(\ltc.frm_counter[13] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0094_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold237 (.A(\ltc.sec_u[0] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold238 (.A(\ltc.frm_counter[16] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0419_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold240 (.A(\ltc.frm_counter[8] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold241 (.A(\ltc.frm_d[0] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold242 (.A(\ltc.frm_counter[12] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold243 (.A(\ltc.frm_counter[9] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold244 (.A(\ltc.frm_counter[7] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold245 (.A(\ltc.frm_counter[14] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0446_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold247 (.A(\ltc.frm_counter[17] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold248 (.A(\ltc.frm_counter[13] ),
    .X(net474));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_4 FILLER_0_28 ();
 sg13g2_fill_1 FILLER_0_32 ();
 sg13g2_fill_2 FILLER_0_49 ();
 sg13g2_fill_1 FILLER_0_51 ();
 sg13g2_fill_1 FILLER_0_69 ();
 sg13g2_decap_8 FILLER_0_74 ();
 sg13g2_decap_4 FILLER_0_81 ();
 sg13g2_decap_8 FILLER_0_89 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_117 ();
 sg13g2_decap_8 FILLER_0_124 ();
 sg13g2_decap_8 FILLER_0_131 ();
 sg13g2_decap_8 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_decap_8 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_fill_1 FILLER_1_60 ();
 sg13g2_decap_8 FILLER_1_93 ();
 sg13g2_fill_1 FILLER_1_100 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_fill_2 FILLER_1_189 ();
 sg13g2_fill_2 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_214 ();
 sg13g2_decap_8 FILLER_1_221 ();
 sg13g2_decap_8 FILLER_1_228 ();
 sg13g2_decap_8 FILLER_1_235 ();
 sg13g2_decap_8 FILLER_1_242 ();
 sg13g2_decap_8 FILLER_1_249 ();
 sg13g2_decap_8 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_305 ();
 sg13g2_decap_8 FILLER_1_312 ();
 sg13g2_decap_8 FILLER_1_319 ();
 sg13g2_decap_8 FILLER_1_326 ();
 sg13g2_decap_8 FILLER_1_333 ();
 sg13g2_decap_8 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_354 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_375 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_4 FILLER_1_403 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_7 ();
 sg13g2_fill_1 FILLER_2_36 ();
 sg13g2_decap_4 FILLER_2_51 ();
 sg13g2_fill_2 FILLER_2_107 ();
 sg13g2_fill_1 FILLER_2_109 ();
 sg13g2_decap_4 FILLER_2_114 ();
 sg13g2_fill_1 FILLER_2_118 ();
 sg13g2_fill_2 FILLER_2_147 ();
 sg13g2_fill_1 FILLER_2_149 ();
 sg13g2_decap_8 FILLER_2_177 ();
 sg13g2_decap_4 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_216 ();
 sg13g2_decap_8 FILLER_2_223 ();
 sg13g2_decap_8 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_237 ();
 sg13g2_decap_8 FILLER_2_244 ();
 sg13g2_decap_8 FILLER_2_251 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_8 FILLER_2_279 ();
 sg13g2_decap_8 FILLER_2_286 ();
 sg13g2_decap_8 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_300 ();
 sg13g2_decap_8 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_12 ();
 sg13g2_decap_8 FILLER_3_17 ();
 sg13g2_decap_4 FILLER_3_24 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_64 ();
 sg13g2_decap_4 FILLER_3_139 ();
 sg13g2_fill_2 FILLER_3_143 ();
 sg13g2_fill_1 FILLER_3_162 ();
 sg13g2_fill_1 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_178 ();
 sg13g2_fill_2 FILLER_3_191 ();
 sg13g2_fill_1 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_236 ();
 sg13g2_decap_8 FILLER_3_243 ();
 sg13g2_decap_8 FILLER_3_250 ();
 sg13g2_decap_8 FILLER_3_257 ();
 sg13g2_decap_8 FILLER_3_264 ();
 sg13g2_decap_8 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_decap_8 FILLER_3_285 ();
 sg13g2_decap_8 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_299 ();
 sg13g2_decap_8 FILLER_3_306 ();
 sg13g2_decap_8 FILLER_3_313 ();
 sg13g2_decap_8 FILLER_3_320 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_decap_8 FILLER_3_334 ();
 sg13g2_decap_8 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_2 ();
 sg13g2_fill_1 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_59 ();
 sg13g2_fill_2 FILLER_4_67 ();
 sg13g2_fill_1 FILLER_4_91 ();
 sg13g2_fill_2 FILLER_4_111 ();
 sg13g2_fill_2 FILLER_4_160 ();
 sg13g2_fill_2 FILLER_4_178 ();
 sg13g2_fill_2 FILLER_4_207 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_decap_8 FILLER_4_232 ();
 sg13g2_decap_8 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_246 ();
 sg13g2_decap_8 FILLER_4_253 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_295 ();
 sg13g2_decap_8 FILLER_4_302 ();
 sg13g2_decap_8 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_21 ();
 sg13g2_fill_2 FILLER_5_49 ();
 sg13g2_fill_1 FILLER_5_56 ();
 sg13g2_fill_2 FILLER_5_75 ();
 sg13g2_fill_2 FILLER_5_119 ();
 sg13g2_fill_1 FILLER_5_152 ();
 sg13g2_decap_4 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_236 ();
 sg13g2_decap_8 FILLER_5_243 ();
 sg13g2_decap_8 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_271 ();
 sg13g2_decap_8 FILLER_5_278 ();
 sg13g2_decap_8 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_5_306 ();
 sg13g2_decap_8 FILLER_5_313 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_334 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_2 ();
 sg13g2_fill_2 FILLER_6_40 ();
 sg13g2_fill_2 FILLER_6_50 ();
 sg13g2_fill_1 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_57 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_fill_2 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_93 ();
 sg13g2_decap_4 FILLER_6_112 ();
 sg13g2_fill_1 FILLER_6_116 ();
 sg13g2_fill_1 FILLER_6_127 ();
 sg13g2_decap_8 FILLER_6_141 ();
 sg13g2_fill_2 FILLER_6_148 ();
 sg13g2_decap_4 FILLER_6_180 ();
 sg13g2_fill_1 FILLER_6_184 ();
 sg13g2_decap_4 FILLER_6_193 ();
 sg13g2_fill_1 FILLER_6_197 ();
 sg13g2_fill_2 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_237 ();
 sg13g2_decap_8 FILLER_6_244 ();
 sg13g2_decap_8 FILLER_6_251 ();
 sg13g2_decap_8 FILLER_6_258 ();
 sg13g2_decap_8 FILLER_6_265 ();
 sg13g2_decap_8 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_27 ();
 sg13g2_fill_1 FILLER_7_97 ();
 sg13g2_fill_2 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_109 ();
 sg13g2_fill_2 FILLER_7_118 ();
 sg13g2_fill_1 FILLER_7_120 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_128 ();
 sg13g2_fill_2 FILLER_7_164 ();
 sg13g2_fill_1 FILLER_7_179 ();
 sg13g2_decap_8 FILLER_7_197 ();
 sg13g2_fill_2 FILLER_7_204 ();
 sg13g2_fill_1 FILLER_7_206 ();
 sg13g2_decap_8 FILLER_7_211 ();
 sg13g2_decap_8 FILLER_7_218 ();
 sg13g2_decap_4 FILLER_7_225 ();
 sg13g2_decap_8 FILLER_7_246 ();
 sg13g2_decap_8 FILLER_7_253 ();
 sg13g2_decap_8 FILLER_7_260 ();
 sg13g2_decap_8 FILLER_7_267 ();
 sg13g2_decap_8 FILLER_7_274 ();
 sg13g2_decap_8 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_288 ();
 sg13g2_decap_8 FILLER_7_295 ();
 sg13g2_decap_8 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_316 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_8 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_2 FILLER_8_30 ();
 sg13g2_fill_1 FILLER_8_32 ();
 sg13g2_fill_1 FILLER_8_47 ();
 sg13g2_fill_2 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_150 ();
 sg13g2_fill_2 FILLER_8_157 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_257 ();
 sg13g2_decap_8 FILLER_8_264 ();
 sg13g2_decap_8 FILLER_8_271 ();
 sg13g2_decap_8 FILLER_8_278 ();
 sg13g2_decap_4 FILLER_8_285 ();
 sg13g2_fill_2 FILLER_8_289 ();
 sg13g2_fill_2 FILLER_8_294 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_decap_4 FILLER_8_313 ();
 sg13g2_decap_8 FILLER_8_320 ();
 sg13g2_decap_8 FILLER_8_327 ();
 sg13g2_decap_8 FILLER_8_334 ();
 sg13g2_decap_8 FILLER_8_341 ();
 sg13g2_decap_8 FILLER_8_348 ();
 sg13g2_decap_8 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_362 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_8 ();
 sg13g2_fill_1 FILLER_9_12 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_fill_1 FILLER_9_50 ();
 sg13g2_fill_2 FILLER_9_64 ();
 sg13g2_fill_2 FILLER_9_79 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_fill_2 FILLER_9_178 ();
 sg13g2_fill_1 FILLER_9_180 ();
 sg13g2_fill_2 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_227 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_4 FILLER_9_280 ();
 sg13g2_fill_1 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_4 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_45 ();
 sg13g2_fill_2 FILLER_10_74 ();
 sg13g2_fill_2 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_101 ();
 sg13g2_decap_8 FILLER_10_111 ();
 sg13g2_fill_2 FILLER_10_118 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_fill_2 FILLER_10_181 ();
 sg13g2_fill_2 FILLER_10_192 ();
 sg13g2_fill_1 FILLER_10_194 ();
 sg13g2_decap_4 FILLER_10_211 ();
 sg13g2_fill_2 FILLER_10_215 ();
 sg13g2_fill_2 FILLER_10_243 ();
 sg13g2_fill_2 FILLER_10_267 ();
 sg13g2_fill_1 FILLER_10_269 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_fill_1 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_fill_1 FILLER_11_16 ();
 sg13g2_fill_1 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_48 ();
 sg13g2_decap_4 FILLER_11_89 ();
 sg13g2_decap_4 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_fill_2 FILLER_11_180 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_209 ();
 sg13g2_fill_2 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_232 ();
 sg13g2_decap_8 FILLER_11_260 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_fill_2 FILLER_11_332 ();
 sg13g2_fill_1 FILLER_11_334 ();
 sg13g2_decap_4 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_2 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_4 FILLER_12_84 ();
 sg13g2_fill_2 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_100 ();
 sg13g2_decap_4 FILLER_12_129 ();
 sg13g2_fill_1 FILLER_12_133 ();
 sg13g2_fill_2 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_fill_1 FILLER_12_199 ();
 sg13g2_fill_2 FILLER_12_219 ();
 sg13g2_fill_1 FILLER_12_221 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_248 ();
 sg13g2_fill_1 FILLER_12_263 ();
 sg13g2_fill_1 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_339 ();
 sg13g2_fill_2 FILLER_12_353 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_29 ();
 sg13g2_fill_2 FILLER_13_73 ();
 sg13g2_fill_1 FILLER_13_75 ();
 sg13g2_fill_2 FILLER_13_84 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_286 ();
 sg13g2_fill_1 FILLER_13_288 ();
 sg13g2_fill_2 FILLER_13_293 ();
 sg13g2_fill_1 FILLER_13_298 ();
 sg13g2_fill_2 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_fill_2 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_2 FILLER_14_87 ();
 sg13g2_fill_1 FILLER_14_89 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_fill_1 FILLER_14_129 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_fill_1 FILLER_14_164 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_decap_4 FILLER_14_203 ();
 sg13g2_fill_2 FILLER_14_211 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_fill_2 FILLER_14_277 ();
 sg13g2_fill_1 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_decap_4 FILLER_14_387 ();
 sg13g2_fill_1 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_33 ();
 sg13g2_fill_1 FILLER_15_44 ();
 sg13g2_decap_4 FILLER_15_81 ();
 sg13g2_fill_2 FILLER_15_112 ();
 sg13g2_fill_2 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_130 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_decap_4 FILLER_15_296 ();
 sg13g2_fill_2 FILLER_15_300 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_decap_4 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_41 ();
 sg13g2_fill_1 FILLER_16_43 ();
 sg13g2_fill_2 FILLER_16_89 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_4 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_decap_8 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_184 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_fill_1 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_4 FILLER_16_228 ();
 sg13g2_fill_1 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_18 ();
 sg13g2_decap_8 FILLER_17_23 ();
 sg13g2_decap_4 FILLER_17_30 ();
 sg13g2_fill_2 FILLER_17_75 ();
 sg13g2_fill_1 FILLER_17_104 ();
 sg13g2_fill_2 FILLER_17_109 ();
 sg13g2_fill_1 FILLER_17_111 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_decap_4 FILLER_17_190 ();
 sg13g2_fill_1 FILLER_17_194 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_247 ();
 sg13g2_decap_4 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_294 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_fill_1 FILLER_17_314 ();
 sg13g2_fill_2 FILLER_17_332 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_4 FILLER_17_386 ();
 sg13g2_fill_1 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_fill_1 FILLER_18_81 ();
 sg13g2_decap_4 FILLER_18_86 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_145 ();
 sg13g2_fill_1 FILLER_18_162 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_4 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_decap_4 FILLER_18_232 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_333 ();
 sg13g2_fill_1 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_23 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_39 ();
 sg13g2_fill_1 FILLER_19_61 ();
 sg13g2_decap_4 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_95 ();
 sg13g2_decap_4 FILLER_19_115 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_decap_4 FILLER_19_188 ();
 sg13g2_decap_4 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_decap_4 FILLER_20_74 ();
 sg13g2_fill_1 FILLER_20_95 ();
 sg13g2_fill_2 FILLER_20_104 ();
 sg13g2_fill_2 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_237 ();
 sg13g2_decap_4 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_4 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_decap_4 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_39 ();
 sg13g2_decap_4 FILLER_21_45 ();
 sg13g2_fill_2 FILLER_21_62 ();
 sg13g2_fill_1 FILLER_21_99 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_decap_4 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_314 ();
 sg13g2_fill_2 FILLER_21_321 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_decap_4 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_25 ();
 sg13g2_fill_1 FILLER_22_46 ();
 sg13g2_fill_2 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_fill_2 FILLER_22_58 ();
 sg13g2_decap_8 FILLER_22_100 ();
 sg13g2_fill_2 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_decap_4 FILLER_22_123 ();
 sg13g2_fill_1 FILLER_22_127 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_decap_8 FILLER_22_268 ();
 sg13g2_fill_2 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_277 ();
 sg13g2_decap_4 FILLER_22_287 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_69 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_82 ();
 sg13g2_decap_8 FILLER_23_87 ();
 sg13g2_decap_8 FILLER_23_94 ();
 sg13g2_fill_1 FILLER_23_101 ();
 sg13g2_decap_4 FILLER_23_106 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_fill_2 FILLER_23_138 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_decap_4 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_decap_8 FILLER_23_222 ();
 sg13g2_decap_8 FILLER_23_229 ();
 sg13g2_fill_2 FILLER_23_293 ();
 sg13g2_decap_4 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_359 ();
 sg13g2_decap_8 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_31 ();
 sg13g2_fill_2 FILLER_24_50 ();
 sg13g2_fill_1 FILLER_24_52 ();
 sg13g2_fill_2 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_155 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_8 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_252 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_160 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_fill_2 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_226 ();
 sg13g2_decap_4 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_fill_2 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_41 ();
 sg13g2_fill_2 FILLER_26_52 ();
 sg13g2_fill_1 FILLER_26_54 ();
 sg13g2_fill_1 FILLER_26_69 ();
 sg13g2_fill_1 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_fill_2 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_295 ();
 sg13g2_decap_4 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_decap_4 FILLER_27_36 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_decap_4 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_107 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_128 ();
 sg13g2_fill_2 FILLER_28_166 ();
 sg13g2_decap_8 FILLER_28_199 ();
 sg13g2_decap_4 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_234 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_decap_4 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_53 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_137 ();
 sg13g2_decap_8 FILLER_29_155 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_fill_1 FILLER_29_193 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_2 FILLER_29_281 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_decap_4 FILLER_29_321 ();
 sg13g2_fill_2 FILLER_29_325 ();
 sg13g2_fill_2 FILLER_29_393 ();
 sg13g2_fill_1 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_4 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_79 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_decap_4 FILLER_30_86 ();
 sg13g2_fill_1 FILLER_30_90 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_236 ();
 sg13g2_fill_2 FILLER_30_268 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_319 ();
 sg13g2_fill_2 FILLER_30_336 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_decap_4 FILLER_31_58 ();
 sg13g2_decap_4 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_decap_4 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_182 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_261 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_fill_2 FILLER_31_277 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_decap_4 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_decap_4 FILLER_31_321 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_26 ();
 sg13g2_fill_2 FILLER_32_30 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_349 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_43 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_fill_1 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_fill_2 FILLER_33_136 ();
 sg13g2_decap_8 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_150 ();
 sg13g2_decap_4 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_decap_4 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_decap_4 FILLER_33_324 ();
 sg13g2_fill_2 FILLER_33_328 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_18 ();
 sg13g2_fill_1 FILLER_34_94 ();
 sg13g2_fill_2 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_114 ();
 sg13g2_fill_2 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_154 ();
 sg13g2_decap_4 FILLER_34_159 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_197 ();
 sg13g2_decap_8 FILLER_34_205 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_2 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_80 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_decap_4 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_2 FILLER_35_240 ();
 sg13g2_fill_1 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_272 ();
 sg13g2_fill_2 FILLER_35_285 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_2 FILLER_35_301 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_25 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_34 ();
 sg13g2_fill_1 FILLER_36_99 ();
 sg13g2_decap_8 FILLER_36_157 ();
 sg13g2_decap_4 FILLER_36_164 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_4 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_78 ();
 sg13g2_fill_2 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_214 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_2 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_93 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_fill_2 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_227 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_fill_1 FILLER_38_331 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net226;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
endmodule
