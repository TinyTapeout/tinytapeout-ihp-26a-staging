module tt_um_corey (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15922_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire _15934_;
 wire _15935_;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire _15945_;
 wire _15946_;
 wire _15947_;
 wire _15948_;
 wire _15949_;
 wire _15950_;
 wire _15951_;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire _15958_;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire _16040_;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire _16052_;
 wire _16053_;
 wire _16054_;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire _16080_;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire _16152_;
 wire _16153_;
 wire _16154_;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16196_;
 wire _16197_;
 wire _16198_;
 wire _16199_;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire _16218_;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire _16264_;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16380_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire _16443_;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire _16458_;
 wire _16459_;
 wire _16460_;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire _16569_;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire _16720_;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire _17813_;
 wire _17814_;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire _18322_;
 wire _18323_;
 wire _18324_;
 wire _18325_;
 wire _18326_;
 wire _18327_;
 wire _18328_;
 wire _18329_;
 wire _18330_;
 wire _18331_;
 wire _18332_;
 wire _18333_;
 wire _18334_;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire _18338_;
 wire _18339_;
 wire _18340_;
 wire _18341_;
 wire _18342_;
 wire _18343_;
 wire _18344_;
 wire _18345_;
 wire _18346_;
 wire _18347_;
 wire _18348_;
 wire _18349_;
 wire _18350_;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire _18354_;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire _18358_;
 wire _18359_;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire _18364_;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire _18368_;
 wire _18369_;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire _18373_;
 wire _18374_;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire _18378_;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire _18398_;
 wire _18399_;
 wire _18400_;
 wire _18401_;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire _18406_;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire _18411_;
 wire _18412_;
 wire _18413_;
 wire _18414_;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire _18420_;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire _18428_;
 wire _18429_;
 wire _18430_;
 wire _18431_;
 wire _18432_;
 wire _18433_;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire _18438_;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire _18443_;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire _18448_;
 wire _18449_;
 wire _18450_;
 wire _18451_;
 wire _18452_;
 wire _18453_;
 wire _18454_;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire _18458_;
 wire _18459_;
 wire _18460_;
 wire _18461_;
 wire _18462_;
 wire _18463_;
 wire _18464_;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire _18468_;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire _18473_;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire _18606_;
 wire _18607_;
 wire _18608_;
 wire _18609_;
 wire _18610_;
 wire _18611_;
 wire _18612_;
 wire _18613_;
 wire _18614_;
 wire _18615_;
 wire _18616_;
 wire _18617_;
 wire _18618_;
 wire _18619_;
 wire _18620_;
 wire _18621_;
 wire _18622_;
 wire _18623_;
 wire _18624_;
 wire _18625_;
 wire _18626_;
 wire _18627_;
 wire _18628_;
 wire _18629_;
 wire _18630_;
 wire _18631_;
 wire _18632_;
 wire _18633_;
 wire _18634_;
 wire _18635_;
 wire _18636_;
 wire _18637_;
 wire _18638_;
 wire _18639_;
 wire _18640_;
 wire _18641_;
 wire _18642_;
 wire _18643_;
 wire _18644_;
 wire _18645_;
 wire _18646_;
 wire _18647_;
 wire _18648_;
 wire _18649_;
 wire _18650_;
 wire _18651_;
 wire _18652_;
 wire _18653_;
 wire _18654_;
 wire _18655_;
 wire _18656_;
 wire _18657_;
 wire _18658_;
 wire _18659_;
 wire _18660_;
 wire _18661_;
 wire _18662_;
 wire _18663_;
 wire _18664_;
 wire _18665_;
 wire _18666_;
 wire _18667_;
 wire _18668_;
 wire _18669_;
 wire _18670_;
 wire _18671_;
 wire _18672_;
 wire _18673_;
 wire _18674_;
 wire _18675_;
 wire _18676_;
 wire _18677_;
 wire _18678_;
 wire _18679_;
 wire _18680_;
 wire _18681_;
 wire _18682_;
 wire _18683_;
 wire _18684_;
 wire _18685_;
 wire _18686_;
 wire _18687_;
 wire _18688_;
 wire _18689_;
 wire _18690_;
 wire _18691_;
 wire _18692_;
 wire _18693_;
 wire _18694_;
 wire _18695_;
 wire _18696_;
 wire _18697_;
 wire _18698_;
 wire _18699_;
 wire _18700_;
 wire _18701_;
 wire _18702_;
 wire _18703_;
 wire _18704_;
 wire _18705_;
 wire _18706_;
 wire _18707_;
 wire _18708_;
 wire _18709_;
 wire _18710_;
 wire _18711_;
 wire _18712_;
 wire _18713_;
 wire _18714_;
 wire _18715_;
 wire _18716_;
 wire _18717_;
 wire _18718_;
 wire _18719_;
 wire _18720_;
 wire _18721_;
 wire _18722_;
 wire _18723_;
 wire _18724_;
 wire _18725_;
 wire _18726_;
 wire _18727_;
 wire _18728_;
 wire _18729_;
 wire _18730_;
 wire _18731_;
 wire _18732_;
 wire _18733_;
 wire _18734_;
 wire _18735_;
 wire _18736_;
 wire _18737_;
 wire _18738_;
 wire _18739_;
 wire _18740_;
 wire _18741_;
 wire _18742_;
 wire _18743_;
 wire _18744_;
 wire _18745_;
 wire _18746_;
 wire _18747_;
 wire _18748_;
 wire _18749_;
 wire _18750_;
 wire _18751_;
 wire _18752_;
 wire _18753_;
 wire _18754_;
 wire _18755_;
 wire _18756_;
 wire _18757_;
 wire _18758_;
 wire _18759_;
 wire _18760_;
 wire _18761_;
 wire _18762_;
 wire _18763_;
 wire _18764_;
 wire _18765_;
 wire _18766_;
 wire _18767_;
 wire _18768_;
 wire _18769_;
 wire _18770_;
 wire _18771_;
 wire _18772_;
 wire _18773_;
 wire _18774_;
 wire _18775_;
 wire _18776_;
 wire _18777_;
 wire _18778_;
 wire _18779_;
 wire _18780_;
 wire _18781_;
 wire _18782_;
 wire _18783_;
 wire _18784_;
 wire _18785_;
 wire _18786_;
 wire _18787_;
 wire _18788_;
 wire _18789_;
 wire _18790_;
 wire _18791_;
 wire _18792_;
 wire _18793_;
 wire _18794_;
 wire _18795_;
 wire _18796_;
 wire _18797_;
 wire _18798_;
 wire _18799_;
 wire _18800_;
 wire _18801_;
 wire _18802_;
 wire _18803_;
 wire _18804_;
 wire _18805_;
 wire _18806_;
 wire _18807_;
 wire _18808_;
 wire _18809_;
 wire _18810_;
 wire _18811_;
 wire _18812_;
 wire _18813_;
 wire _18814_;
 wire _18815_;
 wire _18816_;
 wire _18817_;
 wire _18818_;
 wire _18819_;
 wire _18820_;
 wire _18821_;
 wire _18822_;
 wire _18823_;
 wire _18824_;
 wire _18825_;
 wire _18826_;
 wire _18827_;
 wire _18828_;
 wire _18829_;
 wire _18830_;
 wire _18831_;
 wire _18832_;
 wire _18833_;
 wire _18834_;
 wire _18835_;
 wire _18836_;
 wire _18837_;
 wire _18838_;
 wire _18839_;
 wire _18840_;
 wire _18841_;
 wire _18842_;
 wire _18843_;
 wire _18844_;
 wire _18845_;
 wire _18846_;
 wire _18847_;
 wire _18848_;
 wire _18849_;
 wire _18850_;
 wire _18851_;
 wire _18852_;
 wire _18853_;
 wire _18854_;
 wire _18855_;
 wire _18856_;
 wire _18857_;
 wire _18858_;
 wire _18859_;
 wire _18860_;
 wire _18861_;
 wire _18862_;
 wire _18863_;
 wire _18864_;
 wire _18865_;
 wire _18866_;
 wire _18867_;
 wire _18868_;
 wire _18869_;
 wire _18870_;
 wire _18871_;
 wire _18872_;
 wire _18873_;
 wire _18874_;
 wire _18875_;
 wire _18876_;
 wire _18877_;
 wire _18878_;
 wire _18879_;
 wire _18880_;
 wire _18881_;
 wire _18882_;
 wire _18883_;
 wire _18884_;
 wire _18885_;
 wire _18886_;
 wire _18887_;
 wire _18888_;
 wire _18889_;
 wire _18890_;
 wire _18891_;
 wire _18892_;
 wire _18893_;
 wire _18894_;
 wire _18895_;
 wire _18896_;
 wire _18897_;
 wire _18898_;
 wire _18899_;
 wire _18900_;
 wire _18901_;
 wire _18902_;
 wire _18903_;
 wire _18904_;
 wire _18905_;
 wire _18906_;
 wire _18907_;
 wire _18908_;
 wire _18909_;
 wire _18910_;
 wire _18911_;
 wire _18912_;
 wire _18913_;
 wire _18914_;
 wire _18915_;
 wire _18916_;
 wire _18917_;
 wire _18918_;
 wire _18919_;
 wire _18920_;
 wire _18921_;
 wire _18922_;
 wire _18923_;
 wire _18924_;
 wire _18925_;
 wire _18926_;
 wire _18927_;
 wire _18928_;
 wire _18929_;
 wire _18930_;
 wire _18931_;
 wire _18932_;
 wire _18933_;
 wire _18934_;
 wire _18935_;
 wire _18936_;
 wire _18937_;
 wire _18938_;
 wire _18939_;
 wire _18940_;
 wire _18941_;
 wire _18942_;
 wire _18943_;
 wire _18944_;
 wire _18945_;
 wire _18946_;
 wire _18947_;
 wire _18948_;
 wire _18949_;
 wire _18950_;
 wire _18951_;
 wire _18952_;
 wire _18953_;
 wire _18954_;
 wire _18955_;
 wire _18956_;
 wire _18957_;
 wire _18958_;
 wire _18959_;
 wire _18960_;
 wire _18961_;
 wire _18962_;
 wire _18963_;
 wire _18964_;
 wire _18965_;
 wire _18966_;
 wire _18967_;
 wire _18968_;
 wire _18969_;
 wire _18970_;
 wire _18971_;
 wire _18972_;
 wire _18973_;
 wire _18974_;
 wire _18975_;
 wire _18976_;
 wire _18977_;
 wire _18978_;
 wire _18979_;
 wire _18980_;
 wire _18981_;
 wire _18982_;
 wire _18983_;
 wire _18984_;
 wire _18985_;
 wire _18986_;
 wire _18987_;
 wire _18988_;
 wire _18989_;
 wire _18990_;
 wire _18991_;
 wire _18992_;
 wire _18993_;
 wire _18994_;
 wire _18995_;
 wire _18996_;
 wire _18997_;
 wire _18998_;
 wire _18999_;
 wire _19000_;
 wire _19001_;
 wire _19002_;
 wire _19003_;
 wire _19004_;
 wire _19005_;
 wire _19006_;
 wire _19007_;
 wire _19008_;
 wire _19009_;
 wire _19010_;
 wire _19011_;
 wire _19012_;
 wire _19013_;
 wire _19014_;
 wire _19015_;
 wire _19016_;
 wire _19017_;
 wire _19018_;
 wire _19019_;
 wire _19020_;
 wire _19021_;
 wire _19022_;
 wire _19023_;
 wire _19024_;
 wire _19025_;
 wire _19026_;
 wire _19027_;
 wire _19028_;
 wire _19029_;
 wire _19030_;
 wire _19031_;
 wire _19032_;
 wire _19033_;
 wire _19034_;
 wire _19035_;
 wire _19036_;
 wire _19037_;
 wire _19038_;
 wire _19039_;
 wire _19040_;
 wire _19041_;
 wire _19042_;
 wire _19043_;
 wire _19044_;
 wire _19045_;
 wire _19046_;
 wire _19047_;
 wire _19048_;
 wire _19049_;
 wire _19050_;
 wire _19051_;
 wire _19052_;
 wire _19053_;
 wire _19054_;
 wire _19055_;
 wire _19056_;
 wire _19057_;
 wire _19058_;
 wire _19059_;
 wire _19060_;
 wire _19061_;
 wire _19062_;
 wire _19063_;
 wire _19064_;
 wire _19065_;
 wire _19066_;
 wire _19067_;
 wire _19068_;
 wire _19069_;
 wire _19070_;
 wire _19071_;
 wire _19072_;
 wire _19073_;
 wire _19074_;
 wire _19075_;
 wire _19076_;
 wire _19077_;
 wire _19078_;
 wire _19079_;
 wire _19080_;
 wire _19081_;
 wire _19082_;
 wire _19083_;
 wire _19084_;
 wire _19085_;
 wire _19086_;
 wire _19087_;
 wire _19088_;
 wire _19089_;
 wire _19090_;
 wire _19091_;
 wire _19092_;
 wire _19093_;
 wire _19094_;
 wire _19095_;
 wire _19096_;
 wire _19097_;
 wire _19098_;
 wire _19099_;
 wire _19100_;
 wire _19101_;
 wire _19102_;
 wire _19103_;
 wire _19104_;
 wire _19105_;
 wire _19106_;
 wire _19107_;
 wire _19108_;
 wire _19109_;
 wire _19110_;
 wire _19111_;
 wire _19112_;
 wire _19113_;
 wire _19114_;
 wire _19115_;
 wire _19116_;
 wire _19117_;
 wire _19118_;
 wire _19119_;
 wire _19120_;
 wire _19121_;
 wire _19122_;
 wire _19123_;
 wire _19124_;
 wire _19125_;
 wire _19126_;
 wire _19127_;
 wire _19128_;
 wire _19129_;
 wire _19130_;
 wire _19131_;
 wire _19132_;
 wire _19133_;
 wire _19134_;
 wire _19135_;
 wire _19136_;
 wire _19137_;
 wire _19138_;
 wire _19139_;
 wire _19140_;
 wire _19141_;
 wire _19142_;
 wire _19143_;
 wire _19144_;
 wire _19145_;
 wire _19146_;
 wire _19147_;
 wire _19148_;
 wire _19149_;
 wire _19150_;
 wire _19151_;
 wire _19152_;
 wire _19153_;
 wire _19154_;
 wire _19155_;
 wire _19156_;
 wire _19157_;
 wire _19158_;
 wire _19159_;
 wire _19160_;
 wire _19161_;
 wire _19162_;
 wire _19163_;
 wire _19164_;
 wire _19165_;
 wire _19166_;
 wire _19167_;
 wire _19168_;
 wire _19169_;
 wire _19170_;
 wire _19171_;
 wire _19172_;
 wire _19173_;
 wire _19174_;
 wire _19175_;
 wire _19176_;
 wire _19177_;
 wire _19178_;
 wire _19179_;
 wire _19180_;
 wire _19181_;
 wire _19182_;
 wire _19183_;
 wire _19184_;
 wire _19185_;
 wire _19186_;
 wire _19187_;
 wire _19188_;
 wire _19189_;
 wire _19190_;
 wire _19191_;
 wire _19192_;
 wire _19193_;
 wire _19194_;
 wire _19195_;
 wire _19196_;
 wire _19197_;
 wire _19198_;
 wire _19199_;
 wire _19200_;
 wire _19201_;
 wire _19202_;
 wire _19203_;
 wire _19204_;
 wire _19205_;
 wire _19206_;
 wire _19207_;
 wire _19208_;
 wire _19209_;
 wire _19210_;
 wire _19211_;
 wire _19212_;
 wire _19213_;
 wire _19214_;
 wire _19215_;
 wire _19216_;
 wire _19217_;
 wire _19218_;
 wire _19219_;
 wire _19220_;
 wire _19221_;
 wire _19222_;
 wire _19223_;
 wire _19224_;
 wire _19225_;
 wire _19226_;
 wire _19227_;
 wire _19228_;
 wire _19229_;
 wire _19230_;
 wire _19231_;
 wire _19232_;
 wire _19233_;
 wire _19234_;
 wire _19235_;
 wire _19236_;
 wire _19237_;
 wire _19238_;
 wire _19239_;
 wire _19240_;
 wire _19241_;
 wire _19242_;
 wire _19243_;
 wire _19244_;
 wire _19245_;
 wire _19246_;
 wire _19247_;
 wire _19248_;
 wire _19249_;
 wire _19250_;
 wire _19251_;
 wire _19252_;
 wire _19253_;
 wire _19254_;
 wire _19255_;
 wire _19256_;
 wire _19257_;
 wire _19258_;
 wire _19259_;
 wire _19260_;
 wire _19261_;
 wire _19262_;
 wire _19263_;
 wire _19264_;
 wire _19265_;
 wire _19266_;
 wire _19267_;
 wire _19268_;
 wire _19269_;
 wire _19270_;
 wire _19271_;
 wire _19272_;
 wire _19273_;
 wire _19274_;
 wire _19275_;
 wire _19276_;
 wire _19277_;
 wire _19278_;
 wire _19279_;
 wire _19280_;
 wire _19281_;
 wire _19282_;
 wire _19283_;
 wire _19284_;
 wire _19285_;
 wire _19286_;
 wire _19287_;
 wire _19288_;
 wire _19289_;
 wire _19290_;
 wire _19291_;
 wire _19292_;
 wire _19293_;
 wire _19294_;
 wire _19295_;
 wire _19296_;
 wire _19297_;
 wire _19298_;
 wire _19299_;
 wire _19300_;
 wire _19301_;
 wire _19302_;
 wire _19303_;
 wire _19304_;
 wire _19305_;
 wire _19306_;
 wire _19307_;
 wire _19308_;
 wire _19309_;
 wire _19310_;
 wire _19311_;
 wire _19312_;
 wire _19313_;
 wire _19314_;
 wire _19315_;
 wire _19316_;
 wire _19317_;
 wire _19318_;
 wire _19319_;
 wire _19320_;
 wire _19321_;
 wire _19322_;
 wire _19323_;
 wire _19324_;
 wire _19325_;
 wire _19326_;
 wire _19327_;
 wire _19328_;
 wire _19329_;
 wire _19330_;
 wire _19331_;
 wire _19332_;
 wire _19333_;
 wire _19334_;
 wire _19335_;
 wire _19336_;
 wire _19337_;
 wire _19338_;
 wire _19339_;
 wire _19340_;
 wire _19341_;
 wire _19342_;
 wire _19343_;
 wire _19344_;
 wire _19345_;
 wire _19346_;
 wire _19347_;
 wire _19348_;
 wire _19349_;
 wire _19350_;
 wire _19351_;
 wire _19352_;
 wire _19353_;
 wire _19354_;
 wire _19355_;
 wire _19356_;
 wire _19357_;
 wire _19358_;
 wire _19359_;
 wire _19360_;
 wire _19361_;
 wire _19362_;
 wire _19363_;
 wire _19364_;
 wire _19365_;
 wire _19366_;
 wire _19367_;
 wire _19368_;
 wire _19369_;
 wire _19370_;
 wire _19371_;
 wire _19372_;
 wire _19373_;
 wire _19374_;
 wire _19375_;
 wire _19376_;
 wire _19377_;
 wire _19378_;
 wire _19379_;
 wire _19380_;
 wire _19381_;
 wire _19382_;
 wire _19383_;
 wire _19384_;
 wire _19385_;
 wire _19386_;
 wire _19387_;
 wire _19388_;
 wire _19389_;
 wire _19390_;
 wire _19391_;
 wire _19392_;
 wire _19393_;
 wire _19394_;
 wire _19395_;
 wire _19396_;
 wire _19397_;
 wire _19398_;
 wire _19399_;
 wire _19400_;
 wire _19401_;
 wire _19402_;
 wire _19403_;
 wire _19404_;
 wire _19405_;
 wire _19406_;
 wire _19407_;
 wire _19408_;
 wire _19409_;
 wire _19410_;
 wire _19411_;
 wire _19412_;
 wire _19413_;
 wire _19414_;
 wire _19415_;
 wire _19416_;
 wire _19417_;
 wire _19418_;
 wire _19419_;
 wire _19420_;
 wire _19421_;
 wire _19422_;
 wire _19423_;
 wire _19424_;
 wire _19425_;
 wire _19426_;
 wire _19427_;
 wire _19428_;
 wire _19429_;
 wire _19430_;
 wire _19431_;
 wire _19432_;
 wire _19433_;
 wire _19434_;
 wire _19435_;
 wire _19436_;
 wire _19437_;
 wire _19438_;
 wire _19439_;
 wire _19440_;
 wire _19441_;
 wire _19442_;
 wire _19443_;
 wire _19444_;
 wire _19445_;
 wire _19446_;
 wire _19447_;
 wire _19448_;
 wire _19449_;
 wire _19450_;
 wire _19451_;
 wire _19452_;
 wire _19453_;
 wire _19454_;
 wire _19455_;
 wire _19456_;
 wire _19457_;
 wire _19458_;
 wire _19459_;
 wire _19460_;
 wire _19461_;
 wire _19462_;
 wire _19463_;
 wire _19464_;
 wire _19465_;
 wire _19466_;
 wire _19467_;
 wire _19468_;
 wire _19469_;
 wire _19470_;
 wire _19471_;
 wire _19472_;
 wire _19473_;
 wire _19474_;
 wire _19475_;
 wire _19476_;
 wire _19477_;
 wire _19478_;
 wire _19479_;
 wire _19480_;
 wire _19481_;
 wire _19482_;
 wire _19483_;
 wire _19484_;
 wire _19485_;
 wire _19486_;
 wire _19487_;
 wire _19488_;
 wire _19489_;
 wire _19490_;
 wire _19491_;
 wire _19492_;
 wire _19493_;
 wire _19494_;
 wire _19495_;
 wire _19496_;
 wire _19497_;
 wire _19498_;
 wire _19499_;
 wire _19500_;
 wire _19501_;
 wire _19502_;
 wire _19503_;
 wire _19504_;
 wire _19505_;
 wire _19506_;
 wire _19507_;
 wire _19508_;
 wire _19509_;
 wire _19510_;
 wire _19511_;
 wire _19512_;
 wire _19513_;
 wire _19514_;
 wire _19515_;
 wire _19516_;
 wire _19517_;
 wire _19518_;
 wire _19519_;
 wire _19520_;
 wire _19521_;
 wire _19522_;
 wire _19523_;
 wire _19524_;
 wire _19525_;
 wire _19526_;
 wire _19527_;
 wire _19528_;
 wire _19529_;
 wire _19530_;
 wire _19531_;
 wire _19532_;
 wire _19533_;
 wire _19534_;
 wire _19535_;
 wire _19536_;
 wire _19537_;
 wire _19538_;
 wire _19539_;
 wire _19540_;
 wire _19541_;
 wire _19542_;
 wire _19543_;
 wire _19544_;
 wire _19545_;
 wire _19546_;
 wire _19547_;
 wire _19548_;
 wire _19549_;
 wire _19550_;
 wire _19551_;
 wire _19552_;
 wire _19553_;
 wire _19554_;
 wire _19555_;
 wire _19556_;
 wire _19557_;
 wire _19558_;
 wire _19559_;
 wire _19560_;
 wire _19561_;
 wire _19562_;
 wire _19563_;
 wire _19564_;
 wire _19565_;
 wire _19566_;
 wire _19567_;
 wire _19568_;
 wire _19569_;
 wire _19570_;
 wire _19571_;
 wire _19572_;
 wire _19573_;
 wire _19574_;
 wire _19575_;
 wire _19576_;
 wire _19577_;
 wire _19578_;
 wire _19579_;
 wire _19580_;
 wire _19581_;
 wire _19582_;
 wire _19583_;
 wire _19584_;
 wire _19585_;
 wire _19586_;
 wire _19587_;
 wire _19588_;
 wire _19589_;
 wire _19590_;
 wire _19591_;
 wire _19592_;
 wire _19593_;
 wire _19594_;
 wire _19595_;
 wire _19596_;
 wire _19597_;
 wire _19598_;
 wire _19599_;
 wire _19600_;
 wire _19601_;
 wire _19602_;
 wire _19603_;
 wire _19604_;
 wire _19605_;
 wire _19606_;
 wire _19607_;
 wire _19608_;
 wire _19609_;
 wire _19610_;
 wire _19611_;
 wire _19612_;
 wire _19613_;
 wire _19614_;
 wire _19615_;
 wire _19616_;
 wire _19617_;
 wire _19618_;
 wire _19619_;
 wire _19620_;
 wire _19621_;
 wire _19622_;
 wire _19623_;
 wire _19624_;
 wire _19625_;
 wire _19626_;
 wire _19627_;
 wire _19628_;
 wire _19629_;
 wire _19630_;
 wire _19631_;
 wire _19632_;
 wire _19633_;
 wire _19634_;
 wire _19635_;
 wire _19636_;
 wire _19637_;
 wire _19638_;
 wire _19639_;
 wire _19640_;
 wire _19641_;
 wire _19642_;
 wire _19643_;
 wire _19644_;
 wire _19645_;
 wire _19646_;
 wire _19647_;
 wire _19648_;
 wire _19649_;
 wire _19650_;
 wire _19651_;
 wire _19652_;
 wire _19653_;
 wire _19654_;
 wire _19655_;
 wire _19656_;
 wire _19657_;
 wire _19658_;
 wire _19659_;
 wire _19660_;
 wire _19661_;
 wire _19662_;
 wire _19663_;
 wire _19664_;
 wire _19665_;
 wire _19666_;
 wire _19667_;
 wire _19668_;
 wire _19669_;
 wire _19670_;
 wire _19671_;
 wire _19672_;
 wire _19673_;
 wire _19674_;
 wire _19675_;
 wire _19676_;
 wire _19677_;
 wire _19678_;
 wire _19679_;
 wire _19680_;
 wire _19681_;
 wire _19682_;
 wire _19683_;
 wire _19684_;
 wire _19685_;
 wire _19686_;
 wire _19687_;
 wire _19688_;
 wire _19689_;
 wire _19690_;
 wire _19691_;
 wire _19692_;
 wire _19693_;
 wire _19694_;
 wire _19695_;
 wire _19696_;
 wire _19697_;
 wire _19698_;
 wire _19699_;
 wire _19700_;
 wire _19701_;
 wire _19702_;
 wire _19703_;
 wire _19704_;
 wire _19705_;
 wire _19706_;
 wire _19707_;
 wire _19708_;
 wire _19709_;
 wire _19710_;
 wire _19711_;
 wire _19712_;
 wire _19713_;
 wire _19714_;
 wire _19715_;
 wire _19716_;
 wire _19717_;
 wire _19718_;
 wire _19719_;
 wire _19720_;
 wire _19721_;
 wire _19722_;
 wire _19723_;
 wire _19724_;
 wire _19725_;
 wire _19726_;
 wire _19727_;
 wire _19728_;
 wire _19729_;
 wire _19730_;
 wire _19731_;
 wire _19732_;
 wire _19733_;
 wire _19734_;
 wire _19735_;
 wire _19736_;
 wire _19737_;
 wire _19738_;
 wire _19739_;
 wire _19740_;
 wire _19741_;
 wire _19742_;
 wire _19743_;
 wire _19744_;
 wire _19745_;
 wire _19746_;
 wire _19747_;
 wire _19748_;
 wire _19749_;
 wire _19750_;
 wire _19751_;
 wire _19752_;
 wire _19753_;
 wire _19754_;
 wire _19755_;
 wire _19756_;
 wire _19757_;
 wire _19758_;
 wire _19759_;
 wire _19760_;
 wire _19761_;
 wire _19762_;
 wire _19763_;
 wire _19764_;
 wire _19765_;
 wire _19766_;
 wire _19767_;
 wire _19768_;
 wire _19769_;
 wire _19770_;
 wire _19771_;
 wire _19772_;
 wire _19773_;
 wire _19774_;
 wire _19775_;
 wire _19776_;
 wire _19777_;
 wire _19778_;
 wire _19779_;
 wire _19780_;
 wire _19781_;
 wire _19782_;
 wire _19783_;
 wire _19784_;
 wire _19785_;
 wire _19786_;
 wire _19787_;
 wire _19788_;
 wire _19789_;
 wire _19790_;
 wire _19791_;
 wire _19792_;
 wire _19793_;
 wire _19794_;
 wire _19795_;
 wire _19796_;
 wire _19797_;
 wire _19798_;
 wire _19799_;
 wire _19800_;
 wire _19801_;
 wire _19802_;
 wire _19803_;
 wire _19804_;
 wire _19805_;
 wire _19806_;
 wire _19807_;
 wire _19808_;
 wire _19809_;
 wire _19810_;
 wire _19811_;
 wire _19812_;
 wire _19813_;
 wire _19814_;
 wire _19815_;
 wire _19816_;
 wire _19817_;
 wire _19818_;
 wire _19819_;
 wire _19820_;
 wire _19821_;
 wire _19822_;
 wire _19823_;
 wire _19824_;
 wire _19825_;
 wire _19826_;
 wire _19827_;
 wire _19828_;
 wire _19829_;
 wire _19830_;
 wire _19831_;
 wire _19832_;
 wire _19833_;
 wire _19834_;
 wire _19835_;
 wire _19836_;
 wire _19837_;
 wire _19838_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire accepting;
 wire \byte_cnt[0] ;
 wire \byte_cnt[1] ;
 wire \byte_cnt[2] ;
 wire \byte_cnt[3] ;
 wire \byte_cnt[4] ;
 wire \inv_cycles[0] ;
 wire \inv_cycles[1] ;
 wire \inv_cycles[2] ;
 wire \inv_cycles[3] ;
 wire \inv_cycles[4] ;
 wire \inv_cycles[5] ;
 wire \inv_cycles[6] ;
 wire \inv_cycles[7] ;
 wire \inv_cycles[8] ;
 wire \inv_cycles[9] ;
 wire inv_done;
 wire inv_go;
 wire \inv_result[0] ;
 wire \inv_result[100] ;
 wire \inv_result[101] ;
 wire \inv_result[102] ;
 wire \inv_result[103] ;
 wire \inv_result[104] ;
 wire \inv_result[105] ;
 wire \inv_result[106] ;
 wire \inv_result[107] ;
 wire \inv_result[108] ;
 wire \inv_result[109] ;
 wire \inv_result[10] ;
 wire \inv_result[110] ;
 wire \inv_result[111] ;
 wire \inv_result[112] ;
 wire \inv_result[113] ;
 wire \inv_result[114] ;
 wire \inv_result[115] ;
 wire \inv_result[116] ;
 wire \inv_result[117] ;
 wire \inv_result[118] ;
 wire \inv_result[119] ;
 wire \inv_result[11] ;
 wire \inv_result[120] ;
 wire \inv_result[121] ;
 wire \inv_result[122] ;
 wire \inv_result[123] ;
 wire \inv_result[124] ;
 wire \inv_result[125] ;
 wire \inv_result[126] ;
 wire \inv_result[127] ;
 wire \inv_result[128] ;
 wire \inv_result[129] ;
 wire \inv_result[12] ;
 wire \inv_result[130] ;
 wire \inv_result[131] ;
 wire \inv_result[132] ;
 wire \inv_result[133] ;
 wire \inv_result[134] ;
 wire \inv_result[135] ;
 wire \inv_result[136] ;
 wire \inv_result[137] ;
 wire \inv_result[138] ;
 wire \inv_result[139] ;
 wire \inv_result[13] ;
 wire \inv_result[140] ;
 wire \inv_result[141] ;
 wire \inv_result[142] ;
 wire \inv_result[143] ;
 wire \inv_result[144] ;
 wire \inv_result[145] ;
 wire \inv_result[146] ;
 wire \inv_result[147] ;
 wire \inv_result[148] ;
 wire \inv_result[149] ;
 wire \inv_result[14] ;
 wire \inv_result[150] ;
 wire \inv_result[151] ;
 wire \inv_result[152] ;
 wire \inv_result[153] ;
 wire \inv_result[154] ;
 wire \inv_result[155] ;
 wire \inv_result[156] ;
 wire \inv_result[157] ;
 wire \inv_result[158] ;
 wire \inv_result[159] ;
 wire \inv_result[15] ;
 wire \inv_result[160] ;
 wire \inv_result[161] ;
 wire \inv_result[162] ;
 wire \inv_result[163] ;
 wire \inv_result[164] ;
 wire \inv_result[165] ;
 wire \inv_result[166] ;
 wire \inv_result[167] ;
 wire \inv_result[168] ;
 wire \inv_result[169] ;
 wire \inv_result[16] ;
 wire \inv_result[170] ;
 wire \inv_result[171] ;
 wire \inv_result[172] ;
 wire \inv_result[173] ;
 wire \inv_result[174] ;
 wire \inv_result[175] ;
 wire \inv_result[176] ;
 wire \inv_result[177] ;
 wire \inv_result[178] ;
 wire \inv_result[179] ;
 wire \inv_result[17] ;
 wire \inv_result[180] ;
 wire \inv_result[181] ;
 wire \inv_result[182] ;
 wire \inv_result[183] ;
 wire \inv_result[184] ;
 wire \inv_result[185] ;
 wire \inv_result[186] ;
 wire \inv_result[187] ;
 wire \inv_result[188] ;
 wire \inv_result[189] ;
 wire \inv_result[18] ;
 wire \inv_result[190] ;
 wire \inv_result[191] ;
 wire \inv_result[192] ;
 wire \inv_result[193] ;
 wire \inv_result[194] ;
 wire \inv_result[195] ;
 wire \inv_result[196] ;
 wire \inv_result[197] ;
 wire \inv_result[198] ;
 wire \inv_result[199] ;
 wire \inv_result[19] ;
 wire \inv_result[1] ;
 wire \inv_result[200] ;
 wire \inv_result[201] ;
 wire \inv_result[202] ;
 wire \inv_result[203] ;
 wire \inv_result[204] ;
 wire \inv_result[205] ;
 wire \inv_result[206] ;
 wire \inv_result[207] ;
 wire \inv_result[208] ;
 wire \inv_result[209] ;
 wire \inv_result[20] ;
 wire \inv_result[210] ;
 wire \inv_result[211] ;
 wire \inv_result[212] ;
 wire \inv_result[213] ;
 wire \inv_result[214] ;
 wire \inv_result[215] ;
 wire \inv_result[216] ;
 wire \inv_result[217] ;
 wire \inv_result[218] ;
 wire \inv_result[219] ;
 wire \inv_result[21] ;
 wire \inv_result[220] ;
 wire \inv_result[221] ;
 wire \inv_result[222] ;
 wire \inv_result[223] ;
 wire \inv_result[224] ;
 wire \inv_result[225] ;
 wire \inv_result[226] ;
 wire \inv_result[227] ;
 wire \inv_result[228] ;
 wire \inv_result[229] ;
 wire \inv_result[22] ;
 wire \inv_result[230] ;
 wire \inv_result[231] ;
 wire \inv_result[232] ;
 wire \inv_result[233] ;
 wire \inv_result[234] ;
 wire \inv_result[235] ;
 wire \inv_result[236] ;
 wire \inv_result[237] ;
 wire \inv_result[238] ;
 wire \inv_result[239] ;
 wire \inv_result[23] ;
 wire \inv_result[240] ;
 wire \inv_result[241] ;
 wire \inv_result[242] ;
 wire \inv_result[243] ;
 wire \inv_result[244] ;
 wire \inv_result[245] ;
 wire \inv_result[246] ;
 wire \inv_result[247] ;
 wire \inv_result[248] ;
 wire \inv_result[249] ;
 wire \inv_result[24] ;
 wire \inv_result[250] ;
 wire \inv_result[251] ;
 wire \inv_result[252] ;
 wire \inv_result[253] ;
 wire \inv_result[254] ;
 wire \inv_result[255] ;
 wire \inv_result[25] ;
 wire \inv_result[26] ;
 wire \inv_result[27] ;
 wire \inv_result[28] ;
 wire \inv_result[29] ;
 wire \inv_result[2] ;
 wire \inv_result[30] ;
 wire \inv_result[31] ;
 wire \inv_result[32] ;
 wire \inv_result[33] ;
 wire \inv_result[34] ;
 wire \inv_result[35] ;
 wire \inv_result[36] ;
 wire \inv_result[37] ;
 wire \inv_result[38] ;
 wire \inv_result[39] ;
 wire \inv_result[3] ;
 wire \inv_result[40] ;
 wire \inv_result[41] ;
 wire \inv_result[42] ;
 wire \inv_result[43] ;
 wire \inv_result[44] ;
 wire \inv_result[45] ;
 wire \inv_result[46] ;
 wire \inv_result[47] ;
 wire \inv_result[48] ;
 wire \inv_result[49] ;
 wire \inv_result[4] ;
 wire \inv_result[50] ;
 wire \inv_result[51] ;
 wire \inv_result[52] ;
 wire \inv_result[53] ;
 wire \inv_result[54] ;
 wire \inv_result[55] ;
 wire \inv_result[56] ;
 wire \inv_result[57] ;
 wire \inv_result[58] ;
 wire \inv_result[59] ;
 wire \inv_result[5] ;
 wire \inv_result[60] ;
 wire \inv_result[61] ;
 wire \inv_result[62] ;
 wire \inv_result[63] ;
 wire \inv_result[64] ;
 wire \inv_result[65] ;
 wire \inv_result[66] ;
 wire \inv_result[67] ;
 wire \inv_result[68] ;
 wire \inv_result[69] ;
 wire \inv_result[6] ;
 wire \inv_result[70] ;
 wire \inv_result[71] ;
 wire \inv_result[72] ;
 wire \inv_result[73] ;
 wire \inv_result[74] ;
 wire \inv_result[75] ;
 wire \inv_result[76] ;
 wire \inv_result[77] ;
 wire \inv_result[78] ;
 wire \inv_result[79] ;
 wire \inv_result[7] ;
 wire \inv_result[80] ;
 wire \inv_result[81] ;
 wire \inv_result[82] ;
 wire \inv_result[83] ;
 wire \inv_result[84] ;
 wire \inv_result[85] ;
 wire \inv_result[86] ;
 wire \inv_result[87] ;
 wire \inv_result[88] ;
 wire \inv_result[89] ;
 wire \inv_result[8] ;
 wire \inv_result[90] ;
 wire \inv_result[91] ;
 wire \inv_result[92] ;
 wire \inv_result[93] ;
 wire \inv_result[94] ;
 wire \inv_result[95] ;
 wire \inv_result[96] ;
 wire \inv_result[97] ;
 wire \inv_result[98] ;
 wire \inv_result[99] ;
 wire \inv_result[9] ;
 wire next_loaded;
 wire pipe_pending;
 wire rd_prev;
 wire \shift_reg[0] ;
 wire \shift_reg[100] ;
 wire \shift_reg[101] ;
 wire \shift_reg[102] ;
 wire \shift_reg[103] ;
 wire \shift_reg[104] ;
 wire \shift_reg[105] ;
 wire \shift_reg[106] ;
 wire \shift_reg[107] ;
 wire \shift_reg[108] ;
 wire \shift_reg[109] ;
 wire \shift_reg[10] ;
 wire \shift_reg[110] ;
 wire \shift_reg[111] ;
 wire \shift_reg[112] ;
 wire \shift_reg[113] ;
 wire \shift_reg[114] ;
 wire \shift_reg[115] ;
 wire \shift_reg[116] ;
 wire \shift_reg[117] ;
 wire \shift_reg[118] ;
 wire \shift_reg[119] ;
 wire \shift_reg[11] ;
 wire \shift_reg[120] ;
 wire \shift_reg[121] ;
 wire \shift_reg[122] ;
 wire \shift_reg[123] ;
 wire \shift_reg[124] ;
 wire \shift_reg[125] ;
 wire \shift_reg[126] ;
 wire \shift_reg[127] ;
 wire \shift_reg[128] ;
 wire \shift_reg[129] ;
 wire \shift_reg[12] ;
 wire \shift_reg[130] ;
 wire \shift_reg[131] ;
 wire \shift_reg[132] ;
 wire \shift_reg[133] ;
 wire \shift_reg[134] ;
 wire \shift_reg[135] ;
 wire \shift_reg[136] ;
 wire \shift_reg[137] ;
 wire \shift_reg[138] ;
 wire \shift_reg[139] ;
 wire \shift_reg[13] ;
 wire \shift_reg[140] ;
 wire \shift_reg[141] ;
 wire \shift_reg[142] ;
 wire \shift_reg[143] ;
 wire \shift_reg[144] ;
 wire \shift_reg[145] ;
 wire \shift_reg[146] ;
 wire \shift_reg[147] ;
 wire \shift_reg[148] ;
 wire \shift_reg[149] ;
 wire \shift_reg[14] ;
 wire \shift_reg[150] ;
 wire \shift_reg[151] ;
 wire \shift_reg[152] ;
 wire \shift_reg[153] ;
 wire \shift_reg[154] ;
 wire \shift_reg[155] ;
 wire \shift_reg[156] ;
 wire \shift_reg[157] ;
 wire \shift_reg[158] ;
 wire \shift_reg[159] ;
 wire \shift_reg[15] ;
 wire \shift_reg[160] ;
 wire \shift_reg[161] ;
 wire \shift_reg[162] ;
 wire \shift_reg[163] ;
 wire \shift_reg[164] ;
 wire \shift_reg[165] ;
 wire \shift_reg[166] ;
 wire \shift_reg[167] ;
 wire \shift_reg[168] ;
 wire \shift_reg[169] ;
 wire \shift_reg[16] ;
 wire \shift_reg[170] ;
 wire \shift_reg[171] ;
 wire \shift_reg[172] ;
 wire \shift_reg[173] ;
 wire \shift_reg[174] ;
 wire \shift_reg[175] ;
 wire \shift_reg[176] ;
 wire \shift_reg[177] ;
 wire \shift_reg[178] ;
 wire \shift_reg[179] ;
 wire \shift_reg[17] ;
 wire \shift_reg[180] ;
 wire \shift_reg[181] ;
 wire \shift_reg[182] ;
 wire \shift_reg[183] ;
 wire \shift_reg[184] ;
 wire \shift_reg[185] ;
 wire \shift_reg[186] ;
 wire \shift_reg[187] ;
 wire \shift_reg[188] ;
 wire \shift_reg[189] ;
 wire \shift_reg[18] ;
 wire \shift_reg[190] ;
 wire \shift_reg[191] ;
 wire \shift_reg[192] ;
 wire \shift_reg[193] ;
 wire \shift_reg[194] ;
 wire \shift_reg[195] ;
 wire \shift_reg[196] ;
 wire \shift_reg[197] ;
 wire \shift_reg[198] ;
 wire \shift_reg[199] ;
 wire \shift_reg[19] ;
 wire \shift_reg[1] ;
 wire \shift_reg[200] ;
 wire \shift_reg[201] ;
 wire \shift_reg[202] ;
 wire \shift_reg[203] ;
 wire \shift_reg[204] ;
 wire \shift_reg[205] ;
 wire \shift_reg[206] ;
 wire \shift_reg[207] ;
 wire \shift_reg[208] ;
 wire \shift_reg[209] ;
 wire \shift_reg[20] ;
 wire \shift_reg[210] ;
 wire \shift_reg[211] ;
 wire \shift_reg[212] ;
 wire \shift_reg[213] ;
 wire \shift_reg[214] ;
 wire \shift_reg[215] ;
 wire \shift_reg[216] ;
 wire \shift_reg[217] ;
 wire \shift_reg[218] ;
 wire \shift_reg[219] ;
 wire \shift_reg[21] ;
 wire \shift_reg[220] ;
 wire \shift_reg[221] ;
 wire \shift_reg[222] ;
 wire \shift_reg[223] ;
 wire \shift_reg[224] ;
 wire \shift_reg[225] ;
 wire \shift_reg[226] ;
 wire \shift_reg[227] ;
 wire \shift_reg[228] ;
 wire \shift_reg[229] ;
 wire \shift_reg[22] ;
 wire \shift_reg[230] ;
 wire \shift_reg[231] ;
 wire \shift_reg[232] ;
 wire \shift_reg[233] ;
 wire \shift_reg[234] ;
 wire \shift_reg[235] ;
 wire \shift_reg[236] ;
 wire \shift_reg[237] ;
 wire \shift_reg[238] ;
 wire \shift_reg[239] ;
 wire \shift_reg[23] ;
 wire \shift_reg[240] ;
 wire \shift_reg[241] ;
 wire \shift_reg[242] ;
 wire \shift_reg[243] ;
 wire \shift_reg[244] ;
 wire \shift_reg[245] ;
 wire \shift_reg[246] ;
 wire \shift_reg[247] ;
 wire \shift_reg[248] ;
 wire \shift_reg[249] ;
 wire \shift_reg[24] ;
 wire \shift_reg[250] ;
 wire \shift_reg[251] ;
 wire \shift_reg[252] ;
 wire \shift_reg[253] ;
 wire \shift_reg[254] ;
 wire \shift_reg[255] ;
 wire \shift_reg[256] ;
 wire \shift_reg[257] ;
 wire \shift_reg[258] ;
 wire \shift_reg[259] ;
 wire \shift_reg[25] ;
 wire \shift_reg[260] ;
 wire \shift_reg[261] ;
 wire \shift_reg[262] ;
 wire \shift_reg[263] ;
 wire \shift_reg[264] ;
 wire \shift_reg[265] ;
 wire \shift_reg[266] ;
 wire \shift_reg[267] ;
 wire \shift_reg[268] ;
 wire \shift_reg[269] ;
 wire \shift_reg[26] ;
 wire \shift_reg[270] ;
 wire \shift_reg[271] ;
 wire \shift_reg[27] ;
 wire \shift_reg[28] ;
 wire \shift_reg[29] ;
 wire \shift_reg[2] ;
 wire \shift_reg[30] ;
 wire \shift_reg[31] ;
 wire \shift_reg[32] ;
 wire \shift_reg[33] ;
 wire \shift_reg[34] ;
 wire \shift_reg[35] ;
 wire \shift_reg[36] ;
 wire \shift_reg[37] ;
 wire \shift_reg[38] ;
 wire \shift_reg[39] ;
 wire \shift_reg[3] ;
 wire \shift_reg[40] ;
 wire \shift_reg[41] ;
 wire \shift_reg[42] ;
 wire \shift_reg[43] ;
 wire \shift_reg[44] ;
 wire \shift_reg[45] ;
 wire \shift_reg[46] ;
 wire \shift_reg[47] ;
 wire \shift_reg[48] ;
 wire \shift_reg[49] ;
 wire \shift_reg[4] ;
 wire \shift_reg[50] ;
 wire \shift_reg[51] ;
 wire \shift_reg[52] ;
 wire \shift_reg[53] ;
 wire \shift_reg[54] ;
 wire \shift_reg[55] ;
 wire \shift_reg[56] ;
 wire \shift_reg[57] ;
 wire \shift_reg[58] ;
 wire \shift_reg[59] ;
 wire \shift_reg[5] ;
 wire \shift_reg[60] ;
 wire \shift_reg[61] ;
 wire \shift_reg[62] ;
 wire \shift_reg[63] ;
 wire \shift_reg[64] ;
 wire \shift_reg[65] ;
 wire \shift_reg[66] ;
 wire \shift_reg[67] ;
 wire \shift_reg[68] ;
 wire \shift_reg[69] ;
 wire \shift_reg[6] ;
 wire \shift_reg[70] ;
 wire \shift_reg[71] ;
 wire \shift_reg[72] ;
 wire \shift_reg[73] ;
 wire \shift_reg[74] ;
 wire \shift_reg[75] ;
 wire \shift_reg[76] ;
 wire \shift_reg[77] ;
 wire \shift_reg[78] ;
 wire \shift_reg[79] ;
 wire \shift_reg[7] ;
 wire \shift_reg[80] ;
 wire \shift_reg[81] ;
 wire \shift_reg[82] ;
 wire \shift_reg[83] ;
 wire \shift_reg[84] ;
 wire \shift_reg[85] ;
 wire \shift_reg[86] ;
 wire \shift_reg[87] ;
 wire \shift_reg[88] ;
 wire \shift_reg[89] ;
 wire \shift_reg[8] ;
 wire \shift_reg[90] ;
 wire \shift_reg[91] ;
 wire \shift_reg[92] ;
 wire \shift_reg[93] ;
 wire \shift_reg[94] ;
 wire \shift_reg[95] ;
 wire \shift_reg[96] ;
 wire \shift_reg[97] ;
 wire \shift_reg[98] ;
 wire \shift_reg[99] ;
 wire \shift_reg[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \u_inv.counter[0] ;
 wire \u_inv.counter[1] ;
 wire \u_inv.counter[2] ;
 wire \u_inv.counter[3] ;
 wire \u_inv.counter[4] ;
 wire \u_inv.counter[5] ;
 wire \u_inv.counter[6] ;
 wire \u_inv.counter[7] ;
 wire \u_inv.counter[8] ;
 wire \u_inv.counter[9] ;
 wire \u_inv.d_next[0] ;
 wire \u_inv.d_next[100] ;
 wire \u_inv.d_next[101] ;
 wire \u_inv.d_next[102] ;
 wire \u_inv.d_next[103] ;
 wire \u_inv.d_next[104] ;
 wire \u_inv.d_next[105] ;
 wire \u_inv.d_next[106] ;
 wire \u_inv.d_next[107] ;
 wire \u_inv.d_next[108] ;
 wire \u_inv.d_next[109] ;
 wire \u_inv.d_next[10] ;
 wire \u_inv.d_next[110] ;
 wire \u_inv.d_next[111] ;
 wire \u_inv.d_next[112] ;
 wire \u_inv.d_next[113] ;
 wire \u_inv.d_next[114] ;
 wire \u_inv.d_next[115] ;
 wire \u_inv.d_next[116] ;
 wire \u_inv.d_next[117] ;
 wire \u_inv.d_next[118] ;
 wire \u_inv.d_next[119] ;
 wire \u_inv.d_next[11] ;
 wire \u_inv.d_next[120] ;
 wire \u_inv.d_next[121] ;
 wire \u_inv.d_next[122] ;
 wire \u_inv.d_next[123] ;
 wire \u_inv.d_next[124] ;
 wire \u_inv.d_next[125] ;
 wire \u_inv.d_next[126] ;
 wire \u_inv.d_next[127] ;
 wire \u_inv.d_next[128] ;
 wire \u_inv.d_next[129] ;
 wire \u_inv.d_next[12] ;
 wire \u_inv.d_next[130] ;
 wire \u_inv.d_next[131] ;
 wire \u_inv.d_next[132] ;
 wire \u_inv.d_next[133] ;
 wire \u_inv.d_next[134] ;
 wire \u_inv.d_next[135] ;
 wire \u_inv.d_next[136] ;
 wire \u_inv.d_next[137] ;
 wire \u_inv.d_next[138] ;
 wire \u_inv.d_next[139] ;
 wire \u_inv.d_next[13] ;
 wire \u_inv.d_next[140] ;
 wire \u_inv.d_next[141] ;
 wire \u_inv.d_next[142] ;
 wire \u_inv.d_next[143] ;
 wire \u_inv.d_next[144] ;
 wire \u_inv.d_next[145] ;
 wire \u_inv.d_next[146] ;
 wire \u_inv.d_next[147] ;
 wire \u_inv.d_next[148] ;
 wire \u_inv.d_next[149] ;
 wire \u_inv.d_next[14] ;
 wire \u_inv.d_next[150] ;
 wire \u_inv.d_next[151] ;
 wire \u_inv.d_next[152] ;
 wire \u_inv.d_next[153] ;
 wire \u_inv.d_next[154] ;
 wire \u_inv.d_next[155] ;
 wire \u_inv.d_next[156] ;
 wire \u_inv.d_next[157] ;
 wire \u_inv.d_next[158] ;
 wire \u_inv.d_next[159] ;
 wire \u_inv.d_next[15] ;
 wire \u_inv.d_next[160] ;
 wire \u_inv.d_next[161] ;
 wire \u_inv.d_next[162] ;
 wire \u_inv.d_next[163] ;
 wire \u_inv.d_next[164] ;
 wire \u_inv.d_next[165] ;
 wire \u_inv.d_next[166] ;
 wire \u_inv.d_next[167] ;
 wire \u_inv.d_next[168] ;
 wire \u_inv.d_next[169] ;
 wire \u_inv.d_next[16] ;
 wire \u_inv.d_next[170] ;
 wire \u_inv.d_next[171] ;
 wire \u_inv.d_next[172] ;
 wire \u_inv.d_next[173] ;
 wire \u_inv.d_next[174] ;
 wire \u_inv.d_next[175] ;
 wire \u_inv.d_next[176] ;
 wire \u_inv.d_next[177] ;
 wire \u_inv.d_next[178] ;
 wire \u_inv.d_next[179] ;
 wire \u_inv.d_next[17] ;
 wire \u_inv.d_next[180] ;
 wire \u_inv.d_next[181] ;
 wire \u_inv.d_next[182] ;
 wire \u_inv.d_next[183] ;
 wire \u_inv.d_next[184] ;
 wire \u_inv.d_next[185] ;
 wire \u_inv.d_next[186] ;
 wire \u_inv.d_next[187] ;
 wire \u_inv.d_next[188] ;
 wire \u_inv.d_next[189] ;
 wire \u_inv.d_next[18] ;
 wire \u_inv.d_next[190] ;
 wire \u_inv.d_next[191] ;
 wire \u_inv.d_next[192] ;
 wire \u_inv.d_next[193] ;
 wire \u_inv.d_next[194] ;
 wire \u_inv.d_next[195] ;
 wire \u_inv.d_next[196] ;
 wire \u_inv.d_next[197] ;
 wire \u_inv.d_next[198] ;
 wire \u_inv.d_next[199] ;
 wire \u_inv.d_next[19] ;
 wire \u_inv.d_next[1] ;
 wire \u_inv.d_next[200] ;
 wire \u_inv.d_next[201] ;
 wire \u_inv.d_next[202] ;
 wire \u_inv.d_next[203] ;
 wire \u_inv.d_next[204] ;
 wire \u_inv.d_next[205] ;
 wire \u_inv.d_next[206] ;
 wire \u_inv.d_next[207] ;
 wire \u_inv.d_next[208] ;
 wire \u_inv.d_next[209] ;
 wire \u_inv.d_next[20] ;
 wire \u_inv.d_next[210] ;
 wire \u_inv.d_next[211] ;
 wire \u_inv.d_next[212] ;
 wire \u_inv.d_next[213] ;
 wire \u_inv.d_next[214] ;
 wire \u_inv.d_next[215] ;
 wire \u_inv.d_next[216] ;
 wire \u_inv.d_next[217] ;
 wire \u_inv.d_next[218] ;
 wire \u_inv.d_next[219] ;
 wire \u_inv.d_next[21] ;
 wire \u_inv.d_next[220] ;
 wire \u_inv.d_next[221] ;
 wire \u_inv.d_next[222] ;
 wire \u_inv.d_next[223] ;
 wire \u_inv.d_next[224] ;
 wire \u_inv.d_next[225] ;
 wire \u_inv.d_next[226] ;
 wire \u_inv.d_next[227] ;
 wire \u_inv.d_next[228] ;
 wire \u_inv.d_next[229] ;
 wire \u_inv.d_next[22] ;
 wire \u_inv.d_next[230] ;
 wire \u_inv.d_next[231] ;
 wire \u_inv.d_next[232] ;
 wire \u_inv.d_next[233] ;
 wire \u_inv.d_next[234] ;
 wire \u_inv.d_next[235] ;
 wire \u_inv.d_next[236] ;
 wire \u_inv.d_next[237] ;
 wire \u_inv.d_next[238] ;
 wire \u_inv.d_next[239] ;
 wire \u_inv.d_next[23] ;
 wire \u_inv.d_next[240] ;
 wire \u_inv.d_next[241] ;
 wire \u_inv.d_next[242] ;
 wire \u_inv.d_next[243] ;
 wire \u_inv.d_next[244] ;
 wire \u_inv.d_next[245] ;
 wire \u_inv.d_next[246] ;
 wire \u_inv.d_next[247] ;
 wire \u_inv.d_next[248] ;
 wire \u_inv.d_next[249] ;
 wire \u_inv.d_next[24] ;
 wire \u_inv.d_next[250] ;
 wire \u_inv.d_next[251] ;
 wire \u_inv.d_next[252] ;
 wire \u_inv.d_next[253] ;
 wire \u_inv.d_next[254] ;
 wire \u_inv.d_next[255] ;
 wire \u_inv.d_next[256] ;
 wire \u_inv.d_next[25] ;
 wire \u_inv.d_next[26] ;
 wire \u_inv.d_next[27] ;
 wire \u_inv.d_next[28] ;
 wire \u_inv.d_next[29] ;
 wire \u_inv.d_next[2] ;
 wire \u_inv.d_next[30] ;
 wire \u_inv.d_next[31] ;
 wire \u_inv.d_next[32] ;
 wire \u_inv.d_next[33] ;
 wire \u_inv.d_next[34] ;
 wire \u_inv.d_next[35] ;
 wire \u_inv.d_next[36] ;
 wire \u_inv.d_next[37] ;
 wire \u_inv.d_next[38] ;
 wire \u_inv.d_next[39] ;
 wire \u_inv.d_next[3] ;
 wire \u_inv.d_next[40] ;
 wire \u_inv.d_next[41] ;
 wire \u_inv.d_next[42] ;
 wire \u_inv.d_next[43] ;
 wire \u_inv.d_next[44] ;
 wire \u_inv.d_next[45] ;
 wire \u_inv.d_next[46] ;
 wire \u_inv.d_next[47] ;
 wire \u_inv.d_next[48] ;
 wire \u_inv.d_next[49] ;
 wire \u_inv.d_next[4] ;
 wire \u_inv.d_next[50] ;
 wire \u_inv.d_next[51] ;
 wire \u_inv.d_next[52] ;
 wire \u_inv.d_next[53] ;
 wire \u_inv.d_next[54] ;
 wire \u_inv.d_next[55] ;
 wire \u_inv.d_next[56] ;
 wire \u_inv.d_next[57] ;
 wire \u_inv.d_next[58] ;
 wire \u_inv.d_next[59] ;
 wire \u_inv.d_next[5] ;
 wire \u_inv.d_next[60] ;
 wire \u_inv.d_next[61] ;
 wire \u_inv.d_next[62] ;
 wire \u_inv.d_next[63] ;
 wire \u_inv.d_next[64] ;
 wire \u_inv.d_next[65] ;
 wire \u_inv.d_next[66] ;
 wire \u_inv.d_next[67] ;
 wire \u_inv.d_next[68] ;
 wire \u_inv.d_next[69] ;
 wire \u_inv.d_next[6] ;
 wire \u_inv.d_next[70] ;
 wire \u_inv.d_next[71] ;
 wire \u_inv.d_next[72] ;
 wire \u_inv.d_next[73] ;
 wire \u_inv.d_next[74] ;
 wire \u_inv.d_next[75] ;
 wire \u_inv.d_next[76] ;
 wire \u_inv.d_next[77] ;
 wire \u_inv.d_next[78] ;
 wire \u_inv.d_next[79] ;
 wire \u_inv.d_next[7] ;
 wire \u_inv.d_next[80] ;
 wire \u_inv.d_next[81] ;
 wire \u_inv.d_next[82] ;
 wire \u_inv.d_next[83] ;
 wire \u_inv.d_next[84] ;
 wire \u_inv.d_next[85] ;
 wire \u_inv.d_next[86] ;
 wire \u_inv.d_next[87] ;
 wire \u_inv.d_next[88] ;
 wire \u_inv.d_next[89] ;
 wire \u_inv.d_next[8] ;
 wire \u_inv.d_next[90] ;
 wire \u_inv.d_next[91] ;
 wire \u_inv.d_next[92] ;
 wire \u_inv.d_next[93] ;
 wire \u_inv.d_next[94] ;
 wire \u_inv.d_next[95] ;
 wire \u_inv.d_next[96] ;
 wire \u_inv.d_next[97] ;
 wire \u_inv.d_next[98] ;
 wire \u_inv.d_next[99] ;
 wire \u_inv.d_next[9] ;
 wire \u_inv.d_reg[0] ;
 wire \u_inv.d_reg[100] ;
 wire \u_inv.d_reg[101] ;
 wire \u_inv.d_reg[102] ;
 wire \u_inv.d_reg[103] ;
 wire \u_inv.d_reg[104] ;
 wire \u_inv.d_reg[105] ;
 wire \u_inv.d_reg[106] ;
 wire \u_inv.d_reg[107] ;
 wire \u_inv.d_reg[108] ;
 wire \u_inv.d_reg[109] ;
 wire \u_inv.d_reg[10] ;
 wire \u_inv.d_reg[110] ;
 wire \u_inv.d_reg[111] ;
 wire \u_inv.d_reg[112] ;
 wire \u_inv.d_reg[113] ;
 wire \u_inv.d_reg[114] ;
 wire \u_inv.d_reg[115] ;
 wire \u_inv.d_reg[116] ;
 wire \u_inv.d_reg[117] ;
 wire \u_inv.d_reg[118] ;
 wire \u_inv.d_reg[119] ;
 wire \u_inv.d_reg[11] ;
 wire \u_inv.d_reg[120] ;
 wire \u_inv.d_reg[121] ;
 wire \u_inv.d_reg[122] ;
 wire \u_inv.d_reg[123] ;
 wire \u_inv.d_reg[124] ;
 wire \u_inv.d_reg[125] ;
 wire \u_inv.d_reg[126] ;
 wire \u_inv.d_reg[127] ;
 wire \u_inv.d_reg[128] ;
 wire \u_inv.d_reg[129] ;
 wire \u_inv.d_reg[12] ;
 wire \u_inv.d_reg[130] ;
 wire \u_inv.d_reg[131] ;
 wire \u_inv.d_reg[132] ;
 wire \u_inv.d_reg[133] ;
 wire \u_inv.d_reg[134] ;
 wire \u_inv.d_reg[135] ;
 wire \u_inv.d_reg[136] ;
 wire \u_inv.d_reg[137] ;
 wire \u_inv.d_reg[138] ;
 wire \u_inv.d_reg[139] ;
 wire \u_inv.d_reg[13] ;
 wire \u_inv.d_reg[140] ;
 wire \u_inv.d_reg[141] ;
 wire \u_inv.d_reg[142] ;
 wire \u_inv.d_reg[143] ;
 wire \u_inv.d_reg[144] ;
 wire \u_inv.d_reg[145] ;
 wire \u_inv.d_reg[146] ;
 wire \u_inv.d_reg[147] ;
 wire \u_inv.d_reg[148] ;
 wire \u_inv.d_reg[149] ;
 wire \u_inv.d_reg[14] ;
 wire \u_inv.d_reg[150] ;
 wire \u_inv.d_reg[151] ;
 wire \u_inv.d_reg[152] ;
 wire \u_inv.d_reg[153] ;
 wire \u_inv.d_reg[154] ;
 wire \u_inv.d_reg[155] ;
 wire \u_inv.d_reg[156] ;
 wire \u_inv.d_reg[157] ;
 wire \u_inv.d_reg[158] ;
 wire \u_inv.d_reg[159] ;
 wire \u_inv.d_reg[15] ;
 wire \u_inv.d_reg[160] ;
 wire \u_inv.d_reg[161] ;
 wire \u_inv.d_reg[162] ;
 wire \u_inv.d_reg[163] ;
 wire \u_inv.d_reg[164] ;
 wire \u_inv.d_reg[165] ;
 wire \u_inv.d_reg[166] ;
 wire \u_inv.d_reg[167] ;
 wire \u_inv.d_reg[168] ;
 wire \u_inv.d_reg[169] ;
 wire \u_inv.d_reg[16] ;
 wire \u_inv.d_reg[170] ;
 wire \u_inv.d_reg[171] ;
 wire \u_inv.d_reg[172] ;
 wire \u_inv.d_reg[173] ;
 wire \u_inv.d_reg[174] ;
 wire \u_inv.d_reg[175] ;
 wire \u_inv.d_reg[176] ;
 wire \u_inv.d_reg[177] ;
 wire \u_inv.d_reg[178] ;
 wire \u_inv.d_reg[179] ;
 wire \u_inv.d_reg[17] ;
 wire \u_inv.d_reg[180] ;
 wire \u_inv.d_reg[181] ;
 wire \u_inv.d_reg[182] ;
 wire \u_inv.d_reg[183] ;
 wire \u_inv.d_reg[184] ;
 wire \u_inv.d_reg[185] ;
 wire \u_inv.d_reg[186] ;
 wire \u_inv.d_reg[187] ;
 wire \u_inv.d_reg[188] ;
 wire \u_inv.d_reg[189] ;
 wire \u_inv.d_reg[18] ;
 wire \u_inv.d_reg[190] ;
 wire \u_inv.d_reg[191] ;
 wire \u_inv.d_reg[192] ;
 wire \u_inv.d_reg[193] ;
 wire \u_inv.d_reg[194] ;
 wire \u_inv.d_reg[195] ;
 wire \u_inv.d_reg[196] ;
 wire \u_inv.d_reg[197] ;
 wire \u_inv.d_reg[198] ;
 wire \u_inv.d_reg[199] ;
 wire \u_inv.d_reg[19] ;
 wire \u_inv.d_reg[1] ;
 wire \u_inv.d_reg[200] ;
 wire \u_inv.d_reg[201] ;
 wire \u_inv.d_reg[202] ;
 wire \u_inv.d_reg[203] ;
 wire \u_inv.d_reg[204] ;
 wire \u_inv.d_reg[205] ;
 wire \u_inv.d_reg[206] ;
 wire \u_inv.d_reg[207] ;
 wire \u_inv.d_reg[208] ;
 wire \u_inv.d_reg[209] ;
 wire \u_inv.d_reg[20] ;
 wire \u_inv.d_reg[210] ;
 wire \u_inv.d_reg[211] ;
 wire \u_inv.d_reg[212] ;
 wire \u_inv.d_reg[213] ;
 wire \u_inv.d_reg[214] ;
 wire \u_inv.d_reg[215] ;
 wire \u_inv.d_reg[216] ;
 wire \u_inv.d_reg[217] ;
 wire \u_inv.d_reg[218] ;
 wire \u_inv.d_reg[219] ;
 wire \u_inv.d_reg[21] ;
 wire \u_inv.d_reg[220] ;
 wire \u_inv.d_reg[221] ;
 wire \u_inv.d_reg[222] ;
 wire \u_inv.d_reg[223] ;
 wire \u_inv.d_reg[224] ;
 wire \u_inv.d_reg[225] ;
 wire \u_inv.d_reg[226] ;
 wire \u_inv.d_reg[227] ;
 wire \u_inv.d_reg[228] ;
 wire \u_inv.d_reg[229] ;
 wire \u_inv.d_reg[22] ;
 wire \u_inv.d_reg[230] ;
 wire \u_inv.d_reg[231] ;
 wire \u_inv.d_reg[232] ;
 wire \u_inv.d_reg[233] ;
 wire \u_inv.d_reg[234] ;
 wire \u_inv.d_reg[235] ;
 wire \u_inv.d_reg[236] ;
 wire \u_inv.d_reg[237] ;
 wire \u_inv.d_reg[238] ;
 wire \u_inv.d_reg[239] ;
 wire \u_inv.d_reg[23] ;
 wire \u_inv.d_reg[240] ;
 wire \u_inv.d_reg[241] ;
 wire \u_inv.d_reg[242] ;
 wire \u_inv.d_reg[243] ;
 wire \u_inv.d_reg[244] ;
 wire \u_inv.d_reg[245] ;
 wire \u_inv.d_reg[246] ;
 wire \u_inv.d_reg[247] ;
 wire \u_inv.d_reg[248] ;
 wire \u_inv.d_reg[249] ;
 wire \u_inv.d_reg[24] ;
 wire \u_inv.d_reg[250] ;
 wire \u_inv.d_reg[251] ;
 wire \u_inv.d_reg[252] ;
 wire \u_inv.d_reg[253] ;
 wire \u_inv.d_reg[254] ;
 wire \u_inv.d_reg[255] ;
 wire \u_inv.d_reg[256] ;
 wire \u_inv.d_reg[25] ;
 wire \u_inv.d_reg[26] ;
 wire \u_inv.d_reg[27] ;
 wire \u_inv.d_reg[28] ;
 wire \u_inv.d_reg[29] ;
 wire \u_inv.d_reg[2] ;
 wire \u_inv.d_reg[30] ;
 wire \u_inv.d_reg[31] ;
 wire \u_inv.d_reg[32] ;
 wire \u_inv.d_reg[33] ;
 wire \u_inv.d_reg[34] ;
 wire \u_inv.d_reg[35] ;
 wire \u_inv.d_reg[36] ;
 wire \u_inv.d_reg[37] ;
 wire \u_inv.d_reg[38] ;
 wire \u_inv.d_reg[39] ;
 wire \u_inv.d_reg[3] ;
 wire \u_inv.d_reg[40] ;
 wire \u_inv.d_reg[41] ;
 wire \u_inv.d_reg[42] ;
 wire \u_inv.d_reg[43] ;
 wire \u_inv.d_reg[44] ;
 wire \u_inv.d_reg[45] ;
 wire \u_inv.d_reg[46] ;
 wire \u_inv.d_reg[47] ;
 wire \u_inv.d_reg[48] ;
 wire \u_inv.d_reg[49] ;
 wire \u_inv.d_reg[4] ;
 wire \u_inv.d_reg[50] ;
 wire \u_inv.d_reg[51] ;
 wire \u_inv.d_reg[52] ;
 wire \u_inv.d_reg[53] ;
 wire \u_inv.d_reg[54] ;
 wire \u_inv.d_reg[55] ;
 wire \u_inv.d_reg[56] ;
 wire \u_inv.d_reg[57] ;
 wire \u_inv.d_reg[58] ;
 wire \u_inv.d_reg[59] ;
 wire \u_inv.d_reg[5] ;
 wire \u_inv.d_reg[60] ;
 wire \u_inv.d_reg[61] ;
 wire \u_inv.d_reg[62] ;
 wire \u_inv.d_reg[63] ;
 wire \u_inv.d_reg[64] ;
 wire \u_inv.d_reg[65] ;
 wire \u_inv.d_reg[66] ;
 wire \u_inv.d_reg[67] ;
 wire \u_inv.d_reg[68] ;
 wire \u_inv.d_reg[69] ;
 wire \u_inv.d_reg[6] ;
 wire \u_inv.d_reg[70] ;
 wire \u_inv.d_reg[71] ;
 wire \u_inv.d_reg[72] ;
 wire \u_inv.d_reg[73] ;
 wire \u_inv.d_reg[74] ;
 wire \u_inv.d_reg[75] ;
 wire \u_inv.d_reg[76] ;
 wire \u_inv.d_reg[77] ;
 wire \u_inv.d_reg[78] ;
 wire \u_inv.d_reg[79] ;
 wire \u_inv.d_reg[7] ;
 wire \u_inv.d_reg[80] ;
 wire \u_inv.d_reg[81] ;
 wire \u_inv.d_reg[82] ;
 wire \u_inv.d_reg[83] ;
 wire \u_inv.d_reg[84] ;
 wire \u_inv.d_reg[85] ;
 wire \u_inv.d_reg[86] ;
 wire \u_inv.d_reg[87] ;
 wire \u_inv.d_reg[88] ;
 wire \u_inv.d_reg[89] ;
 wire \u_inv.d_reg[8] ;
 wire \u_inv.d_reg[90] ;
 wire \u_inv.d_reg[91] ;
 wire \u_inv.d_reg[92] ;
 wire \u_inv.d_reg[93] ;
 wire \u_inv.d_reg[94] ;
 wire \u_inv.d_reg[95] ;
 wire \u_inv.d_reg[96] ;
 wire \u_inv.d_reg[97] ;
 wire \u_inv.d_reg[98] ;
 wire \u_inv.d_reg[99] ;
 wire \u_inv.d_reg[9] ;
 wire \u_inv.delta_double[0] ;
 wire \u_inv.delta_reg[1] ;
 wire \u_inv.delta_reg[2] ;
 wire \u_inv.delta_reg[3] ;
 wire \u_inv.delta_reg[4] ;
 wire \u_inv.delta_reg[5] ;
 wire \u_inv.delta_reg[6] ;
 wire \u_inv.delta_reg[7] ;
 wire \u_inv.delta_reg[8] ;
 wire \u_inv.delta_reg[9] ;
 wire \u_inv.f_next[0] ;
 wire \u_inv.f_next[100] ;
 wire \u_inv.f_next[101] ;
 wire \u_inv.f_next[102] ;
 wire \u_inv.f_next[103] ;
 wire \u_inv.f_next[104] ;
 wire \u_inv.f_next[105] ;
 wire \u_inv.f_next[106] ;
 wire \u_inv.f_next[107] ;
 wire \u_inv.f_next[108] ;
 wire \u_inv.f_next[109] ;
 wire \u_inv.f_next[10] ;
 wire \u_inv.f_next[110] ;
 wire \u_inv.f_next[111] ;
 wire \u_inv.f_next[112] ;
 wire \u_inv.f_next[113] ;
 wire \u_inv.f_next[114] ;
 wire \u_inv.f_next[115] ;
 wire \u_inv.f_next[116] ;
 wire \u_inv.f_next[117] ;
 wire \u_inv.f_next[118] ;
 wire \u_inv.f_next[119] ;
 wire \u_inv.f_next[11] ;
 wire \u_inv.f_next[120] ;
 wire \u_inv.f_next[121] ;
 wire \u_inv.f_next[122] ;
 wire \u_inv.f_next[123] ;
 wire \u_inv.f_next[124] ;
 wire \u_inv.f_next[125] ;
 wire \u_inv.f_next[126] ;
 wire \u_inv.f_next[127] ;
 wire \u_inv.f_next[128] ;
 wire \u_inv.f_next[129] ;
 wire \u_inv.f_next[12] ;
 wire \u_inv.f_next[130] ;
 wire \u_inv.f_next[131] ;
 wire \u_inv.f_next[132] ;
 wire \u_inv.f_next[133] ;
 wire \u_inv.f_next[134] ;
 wire \u_inv.f_next[135] ;
 wire \u_inv.f_next[136] ;
 wire \u_inv.f_next[137] ;
 wire \u_inv.f_next[138] ;
 wire \u_inv.f_next[139] ;
 wire \u_inv.f_next[13] ;
 wire \u_inv.f_next[140] ;
 wire \u_inv.f_next[141] ;
 wire \u_inv.f_next[142] ;
 wire \u_inv.f_next[143] ;
 wire \u_inv.f_next[144] ;
 wire \u_inv.f_next[145] ;
 wire \u_inv.f_next[146] ;
 wire \u_inv.f_next[147] ;
 wire \u_inv.f_next[148] ;
 wire \u_inv.f_next[149] ;
 wire \u_inv.f_next[14] ;
 wire \u_inv.f_next[150] ;
 wire \u_inv.f_next[151] ;
 wire \u_inv.f_next[152] ;
 wire \u_inv.f_next[153] ;
 wire \u_inv.f_next[154] ;
 wire \u_inv.f_next[155] ;
 wire \u_inv.f_next[156] ;
 wire \u_inv.f_next[157] ;
 wire \u_inv.f_next[158] ;
 wire \u_inv.f_next[159] ;
 wire \u_inv.f_next[15] ;
 wire \u_inv.f_next[160] ;
 wire \u_inv.f_next[161] ;
 wire \u_inv.f_next[162] ;
 wire \u_inv.f_next[163] ;
 wire \u_inv.f_next[164] ;
 wire \u_inv.f_next[165] ;
 wire \u_inv.f_next[166] ;
 wire \u_inv.f_next[167] ;
 wire \u_inv.f_next[168] ;
 wire \u_inv.f_next[169] ;
 wire \u_inv.f_next[16] ;
 wire \u_inv.f_next[170] ;
 wire \u_inv.f_next[171] ;
 wire \u_inv.f_next[172] ;
 wire \u_inv.f_next[173] ;
 wire \u_inv.f_next[174] ;
 wire \u_inv.f_next[175] ;
 wire \u_inv.f_next[176] ;
 wire \u_inv.f_next[177] ;
 wire \u_inv.f_next[178] ;
 wire \u_inv.f_next[179] ;
 wire \u_inv.f_next[17] ;
 wire \u_inv.f_next[180] ;
 wire \u_inv.f_next[181] ;
 wire \u_inv.f_next[182] ;
 wire \u_inv.f_next[183] ;
 wire \u_inv.f_next[184] ;
 wire \u_inv.f_next[185] ;
 wire \u_inv.f_next[186] ;
 wire \u_inv.f_next[187] ;
 wire \u_inv.f_next[188] ;
 wire \u_inv.f_next[189] ;
 wire \u_inv.f_next[18] ;
 wire \u_inv.f_next[190] ;
 wire \u_inv.f_next[191] ;
 wire \u_inv.f_next[192] ;
 wire \u_inv.f_next[193] ;
 wire \u_inv.f_next[194] ;
 wire \u_inv.f_next[195] ;
 wire \u_inv.f_next[196] ;
 wire \u_inv.f_next[197] ;
 wire \u_inv.f_next[198] ;
 wire \u_inv.f_next[199] ;
 wire \u_inv.f_next[19] ;
 wire \u_inv.f_next[1] ;
 wire \u_inv.f_next[200] ;
 wire \u_inv.f_next[201] ;
 wire \u_inv.f_next[202] ;
 wire \u_inv.f_next[203] ;
 wire \u_inv.f_next[204] ;
 wire \u_inv.f_next[205] ;
 wire \u_inv.f_next[206] ;
 wire \u_inv.f_next[207] ;
 wire \u_inv.f_next[208] ;
 wire \u_inv.f_next[209] ;
 wire \u_inv.f_next[20] ;
 wire \u_inv.f_next[210] ;
 wire \u_inv.f_next[211] ;
 wire \u_inv.f_next[212] ;
 wire \u_inv.f_next[213] ;
 wire \u_inv.f_next[214] ;
 wire \u_inv.f_next[215] ;
 wire \u_inv.f_next[216] ;
 wire \u_inv.f_next[217] ;
 wire \u_inv.f_next[218] ;
 wire \u_inv.f_next[219] ;
 wire \u_inv.f_next[21] ;
 wire \u_inv.f_next[220] ;
 wire \u_inv.f_next[221] ;
 wire \u_inv.f_next[222] ;
 wire \u_inv.f_next[223] ;
 wire \u_inv.f_next[224] ;
 wire \u_inv.f_next[225] ;
 wire \u_inv.f_next[226] ;
 wire \u_inv.f_next[227] ;
 wire \u_inv.f_next[228] ;
 wire \u_inv.f_next[229] ;
 wire \u_inv.f_next[22] ;
 wire \u_inv.f_next[230] ;
 wire \u_inv.f_next[231] ;
 wire \u_inv.f_next[232] ;
 wire \u_inv.f_next[233] ;
 wire \u_inv.f_next[234] ;
 wire \u_inv.f_next[235] ;
 wire \u_inv.f_next[236] ;
 wire \u_inv.f_next[237] ;
 wire \u_inv.f_next[238] ;
 wire \u_inv.f_next[239] ;
 wire \u_inv.f_next[23] ;
 wire \u_inv.f_next[240] ;
 wire \u_inv.f_next[241] ;
 wire \u_inv.f_next[242] ;
 wire \u_inv.f_next[243] ;
 wire \u_inv.f_next[244] ;
 wire \u_inv.f_next[245] ;
 wire \u_inv.f_next[246] ;
 wire \u_inv.f_next[247] ;
 wire \u_inv.f_next[248] ;
 wire \u_inv.f_next[249] ;
 wire \u_inv.f_next[24] ;
 wire \u_inv.f_next[250] ;
 wire \u_inv.f_next[251] ;
 wire \u_inv.f_next[252] ;
 wire \u_inv.f_next[253] ;
 wire \u_inv.f_next[254] ;
 wire \u_inv.f_next[255] ;
 wire \u_inv.f_next[256] ;
 wire \u_inv.f_next[25] ;
 wire \u_inv.f_next[26] ;
 wire \u_inv.f_next[27] ;
 wire \u_inv.f_next[28] ;
 wire \u_inv.f_next[29] ;
 wire \u_inv.f_next[2] ;
 wire \u_inv.f_next[30] ;
 wire \u_inv.f_next[31] ;
 wire \u_inv.f_next[32] ;
 wire \u_inv.f_next[33] ;
 wire \u_inv.f_next[34] ;
 wire \u_inv.f_next[35] ;
 wire \u_inv.f_next[36] ;
 wire \u_inv.f_next[37] ;
 wire \u_inv.f_next[38] ;
 wire \u_inv.f_next[39] ;
 wire \u_inv.f_next[3] ;
 wire \u_inv.f_next[40] ;
 wire \u_inv.f_next[41] ;
 wire \u_inv.f_next[42] ;
 wire \u_inv.f_next[43] ;
 wire \u_inv.f_next[44] ;
 wire \u_inv.f_next[45] ;
 wire \u_inv.f_next[46] ;
 wire \u_inv.f_next[47] ;
 wire \u_inv.f_next[48] ;
 wire \u_inv.f_next[49] ;
 wire \u_inv.f_next[4] ;
 wire \u_inv.f_next[50] ;
 wire \u_inv.f_next[51] ;
 wire \u_inv.f_next[52] ;
 wire \u_inv.f_next[53] ;
 wire \u_inv.f_next[54] ;
 wire \u_inv.f_next[55] ;
 wire \u_inv.f_next[56] ;
 wire \u_inv.f_next[57] ;
 wire \u_inv.f_next[58] ;
 wire \u_inv.f_next[59] ;
 wire \u_inv.f_next[5] ;
 wire \u_inv.f_next[60] ;
 wire \u_inv.f_next[61] ;
 wire \u_inv.f_next[62] ;
 wire \u_inv.f_next[63] ;
 wire \u_inv.f_next[64] ;
 wire \u_inv.f_next[65] ;
 wire \u_inv.f_next[66] ;
 wire \u_inv.f_next[67] ;
 wire \u_inv.f_next[68] ;
 wire \u_inv.f_next[69] ;
 wire \u_inv.f_next[6] ;
 wire \u_inv.f_next[70] ;
 wire \u_inv.f_next[71] ;
 wire \u_inv.f_next[72] ;
 wire \u_inv.f_next[73] ;
 wire \u_inv.f_next[74] ;
 wire \u_inv.f_next[75] ;
 wire \u_inv.f_next[76] ;
 wire \u_inv.f_next[77] ;
 wire \u_inv.f_next[78] ;
 wire \u_inv.f_next[79] ;
 wire \u_inv.f_next[7] ;
 wire \u_inv.f_next[80] ;
 wire \u_inv.f_next[81] ;
 wire \u_inv.f_next[82] ;
 wire \u_inv.f_next[83] ;
 wire \u_inv.f_next[84] ;
 wire \u_inv.f_next[85] ;
 wire \u_inv.f_next[86] ;
 wire \u_inv.f_next[87] ;
 wire \u_inv.f_next[88] ;
 wire \u_inv.f_next[89] ;
 wire \u_inv.f_next[8] ;
 wire \u_inv.f_next[90] ;
 wire \u_inv.f_next[91] ;
 wire \u_inv.f_next[92] ;
 wire \u_inv.f_next[93] ;
 wire \u_inv.f_next[94] ;
 wire \u_inv.f_next[95] ;
 wire \u_inv.f_next[96] ;
 wire \u_inv.f_next[97] ;
 wire \u_inv.f_next[98] ;
 wire \u_inv.f_next[99] ;
 wire \u_inv.f_next[9] ;
 wire \u_inv.f_reg[0] ;
 wire \u_inv.f_reg[100] ;
 wire \u_inv.f_reg[101] ;
 wire \u_inv.f_reg[102] ;
 wire \u_inv.f_reg[103] ;
 wire \u_inv.f_reg[104] ;
 wire \u_inv.f_reg[105] ;
 wire \u_inv.f_reg[106] ;
 wire \u_inv.f_reg[107] ;
 wire \u_inv.f_reg[108] ;
 wire \u_inv.f_reg[109] ;
 wire \u_inv.f_reg[10] ;
 wire \u_inv.f_reg[110] ;
 wire \u_inv.f_reg[111] ;
 wire \u_inv.f_reg[112] ;
 wire \u_inv.f_reg[113] ;
 wire \u_inv.f_reg[114] ;
 wire \u_inv.f_reg[115] ;
 wire \u_inv.f_reg[116] ;
 wire \u_inv.f_reg[117] ;
 wire \u_inv.f_reg[118] ;
 wire \u_inv.f_reg[119] ;
 wire \u_inv.f_reg[11] ;
 wire \u_inv.f_reg[120] ;
 wire \u_inv.f_reg[121] ;
 wire \u_inv.f_reg[122] ;
 wire \u_inv.f_reg[123] ;
 wire \u_inv.f_reg[124] ;
 wire \u_inv.f_reg[125] ;
 wire \u_inv.f_reg[126] ;
 wire \u_inv.f_reg[127] ;
 wire \u_inv.f_reg[128] ;
 wire \u_inv.f_reg[129] ;
 wire \u_inv.f_reg[12] ;
 wire \u_inv.f_reg[130] ;
 wire \u_inv.f_reg[131] ;
 wire \u_inv.f_reg[132] ;
 wire \u_inv.f_reg[133] ;
 wire \u_inv.f_reg[134] ;
 wire \u_inv.f_reg[135] ;
 wire \u_inv.f_reg[136] ;
 wire \u_inv.f_reg[137] ;
 wire \u_inv.f_reg[138] ;
 wire \u_inv.f_reg[139] ;
 wire \u_inv.f_reg[13] ;
 wire \u_inv.f_reg[140] ;
 wire \u_inv.f_reg[141] ;
 wire \u_inv.f_reg[142] ;
 wire \u_inv.f_reg[143] ;
 wire \u_inv.f_reg[144] ;
 wire \u_inv.f_reg[145] ;
 wire \u_inv.f_reg[146] ;
 wire \u_inv.f_reg[147] ;
 wire \u_inv.f_reg[148] ;
 wire \u_inv.f_reg[149] ;
 wire \u_inv.f_reg[14] ;
 wire \u_inv.f_reg[150] ;
 wire \u_inv.f_reg[151] ;
 wire \u_inv.f_reg[152] ;
 wire \u_inv.f_reg[153] ;
 wire \u_inv.f_reg[154] ;
 wire \u_inv.f_reg[155] ;
 wire \u_inv.f_reg[156] ;
 wire \u_inv.f_reg[157] ;
 wire \u_inv.f_reg[158] ;
 wire \u_inv.f_reg[159] ;
 wire \u_inv.f_reg[15] ;
 wire \u_inv.f_reg[160] ;
 wire \u_inv.f_reg[161] ;
 wire \u_inv.f_reg[162] ;
 wire \u_inv.f_reg[163] ;
 wire \u_inv.f_reg[164] ;
 wire \u_inv.f_reg[165] ;
 wire \u_inv.f_reg[166] ;
 wire \u_inv.f_reg[167] ;
 wire \u_inv.f_reg[168] ;
 wire \u_inv.f_reg[169] ;
 wire \u_inv.f_reg[16] ;
 wire \u_inv.f_reg[170] ;
 wire \u_inv.f_reg[171] ;
 wire \u_inv.f_reg[172] ;
 wire \u_inv.f_reg[173] ;
 wire \u_inv.f_reg[174] ;
 wire \u_inv.f_reg[175] ;
 wire \u_inv.f_reg[176] ;
 wire \u_inv.f_reg[177] ;
 wire \u_inv.f_reg[178] ;
 wire \u_inv.f_reg[179] ;
 wire \u_inv.f_reg[17] ;
 wire \u_inv.f_reg[180] ;
 wire \u_inv.f_reg[181] ;
 wire \u_inv.f_reg[182] ;
 wire \u_inv.f_reg[183] ;
 wire \u_inv.f_reg[184] ;
 wire \u_inv.f_reg[185] ;
 wire \u_inv.f_reg[186] ;
 wire \u_inv.f_reg[187] ;
 wire \u_inv.f_reg[188] ;
 wire \u_inv.f_reg[189] ;
 wire \u_inv.f_reg[18] ;
 wire \u_inv.f_reg[190] ;
 wire \u_inv.f_reg[191] ;
 wire \u_inv.f_reg[192] ;
 wire \u_inv.f_reg[193] ;
 wire \u_inv.f_reg[194] ;
 wire \u_inv.f_reg[195] ;
 wire \u_inv.f_reg[196] ;
 wire \u_inv.f_reg[197] ;
 wire \u_inv.f_reg[198] ;
 wire \u_inv.f_reg[199] ;
 wire \u_inv.f_reg[19] ;
 wire \u_inv.f_reg[1] ;
 wire \u_inv.f_reg[200] ;
 wire \u_inv.f_reg[201] ;
 wire \u_inv.f_reg[202] ;
 wire \u_inv.f_reg[203] ;
 wire \u_inv.f_reg[204] ;
 wire \u_inv.f_reg[205] ;
 wire \u_inv.f_reg[206] ;
 wire \u_inv.f_reg[207] ;
 wire \u_inv.f_reg[208] ;
 wire \u_inv.f_reg[209] ;
 wire \u_inv.f_reg[20] ;
 wire \u_inv.f_reg[210] ;
 wire \u_inv.f_reg[211] ;
 wire \u_inv.f_reg[212] ;
 wire \u_inv.f_reg[213] ;
 wire \u_inv.f_reg[214] ;
 wire \u_inv.f_reg[215] ;
 wire \u_inv.f_reg[216] ;
 wire \u_inv.f_reg[217] ;
 wire \u_inv.f_reg[218] ;
 wire \u_inv.f_reg[219] ;
 wire \u_inv.f_reg[21] ;
 wire \u_inv.f_reg[220] ;
 wire \u_inv.f_reg[221] ;
 wire \u_inv.f_reg[222] ;
 wire \u_inv.f_reg[223] ;
 wire \u_inv.f_reg[224] ;
 wire \u_inv.f_reg[225] ;
 wire \u_inv.f_reg[226] ;
 wire \u_inv.f_reg[227] ;
 wire \u_inv.f_reg[228] ;
 wire \u_inv.f_reg[229] ;
 wire \u_inv.f_reg[22] ;
 wire \u_inv.f_reg[230] ;
 wire \u_inv.f_reg[231] ;
 wire \u_inv.f_reg[232] ;
 wire \u_inv.f_reg[233] ;
 wire \u_inv.f_reg[234] ;
 wire \u_inv.f_reg[235] ;
 wire \u_inv.f_reg[236] ;
 wire \u_inv.f_reg[237] ;
 wire \u_inv.f_reg[238] ;
 wire \u_inv.f_reg[239] ;
 wire \u_inv.f_reg[23] ;
 wire \u_inv.f_reg[240] ;
 wire \u_inv.f_reg[241] ;
 wire \u_inv.f_reg[242] ;
 wire \u_inv.f_reg[243] ;
 wire \u_inv.f_reg[244] ;
 wire \u_inv.f_reg[245] ;
 wire \u_inv.f_reg[246] ;
 wire \u_inv.f_reg[247] ;
 wire \u_inv.f_reg[248] ;
 wire \u_inv.f_reg[249] ;
 wire \u_inv.f_reg[24] ;
 wire \u_inv.f_reg[250] ;
 wire \u_inv.f_reg[251] ;
 wire \u_inv.f_reg[252] ;
 wire \u_inv.f_reg[253] ;
 wire \u_inv.f_reg[254] ;
 wire \u_inv.f_reg[255] ;
 wire \u_inv.f_reg[256] ;
 wire \u_inv.f_reg[25] ;
 wire \u_inv.f_reg[26] ;
 wire \u_inv.f_reg[27] ;
 wire \u_inv.f_reg[28] ;
 wire \u_inv.f_reg[29] ;
 wire \u_inv.f_reg[2] ;
 wire \u_inv.f_reg[30] ;
 wire \u_inv.f_reg[31] ;
 wire \u_inv.f_reg[32] ;
 wire \u_inv.f_reg[33] ;
 wire \u_inv.f_reg[34] ;
 wire \u_inv.f_reg[35] ;
 wire \u_inv.f_reg[36] ;
 wire \u_inv.f_reg[37] ;
 wire \u_inv.f_reg[38] ;
 wire \u_inv.f_reg[39] ;
 wire \u_inv.f_reg[3] ;
 wire \u_inv.f_reg[40] ;
 wire \u_inv.f_reg[41] ;
 wire \u_inv.f_reg[42] ;
 wire \u_inv.f_reg[43] ;
 wire \u_inv.f_reg[44] ;
 wire \u_inv.f_reg[45] ;
 wire \u_inv.f_reg[46] ;
 wire \u_inv.f_reg[47] ;
 wire \u_inv.f_reg[48] ;
 wire \u_inv.f_reg[49] ;
 wire \u_inv.f_reg[4] ;
 wire \u_inv.f_reg[50] ;
 wire \u_inv.f_reg[51] ;
 wire \u_inv.f_reg[52] ;
 wire \u_inv.f_reg[53] ;
 wire \u_inv.f_reg[54] ;
 wire \u_inv.f_reg[55] ;
 wire \u_inv.f_reg[56] ;
 wire \u_inv.f_reg[57] ;
 wire \u_inv.f_reg[58] ;
 wire \u_inv.f_reg[59] ;
 wire \u_inv.f_reg[5] ;
 wire \u_inv.f_reg[60] ;
 wire \u_inv.f_reg[61] ;
 wire \u_inv.f_reg[62] ;
 wire \u_inv.f_reg[63] ;
 wire \u_inv.f_reg[64] ;
 wire \u_inv.f_reg[65] ;
 wire \u_inv.f_reg[66] ;
 wire \u_inv.f_reg[67] ;
 wire \u_inv.f_reg[68] ;
 wire \u_inv.f_reg[69] ;
 wire \u_inv.f_reg[6] ;
 wire \u_inv.f_reg[70] ;
 wire \u_inv.f_reg[71] ;
 wire \u_inv.f_reg[72] ;
 wire \u_inv.f_reg[73] ;
 wire \u_inv.f_reg[74] ;
 wire \u_inv.f_reg[75] ;
 wire \u_inv.f_reg[76] ;
 wire \u_inv.f_reg[77] ;
 wire \u_inv.f_reg[78] ;
 wire \u_inv.f_reg[79] ;
 wire \u_inv.f_reg[7] ;
 wire \u_inv.f_reg[80] ;
 wire \u_inv.f_reg[81] ;
 wire \u_inv.f_reg[82] ;
 wire \u_inv.f_reg[83] ;
 wire \u_inv.f_reg[84] ;
 wire \u_inv.f_reg[85] ;
 wire \u_inv.f_reg[86] ;
 wire \u_inv.f_reg[87] ;
 wire \u_inv.f_reg[88] ;
 wire \u_inv.f_reg[89] ;
 wire \u_inv.f_reg[8] ;
 wire \u_inv.f_reg[90] ;
 wire \u_inv.f_reg[91] ;
 wire \u_inv.f_reg[92] ;
 wire \u_inv.f_reg[93] ;
 wire \u_inv.f_reg[94] ;
 wire \u_inv.f_reg[95] ;
 wire \u_inv.f_reg[96] ;
 wire \u_inv.f_reg[97] ;
 wire \u_inv.f_reg[98] ;
 wire \u_inv.f_reg[99] ;
 wire \u_inv.f_reg[9] ;
 wire \u_inv.input_reg[0] ;
 wire \u_inv.input_reg[100] ;
 wire \u_inv.input_reg[101] ;
 wire \u_inv.input_reg[102] ;
 wire \u_inv.input_reg[103] ;
 wire \u_inv.input_reg[104] ;
 wire \u_inv.input_reg[105] ;
 wire \u_inv.input_reg[106] ;
 wire \u_inv.input_reg[107] ;
 wire \u_inv.input_reg[108] ;
 wire \u_inv.input_reg[109] ;
 wire \u_inv.input_reg[10] ;
 wire \u_inv.input_reg[110] ;
 wire \u_inv.input_reg[111] ;
 wire \u_inv.input_reg[112] ;
 wire \u_inv.input_reg[113] ;
 wire \u_inv.input_reg[114] ;
 wire \u_inv.input_reg[115] ;
 wire \u_inv.input_reg[116] ;
 wire \u_inv.input_reg[117] ;
 wire \u_inv.input_reg[118] ;
 wire \u_inv.input_reg[119] ;
 wire \u_inv.input_reg[11] ;
 wire \u_inv.input_reg[120] ;
 wire \u_inv.input_reg[121] ;
 wire \u_inv.input_reg[122] ;
 wire \u_inv.input_reg[123] ;
 wire \u_inv.input_reg[124] ;
 wire \u_inv.input_reg[125] ;
 wire \u_inv.input_reg[126] ;
 wire \u_inv.input_reg[127] ;
 wire \u_inv.input_reg[128] ;
 wire \u_inv.input_reg[129] ;
 wire \u_inv.input_reg[12] ;
 wire \u_inv.input_reg[130] ;
 wire \u_inv.input_reg[131] ;
 wire \u_inv.input_reg[132] ;
 wire \u_inv.input_reg[133] ;
 wire \u_inv.input_reg[134] ;
 wire \u_inv.input_reg[135] ;
 wire \u_inv.input_reg[136] ;
 wire \u_inv.input_reg[137] ;
 wire \u_inv.input_reg[138] ;
 wire \u_inv.input_reg[139] ;
 wire \u_inv.input_reg[13] ;
 wire \u_inv.input_reg[140] ;
 wire \u_inv.input_reg[141] ;
 wire \u_inv.input_reg[142] ;
 wire \u_inv.input_reg[143] ;
 wire \u_inv.input_reg[144] ;
 wire \u_inv.input_reg[145] ;
 wire \u_inv.input_reg[146] ;
 wire \u_inv.input_reg[147] ;
 wire \u_inv.input_reg[148] ;
 wire \u_inv.input_reg[149] ;
 wire \u_inv.input_reg[14] ;
 wire \u_inv.input_reg[150] ;
 wire \u_inv.input_reg[151] ;
 wire \u_inv.input_reg[152] ;
 wire \u_inv.input_reg[153] ;
 wire \u_inv.input_reg[154] ;
 wire \u_inv.input_reg[155] ;
 wire \u_inv.input_reg[156] ;
 wire \u_inv.input_reg[157] ;
 wire \u_inv.input_reg[158] ;
 wire \u_inv.input_reg[159] ;
 wire \u_inv.input_reg[15] ;
 wire \u_inv.input_reg[160] ;
 wire \u_inv.input_reg[161] ;
 wire \u_inv.input_reg[162] ;
 wire \u_inv.input_reg[163] ;
 wire \u_inv.input_reg[164] ;
 wire \u_inv.input_reg[165] ;
 wire \u_inv.input_reg[166] ;
 wire \u_inv.input_reg[167] ;
 wire \u_inv.input_reg[168] ;
 wire \u_inv.input_reg[169] ;
 wire \u_inv.input_reg[16] ;
 wire \u_inv.input_reg[170] ;
 wire \u_inv.input_reg[171] ;
 wire \u_inv.input_reg[172] ;
 wire \u_inv.input_reg[173] ;
 wire \u_inv.input_reg[174] ;
 wire \u_inv.input_reg[175] ;
 wire \u_inv.input_reg[176] ;
 wire \u_inv.input_reg[177] ;
 wire \u_inv.input_reg[178] ;
 wire \u_inv.input_reg[179] ;
 wire \u_inv.input_reg[17] ;
 wire \u_inv.input_reg[180] ;
 wire \u_inv.input_reg[181] ;
 wire \u_inv.input_reg[182] ;
 wire \u_inv.input_reg[183] ;
 wire \u_inv.input_reg[184] ;
 wire \u_inv.input_reg[185] ;
 wire \u_inv.input_reg[186] ;
 wire \u_inv.input_reg[187] ;
 wire \u_inv.input_reg[188] ;
 wire \u_inv.input_reg[189] ;
 wire \u_inv.input_reg[18] ;
 wire \u_inv.input_reg[190] ;
 wire \u_inv.input_reg[191] ;
 wire \u_inv.input_reg[192] ;
 wire \u_inv.input_reg[193] ;
 wire \u_inv.input_reg[194] ;
 wire \u_inv.input_reg[195] ;
 wire \u_inv.input_reg[196] ;
 wire \u_inv.input_reg[197] ;
 wire \u_inv.input_reg[198] ;
 wire \u_inv.input_reg[199] ;
 wire \u_inv.input_reg[19] ;
 wire \u_inv.input_reg[1] ;
 wire \u_inv.input_reg[200] ;
 wire \u_inv.input_reg[201] ;
 wire \u_inv.input_reg[202] ;
 wire \u_inv.input_reg[203] ;
 wire \u_inv.input_reg[204] ;
 wire \u_inv.input_reg[205] ;
 wire \u_inv.input_reg[206] ;
 wire \u_inv.input_reg[207] ;
 wire \u_inv.input_reg[208] ;
 wire \u_inv.input_reg[209] ;
 wire \u_inv.input_reg[20] ;
 wire \u_inv.input_reg[210] ;
 wire \u_inv.input_reg[211] ;
 wire \u_inv.input_reg[212] ;
 wire \u_inv.input_reg[213] ;
 wire \u_inv.input_reg[214] ;
 wire \u_inv.input_reg[215] ;
 wire \u_inv.input_reg[216] ;
 wire \u_inv.input_reg[217] ;
 wire \u_inv.input_reg[218] ;
 wire \u_inv.input_reg[219] ;
 wire \u_inv.input_reg[21] ;
 wire \u_inv.input_reg[220] ;
 wire \u_inv.input_reg[221] ;
 wire \u_inv.input_reg[222] ;
 wire \u_inv.input_reg[223] ;
 wire \u_inv.input_reg[224] ;
 wire \u_inv.input_reg[225] ;
 wire \u_inv.input_reg[226] ;
 wire \u_inv.input_reg[227] ;
 wire \u_inv.input_reg[228] ;
 wire \u_inv.input_reg[229] ;
 wire \u_inv.input_reg[22] ;
 wire \u_inv.input_reg[230] ;
 wire \u_inv.input_reg[231] ;
 wire \u_inv.input_reg[232] ;
 wire \u_inv.input_reg[233] ;
 wire \u_inv.input_reg[234] ;
 wire \u_inv.input_reg[235] ;
 wire \u_inv.input_reg[236] ;
 wire \u_inv.input_reg[237] ;
 wire \u_inv.input_reg[238] ;
 wire \u_inv.input_reg[239] ;
 wire \u_inv.input_reg[23] ;
 wire \u_inv.input_reg[240] ;
 wire \u_inv.input_reg[241] ;
 wire \u_inv.input_reg[242] ;
 wire \u_inv.input_reg[243] ;
 wire \u_inv.input_reg[244] ;
 wire \u_inv.input_reg[245] ;
 wire \u_inv.input_reg[246] ;
 wire \u_inv.input_reg[247] ;
 wire \u_inv.input_reg[248] ;
 wire \u_inv.input_reg[249] ;
 wire \u_inv.input_reg[24] ;
 wire \u_inv.input_reg[250] ;
 wire \u_inv.input_reg[251] ;
 wire \u_inv.input_reg[252] ;
 wire \u_inv.input_reg[253] ;
 wire \u_inv.input_reg[254] ;
 wire \u_inv.input_reg[255] ;
 wire \u_inv.input_reg[25] ;
 wire \u_inv.input_reg[26] ;
 wire \u_inv.input_reg[27] ;
 wire \u_inv.input_reg[28] ;
 wire \u_inv.input_reg[29] ;
 wire \u_inv.input_reg[2] ;
 wire \u_inv.input_reg[30] ;
 wire \u_inv.input_reg[31] ;
 wire \u_inv.input_reg[32] ;
 wire \u_inv.input_reg[33] ;
 wire \u_inv.input_reg[34] ;
 wire \u_inv.input_reg[35] ;
 wire \u_inv.input_reg[36] ;
 wire \u_inv.input_reg[37] ;
 wire \u_inv.input_reg[38] ;
 wire \u_inv.input_reg[39] ;
 wire \u_inv.input_reg[3] ;
 wire \u_inv.input_reg[40] ;
 wire \u_inv.input_reg[41] ;
 wire \u_inv.input_reg[42] ;
 wire \u_inv.input_reg[43] ;
 wire \u_inv.input_reg[44] ;
 wire \u_inv.input_reg[45] ;
 wire \u_inv.input_reg[46] ;
 wire \u_inv.input_reg[47] ;
 wire \u_inv.input_reg[48] ;
 wire \u_inv.input_reg[49] ;
 wire \u_inv.input_reg[4] ;
 wire \u_inv.input_reg[50] ;
 wire \u_inv.input_reg[51] ;
 wire \u_inv.input_reg[52] ;
 wire \u_inv.input_reg[53] ;
 wire \u_inv.input_reg[54] ;
 wire \u_inv.input_reg[55] ;
 wire \u_inv.input_reg[56] ;
 wire \u_inv.input_reg[57] ;
 wire \u_inv.input_reg[58] ;
 wire \u_inv.input_reg[59] ;
 wire \u_inv.input_reg[5] ;
 wire \u_inv.input_reg[60] ;
 wire \u_inv.input_reg[61] ;
 wire \u_inv.input_reg[62] ;
 wire \u_inv.input_reg[63] ;
 wire \u_inv.input_reg[64] ;
 wire \u_inv.input_reg[65] ;
 wire \u_inv.input_reg[66] ;
 wire \u_inv.input_reg[67] ;
 wire \u_inv.input_reg[68] ;
 wire \u_inv.input_reg[69] ;
 wire \u_inv.input_reg[6] ;
 wire \u_inv.input_reg[70] ;
 wire \u_inv.input_reg[71] ;
 wire \u_inv.input_reg[72] ;
 wire \u_inv.input_reg[73] ;
 wire \u_inv.input_reg[74] ;
 wire \u_inv.input_reg[75] ;
 wire \u_inv.input_reg[76] ;
 wire \u_inv.input_reg[77] ;
 wire \u_inv.input_reg[78] ;
 wire \u_inv.input_reg[79] ;
 wire \u_inv.input_reg[7] ;
 wire \u_inv.input_reg[80] ;
 wire \u_inv.input_reg[81] ;
 wire \u_inv.input_reg[82] ;
 wire \u_inv.input_reg[83] ;
 wire \u_inv.input_reg[84] ;
 wire \u_inv.input_reg[85] ;
 wire \u_inv.input_reg[86] ;
 wire \u_inv.input_reg[87] ;
 wire \u_inv.input_reg[88] ;
 wire \u_inv.input_reg[89] ;
 wire \u_inv.input_reg[8] ;
 wire \u_inv.input_reg[90] ;
 wire \u_inv.input_reg[91] ;
 wire \u_inv.input_reg[92] ;
 wire \u_inv.input_reg[93] ;
 wire \u_inv.input_reg[94] ;
 wire \u_inv.input_reg[95] ;
 wire \u_inv.input_reg[96] ;
 wire \u_inv.input_reg[97] ;
 wire \u_inv.input_reg[98] ;
 wire \u_inv.input_reg[99] ;
 wire \u_inv.input_reg[9] ;
 wire \u_inv.input_valid ;
 wire \u_inv.load_input ;
 wire \u_inv.state[0] ;
 wire \u_inv.state[1] ;
 wire net1063;
 wire clknet_leaf_0_clk;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire wr_prev;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_5_0_0_clk;
 wire clknet_5_1_0_clk;
 wire clknet_5_2_0_clk;
 wire clknet_5_3_0_clk;
 wire clknet_5_4_0_clk;
 wire clknet_5_5_0_clk;
 wire clknet_5_6_0_clk;
 wire clknet_5_7_0_clk;
 wire clknet_5_8_0_clk;
 wire clknet_5_9_0_clk;
 wire clknet_5_10_0_clk;
 wire clknet_5_11_0_clk;
 wire clknet_5_12_0_clk;
 wire clknet_5_13_0_clk;
 wire clknet_5_14_0_clk;
 wire clknet_5_15_0_clk;
 wire clknet_5_16_0_clk;
 wire clknet_5_17_0_clk;
 wire clknet_5_18_0_clk;
 wire clknet_5_19_0_clk;
 wire clknet_5_20_0_clk;
 wire clknet_5_21_0_clk;
 wire clknet_5_22_0_clk;
 wire clknet_5_23_0_clk;
 wire clknet_5_24_0_clk;
 wire clknet_5_25_0_clk;
 wire clknet_5_26_0_clk;
 wire clknet_5_27_0_clk;
 wire clknet_5_28_0_clk;
 wire clknet_5_29_0_clk;
 wire clknet_5_30_0_clk;
 wire clknet_5_31_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire [0:0] _20877_;
 wire [0:0] _20878_;

 sg13g2_inv_1 _20879_ (.Y(_13919_),
    .A(net2251));
 sg13g2_inv_1 _20880_ (.Y(_13920_),
    .A(\u_inv.f_next[254] ));
 sg13g2_inv_2 _20881_ (.Y(_13921_),
    .A(net2096));
 sg13g2_inv_2 _20882_ (.Y(_13922_),
    .A(net2368));
 sg13g2_inv_2 _20883_ (.Y(_13923_),
    .A(net2754));
 sg13g2_inv_2 _20884_ (.Y(_13924_),
    .A(net3292));
 sg13g2_inv_2 _20885_ (.Y(_13925_),
    .A(net2711));
 sg13g2_inv_1 _20886_ (.Y(_13926_),
    .A(net3364));
 sg13g2_inv_1 _20887_ (.Y(_13927_),
    .A(net3298));
 sg13g2_inv_2 _20888_ (.Y(_13928_),
    .A(net2873));
 sg13g2_inv_2 _20889_ (.Y(_13929_),
    .A(net2800));
 sg13g2_inv_1 _20890_ (.Y(_13930_),
    .A(net3375));
 sg13g2_inv_1 _20891_ (.Y(_13931_),
    .A(net3036));
 sg13g2_inv_1 _20892_ (.Y(_13932_),
    .A(net3337));
 sg13g2_inv_2 _20893_ (.Y(_13933_),
    .A(net2450));
 sg13g2_inv_2 _20894_ (.Y(_13934_),
    .A(net2069));
 sg13g2_inv_1 _20895_ (.Y(_13935_),
    .A(net3363));
 sg13g2_inv_1 _20896_ (.Y(_13936_),
    .A(net3152));
 sg13g2_inv_1 _20897_ (.Y(_13937_),
    .A(net3312));
 sg13g2_inv_1 _20898_ (.Y(_13938_),
    .A(net3336));
 sg13g2_inv_2 _20899_ (.Y(_13939_),
    .A(net2992));
 sg13g2_inv_1 _20900_ (.Y(_13940_),
    .A(net3365));
 sg13g2_inv_1 _20901_ (.Y(_13941_),
    .A(net3157));
 sg13g2_inv_1 _20902_ (.Y(_13942_),
    .A(net3413));
 sg13g2_inv_1 _20903_ (.Y(_13943_),
    .A(net3258));
 sg13g2_inv_2 _20904_ (.Y(_13944_),
    .A(net3310));
 sg13g2_inv_2 _20905_ (.Y(_13945_),
    .A(net2617));
 sg13g2_inv_1 _20906_ (.Y(_13946_),
    .A(net3359));
 sg13g2_inv_1 _20907_ (.Y(_13947_),
    .A(net3225));
 sg13g2_inv_2 _20908_ (.Y(_13948_),
    .A(net3328));
 sg13g2_inv_2 _20909_ (.Y(_13949_),
    .A(net2729));
 sg13g2_inv_2 _20910_ (.Y(_13950_),
    .A(net2991));
 sg13g2_inv_2 _20911_ (.Y(_13951_),
    .A(net2577));
 sg13g2_inv_1 _20912_ (.Y(_13952_),
    .A(net3283));
 sg13g2_inv_2 _20913_ (.Y(_13953_),
    .A(net2630));
 sg13g2_inv_2 _20914_ (.Y(_13954_),
    .A(net1504));
 sg13g2_inv_1 _20915_ (.Y(_13955_),
    .A(net3391));
 sg13g2_inv_1 _20916_ (.Y(_13956_),
    .A(net3396));
 sg13g2_inv_1 _20917_ (.Y(_13957_),
    .A(net3388));
 sg13g2_inv_1 _20918_ (.Y(_13958_),
    .A(net3424));
 sg13g2_inv_1 _20919_ (.Y(_13959_),
    .A(net3373));
 sg13g2_inv_1 _20920_ (.Y(_13960_),
    .A(net2961));
 sg13g2_inv_2 _20921_ (.Y(_13961_),
    .A(net2540));
 sg13g2_inv_1 _20922_ (.Y(_13962_),
    .A(net2713));
 sg13g2_inv_2 _20923_ (.Y(_13963_),
    .A(net2532));
 sg13g2_inv_2 _20924_ (.Y(_13964_),
    .A(net2481));
 sg13g2_inv_1 _20925_ (.Y(_13965_),
    .A(net3408));
 sg13g2_inv_2 _20926_ (.Y(_13966_),
    .A(net2413));
 sg13g2_inv_1 _20927_ (.Y(_13967_),
    .A(net3406));
 sg13g2_inv_1 _20928_ (.Y(_13968_),
    .A(net3139));
 sg13g2_inv_2 _20929_ (.Y(_13969_),
    .A(net2351));
 sg13g2_inv_2 _20930_ (.Y(_13970_),
    .A(net2281));
 sg13g2_inv_1 _20931_ (.Y(_13971_),
    .A(net3357));
 sg13g2_inv_1 _20932_ (.Y(_13972_),
    .A(net3300));
 sg13g2_inv_1 _20933_ (.Y(_13973_),
    .A(net2954));
 sg13g2_inv_2 _20934_ (.Y(_13974_),
    .A(net3006));
 sg13g2_inv_2 _20935_ (.Y(_13975_),
    .A(net2493));
 sg13g2_inv_1 _20936_ (.Y(_13976_),
    .A(net3314));
 sg13g2_inv_2 _20937_ (.Y(_13977_),
    .A(net2579));
 sg13g2_inv_2 _20938_ (.Y(_13978_),
    .A(net3367));
 sg13g2_inv_2 _20939_ (.Y(_13979_),
    .A(net3267));
 sg13g2_inv_2 _20940_ (.Y(_13980_),
    .A(net3394));
 sg13g2_inv_2 _20941_ (.Y(_13981_),
    .A(net3085));
 sg13g2_inv_1 _20942_ (.Y(_13982_),
    .A(net3266));
 sg13g2_inv_1 _20943_ (.Y(_13983_),
    .A(net3059));
 sg13g2_inv_1 _20944_ (.Y(_13984_),
    .A(net2583));
 sg13g2_inv_1 _20945_ (.Y(_13985_),
    .A(net3366));
 sg13g2_inv_1 _20946_ (.Y(_13986_),
    .A(net3334));
 sg13g2_inv_2 _20947_ (.Y(_13987_),
    .A(net2676));
 sg13g2_inv_2 _20948_ (.Y(_13988_),
    .A(net3099));
 sg13g2_inv_2 _20949_ (.Y(_13989_),
    .A(net2796));
 sg13g2_inv_1 _20950_ (.Y(_13990_),
    .A(net3078));
 sg13g2_inv_2 _20951_ (.Y(_13991_),
    .A(net2735));
 sg13g2_inv_1 _20952_ (.Y(_13992_),
    .A(net3000));
 sg13g2_inv_2 _20953_ (.Y(_13993_),
    .A(net2773));
 sg13g2_inv_1 _20954_ (.Y(_13994_),
    .A(net3318));
 sg13g2_inv_1 _20955_ (.Y(_13995_),
    .A(net3293));
 sg13g2_inv_1 _20956_ (.Y(_13996_),
    .A(net3250));
 sg13g2_inv_2 _20957_ (.Y(_13997_),
    .A(net3025));
 sg13g2_inv_1 _20958_ (.Y(_13998_),
    .A(net3423));
 sg13g2_inv_1 _20959_ (.Y(_13999_),
    .A(net3338));
 sg13g2_inv_1 _20960_ (.Y(_14000_),
    .A(net3330));
 sg13g2_inv_1 _20961_ (.Y(_14001_),
    .A(net3398));
 sg13g2_inv_1 _20962_ (.Y(_14002_),
    .A(net3414));
 sg13g2_inv_1 _20963_ (.Y(_14003_),
    .A(net3397));
 sg13g2_inv_1 _20964_ (.Y(_14004_),
    .A(net3282));
 sg13g2_inv_2 _20965_ (.Y(_14005_),
    .A(net3380));
 sg13g2_inv_1 _20966_ (.Y(_14006_),
    .A(net3421));
 sg13g2_inv_2 _20967_ (.Y(_14007_),
    .A(net3154));
 sg13g2_inv_1 _20968_ (.Y(_14008_),
    .A(net3323));
 sg13g2_inv_2 _20969_ (.Y(_14009_),
    .A(net3339));
 sg13g2_inv_1 _20970_ (.Y(_14010_),
    .A(net3079));
 sg13g2_inv_2 _20971_ (.Y(_14011_),
    .A(net2744));
 sg13g2_inv_1 _20972_ (.Y(_14012_),
    .A(net3256));
 sg13g2_inv_2 _20973_ (.Y(_14013_),
    .A(net2654));
 sg13g2_inv_1 _20974_ (.Y(_14014_),
    .A(net3143));
 sg13g2_inv_1 _20975_ (.Y(_14015_),
    .A(net3100));
 sg13g2_inv_1 _20976_ (.Y(_14016_),
    .A(net3275));
 sg13g2_inv_1 _20977_ (.Y(_14017_),
    .A(net3341));
 sg13g2_inv_2 _20978_ (.Y(_14018_),
    .A(net3168));
 sg13g2_inv_2 _20979_ (.Y(_14019_),
    .A(net3141));
 sg13g2_inv_1 _20980_ (.Y(_14020_),
    .A(net3327));
 sg13g2_inv_1 _20981_ (.Y(_14021_),
    .A(net3401));
 sg13g2_inv_1 _20982_ (.Y(_14022_),
    .A(net2681));
 sg13g2_inv_1 _20983_ (.Y(_14023_),
    .A(net3181));
 sg13g2_inv_2 _20984_ (.Y(_14024_),
    .A(net1925));
 sg13g2_inv_1 _20985_ (.Y(_14025_),
    .A(net2702));
 sg13g2_inv_2 _20986_ (.Y(_14026_),
    .A(net1849));
 sg13g2_inv_1 _20987_ (.Y(_14027_),
    .A(net3430));
 sg13g2_inv_2 _20988_ (.Y(_14028_),
    .A(net2946));
 sg13g2_inv_1 _20989_ (.Y(_14029_),
    .A(net3296));
 sg13g2_inv_1 _20990_ (.Y(_14030_),
    .A(net3403));
 sg13g2_inv_2 _20991_ (.Y(_14031_),
    .A(net3060));
 sg13g2_inv_1 _20992_ (.Y(_14032_),
    .A(net3415));
 sg13g2_inv_2 _20993_ (.Y(_14033_),
    .A(net3383));
 sg13g2_inv_1 _20994_ (.Y(_14034_),
    .A(net3361));
 sg13g2_inv_1 _20995_ (.Y(_14035_),
    .A(net3206));
 sg13g2_inv_1 _20996_ (.Y(_14036_),
    .A(net3171));
 sg13g2_inv_1 _20997_ (.Y(_14037_),
    .A(net3061));
 sg13g2_inv_2 _20998_ (.Y(_14038_),
    .A(net2565));
 sg13g2_inv_2 _20999_ (.Y(_14039_),
    .A(net3405));
 sg13g2_inv_1 _21000_ (.Y(_14040_),
    .A(net3409));
 sg13g2_inv_1 _21001_ (.Y(_14041_),
    .A(net3138));
 sg13g2_inv_1 _21002_ (.Y(_14042_),
    .A(net3024));
 sg13g2_inv_1 _21003_ (.Y(_14043_),
    .A(net3137));
 sg13g2_inv_1 _21004_ (.Y(_14044_),
    .A(net3185));
 sg13g2_inv_2 _21005_ (.Y(_14045_),
    .A(net2665));
 sg13g2_inv_2 _21006_ (.Y(_14046_),
    .A(net2783));
 sg13g2_inv_1 _21007_ (.Y(_14047_),
    .A(net3175));
 sg13g2_inv_1 _21008_ (.Y(_14048_),
    .A(net3201));
 sg13g2_inv_2 _21009_ (.Y(_14049_),
    .A(net2846));
 sg13g2_inv_1 _21010_ (.Y(_14050_),
    .A(net3429));
 sg13g2_inv_2 _21011_ (.Y(_14051_),
    .A(net3156));
 sg13g2_inv_1 _21012_ (.Y(_14052_),
    .A(net3219));
 sg13g2_inv_1 _21013_ (.Y(_14053_),
    .A(net3387));
 sg13g2_inv_1 _21014_ (.Y(_14054_),
    .A(net3426));
 sg13g2_inv_1 _21015_ (.Y(_14055_),
    .A(net3386));
 sg13g2_inv_1 _21016_ (.Y(_14056_),
    .A(net3276));
 sg13g2_inv_2 _21017_ (.Y(_14057_),
    .A(net2554));
 sg13g2_inv_1 _21018_ (.Y(_14058_),
    .A(net3211));
 sg13g2_inv_2 _21019_ (.Y(_14059_),
    .A(net2986));
 sg13g2_inv_1 _21020_ (.Y(_14060_),
    .A(net3404));
 sg13g2_inv_1 _21021_ (.Y(_14061_),
    .A(net3052));
 sg13g2_inv_1 _21022_ (.Y(_14062_),
    .A(net3249));
 sg13g2_inv_2 _21023_ (.Y(_14063_),
    .A(net3111));
 sg13g2_inv_1 _21024_ (.Y(_14064_),
    .A(net3326));
 sg13g2_inv_1 _21025_ (.Y(_14065_),
    .A(net3420));
 sg13g2_inv_2 _21026_ (.Y(_14066_),
    .A(net3252));
 sg13g2_inv_1 _21027_ (.Y(_14067_),
    .A(net3422));
 sg13g2_inv_1 _21028_ (.Y(_14068_),
    .A(net3407));
 sg13g2_inv_1 _21029_ (.Y(_14069_),
    .A(net3317));
 sg13g2_inv_1 _21030_ (.Y(_14070_),
    .A(net3262));
 sg13g2_inv_1 _21031_ (.Y(_14071_),
    .A(net3242));
 sg13g2_inv_1 _21032_ (.Y(_14072_),
    .A(net3416));
 sg13g2_inv_2 _21033_ (.Y(_14073_),
    .A(net3342));
 sg13g2_inv_2 _21034_ (.Y(_14074_),
    .A(net2491));
 sg13g2_inv_1 _21035_ (.Y(_14075_),
    .A(net3129));
 sg13g2_inv_1 _21036_ (.Y(_14076_),
    .A(net3374));
 sg13g2_inv_2 _21037_ (.Y(_14077_),
    .A(net2614));
 sg13g2_inv_2 _21038_ (.Y(_14078_),
    .A(net2978));
 sg13g2_inv_2 _21039_ (.Y(_14079_),
    .A(net3196));
 sg13g2_inv_2 _21040_ (.Y(_14080_),
    .A(net2391));
 sg13g2_inv_1 _21041_ (.Y(_14081_),
    .A(net3382));
 sg13g2_inv_1 _21042_ (.Y(_14082_),
    .A(net3308));
 sg13g2_inv_2 _21043_ (.Y(_14083_),
    .A(net3350));
 sg13g2_inv_1 _21044_ (.Y(_14084_),
    .A(net2858));
 sg13g2_inv_1 _21045_ (.Y(_14085_),
    .A(net2295));
 sg13g2_inv_1 _21046_ (.Y(_14086_),
    .A(net2911));
 sg13g2_inv_1 _21047_ (.Y(_14087_),
    .A(net3186));
 sg13g2_inv_1 _21048_ (.Y(_14088_),
    .A(net2951));
 sg13g2_inv_2 _21049_ (.Y(_14089_),
    .A(net2002));
 sg13g2_inv_1 _21050_ (.Y(_14090_),
    .A(net2673));
 sg13g2_inv_1 _21051_ (.Y(_14091_),
    .A(net3253));
 sg13g2_inv_2 _21052_ (.Y(_14092_),
    .A(net1820));
 sg13g2_inv_2 _21053_ (.Y(_14093_),
    .A(net2825));
 sg13g2_inv_1 _21054_ (.Y(_14094_),
    .A(net3362));
 sg13g2_inv_1 _21055_ (.Y(_14095_),
    .A(net3102));
 sg13g2_inv_1 _21056_ (.Y(_14096_),
    .A(net3199));
 sg13g2_inv_1 _21057_ (.Y(_14097_),
    .A(net3145));
 sg13g2_inv_1 _21058_ (.Y(_14098_),
    .A(net3247));
 sg13g2_inv_1 _21059_ (.Y(_14099_),
    .A(net3037));
 sg13g2_inv_1 _21060_ (.Y(_14100_),
    .A(net3286));
 sg13g2_inv_2 _21061_ (.Y(_14101_),
    .A(net3001));
 sg13g2_inv_1 _21062_ (.Y(_14102_),
    .A(net3307));
 sg13g2_inv_1 _21063_ (.Y(_14103_),
    .A(net3351));
 sg13g2_inv_1 _21064_ (.Y(_14104_),
    .A(net3043));
 sg13g2_inv_2 _21065_ (.Y(_14105_),
    .A(net2758));
 sg13g2_inv_2 _21066_ (.Y(_14106_),
    .A(net3020));
 sg13g2_inv_1 _21067_ (.Y(_14107_),
    .A(net3080));
 sg13g2_inv_1 _21068_ (.Y(_14108_),
    .A(net2823));
 sg13g2_inv_1 _21069_ (.Y(_14109_),
    .A(net2159));
 sg13g2_inv_1 _21070_ (.Y(_14110_),
    .A(net3064));
 sg13g2_inv_2 _21071_ (.Y(_14111_),
    .A(net2709));
 sg13g2_inv_1 _21072_ (.Y(_14112_),
    .A(net3385));
 sg13g2_inv_2 _21073_ (.Y(_14113_),
    .A(net3140));
 sg13g2_inv_1 _21074_ (.Y(_14114_),
    .A(net3233));
 sg13g2_inv_1 _21075_ (.Y(_14115_),
    .A(net3109));
 sg13g2_inv_1 _21076_ (.Y(_14116_),
    .A(net3246));
 sg13g2_inv_1 _21077_ (.Y(_14117_),
    .A(net2848));
 sg13g2_inv_2 _21078_ (.Y(_14118_),
    .A(net2546));
 sg13g2_inv_1 _21079_ (.Y(_14119_),
    .A(net3311));
 sg13g2_inv_1 _21080_ (.Y(_14120_),
    .A(net3335));
 sg13g2_inv_1 _21081_ (.Y(_14121_),
    .A(net3369));
 sg13g2_inv_1 _21082_ (.Y(_14122_),
    .A(net2972));
 sg13g2_inv_2 _21083_ (.Y(_14123_),
    .A(net2559));
 sg13g2_inv_2 _21084_ (.Y(_14124_),
    .A(net2512));
 sg13g2_inv_1 _21085_ (.Y(_14125_),
    .A(net3065));
 sg13g2_inv_1 _21086_ (.Y(_14126_),
    .A(net3041));
 sg13g2_inv_2 _21087_ (.Y(_14127_),
    .A(net2778));
 sg13g2_inv_1 _21088_ (.Y(_14128_),
    .A(net3189));
 sg13g2_inv_2 _21089_ (.Y(_14129_),
    .A(net3005));
 sg13g2_inv_1 _21090_ (.Y(_14130_),
    .A(net2960));
 sg13g2_inv_2 _21091_ (.Y(_14131_),
    .A(net2698));
 sg13g2_inv_1 _21092_ (.Y(_14132_),
    .A(net3136));
 sg13g2_inv_2 _21093_ (.Y(_14133_),
    .A(net3070));
 sg13g2_inv_1 _21094_ (.Y(_14134_),
    .A(net3224));
 sg13g2_inv_1 _21095_ (.Y(_14135_),
    .A(net3358));
 sg13g2_inv_1 _21096_ (.Y(_14136_),
    .A(net3263));
 sg13g2_inv_1 _21097_ (.Y(_14137_),
    .A(net3295));
 sg13g2_inv_1 _21098_ (.Y(_14138_),
    .A(net3402));
 sg13g2_inv_1 _21099_ (.Y(_14139_),
    .A(net3251));
 sg13g2_inv_1 _21100_ (.Y(_14140_),
    .A(net3259));
 sg13g2_inv_2 _21101_ (.Y(_14141_),
    .A(net3053));
 sg13g2_inv_1 _21102_ (.Y(_14142_),
    .A(net1743));
 sg13g2_inv_1 _21103_ (.Y(_14143_),
    .A(net3192));
 sg13g2_inv_1 _21104_ (.Y(_14144_),
    .A(net3306));
 sg13g2_inv_1 _21105_ (.Y(_14145_),
    .A(net3147));
 sg13g2_inv_1 _21106_ (.Y(_14146_),
    .A(net3329));
 sg13g2_inv_1 _21107_ (.Y(_14147_),
    .A(net3234));
 sg13g2_inv_1 _21108_ (.Y(_14148_),
    .A(net3291));
 sg13g2_inv_1 _21109_ (.Y(_14149_),
    .A(net2998));
 sg13g2_inv_1 _21110_ (.Y(_14150_),
    .A(net2851));
 sg13g2_inv_1 _21111_ (.Y(_14151_),
    .A(net2364));
 sg13g2_inv_1 _21112_ (.Y(_14152_),
    .A(\u_inv.f_next[22] ));
 sg13g2_inv_2 _21113_ (.Y(_14153_),
    .A(net1554));
 sg13g2_inv_1 _21114_ (.Y(_14154_),
    .A(net3392));
 sg13g2_inv_2 _21115_ (.Y(_14155_),
    .A(net2980));
 sg13g2_inv_1 _21116_ (.Y(_14156_),
    .A(net3340));
 sg13g2_inv_1 _21117_ (.Y(_14157_),
    .A(net3117));
 sg13g2_inv_1 _21118_ (.Y(_14158_),
    .A(net3395));
 sg13g2_inv_2 _21119_ (.Y(_14159_),
    .A(net3008));
 sg13g2_inv_1 _21120_ (.Y(_14160_),
    .A(net3425));
 sg13g2_inv_1 _21121_ (.Y(_14161_),
    .A(net3273));
 sg13g2_inv_1 _21122_ (.Y(_14162_),
    .A(net3169));
 sg13g2_inv_1 _21123_ (.Y(_14163_),
    .A(net3200));
 sg13g2_inv_1 _21124_ (.Y(_14164_),
    .A(net3207));
 sg13g2_inv_1 _21125_ (.Y(_14165_),
    .A(net2526));
 sg13g2_inv_1 _21126_ (.Y(_14166_),
    .A(net1244));
 sg13g2_inv_1 _21127_ (.Y(_14167_),
    .A(net3352));
 sg13g2_inv_1 _21128_ (.Y(_14168_),
    .A(net3393));
 sg13g2_inv_1 _21129_ (.Y(_14169_),
    .A(net3410));
 sg13g2_inv_1 _21130_ (.Y(_14170_),
    .A(net3360));
 sg13g2_inv_8 _21131_ (.Y(_14171_),
    .A(net5751));
 sg13g2_inv_1 _21132_ (.Y(_14172_),
    .A(\u_inv.d_next[256] ));
 sg13g2_inv_1 _21133_ (.Y(_14173_),
    .A(\u_inv.d_next[246] ));
 sg13g2_inv_1 _21134_ (.Y(_14174_),
    .A(\u_inv.d_next[241] ));
 sg13g2_inv_1 _21135_ (.Y(_14175_),
    .A(\u_inv.d_next[239] ));
 sg13g2_inv_1 _21136_ (.Y(_14176_),
    .A(\u_inv.d_next[233] ));
 sg13g2_inv_1 _21137_ (.Y(_14177_),
    .A(\u_inv.d_next[232] ));
 sg13g2_inv_1 _21138_ (.Y(_14178_),
    .A(\u_inv.d_next[229] ));
 sg13g2_inv_1 _21139_ (.Y(_14179_),
    .A(\u_inv.d_next[227] ));
 sg13g2_inv_1 _21140_ (.Y(_14180_),
    .A(\u_inv.d_next[222] ));
 sg13g2_inv_1 _21141_ (.Y(_14181_),
    .A(\u_inv.d_next[221] ));
 sg13g2_inv_1 _21142_ (.Y(_14182_),
    .A(\u_inv.d_next[217] ));
 sg13g2_inv_1 _21143_ (.Y(_14183_),
    .A(\u_inv.d_next[213] ));
 sg13g2_inv_1 _21144_ (.Y(_14184_),
    .A(\u_inv.d_next[209] ));
 sg13g2_inv_1 _21145_ (.Y(_14185_),
    .A(\u_inv.d_next[207] ));
 sg13g2_inv_1 _21146_ (.Y(_14186_),
    .A(\u_inv.d_next[205] ));
 sg13g2_inv_1 _21147_ (.Y(_14187_),
    .A(\u_inv.d_next[203] ));
 sg13g2_inv_1 _21148_ (.Y(_14188_),
    .A(\u_inv.d_next[199] ));
 sg13g2_inv_1 _21149_ (.Y(_14189_),
    .A(\u_inv.d_next[195] ));
 sg13g2_inv_1 _21150_ (.Y(_14190_),
    .A(\u_inv.d_next[193] ));
 sg13g2_inv_1 _21151_ (.Y(_14191_),
    .A(\u_inv.d_next[190] ));
 sg13g2_inv_1 _21152_ (.Y(_14192_),
    .A(\u_inv.d_next[189] ));
 sg13g2_inv_1 _21153_ (.Y(_14193_),
    .A(\u_inv.d_next[183] ));
 sg13g2_inv_1 _21154_ (.Y(_14194_),
    .A(\u_inv.d_next[181] ));
 sg13g2_inv_1 _21155_ (.Y(_14195_),
    .A(\u_inv.d_next[179] ));
 sg13g2_inv_1 _21156_ (.Y(_14196_),
    .A(\u_inv.d_next[177] ));
 sg13g2_inv_1 _21157_ (.Y(_14197_),
    .A(\u_inv.d_next[175] ));
 sg13g2_inv_1 _21158_ (.Y(_14198_),
    .A(\u_inv.d_next[172] ));
 sg13g2_inv_1 _21159_ (.Y(_14199_),
    .A(\u_inv.d_next[167] ));
 sg13g2_inv_1 _21160_ (.Y(_14200_),
    .A(\u_inv.d_next[159] ));
 sg13g2_inv_1 _21161_ (.Y(_14201_),
    .A(\u_inv.d_next[155] ));
 sg13g2_inv_1 _21162_ (.Y(_14202_),
    .A(\u_inv.d_next[153] ));
 sg13g2_inv_1 _21163_ (.Y(_14203_),
    .A(\u_inv.d_next[149] ));
 sg13g2_inv_1 _21164_ (.Y(_14204_),
    .A(\u_inv.d_next[147] ));
 sg13g2_inv_1 _21165_ (.Y(_14205_),
    .A(net5876));
 sg13g2_inv_1 _21166_ (.Y(_14206_),
    .A(\u_inv.d_next[143] ));
 sg13g2_inv_1 _21167_ (.Y(_14207_),
    .A(\u_inv.d_next[141] ));
 sg13g2_inv_1 _21168_ (.Y(_14208_),
    .A(\u_inv.d_next[139] ));
 sg13g2_inv_1 _21169_ (.Y(_14209_),
    .A(\u_inv.d_next[137] ));
 sg13g2_inv_1 _21170_ (.Y(_14210_),
    .A(\u_inv.d_next[135] ));
 sg13g2_inv_1 _21171_ (.Y(_14211_),
    .A(\u_inv.d_next[133] ));
 sg13g2_inv_1 _21172_ (.Y(_14212_),
    .A(\u_inv.d_next[131] ));
 sg13g2_inv_1 _21173_ (.Y(_14213_),
    .A(\u_inv.d_next[125] ));
 sg13g2_inv_1 _21174_ (.Y(_14214_),
    .A(\u_inv.d_next[119] ));
 sg13g2_inv_1 _21175_ (.Y(_14215_),
    .A(\u_inv.d_next[117] ));
 sg13g2_inv_1 _21176_ (.Y(_14216_),
    .A(\u_inv.d_next[114] ));
 sg13g2_inv_1 _21177_ (.Y(_14217_),
    .A(\u_inv.d_next[105] ));
 sg13g2_inv_1 _21178_ (.Y(_14218_),
    .A(\u_inv.d_next[103] ));
 sg13g2_inv_1 _21179_ (.Y(_14219_),
    .A(\u_inv.d_next[93] ));
 sg13g2_inv_1 _21180_ (.Y(_14220_),
    .A(\u_inv.d_next[90] ));
 sg13g2_inv_1 _21181_ (.Y(_14221_),
    .A(\u_inv.d_next[89] ));
 sg13g2_inv_1 _21182_ (.Y(_14222_),
    .A(\u_inv.d_next[85] ));
 sg13g2_inv_1 _21183_ (.Y(_14223_),
    .A(\u_inv.d_next[83] ));
 sg13g2_inv_1 _21184_ (.Y(_14224_),
    .A(net5877));
 sg13g2_inv_1 _21185_ (.Y(_14225_),
    .A(net5880));
 sg13g2_inv_1 _21186_ (.Y(_14226_),
    .A(\u_inv.d_next[63] ));
 sg13g2_inv_1 _21187_ (.Y(_14227_),
    .A(\u_inv.d_next[58] ));
 sg13g2_inv_1 _21188_ (.Y(_14228_),
    .A(\u_inv.d_next[57] ));
 sg13g2_inv_1 _21189_ (.Y(_14229_),
    .A(\u_inv.d_next[55] ));
 sg13g2_inv_1 _21190_ (.Y(_14230_),
    .A(\u_inv.d_next[53] ));
 sg13g2_inv_1 _21191_ (.Y(_14231_),
    .A(\u_inv.d_next[42] ));
 sg13g2_inv_1 _21192_ (.Y(_14232_),
    .A(\u_inv.d_next[41] ));
 sg13g2_inv_1 _21193_ (.Y(_14233_),
    .A(\u_inv.d_next[37] ));
 sg13g2_inv_1 _21194_ (.Y(_14234_),
    .A(\u_inv.d_next[35] ));
 sg13g2_inv_1 _21195_ (.Y(_14235_),
    .A(\u_inv.d_next[34] ));
 sg13g2_inv_1 _21196_ (.Y(_14236_),
    .A(\u_inv.d_next[23] ));
 sg13g2_inv_1 _21197_ (.Y(_14237_),
    .A(\u_inv.d_next[21] ));
 sg13g2_inv_1 _21198_ (.Y(_14238_),
    .A(\u_inv.d_next[17] ));
 sg13g2_inv_1 _21199_ (.Y(_14239_),
    .A(\u_inv.d_next[15] ));
 sg13g2_inv_1 _21200_ (.Y(_14240_),
    .A(\u_inv.d_next[13] ));
 sg13g2_inv_1 _21201_ (.Y(_14241_),
    .A(\u_inv.d_next[5] ));
 sg13g2_inv_1 _21202_ (.Y(_14242_),
    .A(net1384));
 sg13g2_inv_2 _21203_ (.Y(_14243_),
    .A(net3433));
 sg13g2_inv_1 _21204_ (.Y(_14244_),
    .A(net3368));
 sg13g2_inv_1 _21205_ (.Y(_14245_),
    .A(\u_inv.delta_reg[5] ));
 sg13g2_inv_1 _21206_ (.Y(_14246_),
    .A(net3436));
 sg13g2_inv_1 _21207_ (.Y(_14247_),
    .A(net1153));
 sg13g2_inv_1 _21208_ (.Y(_14248_),
    .A(net5829));
 sg13g2_inv_2 _21209_ (.Y(_14249_),
    .A(net3389));
 sg13g2_inv_1 _21210_ (.Y(_14250_),
    .A(net3371));
 sg13g2_inv_2 _21211_ (.Y(_14251_),
    .A(net3431));
 sg13g2_inv_2 _21212_ (.Y(_14252_),
    .A(net3241));
 sg13g2_inv_1 _21213_ (.Y(_14253_),
    .A(net3072));
 sg13g2_inv_2 _21214_ (.Y(_14254_),
    .A(net3343));
 sg13g2_inv_1 _21215_ (.Y(_14255_),
    .A(net2360));
 sg13g2_inv_1 _21216_ (.Y(_14256_),
    .A(net2253));
 sg13g2_inv_1 _21217_ (.Y(_14257_),
    .A(net2833));
 sg13g2_inv_1 _21218_ (.Y(_14258_),
    .A(\u_inv.f_reg[4] ));
 sg13g2_inv_1 _21219_ (.Y(_14259_),
    .A(net2856));
 sg13g2_inv_1 _21220_ (.Y(_14260_),
    .A(net2163));
 sg13g2_inv_1 _21221_ (.Y(_14261_),
    .A(\u_inv.f_reg[7] ));
 sg13g2_inv_1 _21222_ (.Y(_14262_),
    .A(\u_inv.f_reg[8] ));
 sg13g2_inv_1 _21223_ (.Y(_14263_),
    .A(\u_inv.f_reg[9] ));
 sg13g2_inv_1 _21224_ (.Y(_14264_),
    .A(net2924));
 sg13g2_inv_1 _21225_ (.Y(_14265_),
    .A(net2860));
 sg13g2_inv_1 _21226_ (.Y(_14266_),
    .A(\u_inv.f_reg[12] ));
 sg13g2_inv_1 _21227_ (.Y(_14267_),
    .A(net3349));
 sg13g2_inv_1 _21228_ (.Y(_14268_),
    .A(net2817));
 sg13g2_inv_1 _21229_ (.Y(_14269_),
    .A(net2501));
 sg13g2_inv_1 _21230_ (.Y(_14270_),
    .A(net3089));
 sg13g2_inv_1 _21231_ (.Y(_14271_),
    .A(\u_inv.f_reg[17] ));
 sg13g2_inv_1 _21232_ (.Y(_14272_),
    .A(net3034));
 sg13g2_inv_1 _21233_ (.Y(_14273_),
    .A(\u_inv.f_reg[19] ));
 sg13g2_inv_1 _21234_ (.Y(_14274_),
    .A(net2593));
 sg13g2_inv_1 _21235_ (.Y(_14275_),
    .A(\u_inv.f_reg[21] ));
 sg13g2_inv_1 _21236_ (.Y(_14276_),
    .A(net2670));
 sg13g2_inv_1 _21237_ (.Y(_14277_),
    .A(net2867));
 sg13g2_inv_1 _21238_ (.Y(_14278_),
    .A(\u_inv.f_reg[24] ));
 sg13g2_inv_1 _21239_ (.Y(_14279_),
    .A(\u_inv.f_reg[25] ));
 sg13g2_inv_1 _21240_ (.Y(_14280_),
    .A(net2464));
 sg13g2_inv_1 _21241_ (.Y(_14281_),
    .A(net2760));
 sg13g2_inv_1 _21242_ (.Y(_14282_),
    .A(net3161));
 sg13g2_inv_1 _21243_ (.Y(_14283_),
    .A(\u_inv.f_reg[29] ));
 sg13g2_inv_1 _21244_ (.Y(_14284_),
    .A(net3039));
 sg13g2_inv_1 _21245_ (.Y(_14285_),
    .A(\u_inv.f_reg[31] ));
 sg13g2_inv_2 _21246_ (.Y(_14286_),
    .A(\u_inv.f_reg[32] ));
 sg13g2_inv_1 _21247_ (.Y(_14287_),
    .A(\u_inv.f_reg[33] ));
 sg13g2_inv_1 _21248_ (.Y(_14288_),
    .A(net2892));
 sg13g2_inv_1 _21249_ (.Y(_14289_),
    .A(net3299));
 sg13g2_inv_1 _21250_ (.Y(_14290_),
    .A(net2939));
 sg13g2_inv_1 _21251_ (.Y(_14291_),
    .A(net3284));
 sg13g2_inv_1 _21252_ (.Y(_14292_),
    .A(net2766));
 sg13g2_inv_1 _21253_ (.Y(_14293_),
    .A(net3302));
 sg13g2_inv_1 _21254_ (.Y(_14294_),
    .A(net2890));
 sg13g2_inv_1 _21255_ (.Y(_14295_),
    .A(\u_inv.f_reg[41] ));
 sg13g2_inv_1 _21256_ (.Y(_14296_),
    .A(net2409));
 sg13g2_inv_1 _21257_ (.Y(_14297_),
    .A(\u_inv.f_reg[43] ));
 sg13g2_inv_1 _21258_ (.Y(_14298_),
    .A(net2899));
 sg13g2_inv_1 _21259_ (.Y(_14299_),
    .A(net2684));
 sg13g2_inv_1 _21260_ (.Y(_14300_),
    .A(net2242));
 sg13g2_inv_1 _21261_ (.Y(_14301_),
    .A(\u_inv.f_reg[47] ));
 sg13g2_inv_1 _21262_ (.Y(_14302_),
    .A(\u_inv.f_reg[48] ));
 sg13g2_inv_1 _21263_ (.Y(_14303_),
    .A(net3214));
 sg13g2_inv_1 _21264_ (.Y(_14304_),
    .A(\u_inv.f_reg[50] ));
 sg13g2_inv_1 _21265_ (.Y(_14305_),
    .A(\u_inv.f_reg[51] ));
 sg13g2_inv_1 _21266_ (.Y(_14306_),
    .A(net2301));
 sg13g2_inv_1 _21267_ (.Y(_14307_),
    .A(net3179));
 sg13g2_inv_1 _21268_ (.Y(_14308_),
    .A(net3123));
 sg13g2_inv_1 _21269_ (.Y(_14309_),
    .A(net3132));
 sg13g2_inv_1 _21270_ (.Y(_14310_),
    .A(\u_inv.f_reg[56] ));
 sg13g2_inv_1 _21271_ (.Y(_14311_),
    .A(net3294));
 sg13g2_inv_1 _21272_ (.Y(_14312_),
    .A(net2877));
 sg13g2_inv_1 _21273_ (.Y(_14313_),
    .A(\u_inv.f_reg[59] ));
 sg13g2_inv_1 _21274_ (.Y(_14314_),
    .A(net3257));
 sg13g2_inv_1 _21275_ (.Y(_14315_),
    .A(net2913));
 sg13g2_inv_1 _21276_ (.Y(_14316_),
    .A(net1877));
 sg13g2_inv_1 _21277_ (.Y(_14317_),
    .A(\u_inv.f_reg[63] ));
 sg13g2_inv_1 _21278_ (.Y(_14318_),
    .A(net2967));
 sg13g2_inv_1 _21279_ (.Y(_14319_),
    .A(\u_inv.f_reg[65] ));
 sg13g2_inv_1 _21280_ (.Y(_14320_),
    .A(net2752));
 sg13g2_inv_1 _21281_ (.Y(_14321_),
    .A(\u_inv.f_reg[67] ));
 sg13g2_inv_2 _21282_ (.Y(_14322_),
    .A(net2220));
 sg13g2_inv_1 _21283_ (.Y(_14323_),
    .A(\u_inv.f_reg[69] ));
 sg13g2_inv_1 _21284_ (.Y(_14324_),
    .A(net2466));
 sg13g2_inv_1 _21285_ (.Y(_14325_),
    .A(net3237));
 sg13g2_inv_1 _21286_ (.Y(_14326_),
    .A(net3166));
 sg13g2_inv_1 _21287_ (.Y(_14327_),
    .A(\u_inv.f_reg[73] ));
 sg13g2_inv_1 _21288_ (.Y(_14328_),
    .A(net3057));
 sg13g2_inv_1 _21289_ (.Y(_14329_),
    .A(\u_inv.f_reg[75] ));
 sg13g2_inv_1 _21290_ (.Y(_14330_),
    .A(net2894));
 sg13g2_inv_1 _21291_ (.Y(_14331_),
    .A(\u_inv.f_reg[77] ));
 sg13g2_inv_1 _21292_ (.Y(_14332_),
    .A(net2695));
 sg13g2_inv_1 _21293_ (.Y(_14333_),
    .A(\u_inv.f_reg[79] ));
 sg13g2_inv_1 _21294_ (.Y(_14334_),
    .A(net2771));
 sg13g2_inv_1 _21295_ (.Y(_14335_),
    .A(\u_inv.f_reg[81] ));
 sg13g2_inv_1 _21296_ (.Y(_14336_),
    .A(\u_inv.f_reg[82] ));
 sg13g2_inv_1 _21297_ (.Y(_14337_),
    .A(net2838));
 sg13g2_inv_1 _21298_ (.Y(_14338_),
    .A(\u_inv.f_reg[84] ));
 sg13g2_inv_1 _21299_ (.Y(_14339_),
    .A(\u_inv.f_reg[85] ));
 sg13g2_inv_1 _21300_ (.Y(_14340_),
    .A(net2812));
 sg13g2_inv_1 _21301_ (.Y(_14341_),
    .A(net3399));
 sg13g2_inv_1 _21302_ (.Y(_14342_),
    .A(\u_inv.f_reg[88] ));
 sg13g2_inv_1 _21303_ (.Y(_14343_),
    .A(\u_inv.f_reg[89] ));
 sg13g2_inv_1 _21304_ (.Y(_14344_),
    .A(net3046));
 sg13g2_inv_2 _21305_ (.Y(_14345_),
    .A(net2647));
 sg13g2_inv_1 _21306_ (.Y(_14346_),
    .A(\u_inv.f_reg[92] ));
 sg13g2_inv_1 _21307_ (.Y(_14347_),
    .A(net3260));
 sg13g2_inv_1 _21308_ (.Y(_14348_),
    .A(\u_inv.f_reg[94] ));
 sg13g2_inv_1 _21309_ (.Y(_14349_),
    .A(net2585));
 sg13g2_inv_1 _21310_ (.Y(_14350_),
    .A(net3174));
 sg13g2_inv_1 _21311_ (.Y(_14351_),
    .A(\u_inv.f_reg[97] ));
 sg13g2_inv_1 _21312_ (.Y(_14352_),
    .A(net3208));
 sg13g2_inv_1 _21313_ (.Y(_14353_),
    .A(net3370));
 sg13g2_inv_1 _21314_ (.Y(_14354_),
    .A(\u_inv.f_reg[100] ));
 sg13g2_inv_1 _21315_ (.Y(_14355_),
    .A(net2687));
 sg13g2_inv_1 _21316_ (.Y(_14356_),
    .A(net3134));
 sg13g2_inv_1 _21317_ (.Y(_14357_),
    .A(\u_inv.f_reg[103] ));
 sg13g2_inv_1 _21318_ (.Y(_14358_),
    .A(net2789));
 sg13g2_inv_1 _21319_ (.Y(_14359_),
    .A(net3204));
 sg13g2_inv_1 _21320_ (.Y(_14360_),
    .A(net2915));
 sg13g2_inv_1 _21321_ (.Y(_14361_),
    .A(net3344));
 sg13g2_inv_2 _21322_ (.Y(_14362_),
    .A(net1297));
 sg13g2_inv_2 _21323_ (.Y(_14363_),
    .A(net3150));
 sg13g2_inv_1 _21324_ (.Y(_14364_),
    .A(net2489));
 sg13g2_inv_1 _21325_ (.Y(_14365_),
    .A(\u_inv.f_reg[111] ));
 sg13g2_inv_1 _21326_ (.Y(_14366_),
    .A(net3107));
 sg13g2_inv_1 _21327_ (.Y(_14367_),
    .A(net3319));
 sg13g2_inv_1 _21328_ (.Y(_14368_),
    .A(net2829));
 sg13g2_inv_1 _21329_ (.Y(_14369_),
    .A(\u_inv.f_reg[115] ));
 sg13g2_inv_1 _21330_ (.Y(_14370_),
    .A(net3030));
 sg13g2_inv_1 _21331_ (.Y(_14371_),
    .A(\u_inv.f_reg[117] ));
 sg13g2_inv_1 _21332_ (.Y(_14372_),
    .A(net2050));
 sg13g2_inv_1 _21333_ (.Y(_14373_),
    .A(net3353));
 sg13g2_inv_1 _21334_ (.Y(_14374_),
    .A(net2930));
 sg13g2_inv_1 _21335_ (.Y(_14375_),
    .A(net3202));
 sg13g2_inv_1 _21336_ (.Y(_14376_),
    .A(net2038));
 sg13g2_inv_1 _21337_ (.Y(_14377_),
    .A(net2234));
 sg13g2_inv_1 _21338_ (.Y(_14378_),
    .A(net3113));
 sg13g2_inv_1 _21339_ (.Y(_14379_),
    .A(\u_inv.f_reg[125] ));
 sg13g2_inv_1 _21340_ (.Y(_14380_),
    .A(net2746));
 sg13g2_inv_1 _21341_ (.Y(_14381_),
    .A(\u_inv.f_reg[127] ));
 sg13g2_inv_1 _21342_ (.Y(_14382_),
    .A(\u_inv.f_reg[128] ));
 sg13g2_inv_1 _21343_ (.Y(_14383_),
    .A(\u_inv.f_reg[129] ));
 sg13g2_inv_1 _21344_ (.Y(_14384_),
    .A(net2471));
 sg13g2_inv_1 _21345_ (.Y(_14385_),
    .A(net2499));
 sg13g2_inv_1 _21346_ (.Y(_14386_),
    .A(net2661));
 sg13g2_inv_1 _21347_ (.Y(_14387_),
    .A(net2455));
 sg13g2_inv_1 _21348_ (.Y(_14388_),
    .A(net2958));
 sg13g2_inv_1 _21349_ (.Y(_14389_),
    .A(net3163));
 sg13g2_inv_1 _21350_ (.Y(_14390_),
    .A(\u_inv.f_reg[136] ));
 sg13g2_inv_1 _21351_ (.Y(_14391_),
    .A(net1368));
 sg13g2_inv_1 _21352_ (.Y(_14392_),
    .A(net3279));
 sg13g2_inv_1 _21353_ (.Y(_14393_),
    .A(net3297));
 sg13g2_inv_1 _21354_ (.Y(_14394_),
    .A(net2820));
 sg13g2_inv_1 _21355_ (.Y(_14395_),
    .A(net3212));
 sg13g2_inv_1 _21356_ (.Y(_14396_),
    .A(net3268));
 sg13g2_inv_2 _21357_ (.Y(_14397_),
    .A(net2700));
 sg13g2_inv_2 _21358_ (.Y(_14398_),
    .A(net2805));
 sg13g2_inv_1 _21359_ (.Y(_14399_),
    .A(net2424));
 sg13g2_inv_1 _21360_ (.Y(_14400_),
    .A(\u_inv.f_reg[146] ));
 sg13g2_inv_1 _21361_ (.Y(_14401_),
    .A(net2798));
 sg13g2_inv_1 _21362_ (.Y(_14402_),
    .A(\u_inv.f_reg[148] ));
 sg13g2_inv_1 _21363_ (.Y(_14403_),
    .A(net3051));
 sg13g2_inv_1 _21364_ (.Y(_14404_),
    .A(\u_inv.f_reg[150] ));
 sg13g2_inv_1 _21365_ (.Y(_14405_),
    .A(\u_inv.f_reg[151] ));
 sg13g2_inv_1 _21366_ (.Y(_14406_),
    .A(net3248));
 sg13g2_inv_1 _21367_ (.Y(_14407_),
    .A(net3277));
 sg13g2_inv_1 _21368_ (.Y(_14408_),
    .A(net3014));
 sg13g2_inv_1 _21369_ (.Y(_14409_),
    .A(\u_inv.f_reg[155] ));
 sg13g2_inv_2 _21370_ (.Y(_14410_),
    .A(net2598));
 sg13g2_inv_1 _21371_ (.Y(_14411_),
    .A(net3280));
 sg13g2_inv_1 _21372_ (.Y(_14412_),
    .A(net2982));
 sg13g2_inv_1 _21373_ (.Y(_14413_),
    .A(\u_inv.f_reg[159] ));
 sg13g2_inv_1 _21374_ (.Y(_14414_),
    .A(\u_inv.f_reg[160] ));
 sg13g2_inv_1 _21375_ (.Y(_14415_),
    .A(\u_inv.f_reg[161] ));
 sg13g2_inv_1 _21376_ (.Y(_14416_),
    .A(net2719));
 sg13g2_inv_1 _21377_ (.Y(_14417_),
    .A(\u_inv.f_reg[163] ));
 sg13g2_inv_1 _21378_ (.Y(_14418_),
    .A(net2869));
 sg13g2_inv_1 _21379_ (.Y(_14419_),
    .A(net2854));
 sg13g2_inv_1 _21380_ (.Y(_14420_),
    .A(net1818));
 sg13g2_inv_1 _21381_ (.Y(_14421_),
    .A(\u_inv.f_reg[167] ));
 sg13g2_inv_1 _21382_ (.Y(_14422_),
    .A(net3355));
 sg13g2_inv_1 _21383_ (.Y(_14423_),
    .A(net3194));
 sg13g2_inv_1 _21384_ (.Y(_14424_),
    .A(net2748));
 sg13g2_inv_1 _21385_ (.Y(_14425_),
    .A(net3376));
 sg13g2_inv_1 _21386_ (.Y(_14426_),
    .A(net3062));
 sg13g2_inv_1 _21387_ (.Y(_14427_),
    .A(net3324));
 sg13g2_inv_1 _21388_ (.Y(_14428_),
    .A(net2807));
 sg13g2_inv_1 _21389_ (.Y(_14429_),
    .A(net3244));
 sg13g2_inv_1 _21390_ (.Y(_14430_),
    .A(net3190));
 sg13g2_inv_1 _21391_ (.Y(_14431_),
    .A(\u_inv.f_reg[177] ));
 sg13g2_inv_1 _21392_ (.Y(_14432_),
    .A(net3010));
 sg13g2_inv_1 _21393_ (.Y(_14433_),
    .A(net2714));
 sg13g2_inv_1 _21394_ (.Y(_14434_),
    .A(net3018));
 sg13g2_inv_1 _21395_ (.Y(_14435_),
    .A(\u_inv.f_reg[181] ));
 sg13g2_inv_1 _21396_ (.Y(_14436_),
    .A(net2030));
 sg13g2_inv_1 _21397_ (.Y(_14437_),
    .A(\u_inv.f_reg[183] ));
 sg13g2_inv_1 _21398_ (.Y(_14438_),
    .A(net3016));
 sg13g2_inv_1 _21399_ (.Y(_14439_),
    .A(\u_inv.f_reg[185] ));
 sg13g2_inv_1 _21400_ (.Y(_14440_),
    .A(net2353));
 sg13g2_inv_1 _21401_ (.Y(_14441_),
    .A(\u_inv.f_reg[187] ));
 sg13g2_inv_2 _21402_ (.Y(_14442_),
    .A(net2270));
 sg13g2_inv_1 _21403_ (.Y(_14443_),
    .A(net3321));
 sg13g2_inv_1 _21404_ (.Y(_14444_),
    .A(\u_inv.f_reg[190] ));
 sg13g2_inv_1 _21405_ (.Y(_14445_),
    .A(net3372));
 sg13g2_inv_1 _21406_ (.Y(_14446_),
    .A(net3183));
 sg13g2_inv_1 _21407_ (.Y(_14447_),
    .A(\u_inv.f_reg[193] ));
 sg13g2_inv_1 _21408_ (.Y(_14448_),
    .A(net2793));
 sg13g2_inv_1 _21409_ (.Y(_14449_),
    .A(net3197));
 sg13g2_inv_1 _21410_ (.Y(_14450_),
    .A(net2827));
 sg13g2_inv_1 _21411_ (.Y(_14451_),
    .A(\u_inv.f_reg[197] ));
 sg13g2_inv_1 _21412_ (.Y(_14452_),
    .A(net2652));
 sg13g2_inv_1 _21413_ (.Y(_14453_),
    .A(\u_inv.f_reg[199] ));
 sg13g2_inv_1 _21414_ (.Y(_14454_),
    .A(\u_inv.f_reg[200] ));
 sg13g2_inv_1 _21415_ (.Y(_14455_),
    .A(net3274));
 sg13g2_inv_1 _21416_ (.Y(_14456_),
    .A(net2803));
 sg13g2_inv_1 _21417_ (.Y(_14457_),
    .A(net2255));
 sg13g2_inv_1 _21418_ (.Y(_14458_),
    .A(\u_inv.f_reg[204] ));
 sg13g2_inv_1 _21419_ (.Y(_14459_),
    .A(\u_inv.f_reg[205] ));
 sg13g2_inv_1 _21420_ (.Y(_14460_),
    .A(net2764));
 sg13g2_inv_1 _21421_ (.Y(_14461_),
    .A(net3228));
 sg13g2_inv_1 _21422_ (.Y(_14462_),
    .A(\u_inv.f_reg[208] ));
 sg13g2_inv_1 _21423_ (.Y(_14463_),
    .A(net3239));
 sg13g2_inv_1 _21424_ (.Y(_14464_),
    .A(\u_inv.f_reg[210] ));
 sg13g2_inv_1 _21425_ (.Y(_14465_),
    .A(\u_inv.f_reg[211] ));
 sg13g2_inv_2 _21426_ (.Y(_14466_),
    .A(net2297));
 sg13g2_inv_1 _21427_ (.Y(_14467_),
    .A(\u_inv.f_reg[213] ));
 sg13g2_inv_1 _21428_ (.Y(_14468_),
    .A(net3290));
 sg13g2_inv_1 _21429_ (.Y(_14469_),
    .A(net2956));
 sg13g2_inv_1 _21430_ (.Y(_14470_),
    .A(net3172));
 sg13g2_inv_1 _21431_ (.Y(_14471_),
    .A(net3121));
 sg13g2_inv_1 _21432_ (.Y(_14472_),
    .A(net3032));
 sg13g2_inv_1 _21433_ (.Y(_14473_),
    .A(net3127));
 sg13g2_inv_1 _21434_ (.Y(_14474_),
    .A(\u_inv.f_reg[220] ));
 sg13g2_inv_1 _21435_ (.Y(_14475_),
    .A(net2763));
 sg13g2_inv_1 _21436_ (.Y(_14476_),
    .A(net1678));
 sg13g2_inv_1 _21437_ (.Y(_14477_),
    .A(\u_inv.f_reg[223] ));
 sg13g2_inv_1 _21438_ (.Y(_14478_),
    .A(net2785));
 sg13g2_inv_1 _21439_ (.Y(_14479_),
    .A(\u_inv.f_reg[225] ));
 sg13g2_inv_1 _21440_ (.Y(_14480_),
    .A(net2483));
 sg13g2_inv_1 _21441_ (.Y(_14481_),
    .A(net3119));
 sg13g2_inv_1 _21442_ (.Y(_14482_),
    .A(net3049));
 sg13g2_inv_1 _21443_ (.Y(_14483_),
    .A(\u_inv.f_reg[229] ));
 sg13g2_inv_1 _21444_ (.Y(_14484_),
    .A(net2776));
 sg13g2_inv_1 _21445_ (.Y(_14485_),
    .A(net2733));
 sg13g2_inv_1 _21446_ (.Y(_14486_),
    .A(net3159));
 sg13g2_inv_1 _21447_ (.Y(_14487_),
    .A(\u_inv.f_reg[233] ));
 sg13g2_inv_1 _21448_ (.Y(_14488_),
    .A(net2033));
 sg13g2_inv_1 _21449_ (.Y(_14489_),
    .A(\u_inv.f_reg[235] ));
 sg13g2_inv_1 _21450_ (.Y(_14490_),
    .A(net2365));
 sg13g2_inv_1 _21451_ (.Y(_14491_),
    .A(net3115));
 sg13g2_inv_1 _21452_ (.Y(_14492_),
    .A(net2656));
 sg13g2_inv_1 _21453_ (.Y(_14493_),
    .A(net3347));
 sg13g2_inv_1 _21454_ (.Y(_14494_),
    .A(\u_inv.f_reg[240] ));
 sg13g2_inv_1 _21455_ (.Y(_14495_),
    .A(\u_inv.f_reg[241] ));
 sg13g2_inv_1 _21456_ (.Y(_14496_),
    .A(net1869));
 sg13g2_inv_1 _21457_ (.Y(_14497_),
    .A(net2994));
 sg13g2_inv_1 _21458_ (.Y(_14498_),
    .A(net2717));
 sg13g2_inv_1 _21459_ (.Y(_14499_),
    .A(\u_inv.f_reg[245] ));
 sg13g2_inv_1 _21460_ (.Y(_14500_),
    .A(\u_inv.f_reg[246] ));
 sg13g2_inv_1 _21461_ (.Y(_14501_),
    .A(net3264));
 sg13g2_inv_1 _21462_ (.Y(_14502_),
    .A(net2201));
 sg13g2_inv_1 _21463_ (.Y(_14503_),
    .A(\u_inv.f_reg[249] ));
 sg13g2_inv_1 _21464_ (.Y(_14504_),
    .A(net2768));
 sg13g2_inv_1 _21465_ (.Y(_14505_),
    .A(\u_inv.f_reg[251] ));
 sg13g2_inv_1 _21466_ (.Y(_14506_),
    .A(\u_inv.f_reg[252] ));
 sg13g2_inv_1 _21467_ (.Y(_14507_),
    .A(\u_inv.f_reg[253] ));
 sg13g2_inv_1 _21468_ (.Y(_14508_),
    .A(net2196));
 sg13g2_inv_1 _21469_ (.Y(_14509_),
    .A(\u_inv.f_reg[255] ));
 sg13g2_inv_1 _21470_ (.Y(_14510_),
    .A(net5840));
 sg13g2_inv_1 _21471_ (.Y(_14511_),
    .A(inv_go));
 sg13g2_inv_4 _21472_ (.A(\shift_reg[10] ),
    .Y(_14512_));
 sg13g2_inv_2 _21473_ (.Y(_14513_),
    .A(\shift_reg[11] ));
 sg13g2_inv_1 _21474_ (.Y(_14514_),
    .A(net1837));
 sg13g2_inv_2 _21475_ (.Y(_14515_),
    .A(\shift_reg[12] ));
 sg13g2_inv_2 _21476_ (.Y(_14516_),
    .A(\shift_reg[13] ));
 sg13g2_inv_2 _21477_ (.Y(_14517_),
    .A(\shift_reg[14] ));
 sg13g2_inv_4 _21478_ (.A(net1799),
    .Y(_14518_));
 sg13g2_inv_1 _21479_ (.Y(_14519_),
    .A(net1387));
 sg13g2_inv_1 _21480_ (.Y(_14520_),
    .A(net1185));
 sg13g2_inv_1 _21481_ (.Y(_14521_),
    .A(net1095));
 sg13g2_inv_1 _21482_ (.Y(_14522_),
    .A(net1280));
 sg13g2_inv_1 _21483_ (.Y(_14523_),
    .A(net1112));
 sg13g2_inv_1 _21484_ (.Y(_14524_),
    .A(net1300));
 sg13g2_inv_1 _21485_ (.Y(_14525_),
    .A(net1294));
 sg13g2_inv_1 _21486_ (.Y(_14526_),
    .A(net1252));
 sg13g2_inv_1 _21487_ (.Y(_14527_),
    .A(net1350));
 sg13g2_inv_1 _21488_ (.Y(_14528_),
    .A(net1317));
 sg13g2_inv_1 _21489_ (.Y(_14529_),
    .A(net1382));
 sg13g2_inv_1 _21490_ (.Y(_14530_),
    .A(net1258));
 sg13g2_inv_1 _21491_ (.Y(_14531_),
    .A(net2716));
 sg13g2_inv_1 _21492_ (.Y(_14532_),
    .A(net1236));
 sg13g2_inv_1 _21493_ (.Y(_14533_),
    .A(net1102));
 sg13g2_inv_1 _21494_ (.Y(_14534_),
    .A(net2132));
 sg13g2_inv_1 _21495_ (.Y(_14535_),
    .A(net1109));
 sg13g2_inv_1 _21496_ (.Y(_14536_),
    .A(net1101));
 sg13g2_inv_1 _21497_ (.Y(_14537_),
    .A(net1336));
 sg13g2_inv_1 _21498_ (.Y(_14538_),
    .A(net1269));
 sg13g2_inv_1 _21499_ (.Y(_14539_),
    .A(net1108));
 sg13g2_inv_1 _21500_ (.Y(_14540_),
    .A(net1157));
 sg13g2_inv_1 _21501_ (.Y(_14541_),
    .A(net1347));
 sg13g2_inv_1 _21502_ (.Y(_14542_),
    .A(net1616));
 sg13g2_inv_1 _21503_ (.Y(_14543_),
    .A(net1545));
 sg13g2_inv_1 _21504_ (.Y(_14544_),
    .A(net1103));
 sg13g2_inv_1 _21505_ (.Y(_14545_),
    .A(net1104));
 sg13g2_inv_1 _21506_ (.Y(_14546_),
    .A(net1106));
 sg13g2_inv_1 _21507_ (.Y(_14547_),
    .A(net1099));
 sg13g2_inv_1 _21508_ (.Y(_14548_),
    .A(net1120));
 sg13g2_inv_1 _21509_ (.Y(_14549_),
    .A(net1211));
 sg13g2_inv_1 _21510_ (.Y(_14550_),
    .A(net1119));
 sg13g2_inv_1 _21511_ (.Y(_14551_),
    .A(net1609));
 sg13g2_inv_4 _21512_ (.A(\u_inv.d_reg[0] ),
    .Y(_14552_));
 sg13g2_inv_2 _21513_ (.Y(_14553_),
    .A(net2595));
 sg13g2_inv_1 _21514_ (.Y(_14554_),
    .A(\u_inv.d_reg[255] ));
 sg13g2_inv_2 _21515_ (.Y(_14555_),
    .A(net2966));
 sg13g2_inv_2 _21516_ (.Y(_14556_),
    .A(\u_inv.d_reg[253] ));
 sg13g2_inv_4 _21517_ (.A(\u_inv.d_reg[252] ),
    .Y(_14557_));
 sg13g2_inv_2 _21518_ (.Y(_14558_),
    .A(\u_inv.d_reg[251] ));
 sg13g2_inv_1 _21519_ (.Y(_14559_),
    .A(net2511));
 sg13g2_inv_1 _21520_ (.Y(_14560_),
    .A(\u_inv.d_reg[249] ));
 sg13g2_inv_1 _21521_ (.Y(_14561_),
    .A(\u_inv.d_reg[248] ));
 sg13g2_inv_1 _21522_ (.Y(_14562_),
    .A(\u_inv.d_reg[247] ));
 sg13g2_inv_1 _21523_ (.Y(_14563_),
    .A(net2824));
 sg13g2_inv_1 _21524_ (.Y(_14564_),
    .A(\u_inv.d_reg[245] ));
 sg13g2_inv_2 _21525_ (.Y(_14565_),
    .A(\u_inv.d_reg[244] ));
 sg13g2_inv_2 _21526_ (.Y(_14566_),
    .A(\u_inv.d_reg[243] ));
 sg13g2_inv_2 _21527_ (.Y(_14567_),
    .A(\u_inv.d_reg[242] ));
 sg13g2_inv_1 _21528_ (.Y(_14568_),
    .A(\u_inv.d_reg[241] ));
 sg13g2_inv_1 _21529_ (.Y(_14569_),
    .A(net5865));
 sg13g2_inv_2 _21530_ (.Y(_14570_),
    .A(\u_inv.d_reg[239] ));
 sg13g2_inv_2 _21531_ (.Y(_14571_),
    .A(net2724));
 sg13g2_inv_1 _21532_ (.Y(_14572_),
    .A(net2751));
 sg13g2_inv_2 _21533_ (.Y(_14573_),
    .A(net3289));
 sg13g2_inv_1 _21534_ (.Y(_14574_),
    .A(net2680));
 sg13g2_inv_2 _21535_ (.Y(_14575_),
    .A(\u_inv.d_reg[234] ));
 sg13g2_inv_1 _21536_ (.Y(_14576_),
    .A(\u_inv.d_reg[233] ));
 sg13g2_inv_1 _21537_ (.Y(_14577_),
    .A(\u_inv.d_reg[232] ));
 sg13g2_inv_1 _21538_ (.Y(_14578_),
    .A(\u_inv.d_reg[231] ));
 sg13g2_inv_1 _21539_ (.Y(_14579_),
    .A(net2923));
 sg13g2_inv_2 _21540_ (.Y(_14580_),
    .A(\u_inv.d_reg[229] ));
 sg13g2_inv_1 _21541_ (.Y(_14581_),
    .A(\u_inv.d_reg[228] ));
 sg13g2_inv_4 _21542_ (.A(\u_inv.d_reg[227] ),
    .Y(_14582_));
 sg13g2_inv_1 _21543_ (.Y(_14583_),
    .A(net2227));
 sg13g2_inv_1 _21544_ (.Y(_14584_),
    .A(\u_inv.d_reg[225] ));
 sg13g2_inv_1 _21545_ (.Y(_14585_),
    .A(\u_inv.d_reg[224] ));
 sg13g2_inv_2 _21546_ (.Y(_14586_),
    .A(net3021));
 sg13g2_inv_2 _21547_ (.Y(_14587_),
    .A(\u_inv.d_reg[222] ));
 sg13g2_inv_2 _21548_ (.Y(_14588_),
    .A(\u_inv.d_reg[221] ));
 sg13g2_inv_2 _21549_ (.Y(_14589_),
    .A(\u_inv.d_reg[220] ));
 sg13g2_inv_1 _21550_ (.Y(_14590_),
    .A(\u_inv.d_reg[219] ));
 sg13g2_inv_2 _21551_ (.Y(_14591_),
    .A(\u_inv.d_reg[218] ));
 sg13g2_inv_2 _21552_ (.Y(_14592_),
    .A(\u_inv.d_reg[217] ));
 sg13g2_inv_2 _21553_ (.Y(_14593_),
    .A(\u_inv.d_reg[216] ));
 sg13g2_inv_2 _21554_ (.Y(_14594_),
    .A(\u_inv.d_reg[215] ));
 sg13g2_inv_2 _21555_ (.Y(_14595_),
    .A(net3230));
 sg13g2_inv_2 _21556_ (.Y(_14596_),
    .A(\u_inv.d_reg[213] ));
 sg13g2_inv_1 _21557_ (.Y(_14597_),
    .A(net2153));
 sg13g2_inv_1 _21558_ (.Y(_14598_),
    .A(\u_inv.d_reg[211] ));
 sg13g2_inv_1 _21559_ (.Y(_14599_),
    .A(net2248));
 sg13g2_inv_2 _21560_ (.Y(_14600_),
    .A(\u_inv.d_reg[209] ));
 sg13g2_inv_1 _21561_ (.Y(_14601_),
    .A(\u_inv.d_reg[208] ));
 sg13g2_inv_1 _21562_ (.Y(_14602_),
    .A(\u_inv.d_reg[207] ));
 sg13g2_inv_2 _21563_ (.Y(_14603_),
    .A(\u_inv.d_reg[206] ));
 sg13g2_inv_1 _21564_ (.Y(_14604_),
    .A(\u_inv.d_reg[205] ));
 sg13g2_inv_1 _21565_ (.Y(_14605_),
    .A(\u_inv.d_reg[204] ));
 sg13g2_inv_2 _21566_ (.Y(_14606_),
    .A(\u_inv.d_reg[203] ));
 sg13g2_inv_2 _21567_ (.Y(_14607_),
    .A(net2402));
 sg13g2_inv_2 _21568_ (.Y(_14608_),
    .A(\u_inv.d_reg[201] ));
 sg13g2_inv_2 _21569_ (.Y(_14609_),
    .A(net2495));
 sg13g2_inv_1 _21570_ (.Y(_14610_),
    .A(net2969));
 sg13g2_inv_1 _21571_ (.Y(_14611_),
    .A(net2290));
 sg13g2_inv_1 _21572_ (.Y(_14612_),
    .A(\u_inv.d_reg[197] ));
 sg13g2_inv_1 _21573_ (.Y(_14613_),
    .A(\u_inv.d_reg[196] ));
 sg13g2_inv_2 _21574_ (.Y(_14614_),
    .A(net2390));
 sg13g2_inv_1 _21575_ (.Y(_14615_),
    .A(\u_inv.d_reg[194] ));
 sg13g2_inv_2 _21576_ (.Y(_14616_),
    .A(\u_inv.d_reg[193] ));
 sg13g2_inv_1 _21577_ (.Y(_14617_),
    .A(net2330));
 sg13g2_inv_2 _21578_ (.Y(_14618_),
    .A(\u_inv.d_reg[191] ));
 sg13g2_inv_1 _21579_ (.Y(_14619_),
    .A(\u_inv.d_reg[190] ));
 sg13g2_inv_2 _21580_ (.Y(_14620_),
    .A(\u_inv.d_reg[189] ));
 sg13g2_inv_1 _21581_ (.Y(_14621_),
    .A(\u_inv.d_reg[188] ));
 sg13g2_inv_2 _21582_ (.Y(_14622_),
    .A(\u_inv.d_reg[187] ));
 sg13g2_inv_1 _21583_ (.Y(_14623_),
    .A(\u_inv.d_reg[186] ));
 sg13g2_inv_1 _21584_ (.Y(_14624_),
    .A(net2042));
 sg13g2_inv_1 _21585_ (.Y(_14625_),
    .A(net5866));
 sg13g2_inv_2 _21586_ (.Y(_14626_),
    .A(net2809));
 sg13g2_inv_2 _21587_ (.Y(_14627_),
    .A(net2486));
 sg13g2_inv_2 _21588_ (.Y(_14628_),
    .A(\u_inv.d_reg[181] ));
 sg13g2_inv_2 _21589_ (.Y(_14629_),
    .A(\u_inv.d_reg[180] ));
 sg13g2_inv_1 _21590_ (.Y(_14630_),
    .A(net2173));
 sg13g2_inv_1 _21591_ (.Y(_14631_),
    .A(\u_inv.d_reg[178] ));
 sg13g2_inv_2 _21592_ (.Y(_14632_),
    .A(\u_inv.d_reg[177] ));
 sg13g2_inv_1 _21593_ (.Y(_14633_),
    .A(net2346));
 sg13g2_inv_1 _21594_ (.Y(_14634_),
    .A(\u_inv.d_reg[175] ));
 sg13g2_inv_2 _21595_ (.Y(_14635_),
    .A(\u_inv.d_reg[174] ));
 sg13g2_inv_2 _21596_ (.Y(_14636_),
    .A(net3125));
 sg13g2_inv_2 _21597_ (.Y(_14637_),
    .A(\u_inv.d_reg[172] ));
 sg13g2_inv_1 _21598_ (.Y(_14638_),
    .A(net1812));
 sg13g2_inv_1 _21599_ (.Y(_14639_),
    .A(net2498));
 sg13g2_inv_1 _21600_ (.Y(_14640_),
    .A(net2616));
 sg13g2_inv_1 _21601_ (.Y(_14641_),
    .A(\u_inv.d_reg[168] ));
 sg13g2_inv_2 _21602_ (.Y(_14642_),
    .A(\u_inv.d_reg[167] ));
 sg13g2_inv_1 _21603_ (.Y(_14643_),
    .A(\u_inv.d_reg[166] ));
 sg13g2_inv_1 _21604_ (.Y(_14644_),
    .A(\u_inv.d_reg[165] ));
 sg13g2_inv_1 _21605_ (.Y(_14645_),
    .A(net2725));
 sg13g2_inv_1 _21606_ (.Y(_14646_),
    .A(net3149));
 sg13g2_inv_2 _21607_ (.Y(_14647_),
    .A(\u_inv.d_reg[162] ));
 sg13g2_inv_1 _21608_ (.Y(_14648_),
    .A(\u_inv.d_reg[161] ));
 sg13g2_inv_1 _21609_ (.Y(_14649_),
    .A(net5868));
 sg13g2_inv_1 _21610_ (.Y(_14650_),
    .A(net3412));
 sg13g2_inv_1 _21611_ (.Y(_14651_),
    .A(\u_inv.d_reg[158] ));
 sg13g2_inv_2 _21612_ (.Y(_14652_),
    .A(net3126));
 sg13g2_inv_2 _21613_ (.Y(_14653_),
    .A(net2835));
 sg13g2_inv_1 _21614_ (.Y(_14654_),
    .A(\u_inv.d_reg[155] ));
 sg13g2_inv_2 _21615_ (.Y(_14655_),
    .A(net2429));
 sg13g2_inv_2 _21616_ (.Y(_14656_),
    .A(net2535));
 sg13g2_inv_1 _21617_ (.Y(_14657_),
    .A(\u_inv.d_reg[152] ));
 sg13g2_inv_2 _21618_ (.Y(_14658_),
    .A(\u_inv.d_reg[151] ));
 sg13g2_inv_1 _21619_ (.Y(_14659_),
    .A(\u_inv.d_reg[150] ));
 sg13g2_inv_1 _21620_ (.Y(_14660_),
    .A(\u_inv.d_reg[149] ));
 sg13g2_inv_1 _21621_ (.Y(_14661_),
    .A(\u_inv.d_reg[148] ));
 sg13g2_inv_2 _21622_ (.Y(_14662_),
    .A(net3009));
 sg13g2_inv_2 _21623_ (.Y(_14663_),
    .A(\u_inv.d_reg[146] ));
 sg13g2_inv_2 _21624_ (.Y(_14664_),
    .A(\u_inv.d_reg[145] ));
 sg13g2_inv_2 _21625_ (.Y(_14665_),
    .A(\u_inv.d_reg[144] ));
 sg13g2_inv_1 _21626_ (.Y(_14666_),
    .A(\u_inv.d_reg[143] ));
 sg13g2_inv_1 _21627_ (.Y(_14667_),
    .A(\u_inv.d_reg[142] ));
 sg13g2_inv_2 _21628_ (.Y(_14668_),
    .A(\u_inv.d_reg[141] ));
 sg13g2_inv_2 _21629_ (.Y(_14669_),
    .A(net2557));
 sg13g2_inv_2 _21630_ (.Y(_14670_),
    .A(\u_inv.d_reg[139] ));
 sg13g2_inv_1 _21631_ (.Y(_14671_),
    .A(net2428));
 sg13g2_inv_2 _21632_ (.Y(_14672_),
    .A(\u_inv.d_reg[137] ));
 sg13g2_inv_1 _21633_ (.Y(_14673_),
    .A(\u_inv.d_reg[136] ));
 sg13g2_inv_2 _21634_ (.Y(_14674_),
    .A(\u_inv.d_reg[135] ));
 sg13g2_inv_1 _21635_ (.Y(_14675_),
    .A(net2965));
 sg13g2_inv_1 _21636_ (.Y(_14676_),
    .A(\u_inv.d_reg[133] ));
 sg13g2_inv_1 _21637_ (.Y(_14677_),
    .A(net2703));
 sg13g2_inv_2 _21638_ (.Y(_14678_),
    .A(\u_inv.d_reg[131] ));
 sg13g2_inv_2 _21639_ (.Y(_14679_),
    .A(\u_inv.d_reg[130] ));
 sg13g2_inv_1 _21640_ (.Y(_14680_),
    .A(\u_inv.d_reg[129] ));
 sg13g2_inv_2 _21641_ (.Y(_14681_),
    .A(\u_inv.d_reg[128] ));
 sg13g2_inv_1 _21642_ (.Y(_14682_),
    .A(\u_inv.d_reg[127] ));
 sg13g2_inv_1 _21643_ (.Y(_14683_),
    .A(\u_inv.d_reg[126] ));
 sg13g2_inv_1 _21644_ (.Y(_14684_),
    .A(\u_inv.d_reg[125] ));
 sg13g2_inv_2 _21645_ (.Y(_14685_),
    .A(net2822));
 sg13g2_inv_2 _21646_ (.Y(_14686_),
    .A(\u_inv.d_reg[123] ));
 sg13g2_inv_1 _21647_ (.Y(_14687_),
    .A(net2363));
 sg13g2_inv_1 _21648_ (.Y(_14688_),
    .A(\u_inv.d_reg[121] ));
 sg13g2_inv_1 _21649_ (.Y(_14689_),
    .A(\u_inv.d_reg[120] ));
 sg13g2_inv_1 _21650_ (.Y(_14690_),
    .A(\u_inv.d_reg[119] ));
 sg13g2_inv_2 _21651_ (.Y(_14691_),
    .A(\u_inv.d_reg[118] ));
 sg13g2_inv_2 _21652_ (.Y(_14692_),
    .A(\u_inv.d_reg[117] ));
 sg13g2_inv_1 _21653_ (.Y(_14693_),
    .A(\u_inv.d_reg[116] ));
 sg13g2_inv_2 _21654_ (.Y(_14694_),
    .A(\u_inv.d_reg[115] ));
 sg13g2_inv_2 _21655_ (.Y(_14695_),
    .A(\u_inv.d_reg[114] ));
 sg13g2_inv_2 _21656_ (.Y(_14696_),
    .A(\u_inv.d_reg[113] ));
 sg13g2_inv_2 _21657_ (.Y(_14697_),
    .A(net2706));
 sg13g2_inv_1 _21658_ (.Y(_14698_),
    .A(\u_inv.d_reg[111] ));
 sg13g2_inv_1 _21659_ (.Y(_14699_),
    .A(\u_inv.d_reg[110] ));
 sg13g2_inv_1 _21660_ (.Y(_14700_),
    .A(\u_inv.d_reg[109] ));
 sg13g2_inv_1 _21661_ (.Y(_14701_),
    .A(\u_inv.d_reg[108] ));
 sg13g2_inv_2 _21662_ (.Y(_14702_),
    .A(\u_inv.d_reg[107] ));
 sg13g2_inv_2 _21663_ (.Y(_14703_),
    .A(\u_inv.d_reg[106] ));
 sg13g2_inv_1 _21664_ (.Y(_14704_),
    .A(\u_inv.d_reg[105] ));
 sg13g2_inv_2 _21665_ (.Y(_14705_),
    .A(\u_inv.d_reg[104] ));
 sg13g2_inv_1 _21666_ (.Y(_14706_),
    .A(\u_inv.d_reg[103] ));
 sg13g2_inv_2 _21667_ (.Y(_14707_),
    .A(\u_inv.d_reg[102] ));
 sg13g2_inv_1 _21668_ (.Y(_14708_),
    .A(\u_inv.d_reg[101] ));
 sg13g2_inv_1 _21669_ (.Y(_14709_),
    .A(\u_inv.d_reg[100] ));
 sg13g2_inv_1 _21670_ (.Y(_14710_),
    .A(\u_inv.d_reg[99] ));
 sg13g2_inv_1 _21671_ (.Y(_14711_),
    .A(net2185));
 sg13g2_inv_1 _21672_ (.Y(_14712_),
    .A(\u_inv.d_reg[97] ));
 sg13g2_inv_2 _21673_ (.Y(_14713_),
    .A(\u_inv.d_reg[96] ));
 sg13g2_inv_2 _21674_ (.Y(_14714_),
    .A(\u_inv.d_reg[95] ));
 sg13g2_inv_1 _21675_ (.Y(_14715_),
    .A(\u_inv.d_reg[94] ));
 sg13g2_inv_2 _21676_ (.Y(_14716_),
    .A(\u_inv.d_reg[93] ));
 sg13g2_inv_1 _21677_ (.Y(_14717_),
    .A(\u_inv.d_reg[92] ));
 sg13g2_inv_2 _21678_ (.Y(_14718_),
    .A(\u_inv.d_reg[91] ));
 sg13g2_inv_1 _21679_ (.Y(_14719_),
    .A(net5871));
 sg13g2_inv_2 _21680_ (.Y(_14720_),
    .A(\u_inv.d_reg[89] ));
 sg13g2_inv_2 _21681_ (.Y(_14721_),
    .A(\u_inv.d_reg[88] ));
 sg13g2_inv_1 _21682_ (.Y(_14722_),
    .A(\u_inv.d_reg[87] ));
 sg13g2_inv_2 _21683_ (.Y(_14723_),
    .A(\u_inv.d_reg[86] ));
 sg13g2_inv_1 _21684_ (.Y(_14724_),
    .A(\u_inv.d_reg[85] ));
 sg13g2_inv_2 _21685_ (.Y(_14725_),
    .A(\u_inv.d_reg[84] ));
 sg13g2_inv_1 _21686_ (.Y(_14726_),
    .A(\u_inv.d_reg[83] ));
 sg13g2_inv_1 _21687_ (.Y(_14727_),
    .A(\u_inv.d_reg[82] ));
 sg13g2_inv_1 _21688_ (.Y(_14728_),
    .A(\u_inv.d_reg[81] ));
 sg13g2_inv_1 _21689_ (.Y(_14729_),
    .A(\u_inv.d_reg[80] ));
 sg13g2_inv_2 _21690_ (.Y(_14730_),
    .A(\u_inv.d_reg[79] ));
 sg13g2_inv_1 _21691_ (.Y(_14731_),
    .A(\u_inv.d_reg[78] ));
 sg13g2_inv_1 _21692_ (.Y(_14732_),
    .A(net5872));
 sg13g2_inv_2 _21693_ (.Y(_14733_),
    .A(\u_inv.d_reg[76] ));
 sg13g2_inv_2 _21694_ (.Y(_14734_),
    .A(\u_inv.d_reg[75] ));
 sg13g2_inv_4 _21695_ (.A(\u_inv.d_reg[74] ),
    .Y(_14735_));
 sg13g2_inv_2 _21696_ (.Y(_14736_),
    .A(\u_inv.d_reg[73] ));
 sg13g2_inv_2 _21697_ (.Y(_14737_),
    .A(\u_inv.d_reg[72] ));
 sg13g2_inv_2 _21698_ (.Y(_14738_),
    .A(\u_inv.d_reg[71] ));
 sg13g2_inv_2 _21699_ (.Y(_14739_),
    .A(\u_inv.d_reg[70] ));
 sg13g2_inv_2 _21700_ (.Y(_14740_),
    .A(\u_inv.d_reg[69] ));
 sg13g2_inv_2 _21701_ (.Y(_14741_),
    .A(\u_inv.d_reg[68] ));
 sg13g2_inv_2 _21702_ (.Y(_14742_),
    .A(\u_inv.d_reg[67] ));
 sg13g2_inv_2 _21703_ (.Y(_14743_),
    .A(\u_inv.d_reg[66] ));
 sg13g2_inv_2 _21704_ (.Y(_14744_),
    .A(\u_inv.d_reg[65] ));
 sg13g2_inv_2 _21705_ (.Y(_14745_),
    .A(\u_inv.d_reg[64] ));
 sg13g2_inv_1 _21706_ (.Y(_14746_),
    .A(\u_inv.d_reg[63] ));
 sg13g2_inv_2 _21707_ (.Y(_14747_),
    .A(\u_inv.d_reg[62] ));
 sg13g2_inv_2 _21708_ (.Y(_14748_),
    .A(\u_inv.d_reg[61] ));
 sg13g2_inv_2 _21709_ (.Y(_14749_),
    .A(\u_inv.d_reg[60] ));
 sg13g2_inv_1 _21710_ (.Y(_14750_),
    .A(\u_inv.d_reg[59] ));
 sg13g2_inv_4 _21711_ (.A(\u_inv.d_reg[58] ),
    .Y(_14751_));
 sg13g2_inv_2 _21712_ (.Y(_14752_),
    .A(\u_inv.d_reg[57] ));
 sg13g2_inv_2 _21713_ (.Y(_14753_),
    .A(\u_inv.d_reg[56] ));
 sg13g2_inv_2 _21714_ (.Y(_14754_),
    .A(\u_inv.d_reg[55] ));
 sg13g2_inv_2 _21715_ (.Y(_14755_),
    .A(\u_inv.d_reg[54] ));
 sg13g2_inv_2 _21716_ (.Y(_14756_),
    .A(\u_inv.d_reg[53] ));
 sg13g2_inv_2 _21717_ (.Y(_14757_),
    .A(\u_inv.d_reg[52] ));
 sg13g2_inv_1 _21718_ (.Y(_14758_),
    .A(\u_inv.d_reg[51] ));
 sg13g2_inv_1 _21719_ (.Y(_14759_),
    .A(\u_inv.d_reg[50] ));
 sg13g2_inv_2 _21720_ (.Y(_14760_),
    .A(\u_inv.d_reg[49] ));
 sg13g2_inv_2 _21721_ (.Y(_14761_),
    .A(\u_inv.d_reg[48] ));
 sg13g2_inv_1 _21722_ (.Y(_14762_),
    .A(\u_inv.d_reg[47] ));
 sg13g2_inv_1 _21723_ (.Y(_14763_),
    .A(\u_inv.d_reg[46] ));
 sg13g2_inv_1 _21724_ (.Y(_14764_),
    .A(\u_inv.d_reg[45] ));
 sg13g2_inv_2 _21725_ (.Y(_14765_),
    .A(\u_inv.d_reg[44] ));
 sg13g2_inv_1 _21726_ (.Y(_14766_),
    .A(\u_inv.d_reg[43] ));
 sg13g2_inv_2 _21727_ (.Y(_14767_),
    .A(\u_inv.d_reg[42] ));
 sg13g2_inv_2 _21728_ (.Y(_14768_),
    .A(\u_inv.d_reg[41] ));
 sg13g2_inv_2 _21729_ (.Y(_14769_),
    .A(\u_inv.d_reg[40] ));
 sg13g2_inv_1 _21730_ (.Y(_14770_),
    .A(\u_inv.d_reg[39] ));
 sg13g2_inv_1 _21731_ (.Y(_14771_),
    .A(\u_inv.d_reg[38] ));
 sg13g2_inv_2 _21732_ (.Y(_14772_),
    .A(\u_inv.d_reg[37] ));
 sg13g2_inv_2 _21733_ (.Y(_14773_),
    .A(\u_inv.d_reg[36] ));
 sg13g2_inv_2 _21734_ (.Y(_14774_),
    .A(\u_inv.d_reg[35] ));
 sg13g2_inv_2 _21735_ (.Y(_14775_),
    .A(\u_inv.d_reg[34] ));
 sg13g2_inv_1 _21736_ (.Y(_14776_),
    .A(\u_inv.d_reg[33] ));
 sg13g2_inv_1 _21737_ (.Y(_14777_),
    .A(\u_inv.d_reg[32] ));
 sg13g2_inv_2 _21738_ (.Y(_14778_),
    .A(\u_inv.d_reg[31] ));
 sg13g2_inv_2 _21739_ (.Y(_14779_),
    .A(net2525));
 sg13g2_inv_1 _21740_ (.Y(_14780_),
    .A(\u_inv.d_reg[29] ));
 sg13g2_inv_2 _21741_ (.Y(_14781_),
    .A(\u_inv.d_reg[28] ));
 sg13g2_inv_2 _21742_ (.Y(_14782_),
    .A(\u_inv.d_reg[27] ));
 sg13g2_inv_1 _21743_ (.Y(_14783_),
    .A(\u_inv.d_reg[26] ));
 sg13g2_inv_2 _21744_ (.Y(_14784_),
    .A(\u_inv.d_reg[25] ));
 sg13g2_inv_1 _21745_ (.Y(_14785_),
    .A(\u_inv.d_reg[24] ));
 sg13g2_inv_1 _21746_ (.Y(_14786_),
    .A(\u_inv.d_reg[23] ));
 sg13g2_inv_2 _21747_ (.Y(_14787_),
    .A(net2417));
 sg13g2_inv_2 _21748_ (.Y(_14788_),
    .A(\u_inv.d_reg[21] ));
 sg13g2_inv_1 _21749_ (.Y(_14789_),
    .A(\u_inv.d_reg[20] ));
 sg13g2_inv_2 _21750_ (.Y(_14790_),
    .A(\u_inv.d_reg[19] ));
 sg13g2_inv_1 _21751_ (.Y(_14791_),
    .A(\u_inv.d_reg[18] ));
 sg13g2_inv_2 _21752_ (.Y(_14792_),
    .A(\u_inv.d_reg[17] ));
 sg13g2_inv_1 _21753_ (.Y(_14793_),
    .A(net5873));
 sg13g2_inv_2 _21754_ (.Y(_14794_),
    .A(\u_inv.d_reg[15] ));
 sg13g2_inv_2 _21755_ (.Y(_14795_),
    .A(\u_inv.d_reg[14] ));
 sg13g2_inv_2 _21756_ (.Y(_14796_),
    .A(\u_inv.d_reg[13] ));
 sg13g2_inv_2 _21757_ (.Y(_14797_),
    .A(\u_inv.d_reg[12] ));
 sg13g2_inv_1 _21758_ (.Y(_14798_),
    .A(net5874));
 sg13g2_inv_2 _21759_ (.Y(_14799_),
    .A(\u_inv.d_reg[10] ));
 sg13g2_inv_1 _21760_ (.Y(_14800_),
    .A(\u_inv.d_reg[9] ));
 sg13g2_inv_1 _21761_ (.Y(_14801_),
    .A(\u_inv.d_reg[8] ));
 sg13g2_inv_2 _21762_ (.Y(_14802_),
    .A(\u_inv.d_reg[7] ));
 sg13g2_inv_1 _21763_ (.Y(_14803_),
    .A(\u_inv.d_reg[6] ));
 sg13g2_inv_2 _21764_ (.Y(_14804_),
    .A(\u_inv.d_reg[5] ));
 sg13g2_inv_2 _21765_ (.Y(_14805_),
    .A(net2955));
 sg13g2_inv_1 _21766_ (.Y(_14806_),
    .A(\u_inv.d_reg[3] ));
 sg13g2_inv_1 _21767_ (.Y(_14807_),
    .A(\u_inv.d_reg[2] ));
 sg13g2_inv_2 _21768_ (.Y(_14808_),
    .A(\u_inv.d_reg[1] ));
 sg13g2_nand2b_2 _21769_ (.Y(_14809_),
    .B(net3437),
    .A_N(net5882));
 sg13g2_inv_2 _21770_ (.Y(uio_out[1]),
    .A(_14809_));
 sg13g2_a21oi_1 _21771_ (.A1(net5882),
    .A2(next_loaded),
    .Y(accepting),
    .B1(\state[1] ));
 sg13g2_nor2b_2 _21772_ (.A(\state[1] ),
    .B_N(net5882),
    .Y(_14810_));
 sg13g2_nand2_2 _21773_ (.Y(_14811_),
    .A(_14243_),
    .B(net5882));
 sg13g2_nor2_2 _21774_ (.A(net3417),
    .B(_14811_),
    .Y(_14812_));
 sg13g2_and3_2 _21775_ (.X(_14813_),
    .A(net1181),
    .B(net2548),
    .C(net3313));
 sg13g2_nand3_1 _21776_ (.B(net1153),
    .C(_14813_),
    .A(net2831),
    .Y(_14814_));
 sg13g2_nor2b_2 _21777_ (.A(net1830),
    .B_N(net9),
    .Y(_14815_));
 sg13g2_nand2b_2 _21778_ (.Y(_14816_),
    .B(net9),
    .A_N(net1830));
 sg13g2_nand2b_1 _21779_ (.Y(_14817_),
    .B(_14815_),
    .A_N(next_loaded));
 sg13g2_nand3b_1 _21780_ (.B(_14812_),
    .C(_14815_),
    .Y(_14818_),
    .A_N(next_loaded));
 sg13g2_a22oi_1 _21781_ (.Y(_14819_),
    .B1(_14818_),
    .B2(_14809_),
    .A2(_14814_),
    .A1(_14812_));
 sg13g2_and2_1 _21782_ (.A(_14243_),
    .B(_14819_),
    .X(_14820_));
 sg13g2_nor4_1 _21783_ (.A(net3433),
    .B(net5882),
    .C(_14814_),
    .D(_14816_),
    .Y(_14821_));
 sg13g2_or2_1 _21784_ (.X(_20878_[0]),
    .B(net3434),
    .A(_14820_));
 sg13g2_nand2_1 _21785_ (.Y(_14822_),
    .A(\u_inv.counter[6] ),
    .B(\u_inv.counter[5] ));
 sg13g2_nand3_1 _21786_ (.B(\u_inv.counter[6] ),
    .C(\u_inv.counter[5] ),
    .A(\u_inv.counter[7] ),
    .Y(_14823_));
 sg13g2_nor3_1 _21787_ (.A(net5881),
    .B(\u_inv.counter[3] ),
    .C(\u_inv.counter[4] ),
    .Y(_14824_));
 sg13g2_o21ai_1 _21788_ (.B1(_14254_),
    .Y(_14825_),
    .A1(_14823_),
    .A2(_14824_));
 sg13g2_nand2_1 _21789_ (.Y(_14826_),
    .A(net2633),
    .B(_14825_));
 sg13g2_nor2b_1 _21790_ (.A(\u_inv.state[1] ),
    .B_N(\u_inv.state[0] ),
    .Y(_14827_));
 sg13g2_nand2b_1 _21791_ (.Y(_14828_),
    .B(\u_inv.state[0] ),
    .A_N(\u_inv.state[1] ));
 sg13g2_xnor2_1 _21792_ (.Y(_14829_),
    .A(\u_inv.f_next[251] ),
    .B(\u_inv.f_reg[251] ));
 sg13g2_xnor2_1 _21793_ (.Y(_14830_),
    .A(\u_inv.f_next[250] ),
    .B(\u_inv.f_reg[250] ));
 sg13g2_xor2_1 _21794_ (.B(\u_inv.f_reg[247] ),
    .A(\u_inv.f_next[247] ),
    .X(_14831_));
 sg13g2_xnor2_1 _21795_ (.Y(_14832_),
    .A(\u_inv.f_next[247] ),
    .B(\u_inv.f_reg[247] ));
 sg13g2_nor2_1 _21796_ (.A(_13928_),
    .B(_14500_),
    .Y(_14833_));
 sg13g2_xor2_1 _21797_ (.B(\u_inv.f_reg[246] ),
    .A(\u_inv.f_next[246] ),
    .X(_14834_));
 sg13g2_xnor2_1 _21798_ (.Y(_14835_),
    .A(\u_inv.f_next[246] ),
    .B(\u_inv.f_reg[246] ));
 sg13g2_nand2_1 _21799_ (.Y(_14836_),
    .A(\u_inv.f_next[244] ),
    .B(\u_inv.f_reg[244] ));
 sg13g2_a22oi_1 _21800_ (.Y(_14837_),
    .B1(\u_inv.f_reg[245] ),
    .B2(\u_inv.f_next[245] ),
    .A2(\u_inv.f_reg[244] ),
    .A1(\u_inv.f_next[244] ));
 sg13g2_a21o_1 _21801_ (.A2(_14499_),
    .A1(_13929_),
    .B1(_14837_),
    .X(_14838_));
 sg13g2_nor3_1 _21802_ (.A(_14832_),
    .B(_14835_),
    .C(_14838_),
    .Y(_14839_));
 sg13g2_o21ai_1 _21803_ (.B1(_14833_),
    .Y(_14840_),
    .A1(\u_inv.f_next[247] ),
    .A2(\u_inv.f_reg[247] ));
 sg13g2_a21oi_1 _21804_ (.A1(\u_inv.f_next[247] ),
    .A2(\u_inv.f_reg[247] ),
    .Y(_14841_),
    .B1(_14839_));
 sg13g2_xor2_1 _21805_ (.B(\u_inv.f_reg[245] ),
    .A(\u_inv.f_next[245] ),
    .X(_14842_));
 sg13g2_xor2_1 _21806_ (.B(\u_inv.f_reg[244] ),
    .A(\u_inv.f_next[244] ),
    .X(_14843_));
 sg13g2_xnor2_1 _21807_ (.Y(_14844_),
    .A(\u_inv.f_next[244] ),
    .B(\u_inv.f_reg[244] ));
 sg13g2_nand2_1 _21808_ (.Y(_14845_),
    .A(_14842_),
    .B(_14843_));
 sg13g2_nor3_1 _21809_ (.A(_14832_),
    .B(_14835_),
    .C(_14845_),
    .Y(_14846_));
 sg13g2_nand2_1 _21810_ (.Y(_14847_),
    .A(\u_inv.f_next[222] ),
    .B(\u_inv.f_reg[222] ));
 sg13g2_xnor2_1 _21811_ (.Y(_14848_),
    .A(\u_inv.f_next[222] ),
    .B(\u_inv.f_reg[222] ));
 sg13g2_xnor2_1 _21812_ (.Y(_14849_),
    .A(\u_inv.f_next[223] ),
    .B(\u_inv.f_reg[223] ));
 sg13g2_nor2_1 _21813_ (.A(_14848_),
    .B(_14849_),
    .Y(_14850_));
 sg13g2_xnor2_1 _21814_ (.Y(_14851_),
    .A(\u_inv.f_next[221] ),
    .B(\u_inv.f_reg[221] ));
 sg13g2_nor2_1 _21815_ (.A(_13954_),
    .B(_14474_),
    .Y(_14852_));
 sg13g2_xnor2_1 _21816_ (.Y(_14853_),
    .A(\u_inv.f_next[220] ),
    .B(\u_inv.f_reg[220] ));
 sg13g2_inv_1 _21817_ (.Y(_14854_),
    .A(_14853_));
 sg13g2_nor2_1 _21818_ (.A(_14851_),
    .B(_14853_),
    .Y(_14855_));
 sg13g2_nand2_2 _21819_ (.Y(_14856_),
    .A(_14850_),
    .B(_14855_));
 sg13g2_nand2_1 _21820_ (.Y(_14857_),
    .A(\u_inv.f_next[219] ),
    .B(\u_inv.f_reg[219] ));
 sg13g2_xor2_1 _21821_ (.B(\u_inv.f_reg[219] ),
    .A(\u_inv.f_next[219] ),
    .X(_14858_));
 sg13g2_nand2_1 _21822_ (.Y(_14859_),
    .A(\u_inv.f_next[218] ),
    .B(\u_inv.f_reg[218] ));
 sg13g2_xor2_1 _21823_ (.B(\u_inv.f_reg[218] ),
    .A(\u_inv.f_next[218] ),
    .X(_14860_));
 sg13g2_xnor2_1 _21824_ (.Y(_14861_),
    .A(\u_inv.f_next[218] ),
    .B(\u_inv.f_reg[218] ));
 sg13g2_nand2_2 _21825_ (.Y(_14862_),
    .A(_14858_),
    .B(_14860_));
 sg13g2_nand2_1 _21826_ (.Y(_14863_),
    .A(\u_inv.f_next[216] ),
    .B(\u_inv.f_reg[216] ));
 sg13g2_a22oi_1 _21827_ (.Y(_14864_),
    .B1(\u_inv.f_reg[217] ),
    .B2(\u_inv.f_next[217] ),
    .A2(\u_inv.f_reg[216] ),
    .A1(\u_inv.f_next[216] ));
 sg13g2_a21o_1 _21828_ (.A2(_14471_),
    .A1(_13957_),
    .B1(_14864_),
    .X(_14865_));
 sg13g2_a21oi_1 _21829_ (.A1(_13955_),
    .A2(_14473_),
    .Y(_14866_),
    .B1(_14859_));
 sg13g2_o21ai_1 _21830_ (.B1(_14857_),
    .Y(_14867_),
    .A1(_14862_),
    .A2(_14865_));
 sg13g2_nor2_1 _21831_ (.A(_14866_),
    .B(_14867_),
    .Y(_14868_));
 sg13g2_or2_1 _21832_ (.X(_14869_),
    .B(_14868_),
    .A(_14856_));
 sg13g2_a21oi_1 _21833_ (.A1(_13951_),
    .A2(_14477_),
    .Y(_14870_),
    .B1(_14847_));
 sg13g2_a21oi_1 _21834_ (.A1(\u_inv.f_next[221] ),
    .A2(\u_inv.f_reg[221] ),
    .Y(_14871_),
    .B1(_14852_));
 sg13g2_a21oi_1 _21835_ (.A1(_13953_),
    .A2(_14475_),
    .Y(_14872_),
    .B1(_14871_));
 sg13g2_a221oi_1 _21836_ (.B2(_14872_),
    .C1(_14870_),
    .B1(_14850_),
    .A1(\u_inv.f_next[223] ),
    .Y(_14873_),
    .A2(\u_inv.f_reg[223] ));
 sg13g2_xor2_1 _21837_ (.B(\u_inv.f_reg[216] ),
    .A(\u_inv.f_next[216] ),
    .X(_14874_));
 sg13g2_xnor2_1 _21838_ (.Y(_14875_),
    .A(\u_inv.f_next[216] ),
    .B(\u_inv.f_reg[216] ));
 sg13g2_xor2_1 _21839_ (.B(\u_inv.f_reg[217] ),
    .A(\u_inv.f_next[217] ),
    .X(_14876_));
 sg13g2_and2_1 _21840_ (.A(_14874_),
    .B(_14876_),
    .X(_14877_));
 sg13g2_nand2b_1 _21841_ (.Y(_14878_),
    .B(_14877_),
    .A_N(_14862_));
 sg13g2_nor2_1 _21842_ (.A(_14856_),
    .B(_14878_),
    .Y(_14879_));
 sg13g2_nor2_1 _21843_ (.A(_13960_),
    .B(_14468_),
    .Y(_14880_));
 sg13g2_xor2_1 _21844_ (.B(\u_inv.f_reg[214] ),
    .A(\u_inv.f_next[214] ),
    .X(_14881_));
 sg13g2_xnor2_1 _21845_ (.Y(_14882_),
    .A(\u_inv.f_next[214] ),
    .B(\u_inv.f_reg[214] ));
 sg13g2_nand2_1 _21846_ (.Y(_14883_),
    .A(\u_inv.f_next[215] ),
    .B(\u_inv.f_reg[215] ));
 sg13g2_xor2_1 _21847_ (.B(\u_inv.f_reg[215] ),
    .A(\u_inv.f_next[215] ),
    .X(_14884_));
 sg13g2_xnor2_1 _21848_ (.Y(_14885_),
    .A(\u_inv.f_next[215] ),
    .B(\u_inv.f_reg[215] ));
 sg13g2_xnor2_1 _21849_ (.Y(_14886_),
    .A(\u_inv.f_next[213] ),
    .B(\u_inv.f_reg[213] ));
 sg13g2_nor2_1 _21850_ (.A(_13962_),
    .B(_14466_),
    .Y(_14887_));
 sg13g2_xnor2_1 _21851_ (.Y(_14888_),
    .A(\u_inv.f_next[212] ),
    .B(\u_inv.f_reg[212] ));
 sg13g2_inv_1 _21852_ (.Y(_14889_),
    .A(_14888_));
 sg13g2_nor2_1 _21853_ (.A(_14886_),
    .B(_14888_),
    .Y(_14890_));
 sg13g2_nand3_1 _21854_ (.B(_14884_),
    .C(_14890_),
    .A(_14881_),
    .Y(_14891_));
 sg13g2_xnor2_1 _21855_ (.Y(_14892_),
    .A(\u_inv.f_next[211] ),
    .B(\u_inv.f_reg[211] ));
 sg13g2_nor2_1 _21856_ (.A(_13964_),
    .B(_14464_),
    .Y(_14893_));
 sg13g2_xnor2_1 _21857_ (.Y(_14894_),
    .A(\u_inv.f_next[210] ),
    .B(\u_inv.f_reg[210] ));
 sg13g2_nor2_1 _21858_ (.A(_14892_),
    .B(_14894_),
    .Y(_14895_));
 sg13g2_nor2_1 _21859_ (.A(_13966_),
    .B(_14462_),
    .Y(_14896_));
 sg13g2_a21oi_1 _21860_ (.A1(\u_inv.f_next[209] ),
    .A2(\u_inv.f_reg[209] ),
    .Y(_14897_),
    .B1(_14896_));
 sg13g2_a21o_1 _21861_ (.A2(_14463_),
    .A1(_13965_),
    .B1(_14897_),
    .X(_14898_));
 sg13g2_inv_1 _21862_ (.Y(_14899_),
    .A(_14898_));
 sg13g2_a21oi_1 _21863_ (.A1(\u_inv.f_next[211] ),
    .A2(\u_inv.f_reg[211] ),
    .Y(_14900_),
    .B1(_14893_));
 sg13g2_a21oi_1 _21864_ (.A1(_13963_),
    .A2(_14465_),
    .Y(_14901_),
    .B1(_14900_));
 sg13g2_a21oi_1 _21865_ (.A1(_14895_),
    .A2(_14899_),
    .Y(_14902_),
    .B1(_14901_));
 sg13g2_inv_1 _21866_ (.Y(_14903_),
    .A(_14902_));
 sg13g2_or2_1 _21867_ (.X(_14904_),
    .B(_14902_),
    .A(_14891_));
 sg13g2_o21ai_1 _21868_ (.B1(_14880_),
    .Y(_14905_),
    .A1(\u_inv.f_next[215] ),
    .A2(\u_inv.f_reg[215] ));
 sg13g2_a21oi_1 _21869_ (.A1(\u_inv.f_next[213] ),
    .A2(\u_inv.f_reg[213] ),
    .Y(_14906_),
    .B1(_14887_));
 sg13g2_a21o_1 _21870_ (.A2(_14467_),
    .A1(_13961_),
    .B1(_14906_),
    .X(_14907_));
 sg13g2_or3_1 _21871_ (.A(_14882_),
    .B(_14885_),
    .C(_14907_),
    .X(_14908_));
 sg13g2_nand4_1 _21872_ (.B(_14904_),
    .C(_14905_),
    .A(_14883_),
    .Y(_14909_),
    .D(_14908_));
 sg13g2_nand2_1 _21873_ (.Y(_14910_),
    .A(_14879_),
    .B(_14909_));
 sg13g2_xor2_1 _21874_ (.B(\u_inv.f_reg[209] ),
    .A(\u_inv.f_next[209] ),
    .X(_14911_));
 sg13g2_xnor2_1 _21875_ (.Y(_14912_),
    .A(\u_inv.f_next[209] ),
    .B(\u_inv.f_reg[209] ));
 sg13g2_xor2_1 _21876_ (.B(\u_inv.f_reg[208] ),
    .A(\u_inv.f_next[208] ),
    .X(_14913_));
 sg13g2_xor2_1 _21877_ (.B(\u_inv.f_reg[191] ),
    .A(\u_inv.f_next[191] ),
    .X(_14914_));
 sg13g2_xnor2_1 _21878_ (.Y(_14915_),
    .A(\u_inv.f_next[191] ),
    .B(\u_inv.f_reg[191] ));
 sg13g2_nand2_1 _21879_ (.Y(_14916_),
    .A(\u_inv.f_next[190] ),
    .B(\u_inv.f_reg[190] ));
 sg13g2_xnor2_1 _21880_ (.Y(_14917_),
    .A(\u_inv.f_next[190] ),
    .B(\u_inv.f_reg[190] ));
 sg13g2_inv_1 _21881_ (.Y(_14918_),
    .A(_14917_));
 sg13g2_nor2_1 _21882_ (.A(_14915_),
    .B(_14917_),
    .Y(_14919_));
 sg13g2_nor2_1 _21883_ (.A(_13986_),
    .B(_14442_),
    .Y(_14920_));
 sg13g2_xor2_1 _21884_ (.B(\u_inv.f_reg[188] ),
    .A(\u_inv.f_next[188] ),
    .X(_14921_));
 sg13g2_xor2_1 _21885_ (.B(\u_inv.f_reg[189] ),
    .A(\u_inv.f_next[189] ),
    .X(_14922_));
 sg13g2_xnor2_1 _21886_ (.Y(_14923_),
    .A(\u_inv.f_next[189] ),
    .B(\u_inv.f_reg[189] ));
 sg13g2_and2_1 _21887_ (.A(_14921_),
    .B(_14922_),
    .X(_14924_));
 sg13g2_nand2_1 _21888_ (.Y(_14925_),
    .A(_14919_),
    .B(_14924_));
 sg13g2_xnor2_1 _21889_ (.Y(_14926_),
    .A(\u_inv.f_next[187] ),
    .B(\u_inv.f_reg[187] ));
 sg13g2_xnor2_1 _21890_ (.Y(_14927_),
    .A(\u_inv.f_next[186] ),
    .B(\u_inv.f_reg[186] ));
 sg13g2_nor2_1 _21891_ (.A(net5623),
    .B(net5622),
    .Y(_14928_));
 sg13g2_or2_1 _21892_ (.X(_14929_),
    .B(net5622),
    .A(net5623));
 sg13g2_xor2_1 _21893_ (.B(\u_inv.f_reg[185] ),
    .A(\u_inv.f_next[185] ),
    .X(_14930_));
 sg13g2_nand2_1 _21894_ (.Y(_14931_),
    .A(\u_inv.f_next[184] ),
    .B(\u_inv.f_reg[184] ));
 sg13g2_xor2_1 _21895_ (.B(\u_inv.f_reg[184] ),
    .A(\u_inv.f_next[184] ),
    .X(_14932_));
 sg13g2_and2_1 _21896_ (.A(_14930_),
    .B(_14932_),
    .X(_14933_));
 sg13g2_and4_1 _21897_ (.A(_14919_),
    .B(_14924_),
    .C(_14928_),
    .D(_14933_),
    .X(_14934_));
 sg13g2_xor2_1 _21898_ (.B(\u_inv.f_reg[183] ),
    .A(\u_inv.f_next[183] ),
    .X(_14935_));
 sg13g2_nand2_1 _21899_ (.Y(_14936_),
    .A(\u_inv.f_next[182] ),
    .B(\u_inv.f_reg[182] ));
 sg13g2_xor2_1 _21900_ (.B(\u_inv.f_reg[182] ),
    .A(\u_inv.f_next[182] ),
    .X(_14937_));
 sg13g2_inv_1 _21901_ (.Y(_14938_),
    .A(_14937_));
 sg13g2_nand2_1 _21902_ (.Y(_14939_),
    .A(_14935_),
    .B(_14937_));
 sg13g2_xor2_1 _21903_ (.B(\u_inv.f_reg[181] ),
    .A(\u_inv.f_next[181] ),
    .X(_14940_));
 sg13g2_nand2_1 _21904_ (.Y(_14941_),
    .A(\u_inv.f_next[180] ),
    .B(\u_inv.f_reg[180] ));
 sg13g2_nor2_1 _21905_ (.A(\u_inv.f_next[180] ),
    .B(\u_inv.f_reg[180] ),
    .Y(_14942_));
 sg13g2_xor2_1 _21906_ (.B(\u_inv.f_reg[180] ),
    .A(\u_inv.f_next[180] ),
    .X(_14943_));
 sg13g2_nand2_1 _21907_ (.Y(_14944_),
    .A(_14940_),
    .B(_14943_));
 sg13g2_nor2_1 _21908_ (.A(_14939_),
    .B(_14944_),
    .Y(_14945_));
 sg13g2_nor2_1 _21909_ (.A(\u_inv.f_next[179] ),
    .B(\u_inv.f_reg[179] ),
    .Y(_14946_));
 sg13g2_xor2_1 _21910_ (.B(\u_inv.f_reg[179] ),
    .A(\u_inv.f_next[179] ),
    .X(_14947_));
 sg13g2_nand2_1 _21911_ (.Y(_14948_),
    .A(\u_inv.f_next[178] ),
    .B(\u_inv.f_reg[178] ));
 sg13g2_xor2_1 _21912_ (.B(\u_inv.f_reg[178] ),
    .A(\u_inv.f_next[178] ),
    .X(_14949_));
 sg13g2_xnor2_1 _21913_ (.Y(_14950_),
    .A(\u_inv.f_next[178] ),
    .B(\u_inv.f_reg[178] ));
 sg13g2_nand2_1 _21914_ (.Y(_14951_),
    .A(_14947_),
    .B(_14949_));
 sg13g2_inv_1 _21915_ (.Y(_14952_),
    .A(_14951_));
 sg13g2_nor2_1 _21916_ (.A(_13998_),
    .B(_14430_),
    .Y(_14953_));
 sg13g2_xor2_1 _21917_ (.B(\u_inv.f_reg[176] ),
    .A(\u_inv.f_next[176] ),
    .X(_14954_));
 sg13g2_xnor2_1 _21918_ (.Y(_14955_),
    .A(\u_inv.f_next[176] ),
    .B(\u_inv.f_reg[176] ));
 sg13g2_xor2_1 _21919_ (.B(\u_inv.f_reg[177] ),
    .A(\u_inv.f_next[177] ),
    .X(_14956_));
 sg13g2_xnor2_1 _21920_ (.Y(_14957_),
    .A(\u_inv.f_next[177] ),
    .B(\u_inv.f_reg[177] ));
 sg13g2_nand2_1 _21921_ (.Y(_14958_),
    .A(_14954_),
    .B(_14956_));
 sg13g2_nor4_1 _21922_ (.A(_14939_),
    .B(_14944_),
    .C(_14951_),
    .D(_14958_),
    .Y(_14959_));
 sg13g2_inv_1 _21923_ (.Y(_14960_),
    .A(_14959_));
 sg13g2_nand2_2 _21924_ (.Y(_14961_),
    .A(_14934_),
    .B(_14959_));
 sg13g2_nand2_1 _21925_ (.Y(_14962_),
    .A(\u_inv.f_next[160] ),
    .B(\u_inv.f_reg[160] ));
 sg13g2_a22oi_1 _21926_ (.Y(_14963_),
    .B1(\u_inv.f_reg[161] ),
    .B2(\u_inv.f_next[161] ),
    .A2(\u_inv.f_reg[160] ),
    .A1(\u_inv.f_next[160] ));
 sg13g2_a21oi_1 _21927_ (.A1(_14013_),
    .A2(_14415_),
    .Y(_14964_),
    .B1(_14963_));
 sg13g2_xor2_1 _21928_ (.B(\u_inv.f_reg[167] ),
    .A(\u_inv.f_next[167] ),
    .X(_14965_));
 sg13g2_xnor2_1 _21929_ (.Y(_14966_),
    .A(\u_inv.f_next[167] ),
    .B(\u_inv.f_reg[167] ));
 sg13g2_nand2_1 _21930_ (.Y(_14967_),
    .A(\u_inv.f_next[166] ),
    .B(\u_inv.f_reg[166] ));
 sg13g2_xnor2_1 _21931_ (.Y(_14968_),
    .A(\u_inv.f_next[166] ),
    .B(\u_inv.f_reg[166] ));
 sg13g2_nor2_1 _21932_ (.A(_14966_),
    .B(_14968_),
    .Y(_14969_));
 sg13g2_nor2_1 _21933_ (.A(_14010_),
    .B(_14418_),
    .Y(_14970_));
 sg13g2_xnor2_1 _21934_ (.Y(_14971_),
    .A(\u_inv.f_next[164] ),
    .B(\u_inv.f_reg[164] ));
 sg13g2_xor2_1 _21935_ (.B(\u_inv.f_reg[165] ),
    .A(\u_inv.f_next[165] ),
    .X(_14972_));
 sg13g2_xnor2_1 _21936_ (.Y(_14973_),
    .A(\u_inv.f_next[165] ),
    .B(\u_inv.f_reg[165] ));
 sg13g2_nor2_1 _21937_ (.A(_14971_),
    .B(_14973_),
    .Y(_14974_));
 sg13g2_inv_1 _21938_ (.Y(_14975_),
    .A(_14974_));
 sg13g2_nand2_1 _21939_ (.Y(_14976_),
    .A(_14969_),
    .B(_14974_));
 sg13g2_xor2_1 _21940_ (.B(\u_inv.f_reg[163] ),
    .A(\u_inv.f_next[163] ),
    .X(_14977_));
 sg13g2_nor2_1 _21941_ (.A(_14012_),
    .B(_14416_),
    .Y(_14978_));
 sg13g2_xor2_1 _21942_ (.B(\u_inv.f_reg[162] ),
    .A(\u_inv.f_next[162] ),
    .X(_14979_));
 sg13g2_and2_1 _21943_ (.A(_14977_),
    .B(_14979_),
    .X(_14980_));
 sg13g2_nand3_1 _21944_ (.B(_14974_),
    .C(_14980_),
    .A(_14969_),
    .Y(_14981_));
 sg13g2_a21o_1 _21945_ (.A2(\u_inv.f_reg[165] ),
    .A1(\u_inv.f_next[165] ),
    .B1(_14970_),
    .X(_14982_));
 sg13g2_o21ai_1 _21946_ (.B1(_14982_),
    .Y(_14983_),
    .A1(\u_inv.f_next[165] ),
    .A2(\u_inv.f_reg[165] ));
 sg13g2_inv_1 _21947_ (.Y(_14984_),
    .A(_14983_));
 sg13g2_a21oi_1 _21948_ (.A1(_14007_),
    .A2(_14421_),
    .Y(_14985_),
    .B1(_14967_));
 sg13g2_a221oi_1 _21949_ (.B2(_14984_),
    .C1(_14985_),
    .B1(_14969_),
    .A1(\u_inv.f_next[167] ),
    .Y(_14986_),
    .A2(\u_inv.f_reg[167] ));
 sg13g2_a21oi_1 _21950_ (.A1(\u_inv.f_next[163] ),
    .A2(\u_inv.f_reg[163] ),
    .Y(_14987_),
    .B1(_14978_));
 sg13g2_a21o_2 _21951_ (.A2(_14417_),
    .A1(_14011_),
    .B1(_14987_),
    .X(_14988_));
 sg13g2_nand2_1 _21952_ (.Y(_14989_),
    .A(_14964_),
    .B(_14980_));
 sg13g2_a21oi_1 _21953_ (.A1(_14988_),
    .A2(_14989_),
    .Y(_14990_),
    .B1(_14976_));
 sg13g2_nand2b_2 _21954_ (.Y(_14991_),
    .B(_14986_),
    .A_N(_14990_));
 sg13g2_inv_1 _21955_ (.Y(_14992_),
    .A(_14991_));
 sg13g2_xor2_1 _21956_ (.B(\u_inv.f_reg[175] ),
    .A(\u_inv.f_next[175] ),
    .X(_14993_));
 sg13g2_nand2_1 _21957_ (.Y(_14994_),
    .A(\u_inv.f_next[174] ),
    .B(\u_inv.f_reg[174] ));
 sg13g2_nor2_1 _21958_ (.A(\u_inv.f_next[174] ),
    .B(\u_inv.f_reg[174] ),
    .Y(_14995_));
 sg13g2_xor2_1 _21959_ (.B(\u_inv.f_reg[174] ),
    .A(\u_inv.f_next[174] ),
    .X(_14996_));
 sg13g2_nand2_1 _21960_ (.Y(_14997_),
    .A(_14993_),
    .B(_14996_));
 sg13g2_inv_1 _21961_ (.Y(_14998_),
    .A(_14997_));
 sg13g2_xnor2_1 _21962_ (.Y(_14999_),
    .A(\u_inv.f_next[173] ),
    .B(\u_inv.f_reg[173] ));
 sg13g2_nand2_1 _21963_ (.Y(_15000_),
    .A(\u_inv.f_next[172] ),
    .B(\u_inv.f_reg[172] ));
 sg13g2_xor2_1 _21964_ (.B(\u_inv.f_reg[172] ),
    .A(\u_inv.f_next[172] ),
    .X(_15001_));
 sg13g2_xnor2_1 _21965_ (.Y(_15002_),
    .A(\u_inv.f_next[172] ),
    .B(\u_inv.f_reg[172] ));
 sg13g2_nor2_1 _21966_ (.A(_14999_),
    .B(_15002_),
    .Y(_15003_));
 sg13g2_nand2_1 _21967_ (.Y(_15004_),
    .A(_14998_),
    .B(_15003_));
 sg13g2_xor2_1 _21968_ (.B(\u_inv.f_reg[171] ),
    .A(\u_inv.f_next[171] ),
    .X(_15005_));
 sg13g2_xnor2_1 _21969_ (.Y(_15006_),
    .A(\u_inv.f_next[171] ),
    .B(\u_inv.f_reg[171] ));
 sg13g2_nand2_1 _21970_ (.Y(_15007_),
    .A(\u_inv.f_next[170] ),
    .B(\u_inv.f_reg[170] ));
 sg13g2_xnor2_1 _21971_ (.Y(_15008_),
    .A(\u_inv.f_next[170] ),
    .B(\u_inv.f_reg[170] ));
 sg13g2_nor2_2 _21972_ (.A(_15006_),
    .B(_15008_),
    .Y(_15009_));
 sg13g2_xor2_1 _21973_ (.B(\u_inv.f_reg[169] ),
    .A(\u_inv.f_next[169] ),
    .X(_15010_));
 sg13g2_xnor2_1 _21974_ (.Y(_15011_),
    .A(\u_inv.f_next[169] ),
    .B(\u_inv.f_reg[169] ));
 sg13g2_xor2_1 _21975_ (.B(\u_inv.f_reg[168] ),
    .A(\u_inv.f_next[168] ),
    .X(_15012_));
 sg13g2_xnor2_1 _21976_ (.Y(_15013_),
    .A(\u_inv.f_next[168] ),
    .B(\u_inv.f_reg[168] ));
 sg13g2_nand3_1 _21977_ (.B(_15010_),
    .C(_15012_),
    .A(_15009_),
    .Y(_15014_));
 sg13g2_nor2_1 _21978_ (.A(_15004_),
    .B(_15014_),
    .Y(_15015_));
 sg13g2_a22oi_1 _21979_ (.Y(_15016_),
    .B1(\u_inv.f_reg[173] ),
    .B2(\u_inv.f_next[173] ),
    .A2(\u_inv.f_reg[172] ),
    .A1(\u_inv.f_next[172] ));
 sg13g2_a21oi_1 _21980_ (.A1(_14001_),
    .A2(_14427_),
    .Y(_15017_),
    .B1(_15016_));
 sg13g2_a21oi_1 _21981_ (.A1(_13999_),
    .A2(_14429_),
    .Y(_15018_),
    .B1(_14994_));
 sg13g2_a221oi_1 _21982_ (.B2(_15017_),
    .C1(_15018_),
    .B1(_14998_),
    .A1(\u_inv.f_next[175] ),
    .Y(_15019_),
    .A2(\u_inv.f_reg[175] ));
 sg13g2_a22oi_1 _21983_ (.Y(_15020_),
    .B1(\u_inv.f_reg[171] ),
    .B2(\u_inv.f_next[171] ),
    .A2(\u_inv.f_reg[170] ),
    .A1(\u_inv.f_next[170] ));
 sg13g2_a21oi_1 _21984_ (.A1(_14003_),
    .A2(_14425_),
    .Y(_15021_),
    .B1(_15020_));
 sg13g2_a22oi_1 _21985_ (.Y(_15022_),
    .B1(\u_inv.f_reg[169] ),
    .B2(\u_inv.f_next[169] ),
    .A2(\u_inv.f_reg[168] ),
    .A1(\u_inv.f_next[168] ));
 sg13g2_a21oi_1 _21986_ (.A1(_14005_),
    .A2(_14423_),
    .Y(_15023_),
    .B1(_15022_));
 sg13g2_a21oi_1 _21987_ (.A1(_15009_),
    .A2(_15023_),
    .Y(_15024_),
    .B1(_15021_));
 sg13g2_o21ai_1 _21988_ (.B1(_15019_),
    .Y(_15025_),
    .A1(_15004_),
    .A2(_15024_));
 sg13g2_a21oi_2 _21989_ (.B1(_15025_),
    .Y(_15026_),
    .A2(_15015_),
    .A1(_14991_));
 sg13g2_a22oi_1 _21990_ (.Y(_15027_),
    .B1(\u_inv.f_reg[185] ),
    .B2(\u_inv.f_next[185] ),
    .A2(\u_inv.f_reg[184] ),
    .A1(\u_inv.f_next[184] ));
 sg13g2_a21oi_1 _21991_ (.A1(_13989_),
    .A2(_14439_),
    .Y(_15028_),
    .B1(_15027_));
 sg13g2_inv_1 _21992_ (.Y(_15029_),
    .A(_15028_));
 sg13g2_a22oi_1 _21993_ (.Y(_15030_),
    .B1(\u_inv.f_reg[187] ),
    .B2(\u_inv.f_next[187] ),
    .A2(\u_inv.f_reg[186] ),
    .A1(\u_inv.f_next[186] ));
 sg13g2_a21oi_1 _21994_ (.A1(_13987_),
    .A2(_14441_),
    .Y(_15031_),
    .B1(_15030_));
 sg13g2_a21oi_1 _21995_ (.A1(_14928_),
    .A2(_15028_),
    .Y(_15032_),
    .B1(_15031_));
 sg13g2_a21oi_1 _21996_ (.A1(_13983_),
    .A2(_14445_),
    .Y(_15033_),
    .B1(_14916_));
 sg13g2_a21oi_1 _21997_ (.A1(\u_inv.f_next[189] ),
    .A2(\u_inv.f_reg[189] ),
    .Y(_15034_),
    .B1(_14920_));
 sg13g2_a21oi_1 _21998_ (.A1(_13985_),
    .A2(_14443_),
    .Y(_15035_),
    .B1(_15034_));
 sg13g2_a221oi_1 _21999_ (.B2(_15035_),
    .C1(_15033_),
    .B1(_14919_),
    .A1(\u_inv.f_next[191] ),
    .Y(_15036_),
    .A2(\u_inv.f_reg[191] ));
 sg13g2_o21ai_1 _22000_ (.B1(_15036_),
    .Y(_15037_),
    .A1(_14925_),
    .A2(_15032_));
 sg13g2_a21oi_1 _22001_ (.A1(\u_inv.f_next[177] ),
    .A2(\u_inv.f_reg[177] ),
    .Y(_15038_),
    .B1(_14953_));
 sg13g2_a21oi_1 _22002_ (.A1(_13997_),
    .A2(_14431_),
    .Y(_15039_),
    .B1(_15038_));
 sg13g2_a22oi_1 _22003_ (.Y(_15040_),
    .B1(_14952_),
    .B2(_15039_),
    .A2(\u_inv.f_reg[179] ),
    .A1(\u_inv.f_next[179] ));
 sg13g2_o21ai_1 _22004_ (.B1(_15040_),
    .Y(_15041_),
    .A1(_14946_),
    .A2(_14948_));
 sg13g2_a21oi_1 _22005_ (.A1(_13991_),
    .A2(_14437_),
    .Y(_15042_),
    .B1(_14936_));
 sg13g2_a22oi_1 _22006_ (.Y(_15043_),
    .B1(\u_inv.f_reg[181] ),
    .B2(\u_inv.f_next[181] ),
    .A2(\u_inv.f_reg[180] ),
    .A1(\u_inv.f_next[180] ));
 sg13g2_a21o_1 _22007_ (.A2(_14435_),
    .A1(_13993_),
    .B1(_15043_),
    .X(_15044_));
 sg13g2_a221oi_1 _22008_ (.B2(_15041_),
    .C1(_15042_),
    .B1(_14945_),
    .A1(\u_inv.f_next[183] ),
    .Y(_15045_),
    .A2(\u_inv.f_reg[183] ));
 sg13g2_o21ai_1 _22009_ (.B1(_15045_),
    .Y(_15046_),
    .A1(_14939_),
    .A2(_15044_));
 sg13g2_nand2_1 _22010_ (.Y(_15047_),
    .A(_14934_),
    .B(_15046_));
 sg13g2_o21ai_1 _22011_ (.B1(_15047_),
    .Y(_15048_),
    .A1(_14961_),
    .A2(_15026_));
 sg13g2_nor2_2 _22012_ (.A(_15037_),
    .B(_15048_),
    .Y(_15049_));
 sg13g2_xor2_1 _22013_ (.B(\u_inv.f_reg[159] ),
    .A(\u_inv.f_next[159] ),
    .X(_15050_));
 sg13g2_nand2_1 _22014_ (.Y(_15051_),
    .A(\u_inv.f_next[158] ),
    .B(\u_inv.f_reg[158] ));
 sg13g2_xor2_1 _22015_ (.B(\u_inv.f_reg[158] ),
    .A(\u_inv.f_next[158] ),
    .X(_15052_));
 sg13g2_xnor2_1 _22016_ (.Y(_15053_),
    .A(\u_inv.f_next[158] ),
    .B(\u_inv.f_reg[158] ));
 sg13g2_and2_1 _22017_ (.A(_15050_),
    .B(_15052_),
    .X(_15054_));
 sg13g2_xor2_1 _22018_ (.B(\u_inv.f_reg[157] ),
    .A(\u_inv.f_next[157] ),
    .X(_15055_));
 sg13g2_xnor2_1 _22019_ (.Y(_15056_),
    .A(\u_inv.f_next[157] ),
    .B(\u_inv.f_reg[157] ));
 sg13g2_nor2_1 _22020_ (.A(_14018_),
    .B(_14410_),
    .Y(_15057_));
 sg13g2_xor2_1 _22021_ (.B(\u_inv.f_reg[156] ),
    .A(\u_inv.f_next[156] ),
    .X(_15058_));
 sg13g2_and2_1 _22022_ (.A(_15055_),
    .B(_15058_),
    .X(_15059_));
 sg13g2_and2_1 _22023_ (.A(_15054_),
    .B(_15059_),
    .X(_15060_));
 sg13g2_inv_1 _22024_ (.Y(_15061_),
    .A(_15060_));
 sg13g2_nand2_1 _22025_ (.Y(_15062_),
    .A(\u_inv.f_next[155] ),
    .B(\u_inv.f_reg[155] ));
 sg13g2_xor2_1 _22026_ (.B(\u_inv.f_reg[155] ),
    .A(\u_inv.f_next[155] ),
    .X(_15063_));
 sg13g2_xnor2_1 _22027_ (.Y(_15064_),
    .A(\u_inv.f_next[155] ),
    .B(\u_inv.f_reg[155] ));
 sg13g2_nand2_1 _22028_ (.Y(_15065_),
    .A(\u_inv.f_next[154] ),
    .B(\u_inv.f_reg[154] ));
 sg13g2_xor2_1 _22029_ (.B(\u_inv.f_reg[154] ),
    .A(\u_inv.f_next[154] ),
    .X(_15066_));
 sg13g2_xnor2_1 _22030_ (.Y(_15067_),
    .A(\u_inv.f_next[154] ),
    .B(\u_inv.f_reg[154] ));
 sg13g2_nand2_1 _22031_ (.Y(_15068_),
    .A(_15063_),
    .B(_15066_));
 sg13g2_xor2_1 _22032_ (.B(\u_inv.f_reg[153] ),
    .A(\u_inv.f_next[153] ),
    .X(_15069_));
 sg13g2_xnor2_1 _22033_ (.Y(_15070_),
    .A(\u_inv.f_next[153] ),
    .B(\u_inv.f_reg[153] ));
 sg13g2_nand2_1 _22034_ (.Y(_15071_),
    .A(\u_inv.f_next[152] ),
    .B(\u_inv.f_reg[152] ));
 sg13g2_xnor2_1 _22035_ (.Y(_15072_),
    .A(\u_inv.f_next[152] ),
    .B(\u_inv.f_reg[152] ));
 sg13g2_nor2_1 _22036_ (.A(_15070_),
    .B(_15072_),
    .Y(_15073_));
 sg13g2_inv_1 _22037_ (.Y(_15074_),
    .A(_15073_));
 sg13g2_nand4_1 _22038_ (.B(_15063_),
    .C(_15066_),
    .A(_15060_),
    .Y(_15075_),
    .D(_15073_));
 sg13g2_xor2_1 _22039_ (.B(\u_inv.f_reg[147] ),
    .A(\u_inv.f_next[147] ),
    .X(_15076_));
 sg13g2_xnor2_1 _22040_ (.Y(_15077_),
    .A(\u_inv.f_next[147] ),
    .B(\u_inv.f_reg[147] ));
 sg13g2_nor2_1 _22041_ (.A(_14028_),
    .B(_14400_),
    .Y(_15078_));
 sg13g2_xor2_1 _22042_ (.B(\u_inv.f_reg[146] ),
    .A(\u_inv.f_next[146] ),
    .X(_15079_));
 sg13g2_xnor2_1 _22043_ (.Y(_15080_),
    .A(\u_inv.f_next[146] ),
    .B(\u_inv.f_reg[146] ));
 sg13g2_nor2_1 _22044_ (.A(_15077_),
    .B(_15080_),
    .Y(_15081_));
 sg13g2_nor2_1 _22045_ (.A(\u_inv.f_next[145] ),
    .B(\u_inv.f_reg[145] ),
    .Y(_15082_));
 sg13g2_xnor2_1 _22046_ (.Y(_15083_),
    .A(\u_inv.f_next[145] ),
    .B(\u_inv.f_reg[145] ));
 sg13g2_nand2_1 _22047_ (.Y(_15084_),
    .A(\u_inv.f_next[151] ),
    .B(\u_inv.f_reg[151] ));
 sg13g2_xor2_1 _22048_ (.B(\u_inv.f_reg[151] ),
    .A(\u_inv.f_next[151] ),
    .X(_15085_));
 sg13g2_nand2_1 _22049_ (.Y(_15086_),
    .A(\u_inv.f_next[150] ),
    .B(\u_inv.f_reg[150] ));
 sg13g2_xor2_1 _22050_ (.B(\u_inv.f_reg[150] ),
    .A(\u_inv.f_next[150] ),
    .X(_15087_));
 sg13g2_nand2_1 _22051_ (.Y(_15088_),
    .A(_15085_),
    .B(_15087_));
 sg13g2_xor2_1 _22052_ (.B(\u_inv.f_reg[149] ),
    .A(\u_inv.f_next[149] ),
    .X(_15089_));
 sg13g2_inv_2 _22053_ (.Y(_15090_),
    .A(_15089_));
 sg13g2_nor2_1 _22054_ (.A(_14026_),
    .B(_14402_),
    .Y(_15091_));
 sg13g2_xor2_1 _22055_ (.B(\u_inv.f_reg[148] ),
    .A(\u_inv.f_next[148] ),
    .X(_15092_));
 sg13g2_nand2_1 _22056_ (.Y(_15093_),
    .A(_15089_),
    .B(_15092_));
 sg13g2_nor2_1 _22057_ (.A(_15088_),
    .B(_15093_),
    .Y(_15094_));
 sg13g2_xnor2_1 _22058_ (.Y(_15095_),
    .A(\u_inv.f_next[144] ),
    .B(\u_inv.f_reg[144] ));
 sg13g2_or4_1 _22059_ (.A(_15077_),
    .B(_15080_),
    .C(_15083_),
    .D(_15095_),
    .X(_15096_));
 sg13g2_nor4_1 _22060_ (.A(_15075_),
    .B(_15088_),
    .C(_15093_),
    .D(_15096_),
    .Y(_15097_));
 sg13g2_a22oi_1 _22061_ (.Y(_15098_),
    .B1(\u_inv.f_reg[153] ),
    .B2(\u_inv.f_next[153] ),
    .A2(\u_inv.f_reg[152] ),
    .A1(\u_inv.f_next[152] ));
 sg13g2_a21o_1 _22062_ (.A2(_14407_),
    .A1(_14021_),
    .B1(_15098_),
    .X(_15099_));
 sg13g2_a21oi_1 _22063_ (.A1(_14019_),
    .A2(_14409_),
    .Y(_15100_),
    .B1(_15065_));
 sg13g2_o21ai_1 _22064_ (.B1(_15062_),
    .Y(_15101_),
    .A1(_15068_),
    .A2(_15099_));
 sg13g2_nor2_1 _22065_ (.A(_15100_),
    .B(_15101_),
    .Y(_15102_));
 sg13g2_a21oi_1 _22066_ (.A1(_14015_),
    .A2(_14413_),
    .Y(_15103_),
    .B1(_15051_));
 sg13g2_a21oi_1 _22067_ (.A1(\u_inv.f_next[157] ),
    .A2(\u_inv.f_reg[157] ),
    .Y(_15104_),
    .B1(_15057_));
 sg13g2_a21oi_1 _22068_ (.A1(_14017_),
    .A2(_14411_),
    .Y(_15105_),
    .B1(_15104_));
 sg13g2_a221oi_1 _22069_ (.B2(_15105_),
    .C1(_15103_),
    .B1(_15054_),
    .A1(\u_inv.f_next[159] ),
    .Y(_15106_),
    .A2(\u_inv.f_reg[159] ));
 sg13g2_o21ai_1 _22070_ (.B1(_15106_),
    .Y(_15107_),
    .A1(_15061_),
    .A2(_15102_));
 sg13g2_a21oi_1 _22071_ (.A1(\u_inv.f_next[149] ),
    .A2(\u_inv.f_reg[149] ),
    .Y(_15108_),
    .B1(_15091_));
 sg13g2_a21o_1 _22072_ (.A2(_14403_),
    .A1(_14025_),
    .B1(_15108_),
    .X(_15109_));
 sg13g2_a21oi_1 _22073_ (.A1(_14023_),
    .A2(_14405_),
    .Y(_15110_),
    .B1(_15086_));
 sg13g2_o21ai_1 _22074_ (.B1(_15084_),
    .Y(_15111_),
    .A1(_15088_),
    .A2(_15109_));
 sg13g2_nor2_1 _22075_ (.A(_15110_),
    .B(_15111_),
    .Y(_15112_));
 sg13g2_a22oi_1 _22076_ (.Y(_15113_),
    .B1(\u_inv.f_reg[145] ),
    .B2(\u_inv.f_next[145] ),
    .A2(\u_inv.f_reg[144] ),
    .A1(\u_inv.f_next[144] ));
 sg13g2_nor2_1 _22077_ (.A(_15082_),
    .B(_15113_),
    .Y(_15114_));
 sg13g2_o21ai_1 _22078_ (.B1(_15078_),
    .Y(_15115_),
    .A1(\u_inv.f_next[147] ),
    .A2(\u_inv.f_reg[147] ));
 sg13g2_a22oi_1 _22079_ (.Y(_15116_),
    .B1(_15081_),
    .B2(_15114_),
    .A2(\u_inv.f_reg[147] ),
    .A1(\u_inv.f_next[147] ));
 sg13g2_nand2_2 _22080_ (.Y(_15117_),
    .A(_15115_),
    .B(_15116_));
 sg13g2_nand2_1 _22081_ (.Y(_15118_),
    .A(_15094_),
    .B(_15117_));
 sg13g2_a21oi_1 _22082_ (.A1(_15112_),
    .A2(_15118_),
    .Y(_15119_),
    .B1(_15075_));
 sg13g2_nand2_1 _22083_ (.Y(_15120_),
    .A(\u_inv.f_next[102] ),
    .B(\u_inv.f_reg[102] ));
 sg13g2_a22oi_1 _22084_ (.Y(_15121_),
    .B1(\u_inv.f_reg[103] ),
    .B2(\u_inv.f_next[103] ),
    .A2(\u_inv.f_reg[102] ),
    .A1(\u_inv.f_next[102] ));
 sg13g2_a21oi_1 _22085_ (.A1(_14071_),
    .A2(_14357_),
    .Y(_15122_),
    .B1(_15121_));
 sg13g2_xor2_1 _22086_ (.B(\u_inv.f_reg[103] ),
    .A(\u_inv.f_next[103] ),
    .X(_15123_));
 sg13g2_xor2_1 _22087_ (.B(\u_inv.f_reg[102] ),
    .A(\u_inv.f_next[102] ),
    .X(_15124_));
 sg13g2_xnor2_1 _22088_ (.Y(_15125_),
    .A(\u_inv.f_next[102] ),
    .B(\u_inv.f_reg[102] ));
 sg13g2_nand2_1 _22089_ (.Y(_15126_),
    .A(_15123_),
    .B(_15124_));
 sg13g2_xor2_1 _22090_ (.B(\u_inv.f_reg[101] ),
    .A(\u_inv.f_next[101] ),
    .X(_15127_));
 sg13g2_inv_2 _22091_ (.Y(_15128_),
    .A(_15127_));
 sg13g2_nor2_1 _22092_ (.A(_14074_),
    .B(_14354_),
    .Y(_15129_));
 sg13g2_xor2_1 _22093_ (.B(\u_inv.f_reg[100] ),
    .A(\u_inv.f_next[100] ),
    .X(_15130_));
 sg13g2_and2_1 _22094_ (.A(_15127_),
    .B(_15130_),
    .X(_15131_));
 sg13g2_nand2_1 _22095_ (.Y(_15132_),
    .A(\u_inv.f_next[99] ),
    .B(_14353_));
 sg13g2_xor2_1 _22096_ (.B(\u_inv.f_reg[99] ),
    .A(\u_inv.f_next[99] ),
    .X(_15133_));
 sg13g2_nand2_1 _22097_ (.Y(_15134_),
    .A(\u_inv.f_next[98] ),
    .B(\u_inv.f_reg[98] ));
 sg13g2_xor2_1 _22098_ (.B(\u_inv.f_reg[98] ),
    .A(\u_inv.f_next[98] ),
    .X(_15135_));
 sg13g2_xnor2_1 _22099_ (.Y(_15136_),
    .A(\u_inv.f_next[98] ),
    .B(\u_inv.f_reg[98] ));
 sg13g2_nand2_1 _22100_ (.Y(_15137_),
    .A(_15133_),
    .B(_15135_));
 sg13g2_a22oi_1 _22101_ (.Y(_15138_),
    .B1(\u_inv.f_reg[97] ),
    .B2(\u_inv.f_next[97] ),
    .A2(\u_inv.f_reg[96] ),
    .A1(\u_inv.f_next[96] ));
 sg13g2_a21oi_1 _22102_ (.A1(_14077_),
    .A2(_14351_),
    .Y(_15139_),
    .B1(_15138_));
 sg13g2_nor2b_1 _22103_ (.A(_15137_),
    .B_N(_15139_),
    .Y(_15140_));
 sg13g2_a22oi_1 _22104_ (.Y(_15141_),
    .B1(\u_inv.f_reg[99] ),
    .B2(\u_inv.f_next[99] ),
    .A2(\u_inv.f_reg[98] ),
    .A1(\u_inv.f_next[98] ));
 sg13g2_a21oi_1 _22105_ (.A1(_14075_),
    .A2(_14353_),
    .Y(_15142_),
    .B1(_15141_));
 sg13g2_inv_1 _22106_ (.Y(_15143_),
    .A(_15142_));
 sg13g2_o21ai_1 _22107_ (.B1(_15131_),
    .Y(_15144_),
    .A1(_15140_),
    .A2(_15142_));
 sg13g2_a21oi_1 _22108_ (.A1(\u_inv.f_next[101] ),
    .A2(\u_inv.f_reg[101] ),
    .Y(_15145_),
    .B1(_15129_));
 sg13g2_a21o_1 _22109_ (.A2(_14355_),
    .A1(_14073_),
    .B1(_15145_),
    .X(_15146_));
 sg13g2_inv_1 _22110_ (.Y(_15147_),
    .A(_15146_));
 sg13g2_a21oi_1 _22111_ (.A1(_15144_),
    .A2(_15146_),
    .Y(_15148_),
    .B1(_15126_));
 sg13g2_nor2_2 _22112_ (.A(_15122_),
    .B(_15148_),
    .Y(_15149_));
 sg13g2_xor2_1 _22113_ (.B(\u_inv.f_reg[87] ),
    .A(\u_inv.f_next[87] ),
    .X(_15150_));
 sg13g2_xnor2_1 _22114_ (.Y(_15151_),
    .A(\u_inv.f_next[87] ),
    .B(\u_inv.f_reg[87] ));
 sg13g2_nand2_1 _22115_ (.Y(_15152_),
    .A(\u_inv.f_next[86] ),
    .B(\u_inv.f_reg[86] ));
 sg13g2_xnor2_1 _22116_ (.Y(_15153_),
    .A(\u_inv.f_next[86] ),
    .B(\u_inv.f_reg[86] ));
 sg13g2_nor2_1 _22117_ (.A(_15151_),
    .B(_15153_),
    .Y(_15154_));
 sg13g2_nor2_1 _22118_ (.A(\u_inv.f_next[85] ),
    .B(\u_inv.f_reg[85] ),
    .Y(_15155_));
 sg13g2_nand2_1 _22119_ (.Y(_15156_),
    .A(_14089_),
    .B(_14339_));
 sg13g2_nand2_1 _22120_ (.Y(_15157_),
    .A(\u_inv.f_next[85] ),
    .B(\u_inv.f_reg[85] ));
 sg13g2_nand2_1 _22121_ (.Y(_15158_),
    .A(\u_inv.f_next[84] ),
    .B(\u_inv.f_reg[84] ));
 sg13g2_o21ai_1 _22122_ (.B1(_15157_),
    .Y(_15159_),
    .A1(_15155_),
    .A2(_15158_));
 sg13g2_a21oi_1 _22123_ (.A1(_14087_),
    .A2(_14341_),
    .Y(_15160_),
    .B1(_15152_));
 sg13g2_a221oi_1 _22124_ (.B2(_15159_),
    .C1(_15160_),
    .B1(_15154_),
    .A1(\u_inv.f_next[87] ),
    .Y(_15161_),
    .A2(\u_inv.f_reg[87] ));
 sg13g2_inv_1 _22125_ (.Y(_15162_),
    .A(_15161_));
 sg13g2_nand2_2 _22126_ (.Y(_15163_),
    .A(_15156_),
    .B(_15157_));
 sg13g2_xor2_1 _22127_ (.B(\u_inv.f_reg[84] ),
    .A(\u_inv.f_next[84] ),
    .X(_15164_));
 sg13g2_inv_2 _22128_ (.Y(_15165_),
    .A(_15164_));
 sg13g2_nor2_1 _22129_ (.A(_15163_),
    .B(_15165_),
    .Y(_15166_));
 sg13g2_a21oi_2 _22130_ (.B1(_15162_),
    .Y(_15167_),
    .A2(_15166_),
    .A1(_15154_));
 sg13g2_inv_1 _22131_ (.Y(_15168_),
    .A(_15167_));
 sg13g2_xor2_1 _22132_ (.B(\u_inv.f_reg[71] ),
    .A(\u_inv.f_next[71] ),
    .X(_15169_));
 sg13g2_xnor2_1 _22133_ (.Y(_15170_),
    .A(\u_inv.f_next[71] ),
    .B(\u_inv.f_reg[71] ));
 sg13g2_nand2_1 _22134_ (.Y(_15171_),
    .A(\u_inv.f_next[70] ),
    .B(\u_inv.f_reg[70] ));
 sg13g2_xnor2_1 _22135_ (.Y(_15172_),
    .A(\u_inv.f_next[70] ),
    .B(\u_inv.f_reg[70] ));
 sg13g2_nor2_1 _22136_ (.A(_15170_),
    .B(_15172_),
    .Y(_15173_));
 sg13g2_nor2_1 _22137_ (.A(_14106_),
    .B(_14322_),
    .Y(_15174_));
 sg13g2_nand2_1 _22138_ (.Y(_15175_),
    .A(_14106_),
    .B(_14322_));
 sg13g2_nand2b_2 _22139_ (.Y(_15176_),
    .B(_15175_),
    .A_N(_15174_));
 sg13g2_xor2_1 _22140_ (.B(\u_inv.f_reg[69] ),
    .A(\u_inv.f_next[69] ),
    .X(_15177_));
 sg13g2_nor2b_1 _22141_ (.A(_15176_),
    .B_N(_15177_),
    .Y(_15178_));
 sg13g2_nand2_1 _22142_ (.Y(_15179_),
    .A(_15173_),
    .B(_15178_));
 sg13g2_xor2_1 _22143_ (.B(\u_inv.f_reg[67] ),
    .A(\u_inv.f_next[67] ),
    .X(_15180_));
 sg13g2_xor2_1 _22144_ (.B(\u_inv.f_reg[66] ),
    .A(\u_inv.f_next[66] ),
    .X(_15181_));
 sg13g2_and2_1 _22145_ (.A(_15180_),
    .B(_15181_),
    .X(_15182_));
 sg13g2_nand2_1 _22146_ (.Y(_15183_),
    .A(_15180_),
    .B(_15181_));
 sg13g2_nor2_1 _22147_ (.A(\u_inv.f_next[65] ),
    .B(\u_inv.f_reg[65] ),
    .Y(_15184_));
 sg13g2_nand2_1 _22148_ (.Y(_15185_),
    .A(\u_inv.f_next[65] ),
    .B(\u_inv.f_reg[65] ));
 sg13g2_nand2_1 _22149_ (.Y(_15186_),
    .A(\u_inv.f_next[64] ),
    .B(\u_inv.f_reg[64] ));
 sg13g2_o21ai_1 _22150_ (.B1(_15185_),
    .Y(_15187_),
    .A1(_15184_),
    .A2(_15186_));
 sg13g2_a22oi_1 _22151_ (.Y(_15188_),
    .B1(\u_inv.f_reg[67] ),
    .B2(\u_inv.f_next[67] ),
    .A2(\u_inv.f_reg[66] ),
    .A1(\u_inv.f_next[66] ));
 sg13g2_a21oi_1 _22152_ (.A1(_14107_),
    .A2(_14321_),
    .Y(_15189_),
    .B1(_15188_));
 sg13g2_inv_1 _22153_ (.Y(_15190_),
    .A(_15189_));
 sg13g2_a21oi_1 _22154_ (.A1(_15182_),
    .A2(_15187_),
    .Y(_15191_),
    .B1(_15189_));
 sg13g2_a21oi_1 _22155_ (.A1(_14103_),
    .A2(_14325_),
    .Y(_15192_),
    .B1(_15171_));
 sg13g2_a21oi_1 _22156_ (.A1(\u_inv.f_next[71] ),
    .A2(\u_inv.f_reg[71] ),
    .Y(_15193_),
    .B1(_15192_));
 sg13g2_a21oi_1 _22157_ (.A1(\u_inv.f_next[69] ),
    .A2(\u_inv.f_reg[69] ),
    .Y(_15194_),
    .B1(_15174_));
 sg13g2_a21oi_1 _22158_ (.A1(_14105_),
    .A2(_14323_),
    .Y(_15195_),
    .B1(_15194_));
 sg13g2_o21ai_1 _22159_ (.B1(_15193_),
    .Y(_15196_),
    .A1(_15179_),
    .A2(_15191_));
 sg13g2_a21oi_1 _22160_ (.A1(_15173_),
    .A2(_15195_),
    .Y(_15197_),
    .B1(_15196_));
 sg13g2_xnor2_1 _22161_ (.Y(_15198_),
    .A(\u_inv.f_next[63] ),
    .B(\u_inv.f_reg[63] ));
 sg13g2_nand2_1 _22162_ (.Y(_15199_),
    .A(\u_inv.f_next[62] ),
    .B(\u_inv.f_reg[62] ));
 sg13g2_xnor2_1 _22163_ (.Y(_15200_),
    .A(\u_inv.f_next[62] ),
    .B(\u_inv.f_reg[62] ));
 sg13g2_nor2_1 _22164_ (.A(_15198_),
    .B(_15200_),
    .Y(_15201_));
 sg13g2_nor2_1 _22165_ (.A(_14114_),
    .B(_14314_),
    .Y(_15202_));
 sg13g2_xor2_1 _22166_ (.B(\u_inv.f_reg[60] ),
    .A(\u_inv.f_next[60] ),
    .X(_15203_));
 sg13g2_xnor2_1 _22167_ (.Y(_15204_),
    .A(\u_inv.f_next[60] ),
    .B(\u_inv.f_reg[60] ));
 sg13g2_xnor2_1 _22168_ (.Y(_15205_),
    .A(\u_inv.f_next[61] ),
    .B(\u_inv.f_reg[61] ));
 sg13g2_nor2_1 _22169_ (.A(_15204_),
    .B(_15205_),
    .Y(_15206_));
 sg13g2_nand2_1 _22170_ (.Y(_15207_),
    .A(_15201_),
    .B(_15206_));
 sg13g2_xor2_1 _22171_ (.B(\u_inv.f_reg[59] ),
    .A(\u_inv.f_next[59] ),
    .X(_15208_));
 sg13g2_nand2_1 _22172_ (.Y(_15209_),
    .A(\u_inv.f_next[58] ),
    .B(\u_inv.f_reg[58] ));
 sg13g2_xor2_1 _22173_ (.B(\u_inv.f_reg[58] ),
    .A(\u_inv.f_next[58] ),
    .X(_15210_));
 sg13g2_xnor2_1 _22174_ (.Y(_15211_),
    .A(\u_inv.f_next[58] ),
    .B(\u_inv.f_reg[58] ));
 sg13g2_nand2_1 _22175_ (.Y(_15212_),
    .A(_15208_),
    .B(_15210_));
 sg13g2_nor2_1 _22176_ (.A(_14118_),
    .B(_14310_),
    .Y(_15213_));
 sg13g2_a21oi_1 _22177_ (.A1(\u_inv.f_next[57] ),
    .A2(\u_inv.f_reg[57] ),
    .Y(_15214_),
    .B1(_15213_));
 sg13g2_a21oi_1 _22178_ (.A1(_14117_),
    .A2(_14311_),
    .Y(_15215_),
    .B1(_15214_));
 sg13g2_nor2b_1 _22179_ (.A(_15212_),
    .B_N(_15215_),
    .Y(_15216_));
 sg13g2_a22oi_1 _22180_ (.Y(_15217_),
    .B1(\u_inv.f_reg[59] ),
    .B2(\u_inv.f_next[59] ),
    .A2(\u_inv.f_reg[58] ),
    .A1(\u_inv.f_next[58] ));
 sg13g2_a21oi_1 _22181_ (.A1(_14115_),
    .A2(_14313_),
    .Y(_15218_),
    .B1(_15217_));
 sg13g2_inv_1 _22182_ (.Y(_15219_),
    .A(_15218_));
 sg13g2_nor2_1 _22183_ (.A(_15216_),
    .B(_15218_),
    .Y(_15220_));
 sg13g2_a21oi_1 _22184_ (.A1(_14111_),
    .A2(_14317_),
    .Y(_15221_),
    .B1(_15199_));
 sg13g2_a21oi_1 _22185_ (.A1(\u_inv.f_next[61] ),
    .A2(\u_inv.f_reg[61] ),
    .Y(_15222_),
    .B1(_15202_));
 sg13g2_a21oi_1 _22186_ (.A1(_14113_),
    .A2(_14315_),
    .Y(_15223_),
    .B1(_15222_));
 sg13g2_a221oi_1 _22187_ (.B2(_15223_),
    .C1(_15221_),
    .B1(_15201_),
    .A1(\u_inv.f_next[63] ),
    .Y(_15224_),
    .A2(\u_inv.f_reg[63] ));
 sg13g2_o21ai_1 _22188_ (.B1(_15224_),
    .Y(_15225_),
    .A1(_15207_),
    .A2(_15220_));
 sg13g2_xor2_1 _22189_ (.B(\u_inv.f_reg[39] ),
    .A(\u_inv.f_next[39] ),
    .X(_15226_));
 sg13g2_nand2_1 _22190_ (.Y(_15227_),
    .A(\u_inv.f_next[38] ),
    .B(\u_inv.f_reg[38] ));
 sg13g2_nor2_1 _22191_ (.A(\u_inv.f_next[38] ),
    .B(\u_inv.f_reg[38] ),
    .Y(_15228_));
 sg13g2_xor2_1 _22192_ (.B(\u_inv.f_reg[38] ),
    .A(\u_inv.f_next[38] ),
    .X(_15229_));
 sg13g2_and2_1 _22193_ (.A(_15226_),
    .B(_15229_),
    .X(_15230_));
 sg13g2_nand2_1 _22194_ (.Y(_15231_),
    .A(\u_inv.f_next[36] ),
    .B(\u_inv.f_reg[36] ));
 sg13g2_xor2_1 _22195_ (.B(\u_inv.f_reg[36] ),
    .A(\u_inv.f_next[36] ),
    .X(_15232_));
 sg13g2_xnor2_1 _22196_ (.Y(_15233_),
    .A(\u_inv.f_next[36] ),
    .B(\u_inv.f_reg[36] ));
 sg13g2_xor2_1 _22197_ (.B(\u_inv.f_reg[37] ),
    .A(\u_inv.f_next[37] ),
    .X(_15234_));
 sg13g2_xnor2_1 _22198_ (.Y(_15235_),
    .A(\u_inv.f_next[37] ),
    .B(\u_inv.f_reg[37] ));
 sg13g2_nor2_1 _22199_ (.A(_15233_),
    .B(_15235_),
    .Y(_15236_));
 sg13g2_nand2_1 _22200_ (.Y(_15237_),
    .A(_15230_),
    .B(_15236_));
 sg13g2_xor2_1 _22201_ (.B(\u_inv.f_reg[35] ),
    .A(\u_inv.f_next[35] ),
    .X(_15238_));
 sg13g2_xnor2_1 _22202_ (.Y(_15239_),
    .A(\u_inv.f_next[35] ),
    .B(\u_inv.f_reg[35] ));
 sg13g2_nand2_1 _22203_ (.Y(_15240_),
    .A(\u_inv.f_next[34] ),
    .B(\u_inv.f_reg[34] ));
 sg13g2_xnor2_1 _22204_ (.Y(_15241_),
    .A(\u_inv.f_next[34] ),
    .B(\u_inv.f_reg[34] ));
 sg13g2_nor2_1 _22205_ (.A(_15239_),
    .B(_15241_),
    .Y(_15242_));
 sg13g2_nor2_1 _22206_ (.A(_14142_),
    .B(_14286_),
    .Y(_15243_));
 sg13g2_a21oi_1 _22207_ (.A1(\u_inv.f_next[33] ),
    .A2(\u_inv.f_reg[33] ),
    .Y(_15244_),
    .B1(_15243_));
 sg13g2_a21oi_1 _22208_ (.A1(_14141_),
    .A2(_14287_),
    .Y(_15245_),
    .B1(_15244_));
 sg13g2_a22oi_1 _22209_ (.Y(_15246_),
    .B1(\u_inv.f_reg[35] ),
    .B2(\u_inv.f_next[35] ),
    .A2(\u_inv.f_reg[34] ),
    .A1(\u_inv.f_next[34] ));
 sg13g2_a21oi_1 _22210_ (.A1(_14139_),
    .A2(_14289_),
    .Y(_15247_),
    .B1(_15246_));
 sg13g2_a21oi_1 _22211_ (.A1(_15242_),
    .A2(_15245_),
    .Y(_15248_),
    .B1(_15247_));
 sg13g2_a22oi_1 _22212_ (.Y(_15249_),
    .B1(\u_inv.f_reg[37] ),
    .B2(\u_inv.f_next[37] ),
    .A2(\u_inv.f_reg[36] ),
    .A1(\u_inv.f_next[36] ));
 sg13g2_a21oi_1 _22213_ (.A1(_14137_),
    .A2(_14291_),
    .Y(_15250_),
    .B1(_15249_));
 sg13g2_a21oi_1 _22214_ (.A1(_14135_),
    .A2(_14293_),
    .Y(_15251_),
    .B1(_15227_));
 sg13g2_a221oi_1 _22215_ (.B2(_15250_),
    .C1(_15251_),
    .B1(_15230_),
    .A1(\u_inv.f_next[39] ),
    .Y(_15252_),
    .A2(\u_inv.f_reg[39] ));
 sg13g2_o21ai_1 _22216_ (.B1(_15252_),
    .Y(_15253_),
    .A1(_15237_),
    .A2(_15248_));
 sg13g2_nand2_1 _22217_ (.Y(_15254_),
    .A(\u_inv.f_next[15] ),
    .B(\u_inv.f_reg[15] ));
 sg13g2_nand2_1 _22218_ (.Y(_15255_),
    .A(_14159_),
    .B(_14269_));
 sg13g2_nand2_1 _22219_ (.Y(_15256_),
    .A(\u_inv.f_next[13] ),
    .B(\u_inv.f_reg[13] ));
 sg13g2_nor2_1 _22220_ (.A(\u_inv.f_next[13] ),
    .B(\u_inv.f_reg[13] ),
    .Y(_15257_));
 sg13g2_nand2_1 _22221_ (.Y(_15258_),
    .A(\u_inv.f_next[12] ),
    .B(\u_inv.f_reg[12] ));
 sg13g2_nand2_1 _22222_ (.Y(_15259_),
    .A(_14163_),
    .B(_14265_));
 sg13g2_nand2_2 _22223_ (.Y(_15260_),
    .A(\u_inv.f_next[11] ),
    .B(\u_inv.f_reg[11] ));
 sg13g2_nor2_1 _22224_ (.A(_14164_),
    .B(_14264_),
    .Y(_15261_));
 sg13g2_xor2_1 _22225_ (.B(\u_inv.f_reg[10] ),
    .A(\u_inv.f_next[10] ),
    .X(_15262_));
 sg13g2_inv_1 _22226_ (.Y(_15263_),
    .A(_15262_));
 sg13g2_nor2_1 _22227_ (.A(\u_inv.f_next[9] ),
    .B(\u_inv.f_reg[9] ),
    .Y(_15264_));
 sg13g2_nor2_1 _22228_ (.A(_14166_),
    .B(_14262_),
    .Y(_15265_));
 sg13g2_xor2_1 _22229_ (.B(\u_inv.f_reg[8] ),
    .A(\u_inv.f_next[8] ),
    .X(_15266_));
 sg13g2_nand2_1 _22230_ (.Y(_15267_),
    .A(\u_inv.f_next[7] ),
    .B(\u_inv.f_reg[7] ));
 sg13g2_xnor2_1 _22231_ (.Y(_15268_),
    .A(\u_inv.f_next[7] ),
    .B(\u_inv.f_reg[7] ));
 sg13g2_and2_1 _22232_ (.A(\u_inv.f_next[6] ),
    .B(\u_inv.f_reg[6] ),
    .X(_15269_));
 sg13g2_xor2_1 _22233_ (.B(\u_inv.f_reg[6] ),
    .A(\u_inv.f_next[6] ),
    .X(_15270_));
 sg13g2_nand2_1 _22234_ (.Y(_15271_),
    .A(\u_inv.f_next[5] ),
    .B(\u_inv.f_reg[5] ));
 sg13g2_xnor2_1 _22235_ (.Y(_15272_),
    .A(\u_inv.f_next[5] ),
    .B(\u_inv.f_reg[5] ));
 sg13g2_nand2_1 _22236_ (.Y(_15273_),
    .A(\u_inv.f_next[4] ),
    .B(\u_inv.f_reg[4] ));
 sg13g2_inv_1 _22237_ (.Y(_15274_),
    .A(_15273_));
 sg13g2_xor2_1 _22238_ (.B(\u_inv.f_reg[4] ),
    .A(\u_inv.f_next[4] ),
    .X(_15275_));
 sg13g2_nand2_1 _22239_ (.Y(_15276_),
    .A(\u_inv.f_next[3] ),
    .B(\u_inv.f_reg[3] ));
 sg13g2_xnor2_1 _22240_ (.Y(_15277_),
    .A(\u_inv.f_next[3] ),
    .B(\u_inv.f_reg[3] ));
 sg13g2_nand2_1 _22241_ (.Y(_15278_),
    .A(\u_inv.f_next[2] ),
    .B(\u_inv.f_reg[2] ));
 sg13g2_inv_1 _22242_ (.Y(_15279_),
    .A(_15278_));
 sg13g2_or2_1 _22243_ (.X(_15280_),
    .B(\u_inv.f_reg[2] ),
    .A(\u_inv.f_next[2] ));
 sg13g2_and2_1 _22244_ (.A(_15278_),
    .B(_15280_),
    .X(_15281_));
 sg13g2_nand2_1 _22245_ (.Y(_15282_),
    .A(\u_inv.f_next[1] ),
    .B(\u_inv.f_reg[1] ));
 sg13g2_nor2b_1 _22246_ (.A(\u_inv.f_next[1] ),
    .B_N(\u_inv.f_reg[1] ),
    .Y(_15283_));
 sg13g2_nand2b_1 _22247_ (.Y(_15284_),
    .B(\u_inv.f_next[1] ),
    .A_N(\u_inv.f_reg[1] ));
 sg13g2_xnor2_1 _22248_ (.Y(_15285_),
    .A(\u_inv.f_next[1] ),
    .B(\u_inv.f_reg[1] ));
 sg13g2_nand2_1 _22249_ (.Y(_15286_),
    .A(net5725),
    .B(\u_inv.f_reg[0] ));
 sg13g2_o21ai_1 _22250_ (.B1(_15282_),
    .Y(_15287_),
    .A1(_15285_),
    .A2(_15286_));
 sg13g2_a21oi_1 _22251_ (.A1(_15281_),
    .A2(_15287_),
    .Y(_15288_),
    .B1(_15279_));
 sg13g2_o21ai_1 _22252_ (.B1(_15276_),
    .Y(_15289_),
    .A1(_15277_),
    .A2(_15288_));
 sg13g2_a21oi_1 _22253_ (.A1(_15275_),
    .A2(_15289_),
    .Y(_15290_),
    .B1(_15274_));
 sg13g2_or2_1 _22254_ (.X(_15291_),
    .B(_15290_),
    .A(_15272_));
 sg13g2_o21ai_1 _22255_ (.B1(_15271_),
    .Y(_15292_),
    .A1(_15272_),
    .A2(_15290_));
 sg13g2_and2_1 _22256_ (.A(_15270_),
    .B(_15292_),
    .X(_15293_));
 sg13g2_a21oi_1 _22257_ (.A1(_15270_),
    .A2(_15292_),
    .Y(_15294_),
    .B1(_15269_));
 sg13g2_o21ai_1 _22258_ (.B1(_15267_),
    .Y(_15295_),
    .A1(_15268_),
    .A2(_15294_));
 sg13g2_a21o_1 _22259_ (.A2(_15295_),
    .A1(_15266_),
    .B1(_15265_),
    .X(_15296_));
 sg13g2_a221oi_1 _22260_ (.B2(_15295_),
    .C1(_15265_),
    .B1(_15266_),
    .A1(\u_inv.f_next[9] ),
    .Y(_15297_),
    .A2(\u_inv.f_reg[9] ));
 sg13g2_nor3_1 _22261_ (.A(_15263_),
    .B(_15264_),
    .C(_15297_),
    .Y(_15298_));
 sg13g2_nor2_1 _22262_ (.A(_15261_),
    .B(_15298_),
    .Y(_15299_));
 sg13g2_o21ai_1 _22263_ (.B1(_15259_),
    .Y(_15300_),
    .A1(_15261_),
    .A2(_15298_));
 sg13g2_nand2_1 _22264_ (.Y(_15301_),
    .A(_15260_),
    .B(_15300_));
 sg13g2_xor2_1 _22265_ (.B(\u_inv.f_reg[12] ),
    .A(\u_inv.f_next[12] ),
    .X(_15302_));
 sg13g2_nand2_1 _22266_ (.Y(_15303_),
    .A(_15301_),
    .B(_15302_));
 sg13g2_nand2_1 _22267_ (.Y(_15304_),
    .A(_15258_),
    .B(_15303_));
 sg13g2_o21ai_1 _22268_ (.B1(_15256_),
    .Y(_15305_),
    .A1(_15257_),
    .A2(_15258_));
 sg13g2_xor2_1 _22269_ (.B(\u_inv.f_reg[13] ),
    .A(\u_inv.f_next[13] ),
    .X(_15306_));
 sg13g2_nand2_1 _22270_ (.Y(_15307_),
    .A(_15302_),
    .B(_15306_));
 sg13g2_a21oi_2 _22271_ (.B1(_15307_),
    .Y(_15308_),
    .A2(_15300_),
    .A1(_15260_));
 sg13g2_nor2_1 _22272_ (.A(_15305_),
    .B(_15308_),
    .Y(_15309_));
 sg13g2_xor2_1 _22273_ (.B(\u_inv.f_reg[14] ),
    .A(\u_inv.f_next[14] ),
    .X(_15310_));
 sg13g2_xnor2_1 _22274_ (.Y(_15311_),
    .A(\u_inv.f_next[14] ),
    .B(\u_inv.f_reg[14] ));
 sg13g2_nor2_1 _22275_ (.A(_15309_),
    .B(_15311_),
    .Y(_15312_));
 sg13g2_a21oi_1 _22276_ (.A1(\u_inv.f_next[14] ),
    .A2(\u_inv.f_reg[14] ),
    .Y(_15313_),
    .B1(_15312_));
 sg13g2_nand3_1 _22277_ (.B(\u_inv.f_reg[14] ),
    .C(_15255_),
    .A(\u_inv.f_next[14] ),
    .Y(_15314_));
 sg13g2_nand2_2 _22278_ (.Y(_15315_),
    .A(_15254_),
    .B(_15255_));
 sg13g2_nor2_1 _22279_ (.A(_15311_),
    .B(_15315_),
    .Y(_15316_));
 sg13g2_o21ai_1 _22280_ (.B1(_15316_),
    .Y(_15317_),
    .A1(_15305_),
    .A2(_15308_));
 sg13g2_and3_2 _22281_ (.X(_15318_),
    .A(_15254_),
    .B(_15314_),
    .C(_15317_));
 sg13g2_xor2_1 _22282_ (.B(\u_inv.f_reg[19] ),
    .A(\u_inv.f_next[19] ),
    .X(_15319_));
 sg13g2_xnor2_1 _22283_ (.Y(_15320_),
    .A(\u_inv.f_next[19] ),
    .B(\u_inv.f_reg[19] ));
 sg13g2_nand2_1 _22284_ (.Y(_15321_),
    .A(\u_inv.f_next[18] ),
    .B(\u_inv.f_reg[18] ));
 sg13g2_xor2_1 _22285_ (.B(\u_inv.f_reg[18] ),
    .A(\u_inv.f_next[18] ),
    .X(_15322_));
 sg13g2_xnor2_1 _22286_ (.Y(_15323_),
    .A(\u_inv.f_next[18] ),
    .B(\u_inv.f_reg[18] ));
 sg13g2_nor2_1 _22287_ (.A(_15320_),
    .B(_15323_),
    .Y(_15324_));
 sg13g2_xor2_1 _22288_ (.B(\u_inv.f_reg[17] ),
    .A(\u_inv.f_next[17] ),
    .X(_15325_));
 sg13g2_xor2_1 _22289_ (.B(\u_inv.f_reg[16] ),
    .A(\u_inv.f_next[16] ),
    .X(_15326_));
 sg13g2_xnor2_1 _22290_ (.Y(_15327_),
    .A(\u_inv.f_next[16] ),
    .B(\u_inv.f_reg[16] ));
 sg13g2_nand2_1 _22291_ (.Y(_15328_),
    .A(net5621),
    .B(_15326_));
 sg13g2_nand3_1 _22292_ (.B(net5621),
    .C(_15326_),
    .A(_15324_),
    .Y(_15329_));
 sg13g2_a21oi_1 _22293_ (.A1(_14155_),
    .A2(_14273_),
    .Y(_15330_),
    .B1(_15321_));
 sg13g2_a22oi_1 _22294_ (.Y(_15331_),
    .B1(\u_inv.f_reg[17] ),
    .B2(\u_inv.f_next[17] ),
    .A2(\u_inv.f_reg[16] ),
    .A1(\u_inv.f_next[16] ));
 sg13g2_a21oi_1 _22295_ (.A1(_14157_),
    .A2(_14271_),
    .Y(_15332_),
    .B1(_15331_));
 sg13g2_a221oi_1 _22296_ (.B2(_15332_),
    .C1(_15330_),
    .B1(_15324_),
    .A1(\u_inv.f_next[19] ),
    .Y(_15333_),
    .A2(\u_inv.f_reg[19] ));
 sg13g2_o21ai_1 _22297_ (.B1(_15333_),
    .Y(_15334_),
    .A1(_15318_),
    .A2(_15329_));
 sg13g2_nand2_1 _22298_ (.Y(_15335_),
    .A(\u_inv.f_next[23] ),
    .B(\u_inv.f_reg[23] ));
 sg13g2_nor2_1 _22299_ (.A(\u_inv.f_next[23] ),
    .B(\u_inv.f_reg[23] ),
    .Y(_15336_));
 sg13g2_xor2_1 _22300_ (.B(\u_inv.f_reg[23] ),
    .A(\u_inv.f_next[23] ),
    .X(_15337_));
 sg13g2_nand2_1 _22301_ (.Y(_15338_),
    .A(\u_inv.f_next[22] ),
    .B(\u_inv.f_reg[22] ));
 sg13g2_xor2_1 _22302_ (.B(\u_inv.f_reg[22] ),
    .A(\u_inv.f_next[22] ),
    .X(_15339_));
 sg13g2_xnor2_1 _22303_ (.Y(_15340_),
    .A(\u_inv.f_next[22] ),
    .B(\u_inv.f_reg[22] ));
 sg13g2_nand2_1 _22304_ (.Y(_15341_),
    .A(_14153_),
    .B(_14275_));
 sg13g2_nand2_1 _22305_ (.Y(_15342_),
    .A(\u_inv.f_next[21] ),
    .B(\u_inv.f_reg[21] ));
 sg13g2_and2_1 _22306_ (.A(_15341_),
    .B(_15342_),
    .X(_15343_));
 sg13g2_nand2_2 _22307_ (.Y(_15344_),
    .A(_15341_),
    .B(_15342_));
 sg13g2_nor2_1 _22308_ (.A(_14154_),
    .B(_14274_),
    .Y(_15345_));
 sg13g2_xor2_1 _22309_ (.B(\u_inv.f_reg[20] ),
    .A(\u_inv.f_next[20] ),
    .X(_15346_));
 sg13g2_and2_1 _22310_ (.A(_15343_),
    .B(_15346_),
    .X(_15347_));
 sg13g2_and3_1 _22311_ (.X(_15348_),
    .A(_15337_),
    .B(_15339_),
    .C(_15347_));
 sg13g2_o21ai_1 _22312_ (.B1(_15335_),
    .Y(_15349_),
    .A1(_15336_),
    .A2(_15338_));
 sg13g2_nand2_1 _22313_ (.Y(_15350_),
    .A(_15341_),
    .B(_15345_));
 sg13g2_nand2_1 _22314_ (.Y(_15351_),
    .A(_15342_),
    .B(_15350_));
 sg13g2_and3_1 _22315_ (.X(_15352_),
    .A(_15337_),
    .B(_15339_),
    .C(_15351_));
 sg13g2_or2_1 _22316_ (.X(_15353_),
    .B(_15352_),
    .A(_15349_));
 sg13g2_a21o_2 _22317_ (.A2(_15348_),
    .A1(_15334_),
    .B1(_15353_),
    .X(_15354_));
 sg13g2_nand2_1 _22318_ (.Y(_15355_),
    .A(\u_inv.f_next[27] ),
    .B(\u_inv.f_reg[27] ));
 sg13g2_nor2_1 _22319_ (.A(\u_inv.f_next[27] ),
    .B(\u_inv.f_reg[27] ),
    .Y(_15356_));
 sg13g2_xor2_1 _22320_ (.B(\u_inv.f_reg[27] ),
    .A(\u_inv.f_next[27] ),
    .X(_15357_));
 sg13g2_nand2_1 _22321_ (.Y(_15358_),
    .A(\u_inv.f_next[26] ),
    .B(\u_inv.f_reg[26] ));
 sg13g2_xor2_1 _22322_ (.B(\u_inv.f_reg[26] ),
    .A(\u_inv.f_next[26] ),
    .X(_15359_));
 sg13g2_xnor2_1 _22323_ (.Y(_15360_),
    .A(\u_inv.f_next[26] ),
    .B(\u_inv.f_reg[26] ));
 sg13g2_and2_1 _22324_ (.A(_15357_),
    .B(_15359_),
    .X(_15361_));
 sg13g2_nand2_1 _22325_ (.Y(_15362_),
    .A(\u_inv.f_next[24] ),
    .B(\u_inv.f_reg[24] ));
 sg13g2_inv_1 _22326_ (.Y(_15363_),
    .A(_15362_));
 sg13g2_xor2_1 _22327_ (.B(\u_inv.f_reg[24] ),
    .A(\u_inv.f_next[24] ),
    .X(_15364_));
 sg13g2_xor2_1 _22328_ (.B(\u_inv.f_reg[25] ),
    .A(\u_inv.f_next[25] ),
    .X(_15365_));
 sg13g2_and2_1 _22329_ (.A(_15364_),
    .B(_15365_),
    .X(_15366_));
 sg13g2_and2_1 _22330_ (.A(_15361_),
    .B(_15366_),
    .X(_15367_));
 sg13g2_o21ai_1 _22331_ (.B1(_15355_),
    .Y(_15368_),
    .A1(_15356_),
    .A2(_15358_));
 sg13g2_a21oi_1 _22332_ (.A1(\u_inv.f_next[25] ),
    .A2(\u_inv.f_reg[25] ),
    .Y(_15369_),
    .B1(_15363_));
 sg13g2_a21oi_1 _22333_ (.A1(_14149_),
    .A2(_14279_),
    .Y(_15370_),
    .B1(_15369_));
 sg13g2_a221oi_1 _22334_ (.B2(_15361_),
    .C1(_15368_),
    .B1(_15370_),
    .A1(_15354_),
    .Y(_15371_),
    .A2(_15367_));
 sg13g2_xor2_1 _22335_ (.B(\u_inv.f_reg[31] ),
    .A(\u_inv.f_next[31] ),
    .X(_15372_));
 sg13g2_nand2_1 _22336_ (.Y(_15373_),
    .A(\u_inv.f_next[30] ),
    .B(\u_inv.f_reg[30] ));
 sg13g2_xor2_1 _22337_ (.B(\u_inv.f_reg[30] ),
    .A(\u_inv.f_next[30] ),
    .X(_15374_));
 sg13g2_xnor2_1 _22338_ (.Y(_15375_),
    .A(\u_inv.f_next[30] ),
    .B(\u_inv.f_reg[30] ));
 sg13g2_and2_1 _22339_ (.A(_15372_),
    .B(_15374_),
    .X(_15376_));
 sg13g2_nand2_1 _22340_ (.Y(_15377_),
    .A(\u_inv.f_next[28] ),
    .B(\u_inv.f_reg[28] ));
 sg13g2_xor2_1 _22341_ (.B(\u_inv.f_reg[28] ),
    .A(\u_inv.f_next[28] ),
    .X(_15378_));
 sg13g2_xnor2_1 _22342_ (.Y(_15379_),
    .A(\u_inv.f_next[28] ),
    .B(\u_inv.f_reg[28] ));
 sg13g2_xor2_1 _22343_ (.B(\u_inv.f_reg[29] ),
    .A(\u_inv.f_next[29] ),
    .X(_15380_));
 sg13g2_and2_1 _22344_ (.A(_15378_),
    .B(_15380_),
    .X(_15381_));
 sg13g2_nand2_1 _22345_ (.Y(_15382_),
    .A(_15376_),
    .B(_15381_));
 sg13g2_a21oi_1 _22346_ (.A1(_14143_),
    .A2(_14285_),
    .Y(_15383_),
    .B1(_15373_));
 sg13g2_a22oi_1 _22347_ (.Y(_15384_),
    .B1(\u_inv.f_reg[29] ),
    .B2(\u_inv.f_next[29] ),
    .A2(\u_inv.f_reg[28] ),
    .A1(\u_inv.f_next[28] ));
 sg13g2_a21oi_1 _22348_ (.A1(_14145_),
    .A2(_14283_),
    .Y(_15385_),
    .B1(_15384_));
 sg13g2_a221oi_1 _22349_ (.B2(_15385_),
    .C1(_15383_),
    .B1(_15376_),
    .A1(\u_inv.f_next[31] ),
    .Y(_15386_),
    .A2(\u_inv.f_reg[31] ));
 sg13g2_o21ai_1 _22350_ (.B1(_15386_),
    .Y(_15387_),
    .A1(_15371_),
    .A2(_15382_));
 sg13g2_xor2_1 _22351_ (.B(\u_inv.f_reg[33] ),
    .A(\u_inv.f_next[33] ),
    .X(_15388_));
 sg13g2_xnor2_1 _22352_ (.Y(_15389_),
    .A(\u_inv.f_next[33] ),
    .B(\u_inv.f_reg[33] ));
 sg13g2_xor2_1 _22353_ (.B(\u_inv.f_reg[32] ),
    .A(\u_inv.f_next[32] ),
    .X(_15390_));
 sg13g2_and2_1 _22354_ (.A(_15388_),
    .B(_15390_),
    .X(_15391_));
 sg13g2_and4_1 _22355_ (.A(_15230_),
    .B(_15236_),
    .C(_15242_),
    .D(_15391_),
    .X(_15392_));
 sg13g2_a21oi_2 _22356_ (.B1(_15253_),
    .Y(_15393_),
    .A2(_15392_),
    .A1(_15387_));
 sg13g2_a21o_2 _22357_ (.A2(_15392_),
    .A1(_15387_),
    .B1(_15253_),
    .X(_15394_));
 sg13g2_xnor2_1 _22358_ (.Y(_15395_),
    .A(\u_inv.f_next[47] ),
    .B(\u_inv.f_reg[47] ));
 sg13g2_nand2_1 _22359_ (.Y(_15396_),
    .A(\u_inv.f_next[46] ),
    .B(\u_inv.f_reg[46] ));
 sg13g2_xnor2_1 _22360_ (.Y(_15397_),
    .A(\u_inv.f_next[46] ),
    .B(\u_inv.f_reg[46] ));
 sg13g2_nor2_1 _22361_ (.A(_15395_),
    .B(_15397_),
    .Y(_15398_));
 sg13g2_nand2_1 _22362_ (.Y(_15399_),
    .A(\u_inv.f_next[44] ),
    .B(\u_inv.f_reg[44] ));
 sg13g2_nand2_1 _22363_ (.Y(_15400_),
    .A(_14130_),
    .B(_14298_));
 sg13g2_nand2_2 _22364_ (.Y(_15401_),
    .A(_15399_),
    .B(_15400_));
 sg13g2_xor2_1 _22365_ (.B(\u_inv.f_reg[45] ),
    .A(\u_inv.f_next[45] ),
    .X(_15402_));
 sg13g2_nor2b_1 _22366_ (.A(_15401_),
    .B_N(_15402_),
    .Y(_15403_));
 sg13g2_nand2_1 _22367_ (.Y(_15404_),
    .A(_15398_),
    .B(_15403_));
 sg13g2_xnor2_1 _22368_ (.Y(_15405_),
    .A(\u_inv.f_next[43] ),
    .B(\u_inv.f_reg[43] ));
 sg13g2_nand2_1 _22369_ (.Y(_15406_),
    .A(\u_inv.f_next[42] ),
    .B(\u_inv.f_reg[42] ));
 sg13g2_xnor2_1 _22370_ (.Y(_15407_),
    .A(\u_inv.f_next[42] ),
    .B(\u_inv.f_reg[42] ));
 sg13g2_nor2_1 _22371_ (.A(_15405_),
    .B(net5620),
    .Y(_15408_));
 sg13g2_nand2_1 _22372_ (.Y(_15409_),
    .A(\u_inv.f_next[40] ),
    .B(\u_inv.f_reg[40] ));
 sg13g2_xnor2_1 _22373_ (.Y(_15410_),
    .A(\u_inv.f_next[40] ),
    .B(\u_inv.f_reg[40] ));
 sg13g2_xor2_1 _22374_ (.B(\u_inv.f_reg[41] ),
    .A(\u_inv.f_next[41] ),
    .X(_15411_));
 sg13g2_xnor2_1 _22375_ (.Y(_15412_),
    .A(\u_inv.f_next[41] ),
    .B(\u_inv.f_reg[41] ));
 sg13g2_nand2b_1 _22376_ (.Y(_15413_),
    .B(_15411_),
    .A_N(_15410_));
 sg13g2_inv_1 _22377_ (.Y(_15414_),
    .A(_15413_));
 sg13g2_nor4_1 _22378_ (.A(_15404_),
    .B(_15405_),
    .C(net5620),
    .D(_15413_),
    .Y(_15415_));
 sg13g2_a22oi_1 _22379_ (.Y(_15416_),
    .B1(\u_inv.f_reg[41] ),
    .B2(\u_inv.f_next[41] ),
    .A2(\u_inv.f_reg[40] ),
    .A1(\u_inv.f_next[40] ));
 sg13g2_a21oi_1 _22380_ (.A1(_14133_),
    .A2(_14295_),
    .Y(_15417_),
    .B1(_15416_));
 sg13g2_a22oi_1 _22381_ (.Y(_15418_),
    .B1(\u_inv.f_reg[43] ),
    .B2(\u_inv.f_next[43] ),
    .A2(\u_inv.f_reg[42] ),
    .A1(\u_inv.f_next[42] ));
 sg13g2_a21oi_1 _22382_ (.A1(_14131_),
    .A2(_14297_),
    .Y(_15419_),
    .B1(_15418_));
 sg13g2_a21oi_1 _22383_ (.A1(_15408_),
    .A2(_15417_),
    .Y(_15420_),
    .B1(_15419_));
 sg13g2_a21oi_1 _22384_ (.A1(_14127_),
    .A2(_14301_),
    .Y(_15421_),
    .B1(_15396_));
 sg13g2_a22oi_1 _22385_ (.Y(_15422_),
    .B1(\u_inv.f_reg[45] ),
    .B2(\u_inv.f_next[45] ),
    .A2(\u_inv.f_reg[44] ),
    .A1(\u_inv.f_next[44] ));
 sg13g2_a21oi_1 _22386_ (.A1(_14129_),
    .A2(_14299_),
    .Y(_15423_),
    .B1(_15422_));
 sg13g2_a221oi_1 _22387_ (.B2(_15423_),
    .C1(_15421_),
    .B1(_15398_),
    .A1(\u_inv.f_next[47] ),
    .Y(_15424_),
    .A2(\u_inv.f_reg[47] ));
 sg13g2_o21ai_1 _22388_ (.B1(_15424_),
    .Y(_15425_),
    .A1(_15404_),
    .A2(_15420_));
 sg13g2_a21oi_2 _22389_ (.B1(_15425_),
    .Y(_15426_),
    .A2(_15415_),
    .A1(_15394_));
 sg13g2_nor2_1 _22390_ (.A(\u_inv.f_next[55] ),
    .B(\u_inv.f_reg[55] ),
    .Y(_15427_));
 sg13g2_xor2_1 _22391_ (.B(\u_inv.f_reg[55] ),
    .A(\u_inv.f_next[55] ),
    .X(_15428_));
 sg13g2_xnor2_1 _22392_ (.Y(_15429_),
    .A(\u_inv.f_next[55] ),
    .B(\u_inv.f_reg[55] ));
 sg13g2_nand2_1 _22393_ (.Y(_15430_),
    .A(\u_inv.f_next[54] ),
    .B(\u_inv.f_reg[54] ));
 sg13g2_xor2_1 _22394_ (.B(\u_inv.f_reg[54] ),
    .A(\u_inv.f_next[54] ),
    .X(_15431_));
 sg13g2_xnor2_1 _22395_ (.Y(_15432_),
    .A(\u_inv.f_next[54] ),
    .B(\u_inv.f_reg[54] ));
 sg13g2_nor2_1 _22396_ (.A(_15429_),
    .B(_15432_),
    .Y(_15433_));
 sg13g2_xnor2_1 _22397_ (.Y(_15434_),
    .A(\u_inv.f_next[53] ),
    .B(\u_inv.f_reg[53] ));
 sg13g2_nand2_1 _22398_ (.Y(_15435_),
    .A(\u_inv.f_next[52] ),
    .B(\u_inv.f_reg[52] ));
 sg13g2_xnor2_1 _22399_ (.Y(_15436_),
    .A(\u_inv.f_next[52] ),
    .B(\u_inv.f_reg[52] ));
 sg13g2_nor4_1 _22400_ (.A(_15429_),
    .B(_15432_),
    .C(_15434_),
    .D(_15436_),
    .Y(_15437_));
 sg13g2_nor2_1 _22401_ (.A(_14124_),
    .B(_14304_),
    .Y(_15438_));
 sg13g2_xnor2_1 _22402_ (.Y(_15439_),
    .A(\u_inv.f_next[50] ),
    .B(\u_inv.f_reg[50] ));
 sg13g2_xnor2_1 _22403_ (.Y(_15440_),
    .A(\u_inv.f_next[51] ),
    .B(\u_inv.f_reg[51] ));
 sg13g2_nor2_1 _22404_ (.A(_15439_),
    .B(_15440_),
    .Y(_15441_));
 sg13g2_xnor2_1 _22405_ (.Y(_15442_),
    .A(\u_inv.f_next[49] ),
    .B(\u_inv.f_reg[49] ));
 sg13g2_nand2_1 _22406_ (.Y(_15443_),
    .A(\u_inv.f_next[48] ),
    .B(\u_inv.f_reg[48] ));
 sg13g2_xnor2_1 _22407_ (.Y(_15444_),
    .A(\u_inv.f_next[48] ),
    .B(\u_inv.f_reg[48] ));
 sg13g2_nor2_1 _22408_ (.A(_15442_),
    .B(_15444_),
    .Y(_15445_));
 sg13g2_or2_1 _22409_ (.X(_15446_),
    .B(_15444_),
    .A(_15442_));
 sg13g2_nand3_1 _22410_ (.B(_15441_),
    .C(_15445_),
    .A(_15437_),
    .Y(_15447_));
 sg13g2_a22oi_1 _22411_ (.Y(_15448_),
    .B1(\u_inv.f_reg[55] ),
    .B2(\u_inv.f_next[55] ),
    .A2(\u_inv.f_reg[54] ),
    .A1(\u_inv.f_next[54] ));
 sg13g2_a22oi_1 _22412_ (.Y(_15449_),
    .B1(\u_inv.f_reg[53] ),
    .B2(\u_inv.f_next[53] ),
    .A2(\u_inv.f_reg[52] ),
    .A1(\u_inv.f_next[52] ));
 sg13g2_a21oi_1 _22413_ (.A1(_14121_),
    .A2(_14307_),
    .Y(_15450_),
    .B1(_15449_));
 sg13g2_a22oi_1 _22414_ (.Y(_15451_),
    .B1(\u_inv.f_reg[49] ),
    .B2(\u_inv.f_next[49] ),
    .A2(\u_inv.f_reg[48] ),
    .A1(\u_inv.f_next[48] ));
 sg13g2_a21o_1 _22415_ (.A2(_14303_),
    .A1(_14125_),
    .B1(_15451_),
    .X(_15452_));
 sg13g2_nor3_1 _22416_ (.A(_15439_),
    .B(_15440_),
    .C(_15452_),
    .Y(_15453_));
 sg13g2_a21oi_1 _22417_ (.A1(\u_inv.f_next[51] ),
    .A2(\u_inv.f_reg[51] ),
    .Y(_15454_),
    .B1(_15438_));
 sg13g2_a21oi_1 _22418_ (.A1(_14123_),
    .A2(_14305_),
    .Y(_15455_),
    .B1(_15454_));
 sg13g2_o21ai_1 _22419_ (.B1(_15437_),
    .Y(_15456_),
    .A1(_15453_),
    .A2(_15455_));
 sg13g2_o21ai_1 _22420_ (.B1(_15456_),
    .Y(_15457_),
    .A1(_15427_),
    .A2(_15448_));
 sg13g2_a21oi_1 _22421_ (.A1(_15433_),
    .A2(_15450_),
    .Y(_15458_),
    .B1(_15457_));
 sg13g2_o21ai_1 _22422_ (.B1(_15458_),
    .Y(_15459_),
    .A1(_15426_),
    .A2(_15447_));
 sg13g2_xnor2_1 _22423_ (.Y(_15460_),
    .A(\u_inv.f_next[57] ),
    .B(\u_inv.f_reg[57] ));
 sg13g2_xor2_1 _22424_ (.B(\u_inv.f_reg[56] ),
    .A(\u_inv.f_next[56] ),
    .X(_15461_));
 sg13g2_inv_2 _22425_ (.Y(_15462_),
    .A(_15461_));
 sg13g2_nor2_1 _22426_ (.A(_15460_),
    .B(_15462_),
    .Y(_15463_));
 sg13g2_nor4_1 _22427_ (.A(_15207_),
    .B(_15212_),
    .C(_15460_),
    .D(_15462_),
    .Y(_15464_));
 sg13g2_a21oi_2 _22428_ (.B1(_15225_),
    .Y(_15465_),
    .A2(_15464_),
    .A1(_15459_));
 sg13g2_a21o_2 _22429_ (.A2(_15464_),
    .A1(_15459_),
    .B1(_15225_),
    .X(_15466_));
 sg13g2_xor2_1 _22430_ (.B(\u_inv.f_reg[64] ),
    .A(\u_inv.f_next[64] ),
    .X(_15467_));
 sg13g2_xnor2_1 _22431_ (.Y(_15468_),
    .A(\u_inv.f_next[64] ),
    .B(\u_inv.f_reg[64] ));
 sg13g2_nor2b_2 _22432_ (.A(_15184_),
    .B_N(_15185_),
    .Y(_15469_));
 sg13g2_and2_1 _22433_ (.A(_15467_),
    .B(_15469_),
    .X(_15470_));
 sg13g2_nand4_1 _22434_ (.B(_15178_),
    .C(_15182_),
    .A(_15173_),
    .Y(_15471_),
    .D(_15470_));
 sg13g2_nor2_1 _22435_ (.A(_15465_),
    .B(_15471_),
    .Y(_15472_));
 sg13g2_nor2b_1 _22436_ (.A(_15472_),
    .B_N(_15197_),
    .Y(_15473_));
 sg13g2_o21ai_1 _22437_ (.B1(_15197_),
    .Y(_15474_),
    .A1(_15465_),
    .A2(_15471_));
 sg13g2_xor2_1 _22438_ (.B(\u_inv.f_reg[79] ),
    .A(\u_inv.f_next[79] ),
    .X(_15475_));
 sg13g2_nand2_1 _22439_ (.Y(_15476_),
    .A(\u_inv.f_next[78] ),
    .B(\u_inv.f_reg[78] ));
 sg13g2_nor2_1 _22440_ (.A(\u_inv.f_next[78] ),
    .B(\u_inv.f_reg[78] ),
    .Y(_15477_));
 sg13g2_xor2_1 _22441_ (.B(\u_inv.f_reg[78] ),
    .A(\u_inv.f_next[78] ),
    .X(_15478_));
 sg13g2_and2_1 _22442_ (.A(_15475_),
    .B(_15478_),
    .X(_15479_));
 sg13g2_xnor2_1 _22443_ (.Y(_15480_),
    .A(\u_inv.f_next[77] ),
    .B(\u_inv.f_reg[77] ));
 sg13g2_nand2_1 _22444_ (.Y(_15481_),
    .A(\u_inv.f_next[76] ),
    .B(\u_inv.f_reg[76] ));
 sg13g2_xor2_1 _22445_ (.B(\u_inv.f_reg[76] ),
    .A(\u_inv.f_next[76] ),
    .X(_15482_));
 sg13g2_xnor2_1 _22446_ (.Y(_15483_),
    .A(\u_inv.f_next[76] ),
    .B(\u_inv.f_reg[76] ));
 sg13g2_nor2_1 _22447_ (.A(_15480_),
    .B(_15483_),
    .Y(_15484_));
 sg13g2_nand2_1 _22448_ (.Y(_15485_),
    .A(_15479_),
    .B(_15484_));
 sg13g2_xor2_1 _22449_ (.B(\u_inv.f_reg[75] ),
    .A(\u_inv.f_next[75] ),
    .X(_15486_));
 sg13g2_nand2_1 _22450_ (.Y(_15487_),
    .A(\u_inv.f_next[74] ),
    .B(\u_inv.f_reg[74] ));
 sg13g2_xor2_1 _22451_ (.B(\u_inv.f_reg[74] ),
    .A(\u_inv.f_next[74] ),
    .X(_15488_));
 sg13g2_xnor2_1 _22452_ (.Y(_15489_),
    .A(\u_inv.f_next[74] ),
    .B(\u_inv.f_reg[74] ));
 sg13g2_and2_1 _22453_ (.A(_15486_),
    .B(_15488_),
    .X(_15490_));
 sg13g2_nand2_1 _22454_ (.Y(_15491_),
    .A(_15486_),
    .B(_15488_));
 sg13g2_nand2_1 _22455_ (.Y(_15492_),
    .A(\u_inv.f_next[72] ),
    .B(\u_inv.f_reg[72] ));
 sg13g2_xor2_1 _22456_ (.B(\u_inv.f_reg[72] ),
    .A(\u_inv.f_next[72] ),
    .X(_15493_));
 sg13g2_xnor2_1 _22457_ (.Y(_15494_),
    .A(\u_inv.f_next[72] ),
    .B(\u_inv.f_reg[72] ));
 sg13g2_xor2_1 _22458_ (.B(\u_inv.f_reg[73] ),
    .A(\u_inv.f_next[73] ),
    .X(_15495_));
 sg13g2_xnor2_1 _22459_ (.Y(_15496_),
    .A(\u_inv.f_next[73] ),
    .B(\u_inv.f_reg[73] ));
 sg13g2_nor2_1 _22460_ (.A(_15494_),
    .B(_15496_),
    .Y(_15497_));
 sg13g2_nor4_1 _22461_ (.A(_15485_),
    .B(_15491_),
    .C(_15494_),
    .D(_15496_),
    .Y(_15498_));
 sg13g2_a22oi_1 _22462_ (.Y(_15499_),
    .B1(\u_inv.f_reg[73] ),
    .B2(\u_inv.f_next[73] ),
    .A2(\u_inv.f_reg[72] ),
    .A1(\u_inv.f_next[72] ));
 sg13g2_a21oi_1 _22463_ (.A1(_14101_),
    .A2(_14327_),
    .Y(_15500_),
    .B1(_15499_));
 sg13g2_a22oi_1 _22464_ (.Y(_15501_),
    .B1(\u_inv.f_reg[75] ),
    .B2(\u_inv.f_next[75] ),
    .A2(\u_inv.f_reg[74] ),
    .A1(\u_inv.f_next[74] ));
 sg13g2_a21oi_1 _22465_ (.A1(_14099_),
    .A2(_14329_),
    .Y(_15502_),
    .B1(_15501_));
 sg13g2_a21oi_1 _22466_ (.A1(_15490_),
    .A2(_15500_),
    .Y(_15503_),
    .B1(_15502_));
 sg13g2_a21oi_1 _22467_ (.A1(_14095_),
    .A2(_14333_),
    .Y(_15504_),
    .B1(_15476_));
 sg13g2_a22oi_1 _22468_ (.Y(_15505_),
    .B1(\u_inv.f_reg[77] ),
    .B2(\u_inv.f_next[77] ),
    .A2(\u_inv.f_reg[76] ),
    .A1(\u_inv.f_next[76] ));
 sg13g2_a21oi_1 _22469_ (.A1(_14097_),
    .A2(_14331_),
    .Y(_15506_),
    .B1(_15505_));
 sg13g2_a221oi_1 _22470_ (.B2(_15506_),
    .C1(_15504_),
    .B1(_15479_),
    .A1(\u_inv.f_next[79] ),
    .Y(_15507_),
    .A2(\u_inv.f_reg[79] ));
 sg13g2_o21ai_1 _22471_ (.B1(_15507_),
    .Y(_15508_),
    .A1(_15485_),
    .A2(_15503_));
 sg13g2_a21oi_2 _22472_ (.B1(_15508_),
    .Y(_15509_),
    .A2(_15498_),
    .A1(_15474_));
 sg13g2_xor2_1 _22473_ (.B(\u_inv.f_reg[83] ),
    .A(\u_inv.f_next[83] ),
    .X(_15510_));
 sg13g2_xnor2_1 _22474_ (.Y(_15511_),
    .A(\u_inv.f_next[83] ),
    .B(\u_inv.f_reg[83] ));
 sg13g2_nor2_1 _22475_ (.A(_14092_),
    .B(_14336_),
    .Y(_15512_));
 sg13g2_xor2_1 _22476_ (.B(\u_inv.f_reg[82] ),
    .A(\u_inv.f_next[82] ),
    .X(_15513_));
 sg13g2_and2_1 _22477_ (.A(_15510_),
    .B(_15513_),
    .X(_15514_));
 sg13g2_nand2_1 _22478_ (.Y(_15515_),
    .A(\u_inv.f_next[80] ),
    .B(\u_inv.f_reg[80] ));
 sg13g2_xor2_1 _22479_ (.B(\u_inv.f_reg[80] ),
    .A(\u_inv.f_next[80] ),
    .X(_15516_));
 sg13g2_xnor2_1 _22480_ (.Y(_15517_),
    .A(\u_inv.f_next[80] ),
    .B(\u_inv.f_reg[80] ));
 sg13g2_xor2_1 _22481_ (.B(\u_inv.f_reg[81] ),
    .A(\u_inv.f_next[81] ),
    .X(_15518_));
 sg13g2_xnor2_1 _22482_ (.Y(_15519_),
    .A(\u_inv.f_next[81] ),
    .B(\u_inv.f_reg[81] ));
 sg13g2_nand3_1 _22483_ (.B(_15516_),
    .C(_15518_),
    .A(_15514_),
    .Y(_15520_));
 sg13g2_a22oi_1 _22484_ (.Y(_15521_),
    .B1(\u_inv.f_reg[81] ),
    .B2(\u_inv.f_next[81] ),
    .A2(\u_inv.f_reg[80] ),
    .A1(\u_inv.f_next[80] ));
 sg13g2_a21oi_1 _22485_ (.A1(_14093_),
    .A2(_14335_),
    .Y(_15522_),
    .B1(_15521_));
 sg13g2_o21ai_1 _22486_ (.B1(_15512_),
    .Y(_15523_),
    .A1(\u_inv.f_next[83] ),
    .A2(\u_inv.f_reg[83] ));
 sg13g2_inv_1 _22487_ (.Y(_15524_),
    .A(_15523_));
 sg13g2_a221oi_1 _22488_ (.B2(_15522_),
    .C1(_15524_),
    .B1(_15514_),
    .A1(\u_inv.f_next[83] ),
    .Y(_15525_),
    .A2(\u_inv.f_reg[83] ));
 sg13g2_and2_1 _22489_ (.A(_15161_),
    .B(_15525_),
    .X(_15526_));
 sg13g2_o21ai_1 _22490_ (.B1(_15526_),
    .Y(_15527_),
    .A1(_15509_),
    .A2(_15520_));
 sg13g2_nand2_1 _22491_ (.Y(_15528_),
    .A(_15168_),
    .B(_15527_));
 sg13g2_nand2_1 _22492_ (.Y(_15529_),
    .A(\u_inv.f_next[95] ),
    .B(\u_inv.f_reg[95] ));
 sg13g2_xnor2_1 _22493_ (.Y(_15530_),
    .A(\u_inv.f_next[95] ),
    .B(\u_inv.f_reg[95] ));
 sg13g2_nor2_1 _22494_ (.A(_14080_),
    .B(_14348_),
    .Y(_15531_));
 sg13g2_xnor2_1 _22495_ (.Y(_15532_),
    .A(\u_inv.f_next[94] ),
    .B(\u_inv.f_reg[94] ));
 sg13g2_xor2_1 _22496_ (.B(\u_inv.f_reg[92] ),
    .A(\u_inv.f_next[92] ),
    .X(_15533_));
 sg13g2_xor2_1 _22497_ (.B(\u_inv.f_reg[93] ),
    .A(\u_inv.f_next[93] ),
    .X(_15534_));
 sg13g2_xnor2_1 _22498_ (.Y(_15535_),
    .A(\u_inv.f_next[93] ),
    .B(\u_inv.f_reg[93] ));
 sg13g2_nand2_1 _22499_ (.Y(_15536_),
    .A(_15533_),
    .B(_15534_));
 sg13g2_nor3_1 _22500_ (.A(_15530_),
    .B(_15532_),
    .C(_15536_),
    .Y(_15537_));
 sg13g2_xnor2_1 _22501_ (.Y(_15538_),
    .A(\u_inv.f_next[91] ),
    .B(\u_inv.f_reg[91] ));
 sg13g2_xnor2_1 _22502_ (.Y(_15539_),
    .A(\u_inv.f_next[90] ),
    .B(\u_inv.f_reg[90] ));
 sg13g2_nor2_1 _22503_ (.A(_15538_),
    .B(_15539_),
    .Y(_15540_));
 sg13g2_inv_1 _22504_ (.Y(_15541_),
    .A(_15540_));
 sg13g2_and2_1 _22505_ (.A(_15537_),
    .B(_15540_),
    .X(_15542_));
 sg13g2_nor2_1 _22506_ (.A(\u_inv.f_next[89] ),
    .B(\u_inv.f_reg[89] ),
    .Y(_15543_));
 sg13g2_nand2_1 _22507_ (.Y(_15544_),
    .A(\u_inv.f_next[89] ),
    .B(\u_inv.f_reg[89] ));
 sg13g2_nor2b_2 _22508_ (.A(_15543_),
    .B_N(_15544_),
    .Y(_15545_));
 sg13g2_nand2_1 _22509_ (.Y(_15546_),
    .A(\u_inv.f_next[88] ),
    .B(\u_inv.f_reg[88] ));
 sg13g2_xor2_1 _22510_ (.B(\u_inv.f_reg[88] ),
    .A(\u_inv.f_next[88] ),
    .X(_15547_));
 sg13g2_xnor2_1 _22511_ (.Y(_15548_),
    .A(\u_inv.f_next[88] ),
    .B(\u_inv.f_reg[88] ));
 sg13g2_and2_1 _22512_ (.A(_15545_),
    .B(_15547_),
    .X(_15549_));
 sg13g2_nand4_1 _22513_ (.B(_15527_),
    .C(_15542_),
    .A(_15168_),
    .Y(_15550_),
    .D(_15549_));
 sg13g2_nand2_1 _22514_ (.Y(_15551_),
    .A(_15544_),
    .B(_15546_));
 sg13g2_o21ai_1 _22515_ (.B1(_15544_),
    .Y(_15552_),
    .A1(_15543_),
    .A2(_15546_));
 sg13g2_nand2b_1 _22516_ (.Y(_15553_),
    .B(_15551_),
    .A_N(_15543_));
 sg13g2_a22oi_1 _22517_ (.Y(_15554_),
    .B1(\u_inv.f_reg[93] ),
    .B2(\u_inv.f_next[93] ),
    .A2(\u_inv.f_reg[92] ),
    .A1(\u_inv.f_next[92] ));
 sg13g2_a21o_1 _22518_ (.A2(_14347_),
    .A1(_14081_),
    .B1(_15554_),
    .X(_15555_));
 sg13g2_or3_1 _22519_ (.A(_15530_),
    .B(_15532_),
    .C(_15555_),
    .X(_15556_));
 sg13g2_o21ai_1 _22520_ (.B1(_15531_),
    .Y(_15557_),
    .A1(\u_inv.f_next[95] ),
    .A2(\u_inv.f_reg[95] ));
 sg13g2_nand3_1 _22521_ (.B(_15556_),
    .C(_15557_),
    .A(_15529_),
    .Y(_15558_));
 sg13g2_a22oi_1 _22522_ (.Y(_15559_),
    .B1(\u_inv.f_reg[91] ),
    .B2(\u_inv.f_next[91] ),
    .A2(\u_inv.f_reg[90] ),
    .A1(\u_inv.f_next[90] ));
 sg13g2_a21oi_1 _22523_ (.A1(_14083_),
    .A2(_14345_),
    .Y(_15560_),
    .B1(_15559_));
 sg13g2_a221oi_1 _22524_ (.B2(_15537_),
    .C1(_15558_),
    .B1(_15560_),
    .A1(_15542_),
    .Y(_15561_),
    .A2(_15552_));
 sg13g2_nand2_1 _22525_ (.Y(_15562_),
    .A(_15550_),
    .B(_15561_));
 sg13g2_xor2_1 _22526_ (.B(\u_inv.f_reg[97] ),
    .A(\u_inv.f_next[97] ),
    .X(_15563_));
 sg13g2_xor2_1 _22527_ (.B(\u_inv.f_reg[96] ),
    .A(\u_inv.f_next[96] ),
    .X(_15564_));
 sg13g2_xnor2_1 _22528_ (.Y(_15565_),
    .A(\u_inv.f_next[96] ),
    .B(\u_inv.f_reg[96] ));
 sg13g2_and2_1 _22529_ (.A(_15563_),
    .B(_15564_),
    .X(_15566_));
 sg13g2_nor2b_1 _22530_ (.A(_15126_),
    .B_N(_15566_),
    .Y(_15567_));
 sg13g2_nand4_1 _22531_ (.B(_15133_),
    .C(_15135_),
    .A(_15131_),
    .Y(_15568_),
    .D(_15567_));
 sg13g2_a21o_2 _22532_ (.A2(_15561_),
    .A1(_15550_),
    .B1(_15568_),
    .X(_15569_));
 sg13g2_nand2_2 _22533_ (.Y(_15570_),
    .A(_15149_),
    .B(_15569_));
 sg13g2_xor2_1 _22534_ (.B(\u_inv.f_reg[111] ),
    .A(\u_inv.f_next[111] ),
    .X(_15571_));
 sg13g2_xnor2_1 _22535_ (.Y(_15572_),
    .A(\u_inv.f_next[111] ),
    .B(\u_inv.f_reg[111] ));
 sg13g2_nand2_1 _22536_ (.Y(_15573_),
    .A(\u_inv.f_next[110] ),
    .B(\u_inv.f_reg[110] ));
 sg13g2_nor2_1 _22537_ (.A(\u_inv.f_next[110] ),
    .B(\u_inv.f_reg[110] ),
    .Y(_15574_));
 sg13g2_xor2_1 _22538_ (.B(\u_inv.f_reg[110] ),
    .A(\u_inv.f_next[110] ),
    .X(_15575_));
 sg13g2_and2_1 _22539_ (.A(_15571_),
    .B(_15575_),
    .X(_15576_));
 sg13g2_xor2_1 _22540_ (.B(\u_inv.f_reg[109] ),
    .A(\u_inv.f_next[109] ),
    .X(_15577_));
 sg13g2_xnor2_1 _22541_ (.Y(_15578_),
    .A(\u_inv.f_next[109] ),
    .B(\u_inv.f_reg[109] ));
 sg13g2_nor2_1 _22542_ (.A(_14066_),
    .B(_14362_),
    .Y(_15579_));
 sg13g2_nand2_1 _22543_ (.Y(_15580_),
    .A(_14066_),
    .B(_14362_));
 sg13g2_nand2b_2 _22544_ (.Y(_15581_),
    .B(_15580_),
    .A_N(_15579_));
 sg13g2_nor2_1 _22545_ (.A(_15578_),
    .B(_15581_),
    .Y(_15582_));
 sg13g2_and2_1 _22546_ (.A(_15576_),
    .B(_15582_),
    .X(_15583_));
 sg13g2_xor2_1 _22547_ (.B(\u_inv.f_reg[107] ),
    .A(\u_inv.f_next[107] ),
    .X(_15584_));
 sg13g2_xnor2_1 _22548_ (.Y(_15585_),
    .A(\u_inv.f_next[107] ),
    .B(\u_inv.f_reg[107] ));
 sg13g2_nand2_1 _22549_ (.Y(_15586_),
    .A(\u_inv.f_next[106] ),
    .B(\u_inv.f_reg[106] ));
 sg13g2_xor2_1 _22550_ (.B(\u_inv.f_reg[106] ),
    .A(\u_inv.f_next[106] ),
    .X(_15587_));
 sg13g2_xnor2_1 _22551_ (.Y(_15588_),
    .A(\u_inv.f_next[106] ),
    .B(\u_inv.f_reg[106] ));
 sg13g2_nand2_1 _22552_ (.Y(_15589_),
    .A(_15584_),
    .B(_15587_));
 sg13g2_nor2_1 _22553_ (.A(_14070_),
    .B(_14358_),
    .Y(_15590_));
 sg13g2_xor2_1 _22554_ (.B(\u_inv.f_reg[104] ),
    .A(\u_inv.f_next[104] ),
    .X(_15591_));
 sg13g2_xor2_1 _22555_ (.B(\u_inv.f_reg[105] ),
    .A(\u_inv.f_next[105] ),
    .X(_15592_));
 sg13g2_and2_1 _22556_ (.A(_15591_),
    .B(_15592_),
    .X(_15593_));
 sg13g2_nand4_1 _22557_ (.B(_15584_),
    .C(_15587_),
    .A(_15583_),
    .Y(_15594_),
    .D(_15593_));
 sg13g2_a21oi_2 _22558_ (.B1(_15594_),
    .Y(_15595_),
    .A2(_15569_),
    .A1(_15149_));
 sg13g2_a21o_2 _22559_ (.A2(_15569_),
    .A1(_15149_),
    .B1(_15594_),
    .X(_15596_));
 sg13g2_a21oi_1 _22560_ (.A1(\u_inv.f_next[105] ),
    .A2(\u_inv.f_reg[105] ),
    .Y(_15597_),
    .B1(_15590_));
 sg13g2_a21o_1 _22561_ (.A2(_14359_),
    .A1(_14069_),
    .B1(_15597_),
    .X(_15598_));
 sg13g2_inv_1 _22562_ (.Y(_15599_),
    .A(_15598_));
 sg13g2_a22oi_1 _22563_ (.Y(_15600_),
    .B1(\u_inv.f_reg[107] ),
    .B2(\u_inv.f_next[107] ),
    .A2(\u_inv.f_reg[106] ),
    .A1(\u_inv.f_next[106] ));
 sg13g2_a21o_1 _22564_ (.A2(_14361_),
    .A1(_14067_),
    .B1(_15600_),
    .X(_15601_));
 sg13g2_o21ai_1 _22565_ (.B1(_15601_),
    .Y(_15602_),
    .A1(_15589_),
    .A2(_15598_));
 sg13g2_a21oi_1 _22566_ (.A1(_14063_),
    .A2(_14365_),
    .Y(_15603_),
    .B1(_15573_));
 sg13g2_a21oi_1 _22567_ (.A1(\u_inv.f_next[111] ),
    .A2(\u_inv.f_reg[111] ),
    .Y(_15604_),
    .B1(_15603_));
 sg13g2_a21oi_1 _22568_ (.A1(\u_inv.f_next[109] ),
    .A2(\u_inv.f_reg[109] ),
    .Y(_15605_),
    .B1(_15579_));
 sg13g2_a21oi_1 _22569_ (.A1(_14065_),
    .A2(_14363_),
    .Y(_15606_),
    .B1(_15605_));
 sg13g2_a22oi_1 _22570_ (.Y(_15607_),
    .B1(_15606_),
    .B2(_15576_),
    .A2(_15602_),
    .A1(_15583_));
 sg13g2_nand2_2 _22571_ (.Y(_15608_),
    .A(_15604_),
    .B(_15607_));
 sg13g2_inv_2 _22572_ (.Y(_15609_),
    .A(_15608_));
 sg13g2_nor2_1 _22573_ (.A(_15595_),
    .B(_15608_),
    .Y(_15610_));
 sg13g2_xor2_1 _22574_ (.B(\u_inv.f_reg[127] ),
    .A(\u_inv.f_next[127] ),
    .X(_15611_));
 sg13g2_nand2_1 _22575_ (.Y(_15612_),
    .A(\u_inv.f_next[126] ),
    .B(\u_inv.f_reg[126] ));
 sg13g2_xnor2_1 _22576_ (.Y(_15613_),
    .A(\u_inv.f_next[126] ),
    .B(\u_inv.f_reg[126] ));
 sg13g2_inv_1 _22577_ (.Y(_15614_),
    .A(_15613_));
 sg13g2_and2_1 _22578_ (.A(_15611_),
    .B(_15614_),
    .X(_15615_));
 sg13g2_xor2_1 _22579_ (.B(\u_inv.f_reg[125] ),
    .A(\u_inv.f_next[125] ),
    .X(_15616_));
 sg13g2_nand2_1 _22580_ (.Y(_15617_),
    .A(\u_inv.f_next[124] ),
    .B(\u_inv.f_reg[124] ));
 sg13g2_xor2_1 _22581_ (.B(\u_inv.f_reg[124] ),
    .A(\u_inv.f_next[124] ),
    .X(_15618_));
 sg13g2_xnor2_1 _22582_ (.Y(_15619_),
    .A(\u_inv.f_next[124] ),
    .B(\u_inv.f_reg[124] ));
 sg13g2_nand3_1 _22583_ (.B(_15616_),
    .C(_15618_),
    .A(_15615_),
    .Y(_15620_));
 sg13g2_nor2_1 _22584_ (.A(\u_inv.f_next[123] ),
    .B(\u_inv.f_reg[123] ),
    .Y(_15621_));
 sg13g2_xnor2_1 _22585_ (.Y(_15622_),
    .A(\u_inv.f_next[123] ),
    .B(\u_inv.f_reg[123] ));
 sg13g2_nand2_1 _22586_ (.Y(_15623_),
    .A(\u_inv.f_next[122] ),
    .B(\u_inv.f_reg[122] ));
 sg13g2_xnor2_1 _22587_ (.Y(_15624_),
    .A(\u_inv.f_next[122] ),
    .B(\u_inv.f_reg[122] ));
 sg13g2_nor2_1 _22588_ (.A(_15622_),
    .B(_15624_),
    .Y(_15625_));
 sg13g2_nand2_1 _22589_ (.Y(_15626_),
    .A(\u_inv.f_next[120] ),
    .B(\u_inv.f_reg[120] ));
 sg13g2_xnor2_1 _22590_ (.Y(_15627_),
    .A(\u_inv.f_next[120] ),
    .B(\u_inv.f_reg[120] ));
 sg13g2_xor2_1 _22591_ (.B(\u_inv.f_reg[121] ),
    .A(\u_inv.f_next[121] ),
    .X(_15628_));
 sg13g2_nand2b_1 _22592_ (.Y(_15629_),
    .B(_15628_),
    .A_N(_15627_));
 sg13g2_nor4_2 _22593_ (.A(_15620_),
    .B(_15622_),
    .C(_15624_),
    .Y(_15630_),
    .D(_15629_));
 sg13g2_xnor2_1 _22594_ (.Y(_15631_),
    .A(\u_inv.f_next[119] ),
    .B(\u_inv.f_reg[119] ));
 sg13g2_nand2_1 _22595_ (.Y(_15632_),
    .A(\u_inv.f_next[118] ),
    .B(\u_inv.f_reg[118] ));
 sg13g2_xnor2_1 _22596_ (.Y(_15633_),
    .A(\u_inv.f_next[118] ),
    .B(\u_inv.f_reg[118] ));
 sg13g2_nor2_1 _22597_ (.A(_15631_),
    .B(_15633_),
    .Y(_15634_));
 sg13g2_nand2_1 _22598_ (.Y(_15635_),
    .A(\u_inv.f_next[116] ),
    .B(\u_inv.f_reg[116] ));
 sg13g2_xnor2_1 _22599_ (.Y(_15636_),
    .A(\u_inv.f_next[116] ),
    .B(\u_inv.f_reg[116] ));
 sg13g2_xor2_1 _22600_ (.B(\u_inv.f_reg[117] ),
    .A(\u_inv.f_next[117] ),
    .X(_15637_));
 sg13g2_xnor2_1 _22601_ (.Y(_15638_),
    .A(\u_inv.f_next[117] ),
    .B(\u_inv.f_reg[117] ));
 sg13g2_nor2_1 _22602_ (.A(_15636_),
    .B(_15638_),
    .Y(_15639_));
 sg13g2_nand2_1 _22603_ (.Y(_15640_),
    .A(_15634_),
    .B(_15639_));
 sg13g2_xor2_1 _22604_ (.B(\u_inv.f_reg[115] ),
    .A(\u_inv.f_next[115] ),
    .X(_15641_));
 sg13g2_xnor2_1 _22605_ (.Y(_15642_),
    .A(\u_inv.f_next[115] ),
    .B(\u_inv.f_reg[115] ));
 sg13g2_nand2_1 _22606_ (.Y(_15643_),
    .A(\u_inv.f_next[114] ),
    .B(\u_inv.f_reg[114] ));
 sg13g2_xor2_1 _22607_ (.B(\u_inv.f_reg[114] ),
    .A(\u_inv.f_next[114] ),
    .X(_15644_));
 sg13g2_xnor2_1 _22608_ (.Y(_15645_),
    .A(\u_inv.f_next[114] ),
    .B(\u_inv.f_reg[114] ));
 sg13g2_nand2_1 _22609_ (.Y(_15646_),
    .A(_15641_),
    .B(_15644_));
 sg13g2_inv_1 _22610_ (.Y(_15647_),
    .A(_15646_));
 sg13g2_nand2_1 _22611_ (.Y(_15648_),
    .A(\u_inv.f_next[112] ),
    .B(\u_inv.f_reg[112] ));
 sg13g2_xor2_1 _22612_ (.B(\u_inv.f_reg[112] ),
    .A(\u_inv.f_next[112] ),
    .X(_15649_));
 sg13g2_xnor2_1 _22613_ (.Y(_15650_),
    .A(\u_inv.f_next[112] ),
    .B(\u_inv.f_reg[112] ));
 sg13g2_xor2_1 _22614_ (.B(\u_inv.f_reg[113] ),
    .A(\u_inv.f_next[113] ),
    .X(_15651_));
 sg13g2_xnor2_1 _22615_ (.Y(_15652_),
    .A(\u_inv.f_next[113] ),
    .B(\u_inv.f_reg[113] ));
 sg13g2_nor4_1 _22616_ (.A(_15640_),
    .B(_15646_),
    .C(_15650_),
    .D(_15652_),
    .Y(_15653_));
 sg13g2_nand2_1 _22617_ (.Y(_15654_),
    .A(_15630_),
    .B(_15653_));
 sg13g2_a21oi_2 _22618_ (.B1(_15654_),
    .Y(_15655_),
    .A2(_15609_),
    .A1(_15596_));
 sg13g2_a21o_2 _22619_ (.A2(_15609_),
    .A1(_15596_),
    .B1(_15654_),
    .X(_15656_));
 sg13g2_a22oi_1 _22620_ (.Y(_15657_),
    .B1(\u_inv.f_reg[113] ),
    .B2(\u_inv.f_next[113] ),
    .A2(\u_inv.f_reg[112] ),
    .A1(\u_inv.f_next[112] ));
 sg13g2_a21o_1 _22621_ (.A2(_14367_),
    .A1(_14061_),
    .B1(_15657_),
    .X(_15658_));
 sg13g2_inv_1 _22622_ (.Y(_15659_),
    .A(_15658_));
 sg13g2_a22oi_1 _22623_ (.Y(_15660_),
    .B1(\u_inv.f_reg[115] ),
    .B2(\u_inv.f_next[115] ),
    .A2(\u_inv.f_reg[114] ),
    .A1(\u_inv.f_next[114] ));
 sg13g2_a21oi_1 _22624_ (.A1(_14059_),
    .A2(_14369_),
    .Y(_15661_),
    .B1(_15660_));
 sg13g2_inv_1 _22625_ (.Y(_15662_),
    .A(_15661_));
 sg13g2_a21oi_1 _22626_ (.A1(_15647_),
    .A2(_15659_),
    .Y(_15663_),
    .B1(_15661_));
 sg13g2_a21oi_1 _22627_ (.A1(_14055_),
    .A2(_14373_),
    .Y(_15664_),
    .B1(_15632_));
 sg13g2_a22oi_1 _22628_ (.Y(_15665_),
    .B1(\u_inv.f_reg[117] ),
    .B2(\u_inv.f_next[117] ),
    .A2(\u_inv.f_reg[116] ),
    .A1(\u_inv.f_next[116] ));
 sg13g2_a21oi_1 _22629_ (.A1(_14057_),
    .A2(_14371_),
    .Y(_15666_),
    .B1(_15665_));
 sg13g2_a221oi_1 _22630_ (.B2(_15666_),
    .C1(_15664_),
    .B1(_15634_),
    .A1(\u_inv.f_next[119] ),
    .Y(_15667_),
    .A2(\u_inv.f_reg[119] ));
 sg13g2_o21ai_1 _22631_ (.B1(_15667_),
    .Y(_15668_),
    .A1(_15640_),
    .A2(_15663_));
 sg13g2_inv_1 _22632_ (.Y(_15669_),
    .A(_15668_));
 sg13g2_a22oi_1 _22633_ (.Y(_15670_),
    .B1(\u_inv.f_reg[121] ),
    .B2(\u_inv.f_next[121] ),
    .A2(\u_inv.f_reg[120] ),
    .A1(\u_inv.f_next[120] ));
 sg13g2_a21oi_1 _22634_ (.A1(_14053_),
    .A2(_14375_),
    .Y(_15671_),
    .B1(_15670_));
 sg13g2_a22oi_1 _22635_ (.Y(_15672_),
    .B1(_15625_),
    .B2(_15671_),
    .A2(\u_inv.f_reg[123] ),
    .A1(\u_inv.f_next[123] ));
 sg13g2_o21ai_1 _22636_ (.B1(_15672_),
    .Y(_15673_),
    .A1(_15621_),
    .A2(_15623_));
 sg13g2_nand2b_1 _22637_ (.Y(_15674_),
    .B(_15673_),
    .A_N(_15620_));
 sg13g2_a21oi_1 _22638_ (.A1(_14047_),
    .A2(_14381_),
    .Y(_15675_),
    .B1(_15612_));
 sg13g2_a22oi_1 _22639_ (.Y(_15676_),
    .B1(\u_inv.f_reg[125] ),
    .B2(\u_inv.f_next[125] ),
    .A2(\u_inv.f_reg[124] ),
    .A1(\u_inv.f_next[124] ));
 sg13g2_a21oi_1 _22640_ (.A1(_14049_),
    .A2(_14379_),
    .Y(_15677_),
    .B1(_15676_));
 sg13g2_a221oi_1 _22641_ (.B2(_15677_),
    .C1(_15675_),
    .B1(_15615_),
    .A1(\u_inv.f_next[127] ),
    .Y(_15678_),
    .A2(\u_inv.f_reg[127] ));
 sg13g2_nand2_1 _22642_ (.Y(_15679_),
    .A(_15674_),
    .B(_15678_));
 sg13g2_a21oi_2 _22643_ (.B1(_15679_),
    .Y(_15680_),
    .A2(_15668_),
    .A1(_15630_));
 sg13g2_inv_1 _22644_ (.Y(_15681_),
    .A(_15680_));
 sg13g2_nand2_2 _22645_ (.Y(_15682_),
    .A(_15656_),
    .B(_15680_));
 sg13g2_nand2_1 _22646_ (.Y(_15683_),
    .A(_14031_),
    .B(_14397_));
 sg13g2_nor2_1 _22647_ (.A(_14031_),
    .B(_14397_),
    .Y(_15684_));
 sg13g2_xor2_1 _22648_ (.B(\u_inv.f_reg[143] ),
    .A(\u_inv.f_next[143] ),
    .X(_15685_));
 sg13g2_nor2_1 _22649_ (.A(_14032_),
    .B(_14396_),
    .Y(_15686_));
 sg13g2_xor2_1 _22650_ (.B(\u_inv.f_reg[142] ),
    .A(\u_inv.f_next[142] ),
    .X(_15687_));
 sg13g2_xnor2_1 _22651_ (.Y(_15688_),
    .A(\u_inv.f_next[142] ),
    .B(\u_inv.f_reg[142] ));
 sg13g2_nand2_1 _22652_ (.Y(_15689_),
    .A(_15685_),
    .B(_15687_));
 sg13g2_xor2_1 _22653_ (.B(\u_inv.f_reg[141] ),
    .A(\u_inv.f_next[141] ),
    .X(_15690_));
 sg13g2_xnor2_1 _22654_ (.Y(_15691_),
    .A(\u_inv.f_next[141] ),
    .B(\u_inv.f_reg[141] ));
 sg13g2_nand2_1 _22655_ (.Y(_15692_),
    .A(\u_inv.f_next[140] ),
    .B(\u_inv.f_reg[140] ));
 sg13g2_xnor2_1 _22656_ (.Y(_15693_),
    .A(\u_inv.f_next[140] ),
    .B(\u_inv.f_reg[140] ));
 sg13g2_or2_1 _22657_ (.X(_15694_),
    .B(_15693_),
    .A(_15691_));
 sg13g2_or2_1 _22658_ (.X(_15695_),
    .B(_15694_),
    .A(_15689_));
 sg13g2_nand2_2 _22659_ (.Y(_15696_),
    .A(\u_inv.f_next[136] ),
    .B(\u_inv.f_reg[136] ));
 sg13g2_nand2_1 _22660_ (.Y(_15697_),
    .A(_14038_),
    .B(_14390_));
 sg13g2_and2_1 _22661_ (.A(_15696_),
    .B(_15697_),
    .X(_15698_));
 sg13g2_nand2_1 _22662_ (.Y(_15699_),
    .A(_15696_),
    .B(_15697_));
 sg13g2_nor2_1 _22663_ (.A(\u_inv.f_next[137] ),
    .B(\u_inv.f_reg[137] ),
    .Y(_15700_));
 sg13g2_nand2_1 _22664_ (.Y(_15701_),
    .A(\u_inv.f_next[137] ),
    .B(\u_inv.f_reg[137] ));
 sg13g2_nor2b_2 _22665_ (.A(_15700_),
    .B_N(_15701_),
    .Y(_15702_));
 sg13g2_nand2_1 _22666_ (.Y(_15703_),
    .A(_15698_),
    .B(_15702_));
 sg13g2_xor2_1 _22667_ (.B(\u_inv.f_reg[139] ),
    .A(\u_inv.f_next[139] ),
    .X(_15704_));
 sg13g2_nor2_1 _22668_ (.A(_14036_),
    .B(_14392_),
    .Y(_15705_));
 sg13g2_xor2_1 _22669_ (.B(\u_inv.f_reg[138] ),
    .A(\u_inv.f_next[138] ),
    .X(_15706_));
 sg13g2_xnor2_1 _22670_ (.Y(_15707_),
    .A(\u_inv.f_next[138] ),
    .B(\u_inv.f_reg[138] ));
 sg13g2_and2_1 _22671_ (.A(_15704_),
    .B(_15706_),
    .X(_15708_));
 sg13g2_nand2b_1 _22672_ (.Y(_15709_),
    .B(_15708_),
    .A_N(_15695_));
 sg13g2_nor2_1 _22673_ (.A(_15703_),
    .B(_15709_),
    .Y(_15710_));
 sg13g2_nand2_1 _22674_ (.Y(_15711_),
    .A(\u_inv.f_next[134] ),
    .B(\u_inv.f_reg[134] ));
 sg13g2_xnor2_1 _22675_ (.Y(_15712_),
    .A(\u_inv.f_next[134] ),
    .B(\u_inv.f_reg[134] ));
 sg13g2_xor2_1 _22676_ (.B(\u_inv.f_reg[135] ),
    .A(\u_inv.f_next[135] ),
    .X(_15713_));
 sg13g2_xnor2_1 _22677_ (.Y(_15714_),
    .A(\u_inv.f_next[135] ),
    .B(\u_inv.f_reg[135] ));
 sg13g2_nand2b_1 _22678_ (.Y(_15715_),
    .B(_15713_),
    .A_N(_15712_));
 sg13g2_nand2_1 _22679_ (.Y(_15716_),
    .A(\u_inv.f_next[133] ),
    .B(\u_inv.f_reg[133] ));
 sg13g2_nand2_1 _22680_ (.Y(_15717_),
    .A(_14041_),
    .B(_14387_));
 sg13g2_nand2_2 _22681_ (.Y(_15718_),
    .A(_15716_),
    .B(_15717_));
 sg13g2_nand2_1 _22682_ (.Y(_15719_),
    .A(\u_inv.f_next[132] ),
    .B(\u_inv.f_reg[132] ));
 sg13g2_xnor2_1 _22683_ (.Y(_15720_),
    .A(\u_inv.f_next[132] ),
    .B(\u_inv.f_reg[132] ));
 sg13g2_nor3_1 _22684_ (.A(_15715_),
    .B(_15718_),
    .C(_15720_),
    .Y(_15721_));
 sg13g2_nand2_1 _22685_ (.Y(_15722_),
    .A(\u_inv.f_next[130] ),
    .B(\u_inv.f_reg[130] ));
 sg13g2_xor2_1 _22686_ (.B(\u_inv.f_reg[130] ),
    .A(\u_inv.f_next[130] ),
    .X(_15723_));
 sg13g2_xnor2_1 _22687_ (.Y(_15724_),
    .A(\u_inv.f_next[130] ),
    .B(\u_inv.f_reg[130] ));
 sg13g2_nor2_1 _22688_ (.A(\u_inv.f_next[131] ),
    .B(\u_inv.f_reg[131] ),
    .Y(_15725_));
 sg13g2_xnor2_1 _22689_ (.Y(_15726_),
    .A(\u_inv.f_next[131] ),
    .B(\u_inv.f_reg[131] ));
 sg13g2_nor2_1 _22690_ (.A(_15724_),
    .B(_15726_),
    .Y(_15727_));
 sg13g2_xnor2_1 _22691_ (.Y(_15728_),
    .A(\u_inv.f_next[129] ),
    .B(\u_inv.f_reg[129] ));
 sg13g2_nor2_1 _22692_ (.A(_14046_),
    .B(_14382_),
    .Y(_15729_));
 sg13g2_xor2_1 _22693_ (.B(\u_inv.f_reg[128] ),
    .A(\u_inv.f_next[128] ),
    .X(_15730_));
 sg13g2_xnor2_1 _22694_ (.Y(_15731_),
    .A(\u_inv.f_next[128] ),
    .B(\u_inv.f_reg[128] ));
 sg13g2_nor2_1 _22695_ (.A(_15728_),
    .B(_15731_),
    .Y(_15732_));
 sg13g2_and2_1 _22696_ (.A(_15727_),
    .B(_15732_),
    .X(_15733_));
 sg13g2_inv_1 _22697_ (.Y(_15734_),
    .A(_15733_));
 sg13g2_and3_2 _22698_ (.X(_15735_),
    .A(_15710_),
    .B(_15721_),
    .C(_15733_));
 sg13g2_o21ai_1 _22699_ (.B1(_15735_),
    .Y(_15736_),
    .A1(_15655_),
    .A2(_15681_));
 sg13g2_a21oi_1 _22700_ (.A1(\u_inv.f_next[129] ),
    .A2(\u_inv.f_reg[129] ),
    .Y(_15737_),
    .B1(_15729_));
 sg13g2_a21oi_1 _22701_ (.A1(_14045_),
    .A2(_14383_),
    .Y(_15738_),
    .B1(_15737_));
 sg13g2_a22oi_1 _22702_ (.Y(_15739_),
    .B1(_15727_),
    .B2(_15738_),
    .A2(\u_inv.f_reg[131] ),
    .A1(\u_inv.f_next[131] ));
 sg13g2_o21ai_1 _22703_ (.B1(_15739_),
    .Y(_15740_),
    .A1(_15722_),
    .A2(_15725_));
 sg13g2_nand2_1 _22704_ (.Y(_15741_),
    .A(_15716_),
    .B(_15719_));
 sg13g2_nand2_1 _22705_ (.Y(_15742_),
    .A(_15717_),
    .B(_15741_));
 sg13g2_a21oi_1 _22706_ (.A1(_14039_),
    .A2(_14389_),
    .Y(_15743_),
    .B1(_15711_));
 sg13g2_a221oi_1 _22707_ (.B2(_15740_),
    .C1(_15743_),
    .B1(_15721_),
    .A1(\u_inv.f_next[135] ),
    .Y(_15744_),
    .A2(\u_inv.f_reg[135] ));
 sg13g2_o21ai_1 _22708_ (.B1(_15744_),
    .Y(_15745_),
    .A1(_15715_),
    .A2(_15742_));
 sg13g2_nand2_1 _22709_ (.Y(_15746_),
    .A(_15710_),
    .B(_15745_));
 sg13g2_a22oi_1 _22710_ (.Y(_15747_),
    .B1(\u_inv.f_reg[141] ),
    .B2(\u_inv.f_next[141] ),
    .A2(\u_inv.f_reg[140] ),
    .A1(\u_inv.f_next[140] ));
 sg13g2_a21o_1 _22711_ (.A2(_14395_),
    .A1(_14033_),
    .B1(_15747_),
    .X(_15748_));
 sg13g2_a21oi_1 _22712_ (.A1(_15683_),
    .A2(_15686_),
    .Y(_15749_),
    .B1(_15684_));
 sg13g2_o21ai_1 _22713_ (.B1(_15749_),
    .Y(_15750_),
    .A1(_15689_),
    .A2(_15748_));
 sg13g2_nand2_1 _22714_ (.Y(_15751_),
    .A(_15696_),
    .B(_15701_));
 sg13g2_o21ai_1 _22715_ (.B1(_15701_),
    .Y(_15752_),
    .A1(_15696_),
    .A2(_15700_));
 sg13g2_nand2b_1 _22716_ (.Y(_15753_),
    .B(_15751_),
    .A_N(_15700_));
 sg13g2_o21ai_1 _22717_ (.B1(_15705_),
    .Y(_15754_),
    .A1(\u_inv.f_next[139] ),
    .A2(\u_inv.f_reg[139] ));
 sg13g2_o21ai_1 _22718_ (.B1(_15754_),
    .Y(_15755_),
    .A1(_14035_),
    .A2(_14393_));
 sg13g2_a21oi_1 _22719_ (.A1(_15708_),
    .A2(_15752_),
    .Y(_15756_),
    .B1(_15755_));
 sg13g2_o21ai_1 _22720_ (.B1(_15746_),
    .Y(_15757_),
    .A1(_15695_),
    .A2(_15756_));
 sg13g2_nor2_2 _22721_ (.A(_15750_),
    .B(_15757_),
    .Y(_15758_));
 sg13g2_nor2b_1 _22722_ (.A(_15758_),
    .B_N(_15097_),
    .Y(_15759_));
 sg13g2_nor3_2 _22723_ (.A(_15107_),
    .B(_15119_),
    .C(_15759_),
    .Y(_15760_));
 sg13g2_inv_2 _22724_ (.Y(_15761_),
    .A(_15760_));
 sg13g2_nand2_1 _22725_ (.Y(_15762_),
    .A(_15097_),
    .B(_15735_));
 sg13g2_a21oi_2 _22726_ (.B1(_15762_),
    .Y(_15763_),
    .A2(_15680_),
    .A1(_15656_));
 sg13g2_a21o_2 _22727_ (.A2(_15680_),
    .A1(_15656_),
    .B1(_15762_),
    .X(_15764_));
 sg13g2_nor2_2 _22728_ (.A(_15761_),
    .B(_15763_),
    .Y(_15765_));
 sg13g2_xnor2_1 _22729_ (.Y(_15766_),
    .A(\u_inv.f_next[160] ),
    .B(\u_inv.f_reg[160] ));
 sg13g2_inv_1 _22730_ (.Y(_15767_),
    .A(_15766_));
 sg13g2_xnor2_1 _22731_ (.Y(_15768_),
    .A(\u_inv.f_next[161] ),
    .B(\u_inv.f_reg[161] ));
 sg13g2_or2_1 _22732_ (.X(_15769_),
    .B(_15768_),
    .A(_15766_));
 sg13g2_nor3_1 _22733_ (.A(_14981_),
    .B(_15766_),
    .C(_15768_),
    .Y(_15770_));
 sg13g2_nand2_1 _22734_ (.Y(_15771_),
    .A(_15015_),
    .B(_15770_));
 sg13g2_nor2_1 _22735_ (.A(_14961_),
    .B(_15771_),
    .Y(_15772_));
 sg13g2_o21ai_1 _22736_ (.B1(_15772_),
    .Y(_15773_),
    .A1(_15761_),
    .A2(_15763_));
 sg13g2_nand2_1 _22737_ (.Y(_15774_),
    .A(\u_inv.f_next[198] ),
    .B(\u_inv.f_reg[198] ));
 sg13g2_xor2_1 _22738_ (.B(\u_inv.f_reg[198] ),
    .A(\u_inv.f_next[198] ),
    .X(_15775_));
 sg13g2_xor2_1 _22739_ (.B(\u_inv.f_reg[199] ),
    .A(\u_inv.f_next[199] ),
    .X(_15776_));
 sg13g2_and2_1 _22740_ (.A(_15775_),
    .B(_15776_),
    .X(_15777_));
 sg13g2_xnor2_1 _22741_ (.Y(_15778_),
    .A(\u_inv.f_next[197] ),
    .B(\u_inv.f_reg[197] ));
 sg13g2_nor2_1 _22742_ (.A(_13978_),
    .B(_14450_),
    .Y(_15779_));
 sg13g2_xor2_1 _22743_ (.B(\u_inv.f_reg[196] ),
    .A(\u_inv.f_next[196] ),
    .X(_15780_));
 sg13g2_xnor2_1 _22744_ (.Y(_15781_),
    .A(\u_inv.f_next[196] ),
    .B(\u_inv.f_reg[196] ));
 sg13g2_nor2_1 _22745_ (.A(_15778_),
    .B(_15781_),
    .Y(_15782_));
 sg13g2_nand2_1 _22746_ (.Y(_15783_),
    .A(_15777_),
    .B(_15782_));
 sg13g2_nand2_1 _22747_ (.Y(_15784_),
    .A(\u_inv.f_next[194] ),
    .B(\u_inv.f_reg[194] ));
 sg13g2_xor2_1 _22748_ (.B(\u_inv.f_reg[194] ),
    .A(\u_inv.f_next[194] ),
    .X(_15785_));
 sg13g2_xnor2_1 _22749_ (.Y(_15786_),
    .A(\u_inv.f_next[194] ),
    .B(\u_inv.f_reg[194] ));
 sg13g2_xor2_1 _22750_ (.B(\u_inv.f_reg[195] ),
    .A(\u_inv.f_next[195] ),
    .X(_15787_));
 sg13g2_xnor2_1 _22751_ (.Y(_15788_),
    .A(\u_inv.f_next[195] ),
    .B(\u_inv.f_reg[195] ));
 sg13g2_nor2_1 _22752_ (.A(_15786_),
    .B(_15788_),
    .Y(_15789_));
 sg13g2_nand2_1 _22753_ (.Y(_15790_),
    .A(_15785_),
    .B(_15787_));
 sg13g2_xor2_1 _22754_ (.B(\u_inv.f_reg[193] ),
    .A(\u_inv.f_next[193] ),
    .X(_15791_));
 sg13g2_xnor2_1 _22755_ (.Y(_15792_),
    .A(\u_inv.f_next[193] ),
    .B(\u_inv.f_reg[193] ));
 sg13g2_xor2_1 _22756_ (.B(\u_inv.f_reg[192] ),
    .A(\u_inv.f_next[192] ),
    .X(_15793_));
 sg13g2_xnor2_1 _22757_ (.Y(_15794_),
    .A(\u_inv.f_next[192] ),
    .B(\u_inv.f_reg[192] ));
 sg13g2_nand2_1 _22758_ (.Y(_15795_),
    .A(_15791_),
    .B(_15793_));
 sg13g2_nor3_2 _22759_ (.A(_15783_),
    .B(_15790_),
    .C(_15795_),
    .Y(_15796_));
 sg13g2_inv_1 _22760_ (.Y(_15797_),
    .A(_15796_));
 sg13g2_nand2_1 _22761_ (.Y(_15798_),
    .A(\u_inv.f_next[206] ),
    .B(\u_inv.f_reg[206] ));
 sg13g2_xor2_1 _22762_ (.B(\u_inv.f_reg[206] ),
    .A(\u_inv.f_next[206] ),
    .X(_15799_));
 sg13g2_xnor2_1 _22763_ (.Y(_15800_),
    .A(\u_inv.f_next[206] ),
    .B(\u_inv.f_reg[206] ));
 sg13g2_xor2_1 _22764_ (.B(\u_inv.f_reg[207] ),
    .A(\u_inv.f_next[207] ),
    .X(_15801_));
 sg13g2_and2_1 _22765_ (.A(_15799_),
    .B(_15801_),
    .X(_15802_));
 sg13g2_nor2_1 _22766_ (.A(_13970_),
    .B(_14458_),
    .Y(_15803_));
 sg13g2_xnor2_1 _22767_ (.Y(_15804_),
    .A(\u_inv.f_next[204] ),
    .B(\u_inv.f_reg[204] ));
 sg13g2_inv_1 _22768_ (.Y(_15805_),
    .A(_15804_));
 sg13g2_nand2_1 _22769_ (.Y(_15806_),
    .A(\u_inv.f_next[205] ),
    .B(\u_inv.f_reg[205] ));
 sg13g2_nand2_1 _22770_ (.Y(_15807_),
    .A(_13969_),
    .B(_14459_));
 sg13g2_nand2_2 _22771_ (.Y(_15808_),
    .A(_15806_),
    .B(_15807_));
 sg13g2_nor2_1 _22772_ (.A(_15804_),
    .B(_15808_),
    .Y(_15809_));
 sg13g2_nand2_1 _22773_ (.Y(_15810_),
    .A(_15802_),
    .B(_15809_));
 sg13g2_xor2_1 _22774_ (.B(\u_inv.f_reg[200] ),
    .A(\u_inv.f_next[200] ),
    .X(_15811_));
 sg13g2_xnor2_1 _22775_ (.Y(_15812_),
    .A(\u_inv.f_next[200] ),
    .B(\u_inv.f_reg[200] ));
 sg13g2_xnor2_1 _22776_ (.Y(_15813_),
    .A(\u_inv.f_next[201] ),
    .B(\u_inv.f_reg[201] ));
 sg13g2_nor2_1 _22777_ (.A(_13972_),
    .B(_14456_),
    .Y(_15814_));
 sg13g2_xor2_1 _22778_ (.B(\u_inv.f_reg[202] ),
    .A(\u_inv.f_next[202] ),
    .X(_15815_));
 sg13g2_inv_1 _22779_ (.Y(_15816_),
    .A(_15815_));
 sg13g2_nand2_1 _22780_ (.Y(_15817_),
    .A(\u_inv.f_next[203] ),
    .B(\u_inv.f_reg[203] ));
 sg13g2_xnor2_1 _22781_ (.Y(_15818_),
    .A(\u_inv.f_next[203] ),
    .B(\u_inv.f_reg[203] ));
 sg13g2_or2_1 _22782_ (.X(_15819_),
    .B(_15818_),
    .A(_15816_));
 sg13g2_nor3_1 _22783_ (.A(_15812_),
    .B(_15813_),
    .C(_15819_),
    .Y(_15820_));
 sg13g2_nor2b_1 _22784_ (.A(_15810_),
    .B_N(_15820_),
    .Y(_15821_));
 sg13g2_nand2_2 _22785_ (.Y(_15822_),
    .A(_15796_),
    .B(_15821_));
 sg13g2_a21o_1 _22786_ (.A2(_15773_),
    .A1(_15049_),
    .B1(_15822_),
    .X(_15823_));
 sg13g2_a22oi_1 _22787_ (.Y(_15824_),
    .B1(\u_inv.f_reg[193] ),
    .B2(\u_inv.f_next[193] ),
    .A2(\u_inv.f_reg[192] ),
    .A1(\u_inv.f_next[192] ));
 sg13g2_a21oi_1 _22788_ (.A1(_13981_),
    .A2(_14447_),
    .Y(_15825_),
    .B1(_15824_));
 sg13g2_inv_1 _22789_ (.Y(_15826_),
    .A(_15825_));
 sg13g2_a22oi_1 _22790_ (.Y(_15827_),
    .B1(\u_inv.f_reg[195] ),
    .B2(\u_inv.f_next[195] ),
    .A2(\u_inv.f_reg[194] ),
    .A1(\u_inv.f_next[194] ));
 sg13g2_a21oi_1 _22791_ (.A1(_13979_),
    .A2(_14449_),
    .Y(_15828_),
    .B1(_15827_));
 sg13g2_inv_1 _22792_ (.Y(_15829_),
    .A(_15828_));
 sg13g2_a21oi_1 _22793_ (.A1(_15789_),
    .A2(_15825_),
    .Y(_15830_),
    .B1(_15828_));
 sg13g2_a21oi_1 _22794_ (.A1(_13975_),
    .A2(_14453_),
    .Y(_15831_),
    .B1(_15774_));
 sg13g2_a21oi_1 _22795_ (.A1(\u_inv.f_next[197] ),
    .A2(\u_inv.f_reg[197] ),
    .Y(_15832_),
    .B1(_15779_));
 sg13g2_a21oi_1 _22796_ (.A1(_13977_),
    .A2(_14451_),
    .Y(_15833_),
    .B1(_15832_));
 sg13g2_a221oi_1 _22797_ (.B2(_15833_),
    .C1(_15831_),
    .B1(_15777_),
    .A1(\u_inv.f_next[199] ),
    .Y(_15834_),
    .A2(\u_inv.f_reg[199] ));
 sg13g2_o21ai_1 _22798_ (.B1(_15834_),
    .Y(_15835_),
    .A1(_15783_),
    .A2(_15830_));
 sg13g2_a22oi_1 _22799_ (.Y(_15836_),
    .B1(\u_inv.f_reg[201] ),
    .B2(\u_inv.f_next[201] ),
    .A2(\u_inv.f_reg[200] ),
    .A1(\u_inv.f_next[200] ));
 sg13g2_a21o_1 _22800_ (.A2(_14455_),
    .A1(_13973_),
    .B1(_15836_),
    .X(_15837_));
 sg13g2_o21ai_1 _22801_ (.B1(_15814_),
    .Y(_15838_),
    .A1(\u_inv.f_next[203] ),
    .A2(\u_inv.f_reg[203] ));
 sg13g2_o21ai_1 _22802_ (.B1(_15817_),
    .Y(_15839_),
    .A1(_15819_),
    .A2(_15837_));
 sg13g2_nor2b_2 _22803_ (.A(_15839_),
    .B_N(_15838_),
    .Y(_15840_));
 sg13g2_nand2_1 _22804_ (.Y(_15841_),
    .A(_15803_),
    .B(_15807_));
 sg13g2_nand2_1 _22805_ (.Y(_15842_),
    .A(_15806_),
    .B(_15841_));
 sg13g2_a21oi_1 _22806_ (.A1(_13967_),
    .A2(_14461_),
    .Y(_15843_),
    .B1(_15798_));
 sg13g2_a221oi_1 _22807_ (.B2(_15842_),
    .C1(_15843_),
    .B1(_15802_),
    .A1(\u_inv.f_next[207] ),
    .Y(_15844_),
    .A2(\u_inv.f_reg[207] ));
 sg13g2_o21ai_1 _22808_ (.B1(_15844_),
    .Y(_15845_),
    .A1(_15810_),
    .A2(_15840_));
 sg13g2_a21o_2 _22809_ (.A2(_15835_),
    .A1(_15821_),
    .B1(_15845_),
    .X(_15846_));
 sg13g2_inv_1 _22810_ (.Y(_15847_),
    .A(_15846_));
 sg13g2_nand3_1 _22811_ (.B(_14911_),
    .C(_14913_),
    .A(_14895_),
    .Y(_15848_));
 sg13g2_nor2_1 _22812_ (.A(_14891_),
    .B(_15848_),
    .Y(_15849_));
 sg13g2_inv_1 _22813_ (.Y(_15850_),
    .A(_15849_));
 sg13g2_nand3_1 _22814_ (.B(_15846_),
    .C(_15849_),
    .A(_14879_),
    .Y(_15851_));
 sg13g2_nand4_1 _22815_ (.B(_14873_),
    .C(_14910_),
    .A(_14869_),
    .Y(_15852_),
    .D(_15851_));
 sg13g2_nor4_1 _22816_ (.A(_14856_),
    .B(_14878_),
    .C(_15822_),
    .D(_15850_),
    .Y(_15853_));
 sg13g2_inv_1 _22817_ (.Y(_15854_),
    .A(_15853_));
 sg13g2_a21oi_2 _22818_ (.B1(_15854_),
    .Y(_15855_),
    .A2(_15773_),
    .A1(_15049_));
 sg13g2_xor2_1 _22819_ (.B(\u_inv.f_reg[229] ),
    .A(\u_inv.f_next[229] ),
    .X(_15856_));
 sg13g2_nor2_1 _22820_ (.A(_13946_),
    .B(_14482_),
    .Y(_15857_));
 sg13g2_xor2_1 _22821_ (.B(\u_inv.f_reg[228] ),
    .A(\u_inv.f_next[228] ),
    .X(_15858_));
 sg13g2_xnor2_1 _22822_ (.Y(_15859_),
    .A(\u_inv.f_next[228] ),
    .B(\u_inv.f_reg[228] ));
 sg13g2_and2_1 _22823_ (.A(_15856_),
    .B(_15858_),
    .X(_15860_));
 sg13g2_nand2_1 _22824_ (.Y(_15861_),
    .A(\u_inv.f_next[231] ),
    .B(\u_inv.f_reg[231] ));
 sg13g2_nor2_1 _22825_ (.A(\u_inv.f_next[231] ),
    .B(\u_inv.f_reg[231] ),
    .Y(_15862_));
 sg13g2_xor2_1 _22826_ (.B(\u_inv.f_reg[231] ),
    .A(\u_inv.f_next[231] ),
    .X(_15863_));
 sg13g2_nand2_1 _22827_ (.Y(_15864_),
    .A(\u_inv.f_next[230] ),
    .B(\u_inv.f_reg[230] ));
 sg13g2_xor2_1 _22828_ (.B(\u_inv.f_reg[230] ),
    .A(\u_inv.f_next[230] ),
    .X(_15865_));
 sg13g2_xnor2_1 _22829_ (.Y(_15866_),
    .A(\u_inv.f_next[230] ),
    .B(\u_inv.f_reg[230] ));
 sg13g2_nand3_1 _22830_ (.B(_15863_),
    .C(_15865_),
    .A(_15860_),
    .Y(_15867_));
 sg13g2_nand2_1 _22831_ (.Y(_15868_),
    .A(\u_inv.f_next[227] ),
    .B(\u_inv.f_reg[227] ));
 sg13g2_xor2_1 _22832_ (.B(\u_inv.f_reg[227] ),
    .A(\u_inv.f_next[227] ),
    .X(_15869_));
 sg13g2_nand2_1 _22833_ (.Y(_15870_),
    .A(\u_inv.f_next[226] ),
    .B(\u_inv.f_reg[226] ));
 sg13g2_xor2_1 _22834_ (.B(\u_inv.f_reg[226] ),
    .A(\u_inv.f_next[226] ),
    .X(_15871_));
 sg13g2_xnor2_1 _22835_ (.Y(_15872_),
    .A(\u_inv.f_next[226] ),
    .B(\u_inv.f_reg[226] ));
 sg13g2_nand2_1 _22836_ (.Y(_15873_),
    .A(_15869_),
    .B(_15871_));
 sg13g2_xnor2_1 _22837_ (.Y(_15874_),
    .A(\u_inv.f_next[225] ),
    .B(\u_inv.f_reg[225] ));
 sg13g2_nand2_1 _22838_ (.Y(_15875_),
    .A(\u_inv.f_next[224] ),
    .B(\u_inv.f_reg[224] ));
 sg13g2_xor2_1 _22839_ (.B(\u_inv.f_reg[224] ),
    .A(\u_inv.f_next[224] ),
    .X(_15876_));
 sg13g2_xnor2_1 _22840_ (.Y(_15877_),
    .A(\u_inv.f_next[224] ),
    .B(\u_inv.f_reg[224] ));
 sg13g2_nand2b_1 _22841_ (.Y(_15878_),
    .B(_15876_),
    .A_N(_15874_));
 sg13g2_inv_1 _22842_ (.Y(_15879_),
    .A(_15878_));
 sg13g2_nor3_1 _22843_ (.A(_15867_),
    .B(_15873_),
    .C(_15878_),
    .Y(_15880_));
 sg13g2_xnor2_1 _22844_ (.Y(_15881_),
    .A(\u_inv.f_next[237] ),
    .B(\u_inv.f_reg[237] ));
 sg13g2_nand2_1 _22845_ (.Y(_15882_),
    .A(\u_inv.f_next[236] ),
    .B(\u_inv.f_reg[236] ));
 sg13g2_xnor2_1 _22846_ (.Y(_15883_),
    .A(\u_inv.f_next[236] ),
    .B(\u_inv.f_reg[236] ));
 sg13g2_nor2_1 _22847_ (.A(_15881_),
    .B(_15883_),
    .Y(_15884_));
 sg13g2_xor2_1 _22848_ (.B(\u_inv.f_reg[239] ),
    .A(\u_inv.f_next[239] ),
    .X(_15885_));
 sg13g2_xnor2_1 _22849_ (.Y(_15886_),
    .A(\u_inv.f_next[239] ),
    .B(\u_inv.f_reg[239] ));
 sg13g2_nand2_1 _22850_ (.Y(_15887_),
    .A(\u_inv.f_next[238] ),
    .B(\u_inv.f_reg[238] ));
 sg13g2_xnor2_1 _22851_ (.Y(_15888_),
    .A(\u_inv.f_next[238] ),
    .B(\u_inv.f_reg[238] ));
 sg13g2_nor2_1 _22852_ (.A(_15886_),
    .B(_15888_),
    .Y(_15889_));
 sg13g2_nand2_1 _22853_ (.Y(_15890_),
    .A(_15884_),
    .B(_15889_));
 sg13g2_xnor2_1 _22854_ (.Y(_15891_),
    .A(\u_inv.f_next[233] ),
    .B(\u_inv.f_reg[233] ));
 sg13g2_xnor2_1 _22855_ (.Y(_15892_),
    .A(\u_inv.f_next[232] ),
    .B(\u_inv.f_reg[232] ));
 sg13g2_inv_1 _22856_ (.Y(_15893_),
    .A(_15892_));
 sg13g2_or2_1 _22857_ (.X(_15894_),
    .B(_15892_),
    .A(_15891_));
 sg13g2_nand2_1 _22858_ (.Y(_15895_),
    .A(\u_inv.f_next[234] ),
    .B(\u_inv.f_reg[234] ));
 sg13g2_xor2_1 _22859_ (.B(\u_inv.f_reg[234] ),
    .A(\u_inv.f_next[234] ),
    .X(_15896_));
 sg13g2_xor2_1 _22860_ (.B(\u_inv.f_reg[235] ),
    .A(\u_inv.f_next[235] ),
    .X(_15897_));
 sg13g2_xnor2_1 _22861_ (.Y(_15898_),
    .A(\u_inv.f_next[235] ),
    .B(\u_inv.f_reg[235] ));
 sg13g2_and2_1 _22862_ (.A(_15896_),
    .B(_15897_),
    .X(_15899_));
 sg13g2_nand2b_1 _22863_ (.Y(_15900_),
    .B(_15899_),
    .A_N(_15894_));
 sg13g2_nor2_1 _22864_ (.A(_15890_),
    .B(_15900_),
    .Y(_15901_));
 sg13g2_nand2_1 _22865_ (.Y(_15902_),
    .A(_15880_),
    .B(_15901_));
 sg13g2_inv_1 _22866_ (.Y(_15903_),
    .A(_15902_));
 sg13g2_o21ai_1 _22867_ (.B1(_15903_),
    .Y(_15904_),
    .A1(_15852_),
    .A2(_15855_));
 sg13g2_a22oi_1 _22868_ (.Y(_15905_),
    .B1(\u_inv.f_reg[225] ),
    .B2(\u_inv.f_next[225] ),
    .A2(\u_inv.f_reg[224] ),
    .A1(\u_inv.f_next[224] ));
 sg13g2_a21o_1 _22869_ (.A2(_14479_),
    .A1(_13949_),
    .B1(_15905_),
    .X(_15906_));
 sg13g2_a21oi_1 _22870_ (.A1(_13947_),
    .A2(_14481_),
    .Y(_15907_),
    .B1(_15870_));
 sg13g2_o21ai_1 _22871_ (.B1(_15868_),
    .Y(_15908_),
    .A1(_15873_),
    .A2(_15906_));
 sg13g2_nor2_1 _22872_ (.A(_15907_),
    .B(_15908_),
    .Y(_15909_));
 sg13g2_o21ai_1 _22873_ (.B1(_15861_),
    .Y(_15910_),
    .A1(_15862_),
    .A2(_15864_));
 sg13g2_a21oi_1 _22874_ (.A1(\u_inv.f_next[229] ),
    .A2(\u_inv.f_reg[229] ),
    .Y(_15911_),
    .B1(_15857_));
 sg13g2_a21oi_1 _22875_ (.A1(_13945_),
    .A2(_14483_),
    .Y(_15912_),
    .B1(_15911_));
 sg13g2_nand3_1 _22876_ (.B(_15865_),
    .C(_15912_),
    .A(_15863_),
    .Y(_15913_));
 sg13g2_o21ai_1 _22877_ (.B1(_15913_),
    .Y(_15914_),
    .A1(_15867_),
    .A2(_15909_));
 sg13g2_nor2_2 _22878_ (.A(_15910_),
    .B(_15914_),
    .Y(_15915_));
 sg13g2_nor2b_1 _22879_ (.A(_15915_),
    .B_N(_15901_),
    .Y(_15916_));
 sg13g2_a22oi_1 _22880_ (.Y(_15917_),
    .B1(\u_inv.f_reg[233] ),
    .B2(\u_inv.f_next[233] ),
    .A2(\u_inv.f_reg[232] ),
    .A1(\u_inv.f_next[232] ));
 sg13g2_a21oi_1 _22881_ (.A1(_13941_),
    .A2(_14487_),
    .Y(_15918_),
    .B1(_15917_));
 sg13g2_a21oi_1 _22882_ (.A1(_13939_),
    .A2(_14489_),
    .Y(_15919_),
    .B1(_15895_));
 sg13g2_a221oi_1 _22883_ (.B2(_15918_),
    .C1(_15919_),
    .B1(_15899_),
    .A1(\u_inv.f_next[235] ),
    .Y(_15920_),
    .A2(\u_inv.f_reg[235] ));
 sg13g2_inv_1 _22884_ (.Y(_15921_),
    .A(_15920_));
 sg13g2_a22oi_1 _22885_ (.Y(_15922_),
    .B1(\u_inv.f_reg[237] ),
    .B2(\u_inv.f_next[237] ),
    .A2(\u_inv.f_reg[236] ),
    .A1(\u_inv.f_next[236] ));
 sg13g2_a21oi_1 _22886_ (.A1(_13937_),
    .A2(_14491_),
    .Y(_15923_),
    .B1(_15922_));
 sg13g2_a21oi_1 _22887_ (.A1(_13935_),
    .A2(_14493_),
    .Y(_15924_),
    .B1(_15887_));
 sg13g2_a221oi_1 _22888_ (.B2(_15923_),
    .C1(_15924_),
    .B1(_15889_),
    .A1(\u_inv.f_next[239] ),
    .Y(_15925_),
    .A2(\u_inv.f_reg[239] ));
 sg13g2_o21ai_1 _22889_ (.B1(_15925_),
    .Y(_15926_),
    .A1(_15890_),
    .A2(_15920_));
 sg13g2_nor2_2 _22890_ (.A(_15916_),
    .B(_15926_),
    .Y(_15927_));
 sg13g2_nor2_1 _22891_ (.A(_13934_),
    .B(_14494_),
    .Y(_15928_));
 sg13g2_xnor2_1 _22892_ (.Y(_15929_),
    .A(\u_inv.f_next[240] ),
    .B(\u_inv.f_reg[240] ));
 sg13g2_xnor2_1 _22893_ (.Y(_15930_),
    .A(\u_inv.f_next[241] ),
    .B(\u_inv.f_reg[241] ));
 sg13g2_nor2_1 _22894_ (.A(_15929_),
    .B(_15930_),
    .Y(_15931_));
 sg13g2_inv_1 _22895_ (.Y(_15932_),
    .A(_15931_));
 sg13g2_a21oi_2 _22896_ (.B1(_15932_),
    .Y(_15933_),
    .A2(_15927_),
    .A1(_15904_));
 sg13g2_nand2_1 _22897_ (.Y(_15934_),
    .A(\u_inv.f_next[242] ),
    .B(\u_inv.f_reg[242] ));
 sg13g2_xor2_1 _22898_ (.B(\u_inv.f_reg[242] ),
    .A(\u_inv.f_next[242] ),
    .X(_15935_));
 sg13g2_nor2_1 _22899_ (.A(\u_inv.f_next[243] ),
    .B(\u_inv.f_reg[243] ),
    .Y(_15936_));
 sg13g2_xor2_1 _22900_ (.B(\u_inv.f_reg[243] ),
    .A(\u_inv.f_next[243] ),
    .X(_15937_));
 sg13g2_xnor2_1 _22901_ (.Y(_15938_),
    .A(\u_inv.f_next[243] ),
    .B(\u_inv.f_reg[243] ));
 sg13g2_and2_1 _22902_ (.A(_15935_),
    .B(_15937_),
    .X(_15939_));
 sg13g2_a21oi_1 _22903_ (.A1(\u_inv.f_next[241] ),
    .A2(\u_inv.f_reg[241] ),
    .Y(_15940_),
    .B1(_15928_));
 sg13g2_a21oi_1 _22904_ (.A1(_13933_),
    .A2(_14495_),
    .Y(_15941_),
    .B1(_15940_));
 sg13g2_a22oi_1 _22905_ (.Y(_15942_),
    .B1(_15939_),
    .B2(_15941_),
    .A2(\u_inv.f_reg[243] ),
    .A1(\u_inv.f_next[243] ));
 sg13g2_o21ai_1 _22906_ (.B1(_15942_),
    .Y(_15943_),
    .A1(_15934_),
    .A2(_15936_));
 sg13g2_nand2_1 _22907_ (.Y(_15944_),
    .A(_14846_),
    .B(_15943_));
 sg13g2_nand3_1 _22908_ (.B(_14841_),
    .C(_15944_),
    .A(_14840_),
    .Y(_15945_));
 sg13g2_nand3_1 _22909_ (.B(_15931_),
    .C(_15939_),
    .A(_14846_),
    .Y(_15946_));
 sg13g2_a21oi_1 _22910_ (.A1(_15904_),
    .A2(_15927_),
    .Y(_15947_),
    .B1(_15946_));
 sg13g2_nor2_1 _22911_ (.A(_15945_),
    .B(_15947_),
    .Y(_15948_));
 sg13g2_nand2_1 _22912_ (.Y(_15949_),
    .A(\u_inv.f_next[248] ),
    .B(\u_inv.f_reg[248] ));
 sg13g2_xnor2_1 _22913_ (.Y(_15950_),
    .A(\u_inv.f_next[248] ),
    .B(\u_inv.f_reg[248] ));
 sg13g2_xnor2_1 _22914_ (.Y(_15951_),
    .A(\u_inv.f_next[249] ),
    .B(\u_inv.f_reg[249] ));
 sg13g2_nor2_1 _22915_ (.A(_15950_),
    .B(_15951_),
    .Y(_15952_));
 sg13g2_o21ai_1 _22916_ (.B1(_15952_),
    .Y(_15953_),
    .A1(_15945_),
    .A2(_15947_));
 sg13g2_a22oi_1 _22917_ (.Y(_15954_),
    .B1(\u_inv.f_reg[249] ),
    .B2(\u_inv.f_next[249] ),
    .A2(\u_inv.f_reg[248] ),
    .A1(\u_inv.f_next[248] ));
 sg13g2_a21o_1 _22918_ (.A2(_14503_),
    .A1(_13925_),
    .B1(_15954_),
    .X(_15955_));
 sg13g2_a21oi_1 _22919_ (.A1(_15953_),
    .A2(_15955_),
    .Y(_15956_),
    .B1(_14830_));
 sg13g2_a21oi_1 _22920_ (.A1(\u_inv.f_next[250] ),
    .A2(\u_inv.f_reg[250] ),
    .Y(_15957_),
    .B1(_15956_));
 sg13g2_xnor2_1 _22921_ (.Y(_15958_),
    .A(_14829_),
    .B(_15957_));
 sg13g2_nor2_2 _22922_ (.A(net5714),
    .B(net1224),
    .Y(_15959_));
 sg13g2_or2_1 _22923_ (.X(_15960_),
    .B(\u_inv.delta_reg[2] ),
    .A(\u_inv.delta_reg[1] ));
 sg13g2_nor3_1 _22924_ (.A(\u_inv.delta_reg[3] ),
    .B(\u_inv.delta_reg[4] ),
    .C(_15960_),
    .Y(_15961_));
 sg13g2_nand2_1 _22925_ (.Y(_15962_),
    .A(_14245_),
    .B(_15961_));
 sg13g2_nor2_1 _22926_ (.A(net3441),
    .B(_15962_),
    .Y(_15963_));
 sg13g2_nor3_1 _22927_ (.A(\u_inv.delta_reg[7] ),
    .B(\u_inv.delta_reg[6] ),
    .C(_15962_),
    .Y(_15964_));
 sg13g2_nand2b_1 _22928_ (.Y(_15965_),
    .B(_15964_),
    .A_N(\u_inv.delta_reg[8] ));
 sg13g2_and2_1 _22929_ (.A(_15959_),
    .B(_15965_),
    .X(_15966_));
 sg13g2_nand2_1 _22930_ (.Y(_15967_),
    .A(\u_inv.delta_double[0] ),
    .B(_15959_));
 sg13g2_o21ai_1 _22931_ (.B1(_15959_),
    .Y(_15968_),
    .A1(\u_inv.delta_double[0] ),
    .A2(_15965_));
 sg13g2_nand2b_1 _22932_ (.Y(_15969_),
    .B(_15967_),
    .A_N(_15966_));
 sg13g2_o21ai_1 _22933_ (.B1(net5026),
    .Y(_15970_),
    .A1(\u_inv.f_next[251] ),
    .A2(net5730));
 sg13g2_a21oi_1 _22934_ (.A1(net5730),
    .A2(_15958_),
    .Y(_15971_),
    .B1(_15970_));
 sg13g2_and2_1 _22935_ (.A(_14848_),
    .B(_14849_),
    .X(_15972_));
 sg13g2_and2_1 _22936_ (.A(_14851_),
    .B(_14853_),
    .X(_15973_));
 sg13g2_and2_1 _22937_ (.A(_15972_),
    .B(_15973_),
    .X(_15974_));
 sg13g2_nor2_1 _22938_ (.A(_14874_),
    .B(_14876_),
    .Y(_15975_));
 sg13g2_or2_1 _22939_ (.X(_15976_),
    .B(_14876_),
    .A(_14874_));
 sg13g2_nor2_1 _22940_ (.A(_14858_),
    .B(_14860_),
    .Y(_15977_));
 sg13g2_nand3_1 _22941_ (.B(_15975_),
    .C(_15977_),
    .A(_15974_),
    .Y(_15978_));
 sg13g2_nand2_1 _22942_ (.Y(_15979_),
    .A(_14886_),
    .B(_14888_));
 sg13g2_nor3_1 _22943_ (.A(_14881_),
    .B(_14884_),
    .C(_15979_),
    .Y(_15980_));
 sg13g2_nand2_1 _22944_ (.Y(_15981_),
    .A(_14892_),
    .B(_14894_));
 sg13g2_nor3_1 _22945_ (.A(_14911_),
    .B(_14913_),
    .C(_15981_),
    .Y(_15982_));
 sg13g2_inv_1 _22946_ (.Y(_15983_),
    .A(_15982_));
 sg13g2_nand2_1 _22947_ (.Y(_15984_),
    .A(_15980_),
    .B(_15982_));
 sg13g2_or2_1 _22948_ (.X(_15985_),
    .B(_15984_),
    .A(_15978_));
 sg13g2_nand2_1 _22949_ (.Y(_15986_),
    .A(\u_inv.f_next[219] ),
    .B(_14473_));
 sg13g2_nand2_1 _22950_ (.Y(_15987_),
    .A(\u_inv.f_next[218] ),
    .B(_14472_));
 sg13g2_nand2_1 _22951_ (.Y(_15988_),
    .A(\u_inv.f_next[216] ),
    .B(_14470_));
 sg13g2_nor2_1 _22952_ (.A(_14876_),
    .B(_15988_),
    .Y(_15989_));
 sg13g2_a21o_1 _22953_ (.A2(_14471_),
    .A1(\u_inv.f_next[217] ),
    .B1(_15989_),
    .X(_15990_));
 sg13g2_o21ai_1 _22954_ (.B1(_15986_),
    .Y(_15991_),
    .A1(_14858_),
    .A2(_15987_));
 sg13g2_a21o_1 _22955_ (.A2(_15990_),
    .A1(_15977_),
    .B1(_15991_),
    .X(_15992_));
 sg13g2_and2_1 _22956_ (.A(_15974_),
    .B(_15992_),
    .X(_15993_));
 sg13g2_nor2_1 _22957_ (.A(_13954_),
    .B(\u_inv.f_reg[220] ),
    .Y(_15994_));
 sg13g2_nand2_1 _22958_ (.Y(_15995_),
    .A(_14851_),
    .B(_15994_));
 sg13g2_o21ai_1 _22959_ (.B1(_15995_),
    .Y(_15996_),
    .A1(_13953_),
    .A2(\u_inv.f_reg[221] ));
 sg13g2_nor2_1 _22960_ (.A(_13952_),
    .B(\u_inv.f_reg[222] ),
    .Y(_15997_));
 sg13g2_a22oi_1 _22961_ (.Y(_15998_),
    .B1(_15997_),
    .B2(_14849_),
    .A2(_15996_),
    .A1(_15972_));
 sg13g2_o21ai_1 _22962_ (.B1(_15998_),
    .Y(_15999_),
    .A1(_13951_),
    .A2(\u_inv.f_reg[223] ));
 sg13g2_nor2_1 _22963_ (.A(_13963_),
    .B(\u_inv.f_reg[211] ),
    .Y(_16000_));
 sg13g2_nor2_1 _22964_ (.A(_13964_),
    .B(\u_inv.f_reg[210] ),
    .Y(_16001_));
 sg13g2_nand2_1 _22965_ (.Y(_16002_),
    .A(\u_inv.f_next[209] ),
    .B(_14463_));
 sg13g2_nor2_1 _22966_ (.A(_13966_),
    .B(\u_inv.f_reg[208] ),
    .Y(_16003_));
 sg13g2_nand2_1 _22967_ (.Y(_16004_),
    .A(_14912_),
    .B(_16003_));
 sg13g2_a21oi_1 _22968_ (.A1(_16002_),
    .A2(_16004_),
    .Y(_16005_),
    .B1(_15981_));
 sg13g2_a21oi_1 _22969_ (.A1(_14892_),
    .A2(_16001_),
    .Y(_16006_),
    .B1(_16000_));
 sg13g2_nand2b_1 _22970_ (.Y(_16007_),
    .B(_16006_),
    .A_N(_16005_));
 sg13g2_inv_1 _22971_ (.Y(_16008_),
    .A(_16007_));
 sg13g2_and3_1 _22972_ (.X(_16009_),
    .A(\u_inv.f_next[212] ),
    .B(_14466_),
    .C(_14886_));
 sg13g2_a21oi_1 _22973_ (.A1(\u_inv.f_next[213] ),
    .A2(_14467_),
    .Y(_16010_),
    .B1(_16009_));
 sg13g2_inv_1 _22974_ (.Y(_16011_),
    .A(_16010_));
 sg13g2_nor2_1 _22975_ (.A(_13959_),
    .B(\u_inv.f_reg[215] ),
    .Y(_16012_));
 sg13g2_nand2_1 _22976_ (.Y(_16013_),
    .A(\u_inv.f_next[214] ),
    .B(_14468_));
 sg13g2_o21ai_1 _22977_ (.B1(_16013_),
    .Y(_16014_),
    .A1(_14881_),
    .A2(_16010_));
 sg13g2_a221oi_1 _22978_ (.B2(_14885_),
    .C1(_16012_),
    .B1(_16014_),
    .A1(_15980_),
    .Y(_16015_),
    .A2(_16007_));
 sg13g2_nor2_1 _22979_ (.A(_15978_),
    .B(_16015_),
    .Y(_16016_));
 sg13g2_nand2_1 _22980_ (.Y(_16017_),
    .A(\u_inv.f_next[151] ),
    .B(_14405_));
 sg13g2_nor2_1 _22981_ (.A(_14024_),
    .B(\u_inv.f_reg[150] ),
    .Y(_16018_));
 sg13g2_nand2_1 _22982_ (.Y(_16019_),
    .A(\u_inv.f_next[149] ),
    .B(_14403_));
 sg13g2_nor2_1 _22983_ (.A(_14026_),
    .B(\u_inv.f_reg[148] ),
    .Y(_16020_));
 sg13g2_nand2_1 _22984_ (.Y(_16021_),
    .A(_15090_),
    .B(_16020_));
 sg13g2_a21oi_1 _22985_ (.A1(_16019_),
    .A2(_16021_),
    .Y(_16022_),
    .B1(_15087_));
 sg13g2_nor2_1 _22986_ (.A(_16018_),
    .B(_16022_),
    .Y(_16023_));
 sg13g2_o21ai_1 _22987_ (.B1(_16017_),
    .Y(_16024_),
    .A1(_15085_),
    .A2(_16023_));
 sg13g2_nor4_1 _22988_ (.A(_15085_),
    .B(_15087_),
    .C(_15089_),
    .D(_15092_),
    .Y(_16025_));
 sg13g2_inv_1 _22989_ (.Y(_16026_),
    .A(_16025_));
 sg13g2_nand3_1 _22990_ (.B(_14398_),
    .C(_15083_),
    .A(\u_inv.f_next[144] ),
    .Y(_16027_));
 sg13g2_o21ai_1 _22991_ (.B1(_16027_),
    .Y(_16028_),
    .A1(_14029_),
    .A2(\u_inv.f_reg[145] ));
 sg13g2_nor2_1 _22992_ (.A(_15076_),
    .B(_15079_),
    .Y(_16029_));
 sg13g2_nor2_1 _22993_ (.A(_14027_),
    .B(\u_inv.f_reg[147] ),
    .Y(_16030_));
 sg13g2_nor2_1 _22994_ (.A(_14028_),
    .B(\u_inv.f_reg[146] ),
    .Y(_16031_));
 sg13g2_inv_1 _22995_ (.Y(_16032_),
    .A(_16031_));
 sg13g2_a221oi_1 _22996_ (.B2(_15077_),
    .C1(_16030_),
    .B1(_16031_),
    .A1(_16028_),
    .Y(_16033_),
    .A2(_16029_));
 sg13g2_nor2_1 _22997_ (.A(_16026_),
    .B(_16033_),
    .Y(_16034_));
 sg13g2_or2_1 _22998_ (.X(_16035_),
    .B(_16034_),
    .A(_16024_));
 sg13g2_nor2_1 _22999_ (.A(_15055_),
    .B(_15058_),
    .Y(_16036_));
 sg13g2_nand3b_1 _23000_ (.B(_15053_),
    .C(_16036_),
    .Y(_16037_),
    .A_N(_15050_));
 sg13g2_nand2_1 _23001_ (.Y(_16038_),
    .A(_15064_),
    .B(_15067_));
 sg13g2_and2_1 _23002_ (.A(_15070_),
    .B(_15072_),
    .X(_16039_));
 sg13g2_inv_1 _23003_ (.Y(_16040_),
    .A(_16039_));
 sg13g2_nor3_1 _23004_ (.A(_16037_),
    .B(_16038_),
    .C(_16040_),
    .Y(_16041_));
 sg13g2_nor2_1 _23005_ (.A(_14019_),
    .B(\u_inv.f_reg[155] ),
    .Y(_16042_));
 sg13g2_nand2_1 _23006_ (.Y(_16043_),
    .A(\u_inv.f_next[154] ),
    .B(_14408_));
 sg13g2_nand2_1 _23007_ (.Y(_16044_),
    .A(\u_inv.f_next[152] ),
    .B(_14406_));
 sg13g2_nor2_1 _23008_ (.A(_15069_),
    .B(_16044_),
    .Y(_16045_));
 sg13g2_nand3_1 _23009_ (.B(_14406_),
    .C(_15070_),
    .A(\u_inv.f_next[152] ),
    .Y(_16046_));
 sg13g2_a21oi_1 _23010_ (.A1(\u_inv.f_next[153] ),
    .A2(_14407_),
    .Y(_16047_),
    .B1(_16045_));
 sg13g2_o21ai_1 _23011_ (.B1(_16043_),
    .Y(_16048_),
    .A1(_15066_),
    .A2(_16047_));
 sg13g2_a21oi_1 _23012_ (.A1(_15064_),
    .A2(_16048_),
    .Y(_16049_),
    .B1(_16042_));
 sg13g2_nand2_1 _23013_ (.Y(_16050_),
    .A(\u_inv.f_next[156] ),
    .B(_14410_));
 sg13g2_nor2_1 _23014_ (.A(_15055_),
    .B(_16050_),
    .Y(_16051_));
 sg13g2_nand3_1 _23015_ (.B(_14410_),
    .C(_15056_),
    .A(\u_inv.f_next[156] ),
    .Y(_16052_));
 sg13g2_a21oi_1 _23016_ (.A1(\u_inv.f_next[157] ),
    .A2(_14411_),
    .Y(_16053_),
    .B1(_16051_));
 sg13g2_nor3_1 _23017_ (.A(_15050_),
    .B(_15052_),
    .C(_16053_),
    .Y(_16054_));
 sg13g2_nand2_1 _23018_ (.Y(_16055_),
    .A(\u_inv.f_next[158] ),
    .B(_14412_));
 sg13g2_nor2_1 _23019_ (.A(_15050_),
    .B(_16055_),
    .Y(_16056_));
 sg13g2_nor2_1 _23020_ (.A(_16054_),
    .B(_16056_),
    .Y(_16057_));
 sg13g2_o21ai_1 _23021_ (.B1(_16057_),
    .Y(_16058_),
    .A1(_16037_),
    .A2(_16049_));
 sg13g2_a221oi_1 _23022_ (.B2(_16041_),
    .C1(_16058_),
    .B1(_16035_),
    .A1(\u_inv.f_next[159] ),
    .Y(_16059_),
    .A2(_14413_));
 sg13g2_and2_1 _23023_ (.A(_15083_),
    .B(_15095_),
    .X(_16060_));
 sg13g2_nand2_1 _23024_ (.Y(_16061_),
    .A(_16029_),
    .B(_16060_));
 sg13g2_nand4_1 _23025_ (.B(_16029_),
    .C(_16041_),
    .A(_16025_),
    .Y(_16062_),
    .D(_16060_));
 sg13g2_and2_1 _23026_ (.A(_16059_),
    .B(_16062_),
    .X(_16063_));
 sg13g2_nor2_1 _23027_ (.A(_14155_),
    .B(\u_inv.f_reg[19] ),
    .Y(_16064_));
 sg13g2_nor2_1 _23028_ (.A(_14156_),
    .B(\u_inv.f_reg[18] ),
    .Y(_16065_));
 sg13g2_nand2_1 _23029_ (.Y(_16066_),
    .A(\u_inv.f_next[18] ),
    .B(_14272_));
 sg13g2_and2_1 _23030_ (.A(_15259_),
    .B(_15260_),
    .X(_16067_));
 sg13g2_nand2_1 _23031_ (.Y(_16068_),
    .A(\u_inv.f_next[10] ),
    .B(_14264_));
 sg13g2_nand2_1 _23032_ (.Y(_16069_),
    .A(\u_inv.f_next[9] ),
    .B(_14263_));
 sg13g2_xnor2_1 _23033_ (.Y(_16070_),
    .A(\u_inv.f_next[9] ),
    .B(\u_inv.f_reg[9] ));
 sg13g2_nor2_1 _23034_ (.A(_14166_),
    .B(\u_inv.f_reg[8] ),
    .Y(_16071_));
 sg13g2_nand2_1 _23035_ (.Y(_16072_),
    .A(\u_inv.f_next[7] ),
    .B(_14261_));
 sg13g2_nor2b_1 _23036_ (.A(\u_inv.f_reg[6] ),
    .B_N(\u_inv.f_next[6] ),
    .Y(_16073_));
 sg13g2_nand2_1 _23037_ (.Y(_16074_),
    .A(\u_inv.f_next[5] ),
    .B(_14259_));
 sg13g2_nor2b_1 _23038_ (.A(\u_inv.f_reg[4] ),
    .B_N(\u_inv.f_next[4] ),
    .Y(_16075_));
 sg13g2_nand2_1 _23039_ (.Y(_16076_),
    .A(\u_inv.f_next[3] ),
    .B(_14257_));
 sg13g2_nor2_1 _23040_ (.A(_14169_),
    .B(\u_inv.f_reg[2] ),
    .Y(_16077_));
 sg13g2_nor2b_1 _23041_ (.A(net5725),
    .B_N(\u_inv.f_reg[0] ),
    .Y(_16078_));
 sg13g2_a21oi_1 _23042_ (.A1(_15284_),
    .A2(_16078_),
    .Y(_16079_),
    .B1(_15283_));
 sg13g2_a221oi_1 _23043_ (.B2(_16078_),
    .C1(_15283_),
    .B1(_15284_),
    .A1(_15278_),
    .Y(_16080_),
    .A2(_15280_));
 sg13g2_o21ai_1 _23044_ (.B1(_15277_),
    .Y(_16081_),
    .A1(_16077_),
    .A2(_16080_));
 sg13g2_a21oi_1 _23045_ (.A1(_16076_),
    .A2(_16081_),
    .Y(_16082_),
    .B1(_15275_));
 sg13g2_o21ai_1 _23046_ (.B1(_15272_),
    .Y(_16083_),
    .A1(_16075_),
    .A2(_16082_));
 sg13g2_a21oi_1 _23047_ (.A1(_16074_),
    .A2(_16083_),
    .Y(_16084_),
    .B1(_15270_));
 sg13g2_o21ai_1 _23048_ (.B1(_15268_),
    .Y(_16085_),
    .A1(_16073_),
    .A2(_16084_));
 sg13g2_a21oi_1 _23049_ (.A1(_16072_),
    .A2(_16085_),
    .Y(_16086_),
    .B1(_15266_));
 sg13g2_o21ai_1 _23050_ (.B1(_16070_),
    .Y(_16087_),
    .A1(_16071_),
    .A2(_16086_));
 sg13g2_a21o_1 _23051_ (.A2(_16087_),
    .A1(_16069_),
    .B1(_15262_),
    .X(_16088_));
 sg13g2_a21o_2 _23052_ (.A2(_16088_),
    .A1(_16068_),
    .B1(_16067_),
    .X(_16089_));
 sg13g2_nand2_1 _23053_ (.Y(_16090_),
    .A(\u_inv.f_next[11] ),
    .B(_14265_));
 sg13g2_a21oi_1 _23054_ (.A1(_16089_),
    .A2(_16090_),
    .Y(_16091_),
    .B1(_15302_));
 sg13g2_a21o_1 _23055_ (.A2(_16090_),
    .A1(_16089_),
    .B1(_15302_),
    .X(_16092_));
 sg13g2_a21oi_1 _23056_ (.A1(\u_inv.f_next[12] ),
    .A2(_14266_),
    .Y(_16093_),
    .B1(_16091_));
 sg13g2_a22oi_1 _23057_ (.Y(_16094_),
    .B1(_14267_),
    .B2(\u_inv.f_next[13] ),
    .A2(_14266_),
    .A1(\u_inv.f_next[12] ));
 sg13g2_nand2_1 _23058_ (.Y(_16095_),
    .A(_16092_),
    .B(_16094_));
 sg13g2_o21ai_1 _23059_ (.B1(_16095_),
    .Y(_16096_),
    .A1(\u_inv.f_next[13] ),
    .A2(_14267_));
 sg13g2_nor2_1 _23060_ (.A(_15310_),
    .B(_16096_),
    .Y(_16097_));
 sg13g2_nor2_1 _23061_ (.A(_14160_),
    .B(\u_inv.f_reg[14] ),
    .Y(_16098_));
 sg13g2_nand2_1 _23062_ (.Y(_16099_),
    .A(_15311_),
    .B(_15315_));
 sg13g2_a221oi_1 _23063_ (.B2(_16094_),
    .C1(_16099_),
    .B1(_16092_),
    .A1(_14161_),
    .Y(_16100_),
    .A2(\u_inv.f_reg[13] ));
 sg13g2_nand2_1 _23064_ (.Y(_16101_),
    .A(_15315_),
    .B(_16098_));
 sg13g2_o21ai_1 _23065_ (.B1(_16101_),
    .Y(_16102_),
    .A1(_14159_),
    .A2(\u_inv.f_reg[15] ));
 sg13g2_nor2_1 _23066_ (.A(_16100_),
    .B(_16102_),
    .Y(_16103_));
 sg13g2_o21ai_1 _23067_ (.B1(_15327_),
    .Y(_16104_),
    .A1(_16100_),
    .A2(_16102_));
 sg13g2_nand2_1 _23068_ (.Y(_16105_),
    .A(\u_inv.f_next[16] ),
    .B(_14270_));
 sg13g2_nor2_1 _23069_ (.A(net5621),
    .B(_16105_),
    .Y(_16106_));
 sg13g2_a21oi_1 _23070_ (.A1(\u_inv.f_next[17] ),
    .A2(_14271_),
    .Y(_16107_),
    .B1(_16106_));
 sg13g2_a21o_1 _23071_ (.A2(_16105_),
    .A1(_16104_),
    .B1(net5621),
    .X(_16108_));
 sg13g2_o21ai_1 _23072_ (.B1(_16107_),
    .Y(_16109_),
    .A1(net5621),
    .A2(_16104_));
 sg13g2_nor4_1 _23073_ (.A(_15319_),
    .B(_15322_),
    .C(net5621),
    .D(_15326_),
    .Y(_16110_));
 sg13g2_o21ai_1 _23074_ (.B1(_16110_),
    .Y(_16111_),
    .A1(_16100_),
    .A2(_16102_));
 sg13g2_o21ai_1 _23075_ (.B1(_16066_),
    .Y(_16112_),
    .A1(_15322_),
    .A2(_16107_));
 sg13g2_a21oi_1 _23076_ (.A1(_15320_),
    .A2(_16112_),
    .Y(_16113_),
    .B1(_16064_));
 sg13g2_a21oi_2 _23077_ (.B1(_15346_),
    .Y(_16114_),
    .A2(_16113_),
    .A1(_16111_));
 sg13g2_nand2_1 _23078_ (.Y(_16115_),
    .A(_15344_),
    .B(_16114_));
 sg13g2_or4_1 _23079_ (.A(_15337_),
    .B(_15339_),
    .C(_15343_),
    .D(_15346_),
    .X(_16116_));
 sg13g2_a21o_1 _23080_ (.A2(_16113_),
    .A1(_16111_),
    .B1(_16116_),
    .X(_16117_));
 sg13g2_nor2_1 _23081_ (.A(_14152_),
    .B(\u_inv.f_reg[22] ),
    .Y(_16118_));
 sg13g2_nor2_1 _23082_ (.A(_14154_),
    .B(\u_inv.f_reg[20] ),
    .Y(_16119_));
 sg13g2_nand2_1 _23083_ (.Y(_16120_),
    .A(_15344_),
    .B(_16119_));
 sg13g2_o21ai_1 _23084_ (.B1(_16120_),
    .Y(_16121_),
    .A1(_14153_),
    .A2(\u_inv.f_reg[21] ));
 sg13g2_a21oi_1 _23085_ (.A1(_15340_),
    .A2(_16121_),
    .Y(_16122_),
    .B1(_16118_));
 sg13g2_nor2_1 _23086_ (.A(_15337_),
    .B(_16122_),
    .Y(_16123_));
 sg13g2_a21oi_1 _23087_ (.A1(\u_inv.f_next[23] ),
    .A2(_14277_),
    .Y(_16124_),
    .B1(_16123_));
 sg13g2_and2_1 _23088_ (.A(_16117_),
    .B(_16124_),
    .X(_16125_));
 sg13g2_or4_1 _23089_ (.A(_15357_),
    .B(_15359_),
    .C(_15364_),
    .D(_15365_),
    .X(_16126_));
 sg13g2_a21o_2 _23090_ (.A2(_16124_),
    .A1(_16117_),
    .B1(_16126_),
    .X(_16127_));
 sg13g2_nor2_1 _23091_ (.A(_14148_),
    .B(\u_inv.f_reg[26] ),
    .Y(_16128_));
 sg13g2_nand2_1 _23092_ (.Y(_16129_),
    .A(\u_inv.f_next[25] ),
    .B(_14279_));
 sg13g2_nand2_1 _23093_ (.Y(_16130_),
    .A(\u_inv.f_next[24] ),
    .B(_14278_));
 sg13g2_o21ai_1 _23094_ (.B1(_16129_),
    .Y(_16131_),
    .A1(_15365_),
    .A2(_16130_));
 sg13g2_a21oi_1 _23095_ (.A1(_15360_),
    .A2(_16131_),
    .Y(_16132_),
    .B1(_16128_));
 sg13g2_nor2_1 _23096_ (.A(_15357_),
    .B(_16132_),
    .Y(_16133_));
 sg13g2_a21oi_1 _23097_ (.A1(\u_inv.f_next[27] ),
    .A2(_14281_),
    .Y(_16134_),
    .B1(_16133_));
 sg13g2_nand2_1 _23098_ (.Y(_16135_),
    .A(_16127_),
    .B(_16134_));
 sg13g2_nor4_1 _23099_ (.A(_15372_),
    .B(_15374_),
    .C(_15378_),
    .D(_15380_),
    .Y(_16136_));
 sg13g2_inv_1 _23100_ (.Y(_16137_),
    .A(_16136_));
 sg13g2_a21o_2 _23101_ (.A2(_16134_),
    .A1(_16127_),
    .B1(_16137_),
    .X(_16138_));
 sg13g2_nand2_1 _23102_ (.Y(_16139_),
    .A(\u_inv.f_next[31] ),
    .B(_14285_));
 sg13g2_nand2_1 _23103_ (.Y(_16140_),
    .A(\u_inv.f_next[30] ),
    .B(_14284_));
 sg13g2_nand2_1 _23104_ (.Y(_16141_),
    .A(\u_inv.f_next[29] ),
    .B(_14283_));
 sg13g2_nand2_1 _23105_ (.Y(_16142_),
    .A(\u_inv.f_next[28] ),
    .B(_14282_));
 sg13g2_o21ai_1 _23106_ (.B1(_16141_),
    .Y(_16143_),
    .A1(_15380_),
    .A2(_16142_));
 sg13g2_nand2_1 _23107_ (.Y(_16144_),
    .A(_15375_),
    .B(_16143_));
 sg13g2_and2_1 _23108_ (.A(_16140_),
    .B(_16144_),
    .X(_16145_));
 sg13g2_o21ai_1 _23109_ (.B1(_16139_),
    .Y(_16146_),
    .A1(_15372_),
    .A2(_16145_));
 sg13g2_inv_1 _23110_ (.Y(_16147_),
    .A(_16146_));
 sg13g2_and3_1 _23111_ (.X(_16148_),
    .A(_15239_),
    .B(_15241_),
    .C(_15389_));
 sg13g2_inv_1 _23112_ (.Y(_16149_),
    .A(_16148_));
 sg13g2_nor4_1 _23113_ (.A(_15226_),
    .B(_15229_),
    .C(_15232_),
    .D(_15234_),
    .Y(_16150_));
 sg13g2_nand3b_1 _23114_ (.B(_16148_),
    .C(_16150_),
    .Y(_16151_),
    .A_N(_15390_));
 sg13g2_a21o_2 _23115_ (.A2(_16147_),
    .A1(_16138_),
    .B1(_16151_),
    .X(_16152_));
 sg13g2_nand2_2 _23116_ (.Y(_16153_),
    .A(\u_inv.f_next[32] ),
    .B(_14286_));
 sg13g2_nand2_1 _23117_ (.Y(_16154_),
    .A(\u_inv.f_next[34] ),
    .B(_14288_));
 sg13g2_nor2_1 _23118_ (.A(_14141_),
    .B(\u_inv.f_reg[33] ),
    .Y(_16155_));
 sg13g2_nand2_1 _23119_ (.Y(_16156_),
    .A(_15241_),
    .B(_16155_));
 sg13g2_a21oi_1 _23120_ (.A1(_16154_),
    .A2(_16156_),
    .Y(_16157_),
    .B1(_15238_));
 sg13g2_a21oi_1 _23121_ (.A1(\u_inv.f_next[35] ),
    .A2(_14289_),
    .Y(_16158_),
    .B1(_16157_));
 sg13g2_o21ai_1 _23122_ (.B1(_16158_),
    .Y(_16159_),
    .A1(_16149_),
    .A2(_16153_));
 sg13g2_nand2_1 _23123_ (.Y(_16160_),
    .A(\u_inv.f_next[37] ),
    .B(_14291_));
 sg13g2_nor2_1 _23124_ (.A(_14138_),
    .B(\u_inv.f_reg[36] ),
    .Y(_16161_));
 sg13g2_nand2_1 _23125_ (.Y(_16162_),
    .A(_15235_),
    .B(_16161_));
 sg13g2_nand2_1 _23126_ (.Y(_16163_),
    .A(\u_inv.f_next[38] ),
    .B(_14292_));
 sg13g2_a21o_1 _23127_ (.A2(_16162_),
    .A1(_16160_),
    .B1(_15229_),
    .X(_16164_));
 sg13g2_a21oi_1 _23128_ (.A1(_16163_),
    .A2(_16164_),
    .Y(_16165_),
    .B1(_15226_));
 sg13g2_a221oi_1 _23129_ (.B2(_16159_),
    .C1(_16165_),
    .B1(_16150_),
    .A1(\u_inv.f_next[39] ),
    .Y(_16166_),
    .A2(_14293_));
 sg13g2_nand2_1 _23130_ (.Y(_16167_),
    .A(_16152_),
    .B(_16166_));
 sg13g2_and2_1 _23131_ (.A(_15395_),
    .B(_15397_),
    .X(_16168_));
 sg13g2_nand2b_1 _23132_ (.Y(_16169_),
    .B(_16168_),
    .A_N(_15402_));
 sg13g2_nor2b_1 _23133_ (.A(_16169_),
    .B_N(_15401_),
    .Y(_16170_));
 sg13g2_nand2_1 _23134_ (.Y(_16171_),
    .A(net5620),
    .B(_15412_));
 sg13g2_and4_1 _23135_ (.A(_15405_),
    .B(net5620),
    .C(_15410_),
    .D(_15412_),
    .X(_16172_));
 sg13g2_and2_1 _23136_ (.A(_16170_),
    .B(_16172_),
    .X(_16173_));
 sg13g2_inv_1 _23137_ (.Y(_16174_),
    .A(_16173_));
 sg13g2_a21oi_2 _23138_ (.B1(_16174_),
    .Y(_16175_),
    .A2(_16166_),
    .A1(_16152_));
 sg13g2_nor2_1 _23139_ (.A(_14132_),
    .B(\u_inv.f_reg[42] ),
    .Y(_16176_));
 sg13g2_nor2_1 _23140_ (.A(_14133_),
    .B(\u_inv.f_reg[41] ),
    .Y(_16177_));
 sg13g2_nand2_1 _23141_ (.Y(_16178_),
    .A(\u_inv.f_next[40] ),
    .B(_14294_));
 sg13g2_a21oi_1 _23142_ (.A1(net5620),
    .A2(_16177_),
    .Y(_16179_),
    .B1(_16176_));
 sg13g2_o21ai_1 _23143_ (.B1(_16179_),
    .Y(_16180_),
    .A1(_16171_),
    .A2(_16178_));
 sg13g2_nand2_1 _23144_ (.Y(_16181_),
    .A(_15405_),
    .B(_16180_));
 sg13g2_o21ai_1 _23145_ (.B1(_16181_),
    .Y(_16182_),
    .A1(_14131_),
    .A2(\u_inv.f_reg[43] ));
 sg13g2_nand2_1 _23146_ (.Y(_16183_),
    .A(_16170_),
    .B(_16182_));
 sg13g2_nor2_1 _23147_ (.A(_14129_),
    .B(\u_inv.f_reg[45] ),
    .Y(_16184_));
 sg13g2_nand2_1 _23148_ (.Y(_16185_),
    .A(\u_inv.f_next[44] ),
    .B(_14298_));
 sg13g2_nor2_1 _23149_ (.A(_15402_),
    .B(_16185_),
    .Y(_16186_));
 sg13g2_o21ai_1 _23150_ (.B1(_16168_),
    .Y(_16187_),
    .A1(_16184_),
    .A2(_16186_));
 sg13g2_nor2_1 _23151_ (.A(_14128_),
    .B(\u_inv.f_reg[46] ),
    .Y(_16188_));
 sg13g2_nor2_1 _23152_ (.A(_14127_),
    .B(\u_inv.f_reg[47] ),
    .Y(_16189_));
 sg13g2_a21oi_1 _23153_ (.A1(_15395_),
    .A2(_16188_),
    .Y(_16190_),
    .B1(_16189_));
 sg13g2_nand3_1 _23154_ (.B(_16187_),
    .C(_16190_),
    .A(_16183_),
    .Y(_16191_));
 sg13g2_nand2_1 _23155_ (.Y(_16192_),
    .A(_15434_),
    .B(_15436_));
 sg13g2_nand2_1 _23156_ (.Y(_16193_),
    .A(_15439_),
    .B(_15440_));
 sg13g2_nor2_1 _23157_ (.A(_16192_),
    .B(_16193_),
    .Y(_16194_));
 sg13g2_and2_1 _23158_ (.A(_15442_),
    .B(_15444_),
    .X(_16195_));
 sg13g2_nor2_1 _23159_ (.A(_15428_),
    .B(_15431_),
    .Y(_16196_));
 sg13g2_nand3_1 _23160_ (.B(_16195_),
    .C(_16196_),
    .A(_16194_),
    .Y(_16197_));
 sg13g2_inv_1 _23161_ (.Y(_16198_),
    .A(_16197_));
 sg13g2_o21ai_1 _23162_ (.B1(_16198_),
    .Y(_16199_),
    .A1(_16175_),
    .A2(_16191_));
 sg13g2_nand2_1 _23163_ (.Y(_16200_),
    .A(\u_inv.f_next[48] ),
    .B(_14302_));
 sg13g2_nand3_1 _23164_ (.B(_14302_),
    .C(_15442_),
    .A(\u_inv.f_next[48] ),
    .Y(_16201_));
 sg13g2_nand2_1 _23165_ (.Y(_16202_),
    .A(\u_inv.f_next[49] ),
    .B(_14303_));
 sg13g2_and2_1 _23166_ (.A(_16201_),
    .B(_16202_),
    .X(_16203_));
 sg13g2_nand2b_1 _23167_ (.Y(_16204_),
    .B(_16194_),
    .A_N(_16203_));
 sg13g2_nand2_1 _23168_ (.Y(_16205_),
    .A(\u_inv.f_next[53] ),
    .B(_14307_));
 sg13g2_nor2_1 _23169_ (.A(_14122_),
    .B(\u_inv.f_reg[52] ),
    .Y(_16206_));
 sg13g2_nand2_1 _23170_ (.Y(_16207_),
    .A(_15434_),
    .B(_16206_));
 sg13g2_nand3_1 _23171_ (.B(_14304_),
    .C(_15440_),
    .A(\u_inv.f_next[50] ),
    .Y(_16208_));
 sg13g2_o21ai_1 _23172_ (.B1(_16208_),
    .Y(_16209_),
    .A1(_14123_),
    .A2(\u_inv.f_reg[51] ));
 sg13g2_nand2b_1 _23173_ (.Y(_16210_),
    .B(_16209_),
    .A_N(_16192_));
 sg13g2_nand4_1 _23174_ (.B(_16205_),
    .C(_16207_),
    .A(_16204_),
    .Y(_16211_),
    .D(_16210_));
 sg13g2_nand2_1 _23175_ (.Y(_16212_),
    .A(\u_inv.f_next[54] ),
    .B(_14308_));
 sg13g2_nor2_1 _23176_ (.A(_15428_),
    .B(_16212_),
    .Y(_16213_));
 sg13g2_a221oi_1 _23177_ (.B2(_16211_),
    .C1(_16213_),
    .B1(_16196_),
    .A1(\u_inv.f_next[55] ),
    .Y(_16214_),
    .A2(_14309_));
 sg13g2_nand2_1 _23178_ (.Y(_16215_),
    .A(_16199_),
    .B(_16214_));
 sg13g2_and2_1 _23179_ (.A(_15198_),
    .B(_15200_),
    .X(_16216_));
 sg13g2_nand3_1 _23180_ (.B(_15205_),
    .C(_16216_),
    .A(_15204_),
    .Y(_16217_));
 sg13g2_nor2_1 _23181_ (.A(_15208_),
    .B(_15210_),
    .Y(_16218_));
 sg13g2_nand2_1 _23182_ (.Y(_16219_),
    .A(_15460_),
    .B(_15462_));
 sg13g2_nor4_1 _23183_ (.A(_15208_),
    .B(_15210_),
    .C(_16217_),
    .D(_16219_),
    .Y(_16220_));
 sg13g2_inv_1 _23184_ (.Y(_16221_),
    .A(_16220_));
 sg13g2_a21o_2 _23185_ (.A2(_16214_),
    .A1(_16199_),
    .B1(_16221_),
    .X(_16222_));
 sg13g2_nand2_1 _23186_ (.Y(_16223_),
    .A(\u_inv.f_next[59] ),
    .B(_14313_));
 sg13g2_nor2_1 _23187_ (.A(_14116_),
    .B(\u_inv.f_reg[58] ),
    .Y(_16224_));
 sg13g2_nor2_1 _23188_ (.A(_14118_),
    .B(\u_inv.f_reg[56] ),
    .Y(_16225_));
 sg13g2_and2_1 _23189_ (.A(_15460_),
    .B(_16225_),
    .X(_16226_));
 sg13g2_a21o_1 _23190_ (.A2(_14311_),
    .A1(\u_inv.f_next[57] ),
    .B1(_16226_),
    .X(_16227_));
 sg13g2_a21oi_1 _23191_ (.A1(_15211_),
    .A2(_16227_),
    .Y(_16228_),
    .B1(_16224_));
 sg13g2_o21ai_1 _23192_ (.B1(_16223_),
    .Y(_16229_),
    .A1(_15208_),
    .A2(_16228_));
 sg13g2_nand2b_1 _23193_ (.Y(_16230_),
    .B(_16229_),
    .A_N(_16217_));
 sg13g2_nor2_1 _23194_ (.A(_14113_),
    .B(\u_inv.f_reg[61] ),
    .Y(_16231_));
 sg13g2_nand2_1 _23195_ (.Y(_16232_),
    .A(\u_inv.f_next[60] ),
    .B(_14314_));
 sg13g2_nor2b_1 _23196_ (.A(_16232_),
    .B_N(_15205_),
    .Y(_16233_));
 sg13g2_o21ai_1 _23197_ (.B1(_16216_),
    .Y(_16234_),
    .A1(_16231_),
    .A2(_16233_));
 sg13g2_nor2_1 _23198_ (.A(_14112_),
    .B(\u_inv.f_reg[62] ),
    .Y(_16235_));
 sg13g2_nor2_1 _23199_ (.A(_14111_),
    .B(\u_inv.f_reg[63] ),
    .Y(_16236_));
 sg13g2_a21oi_1 _23200_ (.A1(_15198_),
    .A2(_16235_),
    .Y(_16237_),
    .B1(_16236_));
 sg13g2_and3_2 _23201_ (.X(_16238_),
    .A(_16230_),
    .B(_16234_),
    .C(_16237_));
 sg13g2_nand3_1 _23202_ (.B(_15172_),
    .C(_15176_),
    .A(_15170_),
    .Y(_16239_));
 sg13g2_or2_1 _23203_ (.X(_16240_),
    .B(_16239_),
    .A(_15177_));
 sg13g2_nor2_1 _23204_ (.A(_15180_),
    .B(_15181_),
    .Y(_16241_));
 sg13g2_nand2b_1 _23205_ (.Y(_16242_),
    .B(_16241_),
    .A_N(_15469_));
 sg13g2_or3_1 _23206_ (.A(_15467_),
    .B(_16240_),
    .C(_16242_),
    .X(_16243_));
 sg13g2_a21oi_2 _23207_ (.B1(_16243_),
    .Y(_16244_),
    .A2(_16238_),
    .A1(_16222_));
 sg13g2_nand2_1 _23208_ (.Y(_16245_),
    .A(\u_inv.f_next[66] ),
    .B(_14320_));
 sg13g2_nand2_1 _23209_ (.Y(_16246_),
    .A(\u_inv.f_next[65] ),
    .B(_14319_));
 sg13g2_nand2_1 _23210_ (.Y(_16247_),
    .A(\u_inv.f_next[64] ),
    .B(_14318_));
 sg13g2_o21ai_1 _23211_ (.B1(_16246_),
    .Y(_16248_),
    .A1(_15469_),
    .A2(_16247_));
 sg13g2_nor2_1 _23212_ (.A(_15180_),
    .B(_16245_),
    .Y(_16249_));
 sg13g2_a221oi_1 _23213_ (.B2(_16248_),
    .C1(_16249_),
    .B1(_16241_),
    .A1(\u_inv.f_next[67] ),
    .Y(_16250_),
    .A2(_14321_));
 sg13g2_nand2_1 _23214_ (.Y(_16251_),
    .A(\u_inv.f_next[70] ),
    .B(_14324_));
 sg13g2_nor2_1 _23215_ (.A(_14105_),
    .B(\u_inv.f_reg[69] ),
    .Y(_16252_));
 sg13g2_nor3_1 _23216_ (.A(_14106_),
    .B(\u_inv.f_reg[68] ),
    .C(_15177_),
    .Y(_16253_));
 sg13g2_o21ai_1 _23217_ (.B1(_15172_),
    .Y(_16254_),
    .A1(_16252_),
    .A2(_16253_));
 sg13g2_a21oi_1 _23218_ (.A1(_16251_),
    .A2(_16254_),
    .Y(_16255_),
    .B1(_15169_));
 sg13g2_a21oi_1 _23219_ (.A1(\u_inv.f_next[71] ),
    .A2(_14325_),
    .Y(_16256_),
    .B1(_16255_));
 sg13g2_o21ai_1 _23220_ (.B1(_16256_),
    .Y(_16257_),
    .A1(_16240_),
    .A2(_16250_));
 sg13g2_nor4_1 _23221_ (.A(_15486_),
    .B(_15488_),
    .C(_15493_),
    .D(_15495_),
    .Y(_16258_));
 sg13g2_nor2_1 _23222_ (.A(_15475_),
    .B(_15478_),
    .Y(_16259_));
 sg13g2_nand2_1 _23223_ (.Y(_16260_),
    .A(_15480_),
    .B(_15483_));
 sg13g2_nand4_1 _23224_ (.B(_15483_),
    .C(_16258_),
    .A(_15480_),
    .Y(_16261_),
    .D(_16259_));
 sg13g2_inv_1 _23225_ (.Y(_16262_),
    .A(_16261_));
 sg13g2_o21ai_1 _23226_ (.B1(_16262_),
    .Y(_16263_),
    .A1(_16244_),
    .A2(_16257_));
 sg13g2_nand2_1 _23227_ (.Y(_16264_),
    .A(\u_inv.f_next[78] ),
    .B(_14332_));
 sg13g2_nor2_1 _23228_ (.A(_15475_),
    .B(_16264_),
    .Y(_16265_));
 sg13g2_nand2_1 _23229_ (.Y(_16266_),
    .A(\u_inv.f_next[77] ),
    .B(_14331_));
 sg13g2_nor2_1 _23230_ (.A(_14098_),
    .B(\u_inv.f_reg[76] ),
    .Y(_16267_));
 sg13g2_nand2_1 _23231_ (.Y(_16268_),
    .A(_15480_),
    .B(_16267_));
 sg13g2_and2_1 _23232_ (.A(_16266_),
    .B(_16268_),
    .X(_16269_));
 sg13g2_nand2_1 _23233_ (.Y(_16270_),
    .A(\u_inv.f_next[74] ),
    .B(_14328_));
 sg13g2_nor2_1 _23234_ (.A(_14101_),
    .B(\u_inv.f_reg[73] ),
    .Y(_16271_));
 sg13g2_nand2_1 _23235_ (.Y(_16272_),
    .A(\u_inv.f_next[72] ),
    .B(_14326_));
 sg13g2_nor2_1 _23236_ (.A(_15495_),
    .B(_16272_),
    .Y(_16273_));
 sg13g2_o21ai_1 _23237_ (.B1(_15489_),
    .Y(_16274_),
    .A1(_16271_),
    .A2(_16273_));
 sg13g2_a21oi_1 _23238_ (.A1(_16270_),
    .A2(_16274_),
    .Y(_16275_),
    .B1(_15486_));
 sg13g2_a21oi_1 _23239_ (.A1(\u_inv.f_next[75] ),
    .A2(_14329_),
    .Y(_16276_),
    .B1(_16275_));
 sg13g2_o21ai_1 _23240_ (.B1(_16269_),
    .Y(_16277_),
    .A1(_16260_),
    .A2(_16276_));
 sg13g2_a221oi_1 _23241_ (.B2(_16277_),
    .C1(_16265_),
    .B1(_16259_),
    .A1(\u_inv.f_next[79] ),
    .Y(_16278_),
    .A2(_14333_));
 sg13g2_nor4_1 _23242_ (.A(_15510_),
    .B(_15513_),
    .C(_15516_),
    .D(_15518_),
    .Y(_16279_));
 sg13g2_inv_1 _23243_ (.Y(_16280_),
    .A(_16279_));
 sg13g2_a21oi_2 _23244_ (.B1(_16280_),
    .Y(_16281_),
    .A2(_16278_),
    .A1(_16263_));
 sg13g2_nor2_1 _23245_ (.A(_14092_),
    .B(\u_inv.f_reg[82] ),
    .Y(_16282_));
 sg13g2_nand2_1 _23246_ (.Y(_16283_),
    .A(\u_inv.f_next[81] ),
    .B(_14335_));
 sg13g2_nor2_1 _23247_ (.A(_14094_),
    .B(\u_inv.f_reg[80] ),
    .Y(_16284_));
 sg13g2_nand2_1 _23248_ (.Y(_16285_),
    .A(_15519_),
    .B(_16284_));
 sg13g2_a21oi_1 _23249_ (.A1(_16283_),
    .A2(_16285_),
    .Y(_16286_),
    .B1(_15513_));
 sg13g2_o21ai_1 _23250_ (.B1(_15511_),
    .Y(_16287_),
    .A1(_16282_),
    .A2(_16286_));
 sg13g2_o21ai_1 _23251_ (.B1(_16287_),
    .Y(_16288_),
    .A1(_14091_),
    .A2(\u_inv.f_reg[83] ));
 sg13g2_nand4_1 _23252_ (.B(_15153_),
    .C(_15163_),
    .A(_15151_),
    .Y(_16289_),
    .D(_15165_));
 sg13g2_inv_1 _23253_ (.Y(_16290_),
    .A(_16289_));
 sg13g2_o21ai_1 _23254_ (.B1(_16290_),
    .Y(_16291_),
    .A1(_16281_),
    .A2(_16288_));
 sg13g2_nand2_1 _23255_ (.Y(_16292_),
    .A(\u_inv.f_next[86] ),
    .B(_14340_));
 sg13g2_nand2_1 _23256_ (.Y(_16293_),
    .A(\u_inv.f_next[84] ),
    .B(_14338_));
 sg13g2_nand2b_1 _23257_ (.Y(_16294_),
    .B(_15163_),
    .A_N(_16293_));
 sg13g2_o21ai_1 _23258_ (.B1(_16294_),
    .Y(_16295_),
    .A1(_14089_),
    .A2(\u_inv.f_reg[85] ));
 sg13g2_nand2_1 _23259_ (.Y(_16296_),
    .A(_15153_),
    .B(_16295_));
 sg13g2_a21oi_1 _23260_ (.A1(_16292_),
    .A2(_16296_),
    .Y(_16297_),
    .B1(_15150_));
 sg13g2_a21oi_2 _23261_ (.B1(_16297_),
    .Y(_16298_),
    .A2(_14341_),
    .A1(\u_inv.f_next[87] ));
 sg13g2_nand2_1 _23262_ (.Y(_16299_),
    .A(_16291_),
    .B(_16298_));
 sg13g2_nand2_1 _23263_ (.Y(_16300_),
    .A(_15530_),
    .B(_15532_));
 sg13g2_nor3_1 _23264_ (.A(_15533_),
    .B(_15534_),
    .C(_16300_),
    .Y(_16301_));
 sg13g2_nand2_1 _23265_ (.Y(_16302_),
    .A(_15538_),
    .B(_15539_));
 sg13g2_inv_1 _23266_ (.Y(_16303_),
    .A(_16302_));
 sg13g2_nor2_1 _23267_ (.A(_15545_),
    .B(_15547_),
    .Y(_16304_));
 sg13g2_inv_1 _23268_ (.Y(_16305_),
    .A(_16304_));
 sg13g2_and3_1 _23269_ (.X(_16306_),
    .A(_16301_),
    .B(_16303_),
    .C(_16304_));
 sg13g2_inv_1 _23270_ (.Y(_16307_),
    .A(_16306_));
 sg13g2_a21oi_2 _23271_ (.B1(_16307_),
    .Y(_16308_),
    .A2(_16298_),
    .A1(_16291_));
 sg13g2_nand2_1 _23272_ (.Y(_16309_),
    .A(_16299_),
    .B(_16306_));
 sg13g2_and3_1 _23273_ (.X(_16310_),
    .A(\u_inv.f_next[90] ),
    .B(_14344_),
    .C(_15538_));
 sg13g2_a21oi_1 _23274_ (.A1(\u_inv.f_next[91] ),
    .A2(_14345_),
    .Y(_16311_),
    .B1(_16310_));
 sg13g2_nand2_1 _23275_ (.Y(_16312_),
    .A(\u_inv.f_next[88] ),
    .B(_14342_));
 sg13g2_nor2_1 _23276_ (.A(_15545_),
    .B(_16312_),
    .Y(_16313_));
 sg13g2_a21o_2 _23277_ (.A2(_14343_),
    .A1(\u_inv.f_next[89] ),
    .B1(_16313_),
    .X(_16314_));
 sg13g2_a221oi_1 _23278_ (.B2(_16314_),
    .C1(_16310_),
    .B1(_16303_),
    .A1(\u_inv.f_next[91] ),
    .Y(_16315_),
    .A2(_14345_));
 sg13g2_nand2b_1 _23279_ (.Y(_16316_),
    .B(_16301_),
    .A_N(_16315_));
 sg13g2_nor2_1 _23280_ (.A(_14079_),
    .B(\u_inv.f_reg[95] ),
    .Y(_16317_));
 sg13g2_nor2_1 _23281_ (.A(_14080_),
    .B(\u_inv.f_reg[94] ),
    .Y(_16318_));
 sg13g2_a21oi_1 _23282_ (.A1(_15530_),
    .A2(_16318_),
    .Y(_16319_),
    .B1(_16317_));
 sg13g2_nand2_1 _23283_ (.Y(_16320_),
    .A(\u_inv.f_next[93] ),
    .B(_14347_));
 sg13g2_nand2_1 _23284_ (.Y(_16321_),
    .A(\u_inv.f_next[92] ),
    .B(_14346_));
 sg13g2_o21ai_1 _23285_ (.B1(_16320_),
    .Y(_16322_),
    .A1(_15534_),
    .A2(_16321_));
 sg13g2_nand2b_1 _23286_ (.Y(_16323_),
    .B(_16322_),
    .A_N(_16300_));
 sg13g2_nand3_1 _23287_ (.B(_16319_),
    .C(_16323_),
    .A(_16316_),
    .Y(_16324_));
 sg13g2_inv_1 _23288_ (.Y(_16325_),
    .A(_16324_));
 sg13g2_nor2_1 _23289_ (.A(_15133_),
    .B(_15135_),
    .Y(_16326_));
 sg13g2_nor2_1 _23290_ (.A(_15127_),
    .B(_15130_),
    .Y(_16327_));
 sg13g2_nor2_1 _23291_ (.A(_15123_),
    .B(_15124_),
    .Y(_16328_));
 sg13g2_nor2_1 _23292_ (.A(_15563_),
    .B(_15564_),
    .Y(_16329_));
 sg13g2_and4_1 _23293_ (.A(_16326_),
    .B(_16327_),
    .C(_16328_),
    .D(_16329_),
    .X(_16330_));
 sg13g2_o21ai_1 _23294_ (.B1(_16330_),
    .Y(_16331_),
    .A1(_16308_),
    .A2(_16324_));
 sg13g2_nor2_1 _23295_ (.A(_14074_),
    .B(\u_inv.f_reg[100] ),
    .Y(_16332_));
 sg13g2_nand2_1 _23296_ (.Y(_16333_),
    .A(\u_inv.f_next[98] ),
    .B(_14352_));
 sg13g2_o21ai_1 _23297_ (.B1(_15132_),
    .Y(_16334_),
    .A1(_15133_),
    .A2(_16333_));
 sg13g2_nor2_1 _23298_ (.A(_14073_),
    .B(\u_inv.f_reg[101] ),
    .Y(_16335_));
 sg13g2_nand2_1 _23299_ (.Y(_16336_),
    .A(\u_inv.f_next[96] ),
    .B(_14350_));
 sg13g2_nor2_1 _23300_ (.A(_15563_),
    .B(_16336_),
    .Y(_16337_));
 sg13g2_a21oi_1 _23301_ (.A1(\u_inv.f_next[97] ),
    .A2(_14351_),
    .Y(_16338_),
    .B1(_16337_));
 sg13g2_nor2b_1 _23302_ (.A(_16338_),
    .B_N(_16326_),
    .Y(_16339_));
 sg13g2_o21ai_1 _23303_ (.B1(_16327_),
    .Y(_16340_),
    .A1(_16334_),
    .A2(_16339_));
 sg13g2_a21oi_1 _23304_ (.A1(_15128_),
    .A2(_16332_),
    .Y(_16341_),
    .B1(_16335_));
 sg13g2_nand2_1 _23305_ (.Y(_16342_),
    .A(_16340_),
    .B(_16341_));
 sg13g2_nand2_1 _23306_ (.Y(_16343_),
    .A(\u_inv.f_next[102] ),
    .B(_14356_));
 sg13g2_nor2_1 _23307_ (.A(_15123_),
    .B(_16343_),
    .Y(_16344_));
 sg13g2_a221oi_1 _23308_ (.B2(_16342_),
    .C1(_16344_),
    .B1(_16328_),
    .A1(\u_inv.f_next[103] ),
    .Y(_16345_),
    .A2(_14357_));
 sg13g2_nand2_1 _23309_ (.Y(_16346_),
    .A(_16331_),
    .B(_16345_));
 sg13g2_or4_1 _23310_ (.A(_15584_),
    .B(_15587_),
    .C(_15591_),
    .D(_15592_),
    .X(_16347_));
 sg13g2_nor2_1 _23311_ (.A(_15571_),
    .B(_15575_),
    .Y(_16348_));
 sg13g2_nand2_1 _23312_ (.Y(_16349_),
    .A(_15578_),
    .B(_15581_));
 sg13g2_or4_1 _23313_ (.A(_15571_),
    .B(_15575_),
    .C(_16347_),
    .D(_16349_),
    .X(_16350_));
 sg13g2_a21oi_2 _23314_ (.B1(_16350_),
    .Y(_16351_),
    .A2(_16345_),
    .A1(_16331_));
 sg13g2_a21o_1 _23315_ (.A2(_16345_),
    .A1(_16331_),
    .B1(_16350_),
    .X(_16352_));
 sg13g2_nand2_1 _23316_ (.Y(_16353_),
    .A(\u_inv.f_next[107] ),
    .B(_14361_));
 sg13g2_nor2_1 _23317_ (.A(_14068_),
    .B(\u_inv.f_reg[106] ),
    .Y(_16354_));
 sg13g2_nand2_1 _23318_ (.Y(_16355_),
    .A(\u_inv.f_next[105] ),
    .B(_14359_));
 sg13g2_nand2_1 _23319_ (.Y(_16356_),
    .A(\u_inv.f_next[104] ),
    .B(_14358_));
 sg13g2_o21ai_1 _23320_ (.B1(_16355_),
    .Y(_16357_),
    .A1(_15592_),
    .A2(_16356_));
 sg13g2_a21oi_1 _23321_ (.A1(_15588_),
    .A2(_16357_),
    .Y(_16358_),
    .B1(_16354_));
 sg13g2_o21ai_1 _23322_ (.B1(_16353_),
    .Y(_16359_),
    .A1(_15584_),
    .A2(_16358_));
 sg13g2_nor2b_1 _23323_ (.A(_16349_),
    .B_N(_16359_),
    .Y(_16360_));
 sg13g2_nand2_1 _23324_ (.Y(_16361_),
    .A(\u_inv.f_next[108] ),
    .B(_14362_));
 sg13g2_nand2_1 _23325_ (.Y(_16362_),
    .A(\u_inv.f_next[109] ),
    .B(_14363_));
 sg13g2_o21ai_1 _23326_ (.B1(_16362_),
    .Y(_16363_),
    .A1(_15577_),
    .A2(_16361_));
 sg13g2_o21ai_1 _23327_ (.B1(_16348_),
    .Y(_16364_),
    .A1(_16360_),
    .A2(_16363_));
 sg13g2_nor2_1 _23328_ (.A(_14064_),
    .B(\u_inv.f_reg[110] ),
    .Y(_16365_));
 sg13g2_o21ai_1 _23329_ (.B1(_16364_),
    .Y(_16366_),
    .A1(_14063_),
    .A2(\u_inv.f_reg[111] ));
 sg13g2_a21o_2 _23330_ (.A2(_16365_),
    .A1(_15572_),
    .B1(_16366_),
    .X(_16367_));
 sg13g2_inv_1 _23331_ (.Y(_16368_),
    .A(_16367_));
 sg13g2_nor2_1 _23332_ (.A(_16351_),
    .B(_16367_),
    .Y(_16369_));
 sg13g2_nor4_1 _23333_ (.A(_15611_),
    .B(_15614_),
    .C(_15616_),
    .D(_15618_),
    .Y(_16370_));
 sg13g2_nand3_1 _23334_ (.B(_15624_),
    .C(_15627_),
    .A(_15622_),
    .Y(_16371_));
 sg13g2_nor2_1 _23335_ (.A(_15628_),
    .B(_16371_),
    .Y(_16372_));
 sg13g2_and2_1 _23336_ (.A(_16370_),
    .B(_16372_),
    .X(_16373_));
 sg13g2_nor2_1 _23337_ (.A(_15641_),
    .B(_15644_),
    .Y(_16374_));
 sg13g2_nand3_1 _23338_ (.B(_15652_),
    .C(_16374_),
    .A(_15650_),
    .Y(_16375_));
 sg13g2_and2_1 _23339_ (.A(_15631_),
    .B(_15633_),
    .X(_16376_));
 sg13g2_nand3_1 _23340_ (.B(_15638_),
    .C(_16376_),
    .A(_15636_),
    .Y(_16377_));
 sg13g2_nor2_1 _23341_ (.A(_16375_),
    .B(_16377_),
    .Y(_16378_));
 sg13g2_inv_1 _23342_ (.Y(_16379_),
    .A(_16378_));
 sg13g2_and2_1 _23343_ (.A(_16373_),
    .B(_16378_),
    .X(_16380_));
 sg13g2_o21ai_1 _23344_ (.B1(_16380_),
    .Y(_16381_),
    .A1(_16351_),
    .A2(_16367_));
 sg13g2_nor2_1 _23345_ (.A(_14056_),
    .B(\u_inv.f_reg[118] ),
    .Y(_16382_));
 sg13g2_nor2_1 _23346_ (.A(_14057_),
    .B(\u_inv.f_reg[117] ),
    .Y(_16383_));
 sg13g2_nand2_1 _23347_ (.Y(_16384_),
    .A(\u_inv.f_next[116] ),
    .B(_14370_));
 sg13g2_nor2_1 _23348_ (.A(_15637_),
    .B(_16384_),
    .Y(_16385_));
 sg13g2_or2_1 _23349_ (.X(_16386_),
    .B(_16385_),
    .A(_16383_));
 sg13g2_nor2_1 _23350_ (.A(_14059_),
    .B(\u_inv.f_reg[115] ),
    .Y(_16387_));
 sg13g2_nor2_1 _23351_ (.A(_14060_),
    .B(\u_inv.f_reg[114] ),
    .Y(_16388_));
 sg13g2_nand2_1 _23352_ (.Y(_16389_),
    .A(\u_inv.f_next[113] ),
    .B(_14367_));
 sg13g2_nand2_1 _23353_ (.Y(_16390_),
    .A(\u_inv.f_next[112] ),
    .B(_14366_));
 sg13g2_o21ai_1 _23354_ (.B1(_16389_),
    .Y(_16391_),
    .A1(_15651_),
    .A2(_16390_));
 sg13g2_a221oi_1 _23355_ (.B2(_16374_),
    .C1(_16387_),
    .B1(_16391_),
    .A1(_15642_),
    .Y(_16392_),
    .A2(_16388_));
 sg13g2_inv_1 _23356_ (.Y(_16393_),
    .A(_16392_));
 sg13g2_a22oi_1 _23357_ (.Y(_16394_),
    .B1(_16376_),
    .B2(_16386_),
    .A2(_14373_),
    .A1(\u_inv.f_next[119] ));
 sg13g2_o21ai_1 _23358_ (.B1(_16394_),
    .Y(_16395_),
    .A1(_16377_),
    .A2(_16392_));
 sg13g2_a21oi_1 _23359_ (.A1(_15631_),
    .A2(_16382_),
    .Y(_16396_),
    .B1(_16395_));
 sg13g2_nand2b_1 _23360_ (.Y(_16397_),
    .B(_16373_),
    .A_N(_16396_));
 sg13g2_nor2_1 _23361_ (.A(_14049_),
    .B(\u_inv.f_reg[125] ),
    .Y(_16398_));
 sg13g2_nand2_1 _23362_ (.Y(_16399_),
    .A(\u_inv.f_next[124] ),
    .B(_14378_));
 sg13g2_nor2_1 _23363_ (.A(_15616_),
    .B(_16399_),
    .Y(_16400_));
 sg13g2_nand2_1 _23364_ (.Y(_16401_),
    .A(\u_inv.f_next[126] ),
    .B(_14380_));
 sg13g2_o21ai_1 _23365_ (.B1(_15613_),
    .Y(_16402_),
    .A1(_16398_),
    .A2(_16400_));
 sg13g2_a21oi_1 _23366_ (.A1(_16401_),
    .A2(_16402_),
    .Y(_16403_),
    .B1(_15611_));
 sg13g2_nor2_1 _23367_ (.A(_14052_),
    .B(\u_inv.f_reg[122] ),
    .Y(_16404_));
 sg13g2_nand2_1 _23368_ (.Y(_16405_),
    .A(\u_inv.f_next[121] ),
    .B(_14375_));
 sg13g2_nor2_1 _23369_ (.A(_14054_),
    .B(\u_inv.f_reg[120] ),
    .Y(_16406_));
 sg13g2_nand2_1 _23370_ (.Y(_16407_),
    .A(\u_inv.f_next[120] ),
    .B(_14374_));
 sg13g2_o21ai_1 _23371_ (.B1(_16405_),
    .Y(_16408_),
    .A1(_15628_),
    .A2(_16407_));
 sg13g2_and2_1 _23372_ (.A(_15624_),
    .B(_16408_),
    .X(_16409_));
 sg13g2_o21ai_1 _23373_ (.B1(_15622_),
    .Y(_16410_),
    .A1(_16404_),
    .A2(_16409_));
 sg13g2_o21ai_1 _23374_ (.B1(_16410_),
    .Y(_16411_),
    .A1(_14051_),
    .A2(\u_inv.f_reg[123] ));
 sg13g2_a221oi_1 _23375_ (.B2(_16411_),
    .C1(_16403_),
    .B1(_16370_),
    .A1(\u_inv.f_next[127] ),
    .Y(_16412_),
    .A2(_14381_));
 sg13g2_and2_1 _23376_ (.A(_16397_),
    .B(_16412_),
    .X(_16413_));
 sg13g2_nand2_1 _23377_ (.Y(_16414_),
    .A(_16381_),
    .B(_16413_));
 sg13g2_nand4_1 _23378_ (.B(_15726_),
    .C(_15728_),
    .A(_15724_),
    .Y(_16415_),
    .D(_15731_));
 sg13g2_nand4_1 _23379_ (.B(_15714_),
    .C(_15718_),
    .A(_15712_),
    .Y(_16416_),
    .D(_15720_));
 sg13g2_nor2_1 _23380_ (.A(_16415_),
    .B(_16416_),
    .Y(_16417_));
 sg13g2_nor2_1 _23381_ (.A(_15685_),
    .B(_15687_),
    .Y(_16418_));
 sg13g2_nand3_1 _23382_ (.B(_15693_),
    .C(_16418_),
    .A(_15691_),
    .Y(_16419_));
 sg13g2_or4_1 _23383_ (.A(_15698_),
    .B(_15702_),
    .C(_15704_),
    .D(_15706_),
    .X(_16420_));
 sg13g2_nor2_2 _23384_ (.A(_16419_),
    .B(_16420_),
    .Y(_16421_));
 sg13g2_nand2_1 _23385_ (.Y(_16422_),
    .A(_16417_),
    .B(_16421_));
 sg13g2_a21o_2 _23386_ (.A2(_16413_),
    .A1(_16381_),
    .B1(_16422_),
    .X(_16423_));
 sg13g2_nor2_1 _23387_ (.A(_14046_),
    .B(\u_inv.f_reg[128] ),
    .Y(_16424_));
 sg13g2_nor2_1 _23388_ (.A(_14044_),
    .B(\u_inv.f_reg[130] ),
    .Y(_16425_));
 sg13g2_nand2_1 _23389_ (.Y(_16426_),
    .A(\u_inv.f_next[129] ),
    .B(_14383_));
 sg13g2_nand2_1 _23390_ (.Y(_16427_),
    .A(_15728_),
    .B(_16424_));
 sg13g2_a21oi_1 _23391_ (.A1(_16426_),
    .A2(_16427_),
    .Y(_16428_),
    .B1(_15723_));
 sg13g2_o21ai_1 _23392_ (.B1(_15726_),
    .Y(_16429_),
    .A1(_16425_),
    .A2(_16428_));
 sg13g2_o21ai_1 _23393_ (.B1(_16429_),
    .Y(_16430_),
    .A1(_14043_),
    .A2(\u_inv.f_reg[131] ));
 sg13g2_nand2b_1 _23394_ (.Y(_16431_),
    .B(_16430_),
    .A_N(_16416_));
 sg13g2_nor2_1 _23395_ (.A(_14040_),
    .B(\u_inv.f_reg[134] ),
    .Y(_16432_));
 sg13g2_nand2_1 _23396_ (.Y(_16433_),
    .A(\u_inv.f_next[134] ),
    .B(_14388_));
 sg13g2_nand2_1 _23397_ (.Y(_16434_),
    .A(\u_inv.f_next[132] ),
    .B(_14386_));
 sg13g2_nand2b_1 _23398_ (.Y(_16435_),
    .B(_15718_),
    .A_N(_16434_));
 sg13g2_nand2_1 _23399_ (.Y(_16436_),
    .A(\u_inv.f_next[133] ),
    .B(_14387_));
 sg13g2_and2_1 _23400_ (.A(_16435_),
    .B(_16436_),
    .X(_16437_));
 sg13g2_inv_1 _23401_ (.Y(_16438_),
    .A(_16437_));
 sg13g2_a21o_1 _23402_ (.A2(_16438_),
    .A1(_15712_),
    .B1(_16432_),
    .X(_16439_));
 sg13g2_o21ai_1 _23403_ (.B1(_16431_),
    .Y(_16440_),
    .A1(_14039_),
    .A2(\u_inv.f_reg[135] ));
 sg13g2_a21o_2 _23404_ (.A2(_16439_),
    .A1(_15714_),
    .B1(_16440_),
    .X(_16441_));
 sg13g2_nand2_1 _23405_ (.Y(_16442_),
    .A(\u_inv.f_next[138] ),
    .B(_14392_));
 sg13g2_nor2_1 _23406_ (.A(_14037_),
    .B(\u_inv.f_reg[137] ),
    .Y(_16443_));
 sg13g2_nand2_1 _23407_ (.Y(_16444_),
    .A(\u_inv.f_next[136] ),
    .B(_14390_));
 sg13g2_nor2_1 _23408_ (.A(_15702_),
    .B(_16444_),
    .Y(_16445_));
 sg13g2_o21ai_1 _23409_ (.B1(_15707_),
    .Y(_16446_),
    .A1(_16443_),
    .A2(_16445_));
 sg13g2_a21oi_1 _23410_ (.A1(_16442_),
    .A2(_16446_),
    .Y(_16447_),
    .B1(_15704_));
 sg13g2_a21oi_1 _23411_ (.A1(\u_inv.f_next[139] ),
    .A2(_14393_),
    .Y(_16448_),
    .B1(_16447_));
 sg13g2_nor2_1 _23412_ (.A(_14033_),
    .B(\u_inv.f_reg[141] ),
    .Y(_16449_));
 sg13g2_nand2_1 _23413_ (.Y(_16450_),
    .A(\u_inv.f_next[140] ),
    .B(_14394_));
 sg13g2_nor2_1 _23414_ (.A(_15690_),
    .B(_16450_),
    .Y(_16451_));
 sg13g2_or2_1 _23415_ (.X(_16452_),
    .B(_16451_),
    .A(_16449_));
 sg13g2_nand2_1 _23416_ (.Y(_16453_),
    .A(\u_inv.f_next[142] ),
    .B(_14396_));
 sg13g2_nor2_1 _23417_ (.A(_15685_),
    .B(_16453_),
    .Y(_16454_));
 sg13g2_a221oi_1 _23418_ (.B2(_16452_),
    .C1(_16454_),
    .B1(_16418_),
    .A1(\u_inv.f_next[143] ),
    .Y(_16455_),
    .A2(_14397_));
 sg13g2_o21ai_1 _23419_ (.B1(_16455_),
    .Y(_16456_),
    .A1(_16419_),
    .A2(_16448_));
 sg13g2_a21oi_2 _23420_ (.B1(_16456_),
    .Y(_16457_),
    .A2(_16441_),
    .A1(_16421_));
 sg13g2_and2_1 _23421_ (.A(_16059_),
    .B(_16457_),
    .X(_16458_));
 sg13g2_a21o_2 _23422_ (.A2(_16458_),
    .A1(_16423_),
    .B1(_16063_),
    .X(_16459_));
 sg13g2_nor2_1 _23423_ (.A(_14921_),
    .B(_14922_),
    .Y(_16460_));
 sg13g2_inv_1 _23424_ (.Y(_16461_),
    .A(_16460_));
 sg13g2_nand3_1 _23425_ (.B(_14917_),
    .C(_16460_),
    .A(_14915_),
    .Y(_16462_));
 sg13g2_and2_1 _23426_ (.A(net5623),
    .B(net5622),
    .X(_16463_));
 sg13g2_nand2_1 _23427_ (.Y(_16464_),
    .A(net5623),
    .B(net5622));
 sg13g2_or2_1 _23428_ (.X(_16465_),
    .B(_14932_),
    .A(_14930_));
 sg13g2_nor3_1 _23429_ (.A(_16462_),
    .B(_16464_),
    .C(_16465_),
    .Y(_16466_));
 sg13g2_nor4_1 _23430_ (.A(_14935_),
    .B(_14937_),
    .C(_14940_),
    .D(_14943_),
    .Y(_16467_));
 sg13g2_nor4_1 _23431_ (.A(_14947_),
    .B(_14949_),
    .C(_14954_),
    .D(_14956_),
    .Y(_16468_));
 sg13g2_and2_1 _23432_ (.A(_16467_),
    .B(_16468_),
    .X(_16469_));
 sg13g2_and2_1 _23433_ (.A(_16466_),
    .B(_16469_),
    .X(_16470_));
 sg13g2_nor2_1 _23434_ (.A(_14993_),
    .B(_14996_),
    .Y(_16471_));
 sg13g2_and2_1 _23435_ (.A(_15006_),
    .B(_15008_),
    .X(_16472_));
 sg13g2_nand2_1 _23436_ (.Y(_16473_),
    .A(_15011_),
    .B(_15013_));
 sg13g2_nand4_1 _23437_ (.B(_15002_),
    .C(_16471_),
    .A(_14999_),
    .Y(_16474_),
    .D(_16472_));
 sg13g2_nor2_1 _23438_ (.A(_16473_),
    .B(_16474_),
    .Y(_16475_));
 sg13g2_and2_1 _23439_ (.A(_14966_),
    .B(_14968_),
    .X(_16476_));
 sg13g2_and3_2 _23440_ (.X(_16477_),
    .A(_14971_),
    .B(_14973_),
    .C(_16476_));
 sg13g2_nand2_1 _23441_ (.Y(_16478_),
    .A(_15766_),
    .B(_15768_));
 sg13g2_or3_1 _23442_ (.A(_14977_),
    .B(_14979_),
    .C(_16478_),
    .X(_16479_));
 sg13g2_inv_1 _23443_ (.Y(_16480_),
    .A(_16479_));
 sg13g2_nand3_1 _23444_ (.B(_16477_),
    .C(_16480_),
    .A(_16475_),
    .Y(_16481_));
 sg13g2_nand4_1 _23445_ (.B(_16475_),
    .C(_16477_),
    .A(_16470_),
    .Y(_16482_),
    .D(_16480_));
 sg13g2_a221oi_1 _23446_ (.B2(_16458_),
    .C1(_16482_),
    .B1(_16423_),
    .A1(_16059_),
    .Y(_16483_),
    .A2(_16062_));
 sg13g2_nand2_1 _23447_ (.Y(_16484_),
    .A(\u_inv.f_next[162] ),
    .B(_14416_));
 sg13g2_nand3_1 _23448_ (.B(_14414_),
    .C(_15768_),
    .A(\u_inv.f_next[160] ),
    .Y(_16485_));
 sg13g2_nand2_1 _23449_ (.Y(_16486_),
    .A(\u_inv.f_next[161] ),
    .B(_14415_));
 sg13g2_and2_1 _23450_ (.A(_16485_),
    .B(_16486_),
    .X(_16487_));
 sg13g2_o21ai_1 _23451_ (.B1(_16484_),
    .Y(_16488_),
    .A1(_14979_),
    .A2(_16487_));
 sg13g2_nand2b_1 _23452_ (.Y(_16489_),
    .B(_16488_),
    .A_N(_14977_));
 sg13g2_o21ai_1 _23453_ (.B1(_16489_),
    .Y(_16490_),
    .A1(_14011_),
    .A2(\u_inv.f_reg[163] ));
 sg13g2_nor2_1 _23454_ (.A(_14009_),
    .B(\u_inv.f_reg[165] ),
    .Y(_16491_));
 sg13g2_nand2_1 _23455_ (.Y(_16492_),
    .A(\u_inv.f_next[164] ),
    .B(_14418_));
 sg13g2_nor2_1 _23456_ (.A(_14972_),
    .B(_16492_),
    .Y(_16493_));
 sg13g2_o21ai_1 _23457_ (.B1(_16476_),
    .Y(_16494_),
    .A1(_16491_),
    .A2(_16493_));
 sg13g2_nor2_1 _23458_ (.A(_14008_),
    .B(\u_inv.f_reg[166] ),
    .Y(_16495_));
 sg13g2_nor2_1 _23459_ (.A(_14007_),
    .B(\u_inv.f_reg[167] ),
    .Y(_16496_));
 sg13g2_a221oi_1 _23460_ (.B2(_14966_),
    .C1(_16496_),
    .B1(_16495_),
    .A1(_16477_),
    .Y(_16497_),
    .A2(_16490_));
 sg13g2_nand2_1 _23461_ (.Y(_16498_),
    .A(_16494_),
    .B(_16497_));
 sg13g2_nand2_1 _23462_ (.Y(_16499_),
    .A(_16475_),
    .B(_16498_));
 sg13g2_nand2_1 _23463_ (.Y(_16500_),
    .A(\u_inv.f_next[173] ),
    .B(_14427_));
 sg13g2_nor2_1 _23464_ (.A(_14002_),
    .B(\u_inv.f_reg[172] ),
    .Y(_16501_));
 sg13g2_nand2_1 _23465_ (.Y(_16502_),
    .A(_14999_),
    .B(_16501_));
 sg13g2_nand2_1 _23466_ (.Y(_16503_),
    .A(_16500_),
    .B(_16502_));
 sg13g2_nand2_1 _23467_ (.Y(_16504_),
    .A(\u_inv.f_next[174] ),
    .B(_14428_));
 sg13g2_or2_1 _23468_ (.X(_16505_),
    .B(_16504_),
    .A(_14993_));
 sg13g2_a22oi_1 _23469_ (.Y(_16506_),
    .B1(_16471_),
    .B2(_16503_),
    .A2(_14429_),
    .A1(\u_inv.f_next[175] ));
 sg13g2_nand3_1 _23470_ (.B(_14422_),
    .C(_15011_),
    .A(\u_inv.f_next[168] ),
    .Y(_16507_));
 sg13g2_o21ai_1 _23471_ (.B1(_16507_),
    .Y(_16508_),
    .A1(_14005_),
    .A2(\u_inv.f_reg[169] ));
 sg13g2_nand2_1 _23472_ (.Y(_16509_),
    .A(\u_inv.f_next[170] ),
    .B(_14424_));
 sg13g2_a22oi_1 _23473_ (.Y(_16510_),
    .B1(_16472_),
    .B2(_16508_),
    .A2(_14425_),
    .A1(\u_inv.f_next[171] ));
 sg13g2_o21ai_1 _23474_ (.B1(_16510_),
    .Y(_16511_),
    .A1(_15005_),
    .A2(_16509_));
 sg13g2_inv_1 _23475_ (.Y(_16512_),
    .A(_16511_));
 sg13g2_nand4_1 _23476_ (.B(_15002_),
    .C(_16471_),
    .A(_14999_),
    .Y(_16513_),
    .D(_16511_));
 sg13g2_nand4_1 _23477_ (.B(_16505_),
    .C(_16506_),
    .A(_16499_),
    .Y(_16514_),
    .D(_16513_));
 sg13g2_nor2_1 _23478_ (.A(_13987_),
    .B(\u_inv.f_reg[187] ),
    .Y(_16515_));
 sg13g2_nor2_1 _23479_ (.A(_13988_),
    .B(\u_inv.f_reg[186] ),
    .Y(_16516_));
 sg13g2_nand3b_1 _23480_ (.B(\u_inv.f_next[184] ),
    .C(_14438_),
    .Y(_16517_),
    .A_N(_14930_));
 sg13g2_inv_1 _23481_ (.Y(_16518_),
    .A(_16517_));
 sg13g2_o21ai_1 _23482_ (.B1(_16517_),
    .Y(_16519_),
    .A1(_13989_),
    .A2(\u_inv.f_reg[185] ));
 sg13g2_a21o_1 _23483_ (.A2(_16519_),
    .A1(_14927_),
    .B1(_16516_),
    .X(_16520_));
 sg13g2_a21oi_1 _23484_ (.A1(net5623),
    .A2(_16520_),
    .Y(_16521_),
    .B1(_16515_));
 sg13g2_nand3_1 _23485_ (.B(_14442_),
    .C(_14923_),
    .A(\u_inv.f_next[188] ),
    .Y(_16522_));
 sg13g2_nand2_1 _23486_ (.Y(_16523_),
    .A(\u_inv.f_next[189] ),
    .B(_14443_));
 sg13g2_and2_1 _23487_ (.A(_16522_),
    .B(_16523_),
    .X(_16524_));
 sg13g2_nor3_1 _23488_ (.A(_14914_),
    .B(_14918_),
    .C(_16524_),
    .Y(_16525_));
 sg13g2_nand2_1 _23489_ (.Y(_16526_),
    .A(\u_inv.f_next[190] ),
    .B(_14444_));
 sg13g2_nor2_1 _23490_ (.A(_13992_),
    .B(\u_inv.f_reg[182] ),
    .Y(_16527_));
 sg13g2_nand2_1 _23491_ (.Y(_16528_),
    .A(\u_inv.f_next[180] ),
    .B(_14434_));
 sg13g2_or2_1 _23492_ (.X(_16529_),
    .B(_16528_),
    .A(_14940_));
 sg13g2_o21ai_1 _23493_ (.B1(_16529_),
    .Y(_16530_),
    .A1(_13993_),
    .A2(\u_inv.f_reg[181] ));
 sg13g2_a21oi_1 _23494_ (.A1(_14938_),
    .A2(_16530_),
    .Y(_16531_),
    .B1(_16527_));
 sg13g2_nand2_1 _23495_ (.Y(_16532_),
    .A(\u_inv.f_next[176] ),
    .B(_14430_));
 sg13g2_nand2_1 _23496_ (.Y(_16533_),
    .A(\u_inv.f_next[178] ),
    .B(_14432_));
 sg13g2_nor2_1 _23497_ (.A(_13997_),
    .B(\u_inv.f_reg[177] ),
    .Y(_16534_));
 sg13g2_nor2_1 _23498_ (.A(_14956_),
    .B(_16532_),
    .Y(_16535_));
 sg13g2_o21ai_1 _23499_ (.B1(_14950_),
    .Y(_16536_),
    .A1(_16534_),
    .A2(_16535_));
 sg13g2_a21oi_1 _23500_ (.A1(_16533_),
    .A2(_16536_),
    .Y(_16537_),
    .B1(_14947_));
 sg13g2_a21oi_1 _23501_ (.A1(\u_inv.f_next[179] ),
    .A2(_14433_),
    .Y(_16538_),
    .B1(_16537_));
 sg13g2_nor2b_1 _23502_ (.A(_16538_),
    .B_N(_16467_),
    .Y(_16539_));
 sg13g2_nand2_1 _23503_ (.Y(_16540_),
    .A(\u_inv.f_next[183] ),
    .B(_14437_));
 sg13g2_o21ai_1 _23504_ (.B1(_16540_),
    .Y(_16541_),
    .A1(_14935_),
    .A2(_16531_));
 sg13g2_nor2_2 _23505_ (.A(_16539_),
    .B(_16541_),
    .Y(_16542_));
 sg13g2_inv_1 _23506_ (.Y(_16543_),
    .A(_16542_));
 sg13g2_a21oi_1 _23507_ (.A1(\u_inv.f_next[191] ),
    .A2(_14445_),
    .Y(_16544_),
    .B1(_16525_));
 sg13g2_o21ai_1 _23508_ (.B1(_16544_),
    .Y(_16545_),
    .A1(_16462_),
    .A2(_16521_));
 sg13g2_a221oi_1 _23509_ (.B2(_16466_),
    .C1(_16545_),
    .B1(_16543_),
    .A1(_16470_),
    .Y(_16546_),
    .A2(_16514_));
 sg13g2_o21ai_1 _23510_ (.B1(_16546_),
    .Y(_16547_),
    .A1(_14914_),
    .A2(_16526_));
 sg13g2_nor2_1 _23511_ (.A(_16483_),
    .B(_16547_),
    .Y(_16548_));
 sg13g2_nor2_1 _23512_ (.A(_15785_),
    .B(_15787_),
    .Y(_16549_));
 sg13g2_nand3_1 _23513_ (.B(_15794_),
    .C(_16549_),
    .A(_15792_),
    .Y(_16550_));
 sg13g2_inv_1 _23514_ (.Y(_16551_),
    .A(_16550_));
 sg13g2_or2_1 _23515_ (.X(_16552_),
    .B(_15776_),
    .A(_15775_));
 sg13g2_nand2_1 _23516_ (.Y(_16553_),
    .A(_15778_),
    .B(_15781_));
 sg13g2_nor3_1 _23517_ (.A(_16550_),
    .B(_16552_),
    .C(_16553_),
    .Y(_16554_));
 sg13g2_nand2_1 _23518_ (.Y(_16555_),
    .A(_15804_),
    .B(_15808_));
 sg13g2_or3_1 _23519_ (.A(_15799_),
    .B(_15801_),
    .C(_16555_),
    .X(_16556_));
 sg13g2_nand4_1 _23520_ (.B(_15813_),
    .C(_15816_),
    .A(_15812_),
    .Y(_16557_),
    .D(_15818_));
 sg13g2_nor2_1 _23521_ (.A(_16556_),
    .B(_16557_),
    .Y(_16558_));
 sg13g2_nand2_1 _23522_ (.Y(_16559_),
    .A(_16554_),
    .B(_16558_));
 sg13g2_inv_1 _23523_ (.Y(_16560_),
    .A(_16559_));
 sg13g2_o21ai_1 _23524_ (.B1(_16560_),
    .Y(_16561_),
    .A1(_16483_),
    .A2(_16547_));
 sg13g2_nand2_1 _23525_ (.Y(_16562_),
    .A(\u_inv.f_next[197] ),
    .B(_14451_));
 sg13g2_nor2_1 _23526_ (.A(_13978_),
    .B(\u_inv.f_reg[196] ),
    .Y(_16563_));
 sg13g2_nor2_1 _23527_ (.A(_13979_),
    .B(\u_inv.f_reg[195] ),
    .Y(_16564_));
 sg13g2_nor2_1 _23528_ (.A(_13980_),
    .B(\u_inv.f_reg[194] ),
    .Y(_16565_));
 sg13g2_nor2_1 _23529_ (.A(_13981_),
    .B(\u_inv.f_reg[193] ),
    .Y(_16566_));
 sg13g2_nand2_1 _23530_ (.Y(_16567_),
    .A(\u_inv.f_next[192] ),
    .B(_14446_));
 sg13g2_nor2_1 _23531_ (.A(_15791_),
    .B(_16567_),
    .Y(_16568_));
 sg13g2_or2_1 _23532_ (.X(_16569_),
    .B(_16568_),
    .A(_16566_));
 sg13g2_a221oi_1 _23533_ (.B2(_16549_),
    .C1(_16564_),
    .B1(_16569_),
    .A1(_15788_),
    .Y(_16570_),
    .A2(_16565_));
 sg13g2_nor2_1 _23534_ (.A(_15780_),
    .B(_16570_),
    .Y(_16571_));
 sg13g2_o21ai_1 _23535_ (.B1(_15778_),
    .Y(_16572_),
    .A1(_16563_),
    .A2(_16571_));
 sg13g2_a21oi_1 _23536_ (.A1(_16562_),
    .A2(_16572_),
    .Y(_16573_),
    .B1(_16552_));
 sg13g2_nor3_1 _23537_ (.A(_13976_),
    .B(\u_inv.f_reg[198] ),
    .C(_15776_),
    .Y(_16574_));
 sg13g2_nor2_1 _23538_ (.A(_13975_),
    .B(\u_inv.f_reg[199] ),
    .Y(_16575_));
 sg13g2_nor3_2 _23539_ (.A(_16573_),
    .B(_16574_),
    .C(_16575_),
    .Y(_16576_));
 sg13g2_nor2b_1 _23540_ (.A(_16576_),
    .B_N(_16558_),
    .Y(_16577_));
 sg13g2_nand2_1 _23541_ (.Y(_16578_),
    .A(\u_inv.f_next[204] ),
    .B(_14458_));
 sg13g2_a21oi_1 _23542_ (.A1(_15806_),
    .A2(_15807_),
    .Y(_16579_),
    .B1(_16578_));
 sg13g2_a21oi_1 _23543_ (.A1(\u_inv.f_next[205] ),
    .A2(_14459_),
    .Y(_16580_),
    .B1(_16579_));
 sg13g2_nor2_1 _23544_ (.A(_13968_),
    .B(\u_inv.f_reg[206] ),
    .Y(_16581_));
 sg13g2_nor2_1 _23545_ (.A(_15799_),
    .B(_16580_),
    .Y(_16582_));
 sg13g2_nor2_1 _23546_ (.A(_16581_),
    .B(_16582_),
    .Y(_16583_));
 sg13g2_nor2_1 _23547_ (.A(_15801_),
    .B(_16583_),
    .Y(_16584_));
 sg13g2_a21oi_1 _23548_ (.A1(\u_inv.f_next[207] ),
    .A2(_14461_),
    .Y(_16585_),
    .B1(_16584_));
 sg13g2_nor2_1 _23549_ (.A(_13971_),
    .B(\u_inv.f_reg[203] ),
    .Y(_16586_));
 sg13g2_nand2_1 _23550_ (.Y(_16587_),
    .A(\u_inv.f_next[202] ),
    .B(_14456_));
 sg13g2_nand2_1 _23551_ (.Y(_16588_),
    .A(\u_inv.f_next[201] ),
    .B(_14455_));
 sg13g2_nor2_1 _23552_ (.A(_13974_),
    .B(\u_inv.f_reg[200] ),
    .Y(_16589_));
 sg13g2_nand2_1 _23553_ (.Y(_16590_),
    .A(_15813_),
    .B(_16589_));
 sg13g2_and2_1 _23554_ (.A(_16588_),
    .B(_16590_),
    .X(_16591_));
 sg13g2_o21ai_1 _23555_ (.B1(_16587_),
    .Y(_16592_),
    .A1(_15815_),
    .A2(_16591_));
 sg13g2_a21oi_1 _23556_ (.A1(_15818_),
    .A2(_16592_),
    .Y(_16593_),
    .B1(_16586_));
 sg13g2_o21ai_1 _23557_ (.B1(_16585_),
    .Y(_16594_),
    .A1(_16556_),
    .A2(_16593_));
 sg13g2_nor2_2 _23558_ (.A(_16577_),
    .B(_16594_),
    .Y(_16595_));
 sg13g2_nor2_1 _23559_ (.A(_15985_),
    .B(_16559_),
    .Y(_16596_));
 sg13g2_o21ai_1 _23560_ (.B1(_16596_),
    .Y(_16597_),
    .A1(_16483_),
    .A2(_16547_));
 sg13g2_nor2_1 _23561_ (.A(_15985_),
    .B(_16595_),
    .Y(_16598_));
 sg13g2_nor4_2 _23562_ (.A(_15993_),
    .B(_15999_),
    .C(_16016_),
    .Y(_16599_),
    .D(_16598_));
 sg13g2_nor4_1 _23563_ (.A(_15856_),
    .B(_15858_),
    .C(_15863_),
    .D(_15865_),
    .Y(_16600_));
 sg13g2_nor2_1 _23564_ (.A(_15869_),
    .B(_15871_),
    .Y(_16601_));
 sg13g2_nand2_1 _23565_ (.Y(_16602_),
    .A(_15874_),
    .B(_15877_));
 sg13g2_nand4_1 _23566_ (.B(_15877_),
    .C(_16600_),
    .A(_15874_),
    .Y(_16603_),
    .D(_16601_));
 sg13g2_and2_1 _23567_ (.A(_15891_),
    .B(_15892_),
    .X(_16604_));
 sg13g2_nand3b_1 _23568_ (.B(_15898_),
    .C(_16604_),
    .Y(_16605_),
    .A_N(_15896_));
 sg13g2_nand2_1 _23569_ (.Y(_16606_),
    .A(_15881_),
    .B(_15883_));
 sg13g2_and2_1 _23570_ (.A(_15886_),
    .B(_15888_),
    .X(_16607_));
 sg13g2_nand2b_1 _23571_ (.Y(_16608_),
    .B(_16607_),
    .A_N(_16606_));
 sg13g2_nor2_1 _23572_ (.A(_16605_),
    .B(_16608_),
    .Y(_16609_));
 sg13g2_nand2b_1 _23573_ (.Y(_16610_),
    .B(_16609_),
    .A_N(_16603_));
 sg13g2_a21oi_2 _23574_ (.B1(_16610_),
    .Y(_16611_),
    .A2(_16599_),
    .A1(_16597_));
 sg13g2_nand2_1 _23575_ (.Y(_16612_),
    .A(\u_inv.f_next[227] ),
    .B(_14481_));
 sg13g2_nor2_1 _23576_ (.A(_13948_),
    .B(\u_inv.f_reg[226] ),
    .Y(_16613_));
 sg13g2_inv_1 _23577_ (.Y(_16614_),
    .A(_16613_));
 sg13g2_nor2_1 _23578_ (.A(_13950_),
    .B(\u_inv.f_reg[224] ),
    .Y(_16615_));
 sg13g2_nand2_1 _23579_ (.Y(_16616_),
    .A(_15874_),
    .B(_16615_));
 sg13g2_o21ai_1 _23580_ (.B1(_16616_),
    .Y(_16617_),
    .A1(_13949_),
    .A2(\u_inv.f_reg[225] ));
 sg13g2_a21oi_1 _23581_ (.A1(_15872_),
    .A2(_16617_),
    .Y(_16618_),
    .B1(_16613_));
 sg13g2_o21ai_1 _23582_ (.B1(_16612_),
    .Y(_16619_),
    .A1(_15869_),
    .A2(_16618_));
 sg13g2_nor2_1 _23583_ (.A(_13944_),
    .B(\u_inv.f_reg[230] ),
    .Y(_16620_));
 sg13g2_nand2_1 _23584_ (.Y(_16621_),
    .A(\u_inv.f_next[228] ),
    .B(_14482_));
 sg13g2_nor2_1 _23585_ (.A(_15856_),
    .B(_16621_),
    .Y(_16622_));
 sg13g2_a21oi_1 _23586_ (.A1(\u_inv.f_next[229] ),
    .A2(_14483_),
    .Y(_16623_),
    .B1(_16622_));
 sg13g2_nor3_1 _23587_ (.A(_15863_),
    .B(_15865_),
    .C(_16623_),
    .Y(_16624_));
 sg13g2_nor3_1 _23588_ (.A(_13944_),
    .B(\u_inv.f_reg[230] ),
    .C(_15863_),
    .Y(_16625_));
 sg13g2_a221oi_1 _23589_ (.B2(_16619_),
    .C1(_16625_),
    .B1(_16600_),
    .A1(\u_inv.f_next[231] ),
    .Y(_16626_),
    .A2(_14485_));
 sg13g2_nand2b_2 _23590_ (.Y(_16627_),
    .B(_16626_),
    .A_N(_16624_));
 sg13g2_nor2_1 _23591_ (.A(_13939_),
    .B(\u_inv.f_reg[235] ),
    .Y(_16628_));
 sg13g2_nor2_1 _23592_ (.A(_13940_),
    .B(\u_inv.f_reg[234] ),
    .Y(_16629_));
 sg13g2_inv_1 _23593_ (.Y(_16630_),
    .A(_16629_));
 sg13g2_nand3_1 _23594_ (.B(_14486_),
    .C(_15891_),
    .A(\u_inv.f_next[232] ),
    .Y(_16631_));
 sg13g2_nand2_1 _23595_ (.Y(_16632_),
    .A(\u_inv.f_next[233] ),
    .B(_14487_));
 sg13g2_and2_1 _23596_ (.A(_16631_),
    .B(_16632_),
    .X(_16633_));
 sg13g2_o21ai_1 _23597_ (.B1(_16630_),
    .Y(_16634_),
    .A1(_15896_),
    .A2(_16633_));
 sg13g2_a21oi_1 _23598_ (.A1(_15898_),
    .A2(_16634_),
    .Y(_16635_),
    .B1(_16628_));
 sg13g2_nor2_1 _23599_ (.A(_13938_),
    .B(\u_inv.f_reg[236] ),
    .Y(_16636_));
 sg13g2_and2_1 _23600_ (.A(_15881_),
    .B(_16636_),
    .X(_16637_));
 sg13g2_a21o_1 _23601_ (.A2(_14491_),
    .A1(\u_inv.f_next[237] ),
    .B1(_16637_),
    .X(_16638_));
 sg13g2_nand2_1 _23602_ (.Y(_16639_),
    .A(\u_inv.f_next[238] ),
    .B(_14492_));
 sg13g2_nor2_1 _23603_ (.A(_15885_),
    .B(_16639_),
    .Y(_16640_));
 sg13g2_a221oi_1 _23604_ (.B2(_16638_),
    .C1(_16640_),
    .B1(_16607_),
    .A1(\u_inv.f_next[239] ),
    .Y(_16641_),
    .A2(_14493_));
 sg13g2_o21ai_1 _23605_ (.B1(_16641_),
    .Y(_16642_),
    .A1(_16608_),
    .A2(_16635_));
 sg13g2_a21oi_1 _23606_ (.A1(_16609_),
    .A2(_16627_),
    .Y(_16643_),
    .B1(_16642_));
 sg13g2_inv_1 _23607_ (.Y(_16644_),
    .A(_16643_));
 sg13g2_nor2_1 _23608_ (.A(_16611_),
    .B(_16644_),
    .Y(_16645_));
 sg13g2_nand2b_1 _23609_ (.Y(_16646_),
    .B(_16643_),
    .A_N(_16611_));
 sg13g2_and2_1 _23610_ (.A(_15929_),
    .B(_15930_),
    .X(_16647_));
 sg13g2_nor2_1 _23611_ (.A(_15935_),
    .B(_15937_),
    .Y(_16648_));
 sg13g2_nand2_1 _23612_ (.Y(_16649_),
    .A(_16647_),
    .B(_16648_));
 sg13g2_nor2_1 _23613_ (.A(_14842_),
    .B(_14843_),
    .Y(_16650_));
 sg13g2_nor2_1 _23614_ (.A(_14831_),
    .B(_14834_),
    .Y(_16651_));
 sg13g2_nand2_1 _23615_ (.Y(_16652_),
    .A(_16650_),
    .B(_16651_));
 sg13g2_nor2_1 _23616_ (.A(_16649_),
    .B(_16652_),
    .Y(_16653_));
 sg13g2_o21ai_1 _23617_ (.B1(_16653_),
    .Y(_16654_),
    .A1(_16611_),
    .A2(_16644_));
 sg13g2_nor2_1 _23618_ (.A(_13931_),
    .B(\u_inv.f_reg[243] ),
    .Y(_16655_));
 sg13g2_nor2_1 _23619_ (.A(_13932_),
    .B(\u_inv.f_reg[242] ),
    .Y(_16656_));
 sg13g2_nor2_1 _23620_ (.A(_13934_),
    .B(\u_inv.f_reg[240] ),
    .Y(_16657_));
 sg13g2_nand2_1 _23621_ (.Y(_16658_),
    .A(_15930_),
    .B(_16657_));
 sg13g2_o21ai_1 _23622_ (.B1(_16658_),
    .Y(_16659_),
    .A1(_13933_),
    .A2(\u_inv.f_reg[241] ));
 sg13g2_inv_1 _23623_ (.Y(_16660_),
    .A(_16659_));
 sg13g2_a221oi_1 _23624_ (.B2(_16648_),
    .C1(_16655_),
    .B1(_16659_),
    .A1(_15938_),
    .Y(_16661_),
    .A2(_16656_));
 sg13g2_nor2_1 _23625_ (.A(_16652_),
    .B(_16661_),
    .Y(_16662_));
 sg13g2_nor2_1 _23626_ (.A(_13930_),
    .B(\u_inv.f_reg[244] ),
    .Y(_16663_));
 sg13g2_nand2b_1 _23627_ (.Y(_16664_),
    .B(_16663_),
    .A_N(_14842_));
 sg13g2_o21ai_1 _23628_ (.B1(_16664_),
    .Y(_16665_),
    .A1(_13929_),
    .A2(\u_inv.f_reg[245] ));
 sg13g2_nand2_1 _23629_ (.Y(_16666_),
    .A(\u_inv.f_next[246] ),
    .B(_14500_));
 sg13g2_nor2_1 _23630_ (.A(_14831_),
    .B(_16666_),
    .Y(_16667_));
 sg13g2_a221oi_1 _23631_ (.B2(_16665_),
    .C1(_16667_),
    .B1(_16651_),
    .A1(\u_inv.f_next[247] ),
    .Y(_16668_),
    .A2(_14501_));
 sg13g2_nor2b_1 _23632_ (.A(_16662_),
    .B_N(_16668_),
    .Y(_16669_));
 sg13g2_nand2_1 _23633_ (.Y(_16670_),
    .A(_16654_),
    .B(_16669_));
 sg13g2_nand2_1 _23634_ (.Y(_16671_),
    .A(_15950_),
    .B(_15951_));
 sg13g2_a21oi_1 _23635_ (.A1(_16654_),
    .A2(_16669_),
    .Y(_16672_),
    .B1(_16671_));
 sg13g2_nor2_1 _23636_ (.A(_13926_),
    .B(\u_inv.f_reg[248] ),
    .Y(_16673_));
 sg13g2_nand2_1 _23637_ (.Y(_16674_),
    .A(_15951_),
    .B(_16673_));
 sg13g2_o21ai_1 _23638_ (.B1(_16674_),
    .Y(_16675_),
    .A1(_13925_),
    .A2(\u_inv.f_reg[249] ));
 sg13g2_o21ai_1 _23639_ (.B1(_14830_),
    .Y(_16676_),
    .A1(_16672_),
    .A2(_16675_));
 sg13g2_nor2_1 _23640_ (.A(_13924_),
    .B(\u_inv.f_reg[250] ),
    .Y(_16677_));
 sg13g2_o21ai_1 _23641_ (.B1(_16676_),
    .Y(_16678_),
    .A1(_13924_),
    .A2(\u_inv.f_reg[250] ));
 sg13g2_a21oi_1 _23642_ (.A1(_14829_),
    .A2(_16678_),
    .Y(_16679_),
    .B1(net5026));
 sg13g2_o21ai_1 _23643_ (.B1(_16679_),
    .Y(_16680_),
    .A1(_14829_),
    .A2(_16678_));
 sg13g2_nand2b_2 _23644_ (.Y(_16681_),
    .B(_16680_),
    .A_N(_15971_));
 sg13g2_a21oi_1 _23645_ (.A1(_16597_),
    .A2(_16599_),
    .Y(_16682_),
    .B1(_16603_));
 sg13g2_nor2_1 _23646_ (.A(_16627_),
    .B(_16682_),
    .Y(_16683_));
 sg13g2_or2_1 _23647_ (.X(_16684_),
    .B(_16683_),
    .A(_16605_));
 sg13g2_nand2_1 _23648_ (.Y(_16685_),
    .A(_16635_),
    .B(_16684_));
 sg13g2_a21oi_1 _23649_ (.A1(_16635_),
    .A2(_16684_),
    .Y(_16686_),
    .B1(_16606_));
 sg13g2_o21ai_1 _23650_ (.B1(_15888_),
    .Y(_16687_),
    .A1(_16638_),
    .A2(_16686_));
 sg13g2_and2_1 _23651_ (.A(_16639_),
    .B(_16687_),
    .X(_16688_));
 sg13g2_a21oi_1 _23652_ (.A1(_15885_),
    .A2(_16688_),
    .Y(_16689_),
    .B1(net5034));
 sg13g2_o21ai_1 _23653_ (.B1(_16689_),
    .Y(_16690_),
    .A1(_15885_),
    .A2(_16688_));
 sg13g2_o21ai_1 _23654_ (.B1(_15880_),
    .Y(_16691_),
    .A1(_15852_),
    .A2(_15855_));
 sg13g2_a21oi_2 _23655_ (.B1(_15894_),
    .Y(_16692_),
    .A2(_16691_),
    .A1(_15915_));
 sg13g2_a21oi_1 _23656_ (.A1(_15899_),
    .A2(_16692_),
    .Y(_16693_),
    .B1(_15921_));
 sg13g2_a21o_1 _23657_ (.A2(_16692_),
    .A1(_15899_),
    .B1(_15921_),
    .X(_16694_));
 sg13g2_a21oi_1 _23658_ (.A1(_15884_),
    .A2(_16694_),
    .Y(_16695_),
    .B1(_15923_));
 sg13g2_or2_1 _23659_ (.X(_16696_),
    .B(_16695_),
    .A(_15888_));
 sg13g2_nand2_1 _23660_ (.Y(_16697_),
    .A(_15887_),
    .B(_16696_));
 sg13g2_o21ai_1 _23661_ (.B1(net5738),
    .Y(_16698_),
    .A1(_15886_),
    .A2(_16697_));
 sg13g2_a21oi_1 _23662_ (.A1(_15886_),
    .A2(_16697_),
    .Y(_16699_),
    .B1(_16698_));
 sg13g2_o21ai_1 _23663_ (.B1(net5034),
    .Y(_16700_),
    .A1(\u_inv.f_next[239] ),
    .A2(net5738));
 sg13g2_o21ai_1 _23664_ (.B1(_16690_),
    .Y(_16701_),
    .A1(_16699_),
    .A2(_16700_));
 sg13g2_a21o_2 _23665_ (.A2(_16595_),
    .A1(_16561_),
    .B1(_15984_),
    .X(_16702_));
 sg13g2_and2_1 _23666_ (.A(_16015_),
    .B(_16702_),
    .X(_16703_));
 sg13g2_or2_1 _23667_ (.X(_16704_),
    .B(_16703_),
    .A(_14874_));
 sg13g2_a21oi_2 _23668_ (.B1(_15976_),
    .Y(_16705_),
    .A2(_16702_),
    .A1(_16015_));
 sg13g2_a21o_2 _23669_ (.A2(_16705_),
    .A1(_15977_),
    .B1(_15992_),
    .X(_16706_));
 sg13g2_and2_1 _23670_ (.A(_15973_),
    .B(_16706_),
    .X(_16707_));
 sg13g2_o21ai_1 _23671_ (.B1(_14848_),
    .Y(_16708_),
    .A1(_15996_),
    .A2(_16707_));
 sg13g2_nand2b_1 _23672_ (.Y(_16709_),
    .B(_16708_),
    .A_N(_15997_));
 sg13g2_a21oi_1 _23673_ (.A1(_14849_),
    .A2(_16709_),
    .Y(_16710_),
    .B1(net5041));
 sg13g2_o21ai_1 _23674_ (.B1(_16710_),
    .Y(_16711_),
    .A1(_14849_),
    .A2(_16709_));
 sg13g2_nand2_2 _23675_ (.Y(_16712_),
    .A(_15823_),
    .B(_15847_));
 sg13g2_nand3_1 _23676_ (.B(_14913_),
    .C(_16712_),
    .A(_14911_),
    .Y(_16713_));
 sg13g2_a21oi_1 _23677_ (.A1(_15823_),
    .A2(_15847_),
    .Y(_16714_),
    .B1(_15848_));
 sg13g2_a21oi_1 _23678_ (.A1(_15823_),
    .A2(_15847_),
    .Y(_16715_),
    .B1(_15850_));
 sg13g2_nor2_1 _23679_ (.A(_14909_),
    .B(_16715_),
    .Y(_16716_));
 sg13g2_o21ai_1 _23680_ (.B1(_14877_),
    .Y(_16717_),
    .A1(_14909_),
    .A2(_16715_));
 sg13g2_o21ai_1 _23681_ (.B1(_14868_),
    .Y(_16718_),
    .A1(_14862_),
    .A2(_16717_));
 sg13g2_a21oi_1 _23682_ (.A1(_14855_),
    .A2(_16718_),
    .Y(_16719_),
    .B1(_14872_));
 sg13g2_o21ai_1 _23683_ (.B1(_14847_),
    .Y(_16720_),
    .A1(_14848_),
    .A2(_16719_));
 sg13g2_xnor2_1 _23684_ (.Y(_16721_),
    .A(_14849_),
    .B(_16720_));
 sg13g2_nor2_1 _23685_ (.A(\u_inv.f_next[223] ),
    .B(net5751),
    .Y(_16722_));
 sg13g2_o21ai_1 _23686_ (.B1(net5041),
    .Y(_16723_),
    .A1(net5674),
    .A2(_16721_));
 sg13g2_o21ai_1 _23687_ (.B1(_16711_),
    .Y(_16724_),
    .A1(_16722_),
    .A2(_16723_));
 sg13g2_a21oi_2 _23688_ (.B1(_16602_),
    .Y(_16725_),
    .A2(_16599_),
    .A1(_16597_));
 sg13g2_a21o_1 _23689_ (.A2(_16725_),
    .A1(_16601_),
    .B1(_16619_),
    .X(_16726_));
 sg13g2_nand2_2 _23690_ (.Y(_16727_),
    .A(_15859_),
    .B(_16726_));
 sg13g2_nor2_1 _23691_ (.A(_15856_),
    .B(_16727_),
    .Y(_16728_));
 sg13g2_o21ai_1 _23692_ (.B1(_16623_),
    .Y(_16729_),
    .A1(_15856_),
    .A2(_16727_));
 sg13g2_a21oi_1 _23693_ (.A1(_15866_),
    .A2(_16729_),
    .Y(_16730_),
    .B1(_16620_));
 sg13g2_a21oi_1 _23694_ (.A1(_15863_),
    .A2(_16730_),
    .Y(_16731_),
    .B1(net5035));
 sg13g2_o21ai_1 _23695_ (.B1(_16731_),
    .Y(_16732_),
    .A1(_15863_),
    .A2(_16730_));
 sg13g2_o21ai_1 _23696_ (.B1(_15876_),
    .Y(_16733_),
    .A1(_15852_),
    .A2(_15855_));
 sg13g2_o21ai_1 _23697_ (.B1(_15879_),
    .Y(_16734_),
    .A1(_15852_),
    .A2(_15855_));
 sg13g2_o21ai_1 _23698_ (.B1(_15909_),
    .Y(_16735_),
    .A1(_15873_),
    .A2(_16734_));
 sg13g2_a21oi_1 _23699_ (.A1(_15860_),
    .A2(_16735_),
    .Y(_16736_),
    .B1(_15912_));
 sg13g2_o21ai_1 _23700_ (.B1(_15864_),
    .Y(_16737_),
    .A1(_15866_),
    .A2(_16736_));
 sg13g2_xnor2_1 _23701_ (.Y(_16738_),
    .A(_15863_),
    .B(_16737_));
 sg13g2_a21oi_1 _23702_ (.A1(net5739),
    .A2(_16738_),
    .Y(_16739_),
    .B1(net4942));
 sg13g2_o21ai_1 _23703_ (.B1(_16739_),
    .Y(_16740_),
    .A1(net3258),
    .A2(net5739));
 sg13g2_nand2_1 _23704_ (.Y(_16741_),
    .A(_16732_),
    .B(_16740_));
 sg13g2_and3_1 _23705_ (.X(_16742_),
    .A(_14830_),
    .B(_15953_),
    .C(_15955_));
 sg13g2_o21ai_1 _23706_ (.B1(net5730),
    .Y(_16743_),
    .A1(_15956_),
    .A2(_16742_));
 sg13g2_o21ai_1 _23707_ (.B1(_16743_),
    .Y(_16744_),
    .A1(\u_inv.f_next[250] ),
    .A2(net5730));
 sg13g2_nor3_1 _23708_ (.A(_14830_),
    .B(_16672_),
    .C(_16675_),
    .Y(_16745_));
 sg13g2_nor2_1 _23709_ (.A(net5026),
    .B(_16745_),
    .Y(_16746_));
 sg13g2_nand2_1 _23710_ (.Y(_16747_),
    .A(_16676_),
    .B(_16746_));
 sg13g2_o21ai_1 _23711_ (.B1(_16747_),
    .Y(_16748_),
    .A1(net4928),
    .A2(_16744_));
 sg13g2_a21oi_2 _23712_ (.B1(_15943_),
    .Y(_16749_),
    .A2(_15939_),
    .A1(_15933_));
 sg13g2_o21ai_1 _23713_ (.B1(_14838_),
    .Y(_16750_),
    .A1(_14845_),
    .A2(_16749_));
 sg13g2_xnor2_1 _23714_ (.Y(_16751_),
    .A(_14834_),
    .B(_16750_));
 sg13g2_nand2_1 _23715_ (.Y(_16752_),
    .A(net5735),
    .B(_16751_));
 sg13g2_a21oi_1 _23716_ (.A1(_13928_),
    .A2(net5663),
    .Y(_16753_),
    .B1(net4938));
 sg13g2_o21ai_1 _23717_ (.B1(_16661_),
    .Y(_16754_),
    .A1(_16645_),
    .A2(_16649_));
 sg13g2_a21oi_1 _23718_ (.A1(_16650_),
    .A2(_16754_),
    .Y(_16755_),
    .B1(_16665_));
 sg13g2_nand2_1 _23719_ (.Y(_16756_),
    .A(_14834_),
    .B(_16755_));
 sg13g2_nor2_1 _23720_ (.A(_14834_),
    .B(_16755_),
    .Y(_16757_));
 sg13g2_nor2_1 _23721_ (.A(net5031),
    .B(_16757_),
    .Y(_16758_));
 sg13g2_and2_1 _23722_ (.A(_16756_),
    .B(_16758_),
    .X(_16759_));
 sg13g2_a22oi_1 _23723_ (.Y(_16760_),
    .B1(_16756_),
    .B2(_16758_),
    .A2(_16753_),
    .A1(_16752_));
 sg13g2_a21o_1 _23724_ (.A2(_16753_),
    .A1(_16752_),
    .B1(_16759_),
    .X(_16761_));
 sg13g2_o21ai_1 _23725_ (.B1(_15896_),
    .Y(_16762_),
    .A1(_15918_),
    .A2(_16692_));
 sg13g2_nand2_1 _23726_ (.Y(_16763_),
    .A(_15895_),
    .B(_16762_));
 sg13g2_xnor2_1 _23727_ (.Y(_16764_),
    .A(_15897_),
    .B(_16763_));
 sg13g2_o21ai_1 _23728_ (.B1(net5035),
    .Y(_16765_),
    .A1(\u_inv.f_next[235] ),
    .A2(net5738));
 sg13g2_a21oi_1 _23729_ (.A1(net5738),
    .A2(_16764_),
    .Y(_16766_),
    .B1(_16765_));
 sg13g2_o21ai_1 _23730_ (.B1(_16604_),
    .Y(_16767_),
    .A1(_16627_),
    .A2(_16682_));
 sg13g2_a21oi_1 _23731_ (.A1(_16633_),
    .A2(_16767_),
    .Y(_16768_),
    .B1(_15896_));
 sg13g2_nor2_1 _23732_ (.A(_16629_),
    .B(_16768_),
    .Y(_16769_));
 sg13g2_o21ai_1 _23733_ (.B1(net4941),
    .Y(_16770_),
    .A1(_15897_),
    .A2(_16769_));
 sg13g2_a21oi_1 _23734_ (.A1(_15897_),
    .A2(_16769_),
    .Y(_16771_),
    .B1(_16770_));
 sg13g2_or2_1 _23735_ (.X(_16772_),
    .B(_16771_),
    .A(_16766_));
 sg13g2_o21ai_1 _23736_ (.B1(_15935_),
    .Y(_16773_),
    .A1(_15933_),
    .A2(_15941_));
 sg13g2_a21oi_1 _23737_ (.A1(_15934_),
    .A2(_16773_),
    .Y(_16774_),
    .B1(_15937_));
 sg13g2_and3_1 _23738_ (.X(_16775_),
    .A(_15934_),
    .B(_15937_),
    .C(_16773_));
 sg13g2_nor3_1 _23739_ (.A(net5664),
    .B(_16774_),
    .C(_16775_),
    .Y(_16776_));
 sg13g2_o21ai_1 _23740_ (.B1(net5032),
    .Y(_16777_),
    .A1(\u_inv.f_next[243] ),
    .A2(net5735));
 sg13g2_o21ai_1 _23741_ (.B1(_16647_),
    .Y(_16778_),
    .A1(_16611_),
    .A2(_16644_));
 sg13g2_a21oi_1 _23742_ (.A1(_16660_),
    .A2(_16778_),
    .Y(_16779_),
    .B1(_15935_));
 sg13g2_or3_1 _23743_ (.A(_15938_),
    .B(_16656_),
    .C(_16779_),
    .X(_16780_));
 sg13g2_o21ai_1 _23744_ (.B1(_15938_),
    .Y(_16781_),
    .A1(_16656_),
    .A2(_16779_));
 sg13g2_nand3_1 _23745_ (.B(_16780_),
    .C(_16781_),
    .A(net4938),
    .Y(_16782_));
 sg13g2_o21ai_1 _23746_ (.B1(_16782_),
    .Y(_16783_),
    .A1(_16776_),
    .A2(_16777_));
 sg13g2_xnor2_1 _23747_ (.Y(_16784_),
    .A(_14843_),
    .B(_16749_));
 sg13g2_nor2_1 _23748_ (.A(\u_inv.f_next[244] ),
    .B(net5735),
    .Y(_16785_));
 sg13g2_o21ai_1 _23749_ (.B1(net5037),
    .Y(_16786_),
    .A1(net5664),
    .A2(_16784_));
 sg13g2_nand2_1 _23750_ (.Y(_16787_),
    .A(_14844_),
    .B(_16754_));
 sg13g2_o21ai_1 _23751_ (.B1(net4939),
    .Y(_16788_),
    .A1(_14844_),
    .A2(_16754_));
 sg13g2_nand2b_1 _23752_ (.Y(_16789_),
    .B(_16787_),
    .A_N(_16788_));
 sg13g2_o21ai_1 _23753_ (.B1(_16789_),
    .Y(_16790_),
    .A1(_16785_),
    .A2(_16786_));
 sg13g2_nor2b_1 _23754_ (.A(_16663_),
    .B_N(_14842_),
    .Y(_16791_));
 sg13g2_nand2_1 _23755_ (.Y(_16792_),
    .A(net4939),
    .B(_16664_));
 sg13g2_a221oi_1 _23756_ (.B2(_16791_),
    .C1(_16792_),
    .B1(_16787_),
    .A1(_16650_),
    .Y(_16793_),
    .A2(_16754_));
 sg13g2_o21ai_1 _23757_ (.B1(_14836_),
    .Y(_16794_),
    .A1(_14844_),
    .A2(_16749_));
 sg13g2_xnor2_1 _23758_ (.Y(_16795_),
    .A(_14842_),
    .B(_16794_));
 sg13g2_o21ai_1 _23759_ (.B1(net5037),
    .Y(_16796_),
    .A1(\u_inv.f_next[245] ),
    .A2(net5735));
 sg13g2_a21oi_1 _23760_ (.A1(net5735),
    .A2(_16795_),
    .Y(_16797_),
    .B1(_16796_));
 sg13g2_nor2_2 _23761_ (.A(_16793_),
    .B(_16797_),
    .Y(_16798_));
 sg13g2_or2_1 _23762_ (.X(_16799_),
    .B(_16797_),
    .A(_16793_));
 sg13g2_xnor2_1 _23763_ (.Y(_16800_),
    .A(_14853_),
    .B(_16706_));
 sg13g2_o21ai_1 _23764_ (.B1(net5752),
    .Y(_16801_),
    .A1(_14854_),
    .A2(_16718_));
 sg13g2_a21o_1 _23765_ (.A2(_16718_),
    .A1(_14854_),
    .B1(_16801_),
    .X(_16802_));
 sg13g2_a21oi_1 _23766_ (.A1(\u_inv.f_next[220] ),
    .A2(net5674),
    .Y(_16803_),
    .B1(net4951));
 sg13g2_a22oi_1 _23767_ (.Y(_16804_),
    .B1(_16802_),
    .B2(_16803_),
    .A2(_16800_),
    .A1(net4952));
 sg13g2_or2_1 _23768_ (.X(_16805_),
    .B(_16636_),
    .A(_15881_));
 sg13g2_a21oi_1 _23769_ (.A1(_15883_),
    .A2(_16685_),
    .Y(_16806_),
    .B1(_16805_));
 sg13g2_nor4_1 _23770_ (.A(net5034),
    .B(_16637_),
    .C(_16686_),
    .D(_16806_),
    .Y(_16807_));
 sg13g2_o21ai_1 _23771_ (.B1(_15882_),
    .Y(_16808_),
    .A1(_15883_),
    .A2(_16693_));
 sg13g2_xor2_1 _23772_ (.B(_16808_),
    .A(_15881_),
    .X(_16809_));
 sg13g2_o21ai_1 _23773_ (.B1(net5034),
    .Y(_16810_),
    .A1(\u_inv.f_next[237] ),
    .A2(net5738));
 sg13g2_a21oi_1 _23774_ (.A1(net5738),
    .A2(_16809_),
    .Y(_16811_),
    .B1(_16810_));
 sg13g2_nor2_1 _23775_ (.A(_16807_),
    .B(_16811_),
    .Y(_16812_));
 sg13g2_inv_1 _23776_ (.Y(_16813_),
    .A(_16812_));
 sg13g2_or3_1 _23777_ (.A(_15933_),
    .B(_15935_),
    .C(_15941_),
    .X(_16814_));
 sg13g2_nand2_1 _23778_ (.Y(_16815_),
    .A(_16773_),
    .B(_16814_));
 sg13g2_nor2_1 _23779_ (.A(\u_inv.f_next[242] ),
    .B(net5737),
    .Y(_16816_));
 sg13g2_a21oi_1 _23780_ (.A1(net5735),
    .A2(_16815_),
    .Y(_16817_),
    .B1(_16816_));
 sg13g2_nand3_1 _23781_ (.B(_16660_),
    .C(_16778_),
    .A(_15935_),
    .Y(_16818_));
 sg13g2_nor2_1 _23782_ (.A(net5032),
    .B(_16779_),
    .Y(_16819_));
 sg13g2_a22oi_1 _23783_ (.Y(_16820_),
    .B1(_16818_),
    .B2(_16819_),
    .A2(_16817_),
    .A1(net5032));
 sg13g2_inv_1 _23784_ (.Y(_16821_),
    .A(_16820_));
 sg13g2_o21ai_1 _23785_ (.B1(_15872_),
    .Y(_16822_),
    .A1(_16617_),
    .A2(_16725_));
 sg13g2_nand3_1 _23786_ (.B(_16614_),
    .C(_16822_),
    .A(_15869_),
    .Y(_16823_));
 sg13g2_a21o_1 _23787_ (.A2(_16822_),
    .A1(_16614_),
    .B1(_15869_),
    .X(_16824_));
 sg13g2_nand3_1 _23788_ (.B(_16823_),
    .C(_16824_),
    .A(net4941),
    .Y(_16825_));
 sg13g2_a21o_1 _23789_ (.A2(_16734_),
    .A1(_15906_),
    .B1(_15872_),
    .X(_16826_));
 sg13g2_and3_1 _23790_ (.X(_16827_),
    .A(_15869_),
    .B(_15870_),
    .C(_16826_));
 sg13g2_a21oi_1 _23791_ (.A1(_15870_),
    .A2(_16826_),
    .Y(_16828_),
    .B1(_15869_));
 sg13g2_nor3_1 _23792_ (.A(net5666),
    .B(_16827_),
    .C(_16828_),
    .Y(_16829_));
 sg13g2_o21ai_1 _23793_ (.B1(net5035),
    .Y(_16830_),
    .A1(\u_inv.f_next[227] ),
    .A2(net5739));
 sg13g2_o21ai_1 _23794_ (.B1(_16825_),
    .Y(_16831_),
    .A1(_16829_),
    .A2(_16830_));
 sg13g2_xnor2_1 _23795_ (.Y(_16832_),
    .A(_15948_),
    .B(_15950_));
 sg13g2_o21ai_1 _23796_ (.B1(net5032),
    .Y(_16833_),
    .A1(\u_inv.f_next[248] ),
    .A2(net5736));
 sg13g2_a21oi_1 _23797_ (.A1(net5736),
    .A2(_16832_),
    .Y(_16834_),
    .B1(_16833_));
 sg13g2_xor2_1 _23798_ (.B(_16670_),
    .A(_15950_),
    .X(_16835_));
 sg13g2_a21o_2 _23799_ (.A2(_16835_),
    .A1(net4938),
    .B1(_16834_),
    .X(_16836_));
 sg13g2_o21ai_1 _23800_ (.B1(_15949_),
    .Y(_16837_),
    .A1(_15948_),
    .A2(_15950_));
 sg13g2_xor2_1 _23801_ (.B(_16837_),
    .A(_15951_),
    .X(_16838_));
 sg13g2_o21ai_1 _23802_ (.B1(net5026),
    .Y(_16839_),
    .A1(\u_inv.f_next[249] ),
    .A2(net5730));
 sg13g2_a21oi_1 _23803_ (.A1(net5736),
    .A2(_16838_),
    .Y(_16840_),
    .B1(_16839_));
 sg13g2_a21o_1 _23804_ (.A2(_16670_),
    .A1(_15950_),
    .B1(_16673_),
    .X(_16841_));
 sg13g2_o21ai_1 _23805_ (.B1(net4938),
    .Y(_16842_),
    .A1(_15951_),
    .A2(_16841_));
 sg13g2_a21o_1 _23806_ (.A2(_16841_),
    .A1(_15951_),
    .B1(_16842_),
    .X(_16843_));
 sg13g2_nand2b_2 _23807_ (.Y(_16844_),
    .B(_16843_),
    .A_N(_16840_));
 sg13g2_xnor2_1 _23808_ (.Y(_16845_),
    .A(_14848_),
    .B(_16719_));
 sg13g2_o21ai_1 _23809_ (.B1(net5041),
    .Y(_16846_),
    .A1(\u_inv.f_next[222] ),
    .A2(net5751));
 sg13g2_a21o_1 _23810_ (.A2(_16845_),
    .A1(net5751),
    .B1(_16846_),
    .X(_16847_));
 sg13g2_nor3_1 _23811_ (.A(_14848_),
    .B(_15996_),
    .C(_16707_),
    .Y(_16848_));
 sg13g2_nand2_1 _23812_ (.Y(_16849_),
    .A(net4951),
    .B(_16708_));
 sg13g2_o21ai_1 _23813_ (.B1(_16847_),
    .Y(_16850_),
    .A1(_16848_),
    .A2(_16849_));
 sg13g2_a21o_2 _23814_ (.A2(_15764_),
    .A1(_15760_),
    .B1(_15771_),
    .X(_16851_));
 sg13g2_a21oi_1 _23815_ (.A1(_15026_),
    .A2(_16851_),
    .Y(_16852_),
    .B1(_14960_));
 sg13g2_o21ai_1 _23816_ (.B1(_14932_),
    .Y(_16853_),
    .A1(_15046_),
    .A2(_16852_));
 sg13g2_o21ai_1 _23817_ (.B1(_14933_),
    .Y(_16854_),
    .A1(_15046_),
    .A2(_16852_));
 sg13g2_o21ai_1 _23818_ (.B1(_15032_),
    .Y(_16855_),
    .A1(_14929_),
    .A2(_16854_));
 sg13g2_a21oi_1 _23819_ (.A1(_14924_),
    .A2(_16855_),
    .Y(_16856_),
    .B1(_15035_));
 sg13g2_xnor2_1 _23820_ (.Y(_16857_),
    .A(_14917_),
    .B(_16856_));
 sg13g2_nor2_1 _23821_ (.A(\u_inv.f_next[190] ),
    .B(net5766),
    .Y(_16858_));
 sg13g2_a21oi_1 _23822_ (.A1(net5766),
    .A2(_16857_),
    .Y(_16859_),
    .B1(_16858_));
 sg13g2_a221oi_1 _23823_ (.B2(_16458_),
    .C1(_16481_),
    .B1(_16423_),
    .A1(_16059_),
    .Y(_16860_),
    .A2(_16062_));
 sg13g2_o21ai_1 _23824_ (.B1(_16469_),
    .Y(_16861_),
    .A1(_16514_),
    .A2(_16860_));
 sg13g2_a21oi_2 _23825_ (.B1(_16465_),
    .Y(_16862_),
    .A2(_16861_),
    .A1(_16542_));
 sg13g2_a221oi_1 _23826_ (.B2(_16463_),
    .C1(_16515_),
    .B1(_16862_),
    .A1(net5623),
    .Y(_16863_),
    .A2(_16520_));
 sg13g2_nand2b_1 _23827_ (.Y(_16864_),
    .B(_16460_),
    .A_N(_16863_));
 sg13g2_o21ai_1 _23828_ (.B1(_16524_),
    .Y(_16865_),
    .A1(_16461_),
    .A2(_16863_));
 sg13g2_nor2_1 _23829_ (.A(_14917_),
    .B(_16865_),
    .Y(_16866_));
 sg13g2_nand2_1 _23830_ (.Y(_16867_),
    .A(_14917_),
    .B(_16865_));
 sg13g2_nor2_1 _23831_ (.A(net5055),
    .B(_16866_),
    .Y(_16868_));
 sg13g2_a22oi_1 _23832_ (.Y(_16869_),
    .B1(_16867_),
    .B2(_16868_),
    .A2(_16859_),
    .A1(net5055));
 sg13g2_inv_1 _23833_ (.Y(_16870_),
    .A(_16869_));
 sg13g2_or3_1 _23834_ (.A(_15896_),
    .B(_15918_),
    .C(_16692_),
    .X(_16871_));
 sg13g2_a21o_1 _23835_ (.A2(_16871_),
    .A1(_16762_),
    .B1(net5665),
    .X(_16872_));
 sg13g2_nor2_1 _23836_ (.A(\u_inv.f_next[234] ),
    .B(net5739),
    .Y(_16873_));
 sg13g2_nor2_1 _23837_ (.A(net4941),
    .B(_16873_),
    .Y(_16874_));
 sg13g2_nand2_1 _23838_ (.Y(_16875_),
    .A(net5035),
    .B(_16872_));
 sg13g2_nand3_1 _23839_ (.B(_16633_),
    .C(_16767_),
    .A(_15896_),
    .Y(_16876_));
 sg13g2_nor2_1 _23840_ (.A(net5034),
    .B(_16768_),
    .Y(_16877_));
 sg13g2_nand2_1 _23841_ (.Y(_16878_),
    .A(_16876_),
    .B(_16877_));
 sg13g2_a22oi_1 _23842_ (.Y(_16879_),
    .B1(_16876_),
    .B2(_16877_),
    .A2(_16874_),
    .A1(_16872_));
 sg13g2_o21ai_1 _23843_ (.B1(_16878_),
    .Y(_16880_),
    .A1(_16873_),
    .A2(_16875_));
 sg13g2_a21o_1 _23844_ (.A2(_16706_),
    .A1(_14853_),
    .B1(_15994_),
    .X(_16881_));
 sg13g2_a21oi_1 _23845_ (.A1(_14851_),
    .A2(_16881_),
    .Y(_16882_),
    .B1(net5042));
 sg13g2_o21ai_1 _23846_ (.B1(_16882_),
    .Y(_16883_),
    .A1(_14851_),
    .A2(_16881_));
 sg13g2_a21oi_1 _23847_ (.A1(_14854_),
    .A2(_16718_),
    .Y(_16884_),
    .B1(_14852_));
 sg13g2_xnor2_1 _23848_ (.Y(_16885_),
    .A(_14851_),
    .B(_16884_));
 sg13g2_mux2_1 _23849_ (.A0(_13953_),
    .A1(_16885_),
    .S(net5752),
    .X(_16886_));
 sg13g2_o21ai_1 _23850_ (.B1(_16883_),
    .Y(_16887_),
    .A1(net4952),
    .A2(_16886_));
 sg13g2_a21oi_1 _23851_ (.A1(_14834_),
    .A2(_16750_),
    .Y(_16888_),
    .B1(_14833_));
 sg13g2_or2_1 _23852_ (.X(_16889_),
    .B(_16888_),
    .A(_14831_));
 sg13g2_a21oi_1 _23853_ (.A1(_14831_),
    .A2(_16888_),
    .Y(_16890_),
    .B1(net5663));
 sg13g2_o21ai_1 _23854_ (.B1(net5032),
    .Y(_16891_),
    .A1(\u_inv.f_next[247] ),
    .A2(net5736));
 sg13g2_a21o_1 _23855_ (.A2(_16890_),
    .A1(_16889_),
    .B1(_16891_),
    .X(_16892_));
 sg13g2_o21ai_1 _23856_ (.B1(_16666_),
    .Y(_16893_),
    .A1(_14834_),
    .A2(_16755_));
 sg13g2_and2_1 _23857_ (.A(_14832_),
    .B(_16893_),
    .X(_16894_));
 sg13g2_o21ai_1 _23858_ (.B1(net4938),
    .Y(_16895_),
    .A1(_14832_),
    .A2(_16893_));
 sg13g2_o21ai_1 _23859_ (.B1(_16892_),
    .Y(_16896_),
    .A1(_16894_),
    .A2(_16895_));
 sg13g2_a21oi_1 _23860_ (.A1(_16526_),
    .A2(_16867_),
    .Y(_16897_),
    .B1(_14914_));
 sg13g2_nand3_1 _23861_ (.B(_16526_),
    .C(_16867_),
    .A(_14914_),
    .Y(_16898_));
 sg13g2_nor2_1 _23862_ (.A(net5055),
    .B(_16897_),
    .Y(_16899_));
 sg13g2_o21ai_1 _23863_ (.B1(_14916_),
    .Y(_16900_),
    .A1(_14917_),
    .A2(_16856_));
 sg13g2_xnor2_1 _23864_ (.Y(_16901_),
    .A(_14914_),
    .B(_16900_));
 sg13g2_o21ai_1 _23865_ (.B1(net5055),
    .Y(_16902_),
    .A1(\u_inv.f_next[191] ),
    .A2(net5766));
 sg13g2_a21oi_1 _23866_ (.A1(net5766),
    .A2(_16901_),
    .Y(_16903_),
    .B1(_16902_));
 sg13g2_a21o_2 _23867_ (.A2(_16899_),
    .A1(_16898_),
    .B1(_16903_),
    .X(_16904_));
 sg13g2_xnor2_1 _23868_ (.Y(_16905_),
    .A(_15866_),
    .B(_16736_));
 sg13g2_o21ai_1 _23869_ (.B1(net5035),
    .Y(_16906_),
    .A1(\u_inv.f_next[230] ),
    .A2(net5739));
 sg13g2_a21o_1 _23870_ (.A2(_16905_),
    .A1(net5739),
    .B1(_16906_),
    .X(_16907_));
 sg13g2_xnor2_1 _23871_ (.Y(_16908_),
    .A(_15866_),
    .B(_16729_));
 sg13g2_o21ai_1 _23872_ (.B1(_16907_),
    .Y(_16909_),
    .A1(net5035),
    .A2(_16908_));
 sg13g2_a21oi_1 _23873_ (.A1(_15888_),
    .A2(_16695_),
    .Y(_16910_),
    .B1(net5665));
 sg13g2_a22oi_1 _23874_ (.Y(_16911_),
    .B1(_16696_),
    .B2(_16910_),
    .A2(net5665),
    .A1(\u_inv.f_next[238] ));
 sg13g2_or3_1 _23875_ (.A(_15888_),
    .B(_16638_),
    .C(_16686_),
    .X(_16912_));
 sg13g2_a21oi_1 _23876_ (.A1(_16687_),
    .A2(_16912_),
    .Y(_16913_),
    .B1(net5034));
 sg13g2_a21o_2 _23877_ (.A2(_16911_),
    .A1(net5034),
    .B1(_16913_),
    .X(_16914_));
 sg13g2_inv_1 _23878_ (.Y(_16915_),
    .A(_16914_));
 sg13g2_nor2_1 _23879_ (.A(_13922_),
    .B(_14506_),
    .Y(_16916_));
 sg13g2_xnor2_1 _23880_ (.Y(_16917_),
    .A(\u_inv.f_next[252] ),
    .B(\u_inv.f_reg[252] ));
 sg13g2_inv_1 _23881_ (.Y(_16918_),
    .A(_16917_));
 sg13g2_a22oi_1 _23882_ (.Y(_16919_),
    .B1(\u_inv.f_reg[251] ),
    .B2(\u_inv.f_next[251] ),
    .A2(\u_inv.f_reg[250] ),
    .A1(\u_inv.f_next[250] ));
 sg13g2_a21o_1 _23883_ (.A2(_14505_),
    .A1(_13923_),
    .B1(_16919_),
    .X(_16920_));
 sg13g2_and2_1 _23884_ (.A(_15955_),
    .B(_16920_),
    .X(_16921_));
 sg13g2_or2_1 _23885_ (.X(_16922_),
    .B(_14830_),
    .A(_14829_));
 sg13g2_a22oi_1 _23886_ (.Y(_16923_),
    .B1(_16922_),
    .B2(_16920_),
    .A2(_16921_),
    .A1(_15953_));
 sg13g2_o21ai_1 _23887_ (.B1(net5736),
    .Y(_16924_),
    .A1(_16918_),
    .A2(_16923_));
 sg13g2_a21oi_1 _23888_ (.A1(_16918_),
    .A2(_16923_),
    .Y(_16925_),
    .B1(_16924_));
 sg13g2_a21oi_1 _23889_ (.A1(\u_inv.f_next[252] ),
    .A2(net5663),
    .Y(_16926_),
    .B1(_16925_));
 sg13g2_nand4_1 _23890_ (.B(_14830_),
    .C(_15950_),
    .A(_14829_),
    .Y(_16927_),
    .D(_15951_));
 sg13g2_a21oi_1 _23891_ (.A1(_16654_),
    .A2(_16669_),
    .Y(_16928_),
    .B1(_16927_));
 sg13g2_and2_1 _23892_ (.A(_14830_),
    .B(_16675_),
    .X(_16929_));
 sg13g2_o21ai_1 _23893_ (.B1(_14829_),
    .Y(_16930_),
    .A1(_16677_),
    .A2(_16929_));
 sg13g2_o21ai_1 _23894_ (.B1(_16930_),
    .Y(_16931_),
    .A1(_13923_),
    .A2(\u_inv.f_reg[251] ));
 sg13g2_or2_1 _23895_ (.X(_16932_),
    .B(_16931_),
    .A(_16928_));
 sg13g2_a21oi_1 _23896_ (.A1(_16917_),
    .A2(_16932_),
    .Y(_16933_),
    .B1(net5031));
 sg13g2_o21ai_1 _23897_ (.B1(_16933_),
    .Y(_16934_),
    .A1(_16917_),
    .A2(_16932_));
 sg13g2_o21ai_1 _23898_ (.B1(_16934_),
    .Y(_16935_),
    .A1(net4938),
    .A2(_16926_));
 sg13g2_xnor2_1 _23899_ (.Y(_16936_),
    .A(\u_inv.f_next[253] ),
    .B(\u_inv.f_reg[253] ));
 sg13g2_nor2_1 _23900_ (.A(_13922_),
    .B(\u_inv.f_reg[252] ),
    .Y(_16937_));
 sg13g2_a21o_1 _23901_ (.A2(_16932_),
    .A1(_16917_),
    .B1(_16937_),
    .X(_16938_));
 sg13g2_and2_1 _23902_ (.A(_16917_),
    .B(_16936_),
    .X(_16939_));
 sg13g2_nand2_1 _23903_ (.Y(_16940_),
    .A(_16917_),
    .B(_16936_));
 sg13g2_o21ai_1 _23904_ (.B1(_16939_),
    .Y(_16941_),
    .A1(_16928_),
    .A2(_16931_));
 sg13g2_o21ai_1 _23905_ (.B1(net4938),
    .Y(_16942_),
    .A1(_16936_),
    .A2(_16938_));
 sg13g2_a21o_1 _23906_ (.A2(_16938_),
    .A1(_16936_),
    .B1(_16942_),
    .X(_16943_));
 sg13g2_a21oi_1 _23907_ (.A1(_16918_),
    .A2(_16923_),
    .Y(_16944_),
    .B1(_16916_));
 sg13g2_xor2_1 _23908_ (.B(_16944_),
    .A(_16936_),
    .X(_16945_));
 sg13g2_nor2_1 _23909_ (.A(net5663),
    .B(_16945_),
    .Y(_16946_));
 sg13g2_o21ai_1 _23910_ (.B1(net5027),
    .Y(_16947_),
    .A1(\u_inv.f_next[253] ),
    .A2(net5736));
 sg13g2_o21ai_1 _23911_ (.B1(_16943_),
    .Y(_16948_),
    .A1(_16946_),
    .A2(_16947_));
 sg13g2_a221oi_1 _23912_ (.B2(_16458_),
    .C1(_16479_),
    .B1(_16423_),
    .A1(_16059_),
    .Y(_16949_),
    .A2(_16062_));
 sg13g2_a21oi_1 _23913_ (.A1(_16477_),
    .A2(_16949_),
    .Y(_16950_),
    .B1(_16498_));
 sg13g2_a21o_1 _23914_ (.A2(_16949_),
    .A1(_16477_),
    .B1(_16498_),
    .X(_16951_));
 sg13g2_nor2_1 _23915_ (.A(_16473_),
    .B(_16950_),
    .Y(_16952_));
 sg13g2_inv_1 _23916_ (.Y(_16953_),
    .A(_16952_));
 sg13g2_nand4_1 _23917_ (.B(_15013_),
    .C(_16472_),
    .A(_15011_),
    .Y(_16954_),
    .D(_16951_));
 sg13g2_and2_1 _23918_ (.A(_16512_),
    .B(_16954_),
    .X(_16955_));
 sg13g2_a21oi_1 _23919_ (.A1(_16512_),
    .A2(_16954_),
    .Y(_16956_),
    .B1(_15001_));
 sg13g2_o21ai_1 _23920_ (.B1(_14999_),
    .Y(_16957_),
    .A1(_16501_),
    .A2(_16956_));
 sg13g2_a21o_1 _23921_ (.A2(_16957_),
    .A1(_16500_),
    .B1(_14996_),
    .X(_16958_));
 sg13g2_a21oi_1 _23922_ (.A1(_16504_),
    .A2(_16958_),
    .Y(_16959_),
    .B1(_14993_));
 sg13g2_nand3_1 _23923_ (.B(_16504_),
    .C(_16958_),
    .A(_14993_),
    .Y(_16960_));
 sg13g2_nor2_1 _23924_ (.A(net5066),
    .B(_16959_),
    .Y(_16961_));
 sg13g2_a21oi_1 _23925_ (.A1(_15760_),
    .A2(_15764_),
    .Y(_16962_),
    .B1(_15769_));
 sg13g2_or2_1 _23926_ (.X(_16963_),
    .B(_16962_),
    .A(_14964_));
 sg13g2_o21ai_1 _23927_ (.B1(_15770_),
    .Y(_16964_),
    .A1(_15761_),
    .A2(_15763_));
 sg13g2_a21oi_2 _23928_ (.B1(_15013_),
    .Y(_16965_),
    .A2(_16964_),
    .A1(_14992_));
 sg13g2_a21oi_1 _23929_ (.A1(_15010_),
    .A2(_16965_),
    .Y(_16966_),
    .B1(_15023_));
 sg13g2_a21o_1 _23930_ (.A2(_16965_),
    .A1(_15010_),
    .B1(_15023_),
    .X(_16967_));
 sg13g2_a21oi_1 _23931_ (.A1(_15009_),
    .A2(_16967_),
    .Y(_16968_),
    .B1(_15021_));
 sg13g2_a21o_1 _23932_ (.A2(_16967_),
    .A1(_15009_),
    .B1(_15021_),
    .X(_16969_));
 sg13g2_a21oi_1 _23933_ (.A1(_15003_),
    .A2(_16969_),
    .Y(_16970_),
    .B1(_15017_));
 sg13g2_o21ai_1 _23934_ (.B1(_14994_),
    .Y(_16971_),
    .A1(_14995_),
    .A2(_16970_));
 sg13g2_xnor2_1 _23935_ (.Y(_16972_),
    .A(_14993_),
    .B(_16971_));
 sg13g2_o21ai_1 _23936_ (.B1(net5066),
    .Y(_16973_),
    .A1(\u_inv.f_next[175] ),
    .A2(net5777));
 sg13g2_a21oi_1 _23937_ (.A1(net5778),
    .A2(_16972_),
    .Y(_16974_),
    .B1(_16973_));
 sg13g2_a21o_2 _23938_ (.A2(_16961_),
    .A1(_16960_),
    .B1(_16974_),
    .X(_16975_));
 sg13g2_a21o_1 _23939_ (.A2(_16717_),
    .A1(_14865_),
    .B1(_14861_),
    .X(_16976_));
 sg13g2_nand3_1 _23940_ (.B(_14865_),
    .C(_16717_),
    .A(_14861_),
    .Y(_16977_));
 sg13g2_a21oi_1 _23941_ (.A1(_16976_),
    .A2(_16977_),
    .Y(_16978_),
    .B1(net5674));
 sg13g2_o21ai_1 _23942_ (.B1(net5042),
    .Y(_16979_),
    .A1(\u_inv.f_next[218] ),
    .A2(net5752));
 sg13g2_nor3_1 _23943_ (.A(_14861_),
    .B(_15990_),
    .C(_16705_),
    .Y(_16980_));
 sg13g2_o21ai_1 _23944_ (.B1(_14861_),
    .Y(_16981_),
    .A1(_15990_),
    .A2(_16705_));
 sg13g2_nor2_1 _23945_ (.A(net5042),
    .B(_16980_),
    .Y(_16982_));
 sg13g2_nand2_1 _23946_ (.Y(_16983_),
    .A(_16981_),
    .B(_16982_));
 sg13g2_o21ai_1 _23947_ (.B1(_16983_),
    .Y(_16984_),
    .A1(_16978_),
    .A2(_16979_));
 sg13g2_xnor2_1 _23948_ (.Y(_16985_),
    .A(_15858_),
    .B(_16735_));
 sg13g2_a21oi_1 _23949_ (.A1(net5751),
    .A2(_16985_),
    .Y(_16986_),
    .B1(net4941));
 sg13g2_o21ai_1 _23950_ (.B1(_16986_),
    .Y(_16987_),
    .A1(\u_inv.f_next[228] ),
    .A2(net5752));
 sg13g2_nor2_1 _23951_ (.A(_15859_),
    .B(_16726_),
    .Y(_16988_));
 sg13g2_nand2_1 _23952_ (.Y(_16989_),
    .A(net4942),
    .B(_16727_));
 sg13g2_o21ai_1 _23953_ (.B1(_16987_),
    .Y(_16990_),
    .A1(_16988_),
    .A2(_16989_));
 sg13g2_a21oi_1 _23954_ (.A1(_15026_),
    .A2(_16851_),
    .Y(_16991_),
    .B1(_14955_));
 sg13g2_a21oi_1 _23955_ (.A1(_15026_),
    .A2(_16851_),
    .Y(_16992_),
    .B1(_14958_));
 sg13g2_nor2_1 _23956_ (.A(_15039_),
    .B(_16992_),
    .Y(_16993_));
 sg13g2_a21oi_2 _23957_ (.B1(_15041_),
    .Y(_16994_),
    .A2(_16992_),
    .A1(_14952_));
 sg13g2_o21ai_1 _23958_ (.B1(_15044_),
    .Y(_16995_),
    .A1(_14944_),
    .A2(_16994_));
 sg13g2_nand2_1 _23959_ (.Y(_16996_),
    .A(_14937_),
    .B(_16995_));
 sg13g2_and2_1 _23960_ (.A(_14936_),
    .B(_16996_),
    .X(_16997_));
 sg13g2_a21oi_1 _23961_ (.A1(_14935_),
    .A2(_16997_),
    .Y(_16998_),
    .B1(net5680));
 sg13g2_o21ai_1 _23962_ (.B1(_16998_),
    .Y(_16999_),
    .A1(_14935_),
    .A2(_16997_));
 sg13g2_a21oi_1 _23963_ (.A1(_13991_),
    .A2(net5680),
    .Y(_17000_),
    .B1(net4963));
 sg13g2_o21ai_1 _23964_ (.B1(_16468_),
    .Y(_17001_),
    .A1(_16514_),
    .A2(_16860_));
 sg13g2_a21oi_1 _23965_ (.A1(_16538_),
    .A2(_17001_),
    .Y(_17002_),
    .B1(_14943_));
 sg13g2_nand2b_1 _23966_ (.Y(_17003_),
    .B(_17002_),
    .A_N(_14940_));
 sg13g2_nand2b_1 _23967_ (.Y(_17004_),
    .B(_17003_),
    .A_N(_16530_));
 sg13g2_a21oi_1 _23968_ (.A1(_14938_),
    .A2(_17004_),
    .Y(_17005_),
    .B1(_16527_));
 sg13g2_nor2_1 _23969_ (.A(_14935_),
    .B(_17005_),
    .Y(_17006_));
 sg13g2_nand2_1 _23970_ (.Y(_17007_),
    .A(_14935_),
    .B(_17005_));
 sg13g2_nor2_1 _23971_ (.A(net5056),
    .B(_17006_),
    .Y(_17008_));
 sg13g2_and2_1 _23972_ (.A(_17007_),
    .B(_17008_),
    .X(_17009_));
 sg13g2_a22oi_1 _23973_ (.Y(_17010_),
    .B1(_17007_),
    .B2(_17008_),
    .A2(_17000_),
    .A1(_16999_));
 sg13g2_a21o_1 _23974_ (.A2(_17000_),
    .A1(_16999_),
    .B1(_17009_),
    .X(_17011_));
 sg13g2_nand2b_1 _23975_ (.Y(_17012_),
    .B(_14902_),
    .A_N(_16714_));
 sg13g2_o21ai_1 _23976_ (.B1(_14890_),
    .Y(_17013_),
    .A1(_14903_),
    .A2(_16714_));
 sg13g2_a21oi_1 _23977_ (.A1(_14907_),
    .A2(_17013_),
    .Y(_17014_),
    .B1(_14882_));
 sg13g2_nand3_1 _23978_ (.B(_14907_),
    .C(_17013_),
    .A(_14882_),
    .Y(_17015_));
 sg13g2_nor2b_1 _23979_ (.A(_17014_),
    .B_N(_17015_),
    .Y(_17016_));
 sg13g2_nor2_1 _23980_ (.A(\u_inv.f_next[214] ),
    .B(net5754),
    .Y(_17017_));
 sg13g2_o21ai_1 _23981_ (.B1(net5044),
    .Y(_17018_),
    .A1(net5672),
    .A2(_17016_));
 sg13g2_a21o_1 _23982_ (.A2(_16595_),
    .A1(_16561_),
    .B1(_15983_),
    .X(_17019_));
 sg13g2_and2_1 _23983_ (.A(_16008_),
    .B(_17019_),
    .X(_17020_));
 sg13g2_a21oi_1 _23984_ (.A1(_16008_),
    .A2(_17019_),
    .Y(_17021_),
    .B1(_15979_));
 sg13g2_nand3b_1 _23985_ (.B(_16010_),
    .C(_14881_),
    .Y(_17022_),
    .A_N(_17021_));
 sg13g2_o21ai_1 _23986_ (.B1(_14882_),
    .Y(_17023_),
    .A1(_16011_),
    .A2(_17021_));
 sg13g2_nand3_1 _23987_ (.B(_17022_),
    .C(_17023_),
    .A(net4953),
    .Y(_17024_));
 sg13g2_o21ai_1 _23988_ (.B1(_17024_),
    .Y(_17025_),
    .A1(_17017_),
    .A2(_17018_));
 sg13g2_o21ai_1 _23989_ (.B1(_15794_),
    .Y(_17026_),
    .A1(_16483_),
    .A2(_16547_));
 sg13g2_a21oi_1 _23990_ (.A1(_16567_),
    .A2(_17026_),
    .Y(_17027_),
    .B1(_15791_));
 sg13g2_o21ai_1 _23991_ (.B1(_15786_),
    .Y(_17028_),
    .A1(_16566_),
    .A2(_17027_));
 sg13g2_nor2b_1 _23992_ (.A(_16565_),
    .B_N(_17028_),
    .Y(_17029_));
 sg13g2_a21oi_1 _23993_ (.A1(_15787_),
    .A2(_17029_),
    .Y(_17030_),
    .B1(net5053));
 sg13g2_o21ai_1 _23994_ (.B1(_17030_),
    .Y(_17031_),
    .A1(_15787_),
    .A2(_17029_));
 sg13g2_a21oi_1 _23995_ (.A1(_15049_),
    .A2(_15773_),
    .Y(_17032_),
    .B1(_15794_));
 sg13g2_a21o_1 _23996_ (.A2(_15773_),
    .A1(_15049_),
    .B1(_15795_),
    .X(_17033_));
 sg13g2_and2_1 _23997_ (.A(_15826_),
    .B(_17033_),
    .X(_17034_));
 sg13g2_o21ai_1 _23998_ (.B1(_15784_),
    .Y(_17035_),
    .A1(_15786_),
    .A2(_17034_));
 sg13g2_xnor2_1 _23999_ (.Y(_17036_),
    .A(_15787_),
    .B(_17035_));
 sg13g2_a21oi_1 _24000_ (.A1(net5763),
    .A2(_17036_),
    .Y(_17037_),
    .B1(net4961));
 sg13g2_o21ai_1 _24001_ (.B1(_17037_),
    .Y(_17038_),
    .A1(\u_inv.f_next[195] ),
    .A2(net5763));
 sg13g2_nand2_2 _24002_ (.Y(_17039_),
    .A(_17031_),
    .B(_17038_));
 sg13g2_a21oi_1 _24003_ (.A1(_15826_),
    .A2(_17033_),
    .Y(_17040_),
    .B1(_15790_));
 sg13g2_a21o_1 _24004_ (.A2(_17033_),
    .A1(_15826_),
    .B1(_15790_),
    .X(_17041_));
 sg13g2_nand2_1 _24005_ (.Y(_17042_),
    .A(_15829_),
    .B(_17041_));
 sg13g2_a21oi_1 _24006_ (.A1(_15829_),
    .A2(_17041_),
    .Y(_17043_),
    .B1(_15781_));
 sg13g2_o21ai_1 _24007_ (.B1(_15778_),
    .Y(_17044_),
    .A1(_15779_),
    .A2(_17043_));
 sg13g2_nor3_1 _24008_ (.A(_15778_),
    .B(_15779_),
    .C(_17043_),
    .Y(_17045_));
 sg13g2_nand3b_1 _24009_ (.B(net5762),
    .C(_17044_),
    .Y(_17046_),
    .A_N(_17045_));
 sg13g2_a21oi_1 _24010_ (.A1(_13977_),
    .A2(net5681),
    .Y(_17047_),
    .B1(net4961));
 sg13g2_o21ai_1 _24011_ (.B1(_16551_),
    .Y(_17048_),
    .A1(_16483_),
    .A2(_16547_));
 sg13g2_a21oi_1 _24012_ (.A1(_16570_),
    .A2(_17048_),
    .Y(_17049_),
    .B1(_15780_));
 sg13g2_or3_1 _24013_ (.A(_15778_),
    .B(_16563_),
    .C(_17049_),
    .X(_17050_));
 sg13g2_o21ai_1 _24014_ (.B1(_15778_),
    .Y(_17051_),
    .A1(_16563_),
    .A2(_17049_));
 sg13g2_and2_1 _24015_ (.A(net4965),
    .B(_17051_),
    .X(_17052_));
 sg13g2_a22oi_1 _24016_ (.Y(_17053_),
    .B1(_17050_),
    .B2(_17052_),
    .A2(_17047_),
    .A1(_17046_));
 sg13g2_inv_1 _24017_ (.Y(_17054_),
    .A(_17053_));
 sg13g2_a21oi_1 _24018_ (.A1(_15049_),
    .A2(_15773_),
    .Y(_17055_),
    .B1(_15797_));
 sg13g2_nor2_1 _24019_ (.A(_15835_),
    .B(_17055_),
    .Y(_17056_));
 sg13g2_o21ai_1 _24020_ (.B1(_15811_),
    .Y(_17057_),
    .A1(_15835_),
    .A2(_17055_));
 sg13g2_o21ai_1 _24021_ (.B1(_17057_),
    .Y(_17058_),
    .A1(_13974_),
    .A2(_14454_));
 sg13g2_xor2_1 _24022_ (.B(_17058_),
    .A(_15813_),
    .X(_17059_));
 sg13g2_o21ai_1 _24023_ (.B1(net5052),
    .Y(_17060_),
    .A1(\u_inv.f_next[201] ),
    .A2(net5762));
 sg13g2_a21oi_1 _24024_ (.A1(net5762),
    .A2(_17059_),
    .Y(_17061_),
    .B1(_17060_));
 sg13g2_o21ai_1 _24025_ (.B1(_16554_),
    .Y(_17062_),
    .A1(_16483_),
    .A2(_16547_));
 sg13g2_a21oi_1 _24026_ (.A1(_16576_),
    .A2(_17062_),
    .Y(_17063_),
    .B1(_15811_));
 sg13g2_nor3_1 _24027_ (.A(_15813_),
    .B(_16589_),
    .C(_17063_),
    .Y(_17064_));
 sg13g2_o21ai_1 _24028_ (.B1(_15813_),
    .Y(_17065_),
    .A1(_16589_),
    .A2(_17063_));
 sg13g2_nor2_1 _24029_ (.A(net5052),
    .B(_17064_),
    .Y(_17066_));
 sg13g2_a21oi_1 _24030_ (.A1(_17065_),
    .A2(_17066_),
    .Y(_17067_),
    .B1(_17061_));
 sg13g2_nand2_2 _24031_ (.Y(_17068_),
    .A(_16423_),
    .B(_16457_));
 sg13g2_a21o_1 _24032_ (.A2(_16457_),
    .A1(_16423_),
    .B1(_16061_),
    .X(_17069_));
 sg13g2_a21oi_1 _24033_ (.A1(_16033_),
    .A2(_17069_),
    .Y(_17070_),
    .B1(_16026_));
 sg13g2_o21ai_1 _24034_ (.B1(_15072_),
    .Y(_17071_),
    .A1(_16024_),
    .A2(_17070_));
 sg13g2_o21ai_1 _24035_ (.B1(_16039_),
    .Y(_17072_),
    .A1(_16024_),
    .A2(_17070_));
 sg13g2_o21ai_1 _24036_ (.B1(_16049_),
    .Y(_17073_),
    .A1(_16038_),
    .A2(_17072_));
 sg13g2_nand2b_1 _24037_ (.Y(_17074_),
    .B(_17073_),
    .A_N(_15058_));
 sg13g2_xor2_1 _24038_ (.B(_17073_),
    .A(_15058_),
    .X(_17075_));
 sg13g2_a21o_1 _24039_ (.A2(_15758_),
    .A1(_15736_),
    .B1(_15095_),
    .X(_17076_));
 sg13g2_a21oi_1 _24040_ (.A1(_15736_),
    .A2(_15758_),
    .Y(_17077_),
    .B1(_15096_));
 sg13g2_nor2_1 _24041_ (.A(_15117_),
    .B(_17077_),
    .Y(_17078_));
 sg13g2_or2_1 _24042_ (.X(_17079_),
    .B(_17077_),
    .A(_15117_));
 sg13g2_o21ai_1 _24043_ (.B1(_15094_),
    .Y(_17080_),
    .A1(_15117_),
    .A2(_17077_));
 sg13g2_a21o_1 _24044_ (.A2(_17080_),
    .A1(_15112_),
    .B1(_15072_),
    .X(_17081_));
 sg13g2_a21o_2 _24045_ (.A2(_17080_),
    .A1(_15112_),
    .B1(_15074_),
    .X(_17082_));
 sg13g2_o21ai_1 _24046_ (.B1(_15102_),
    .Y(_17083_),
    .A1(_15068_),
    .A2(_17082_));
 sg13g2_xor2_1 _24047_ (.B(_17083_),
    .A(_15058_),
    .X(_17084_));
 sg13g2_o21ai_1 _24048_ (.B1(net5068),
    .Y(_17085_),
    .A1(_14018_),
    .A2(net5783));
 sg13g2_a21oi_1 _24049_ (.A1(net5783),
    .A2(_17084_),
    .Y(_17086_),
    .B1(_17085_));
 sg13g2_a21oi_2 _24050_ (.B1(_17086_),
    .Y(_17087_),
    .A2(_17075_),
    .A1(net4978));
 sg13g2_o21ai_1 _24051_ (.B1(_14955_),
    .Y(_17088_),
    .A1(_16514_),
    .A2(_16860_));
 sg13g2_a21oi_1 _24052_ (.A1(_16532_),
    .A2(_17088_),
    .Y(_17089_),
    .B1(_14956_));
 sg13g2_o21ai_1 _24053_ (.B1(_14950_),
    .Y(_17090_),
    .A1(_16534_),
    .A2(_17089_));
 sg13g2_a21o_1 _24054_ (.A2(_17090_),
    .A1(_16533_),
    .B1(_14947_),
    .X(_17091_));
 sg13g2_nand3_1 _24055_ (.B(_16533_),
    .C(_17090_),
    .A(_14947_),
    .Y(_17092_));
 sg13g2_nand3_1 _24056_ (.B(_17091_),
    .C(_17092_),
    .A(net4975),
    .Y(_17093_));
 sg13g2_o21ai_1 _24057_ (.B1(_14948_),
    .Y(_17094_),
    .A1(_14950_),
    .A2(_16993_));
 sg13g2_xor2_1 _24058_ (.B(_17094_),
    .A(_14947_),
    .X(_17095_));
 sg13g2_nor2_1 _24059_ (.A(net5689),
    .B(_17095_),
    .Y(_17096_));
 sg13g2_o21ai_1 _24060_ (.B1(net5056),
    .Y(_17097_),
    .A1(\u_inv.f_next[179] ),
    .A2(net5777));
 sg13g2_o21ai_1 _24061_ (.B1(_17093_),
    .Y(_17098_),
    .A1(_17096_),
    .A2(_17097_));
 sg13g2_nor2_1 _24062_ (.A(_16519_),
    .B(_16862_),
    .Y(_17099_));
 sg13g2_o21ai_1 _24063_ (.B1(net5622),
    .Y(_17100_),
    .A1(_16519_),
    .A2(_16862_));
 sg13g2_nand2b_1 _24064_ (.Y(_17101_),
    .B(_17100_),
    .A_N(_16516_));
 sg13g2_a21oi_1 _24065_ (.A1(net5623),
    .A2(_17101_),
    .Y(_17102_),
    .B1(net5055));
 sg13g2_o21ai_1 _24066_ (.B1(_17102_),
    .Y(_17103_),
    .A1(net5623),
    .A2(_17101_));
 sg13g2_a21oi_1 _24067_ (.A1(_15029_),
    .A2(_16854_),
    .Y(_17104_),
    .B1(net5622));
 sg13g2_a21oi_1 _24068_ (.A1(\u_inv.f_next[186] ),
    .A2(\u_inv.f_reg[186] ),
    .Y(_17105_),
    .B1(_17104_));
 sg13g2_xor2_1 _24069_ (.B(_17105_),
    .A(_14926_),
    .X(_17106_));
 sg13g2_nor2_1 _24070_ (.A(net5682),
    .B(_17106_),
    .Y(_17107_));
 sg13g2_o21ai_1 _24071_ (.B1(net5055),
    .Y(_17108_),
    .A1(\u_inv.f_next[187] ),
    .A2(net5766));
 sg13g2_o21ai_1 _24072_ (.B1(_17103_),
    .Y(_17109_),
    .A1(_17107_),
    .A2(_17108_));
 sg13g2_a21oi_1 _24073_ (.A1(_15059_),
    .A2(_17083_),
    .Y(_17110_),
    .B1(_15105_));
 sg13g2_xnor2_1 _24074_ (.Y(_17111_),
    .A(_15052_),
    .B(_17110_));
 sg13g2_nor2_1 _24075_ (.A(\u_inv.f_next[158] ),
    .B(net5783),
    .Y(_17112_));
 sg13g2_o21ai_1 _24076_ (.B1(net5068),
    .Y(_17113_),
    .A1(net5698),
    .A2(_17111_));
 sg13g2_nand2_1 _24077_ (.Y(_17114_),
    .A(_16036_),
    .B(_17073_));
 sg13g2_nand3_1 _24078_ (.B(_16053_),
    .C(_17114_),
    .A(_15052_),
    .Y(_17115_));
 sg13g2_a21o_1 _24079_ (.A2(_17114_),
    .A1(_16053_),
    .B1(_15052_),
    .X(_17116_));
 sg13g2_nand3_1 _24080_ (.B(_17115_),
    .C(_17116_),
    .A(net4978),
    .Y(_17117_));
 sg13g2_o21ai_1 _24081_ (.B1(_17117_),
    .Y(_17118_),
    .A1(_17112_),
    .A2(_17113_));
 sg13g2_o21ai_1 _24082_ (.B1(_15000_),
    .Y(_17119_),
    .A1(_15002_),
    .A2(_16968_));
 sg13g2_xor2_1 _24083_ (.B(_17119_),
    .A(_14999_),
    .X(_17120_));
 sg13g2_o21ai_1 _24084_ (.B1(net5066),
    .Y(_17121_),
    .A1(\u_inv.f_next[173] ),
    .A2(net5778));
 sg13g2_a21oi_1 _24085_ (.A1(net5778),
    .A2(_17120_),
    .Y(_17122_),
    .B1(_17121_));
 sg13g2_nor3_1 _24086_ (.A(_14999_),
    .B(_16501_),
    .C(_16956_),
    .Y(_17123_));
 sg13g2_nor2_1 _24087_ (.A(net5066),
    .B(_17123_),
    .Y(_17124_));
 sg13g2_a21o_2 _24088_ (.A2(_17124_),
    .A1(_16957_),
    .B1(_17122_),
    .X(_17125_));
 sg13g2_o21ai_1 _24089_ (.B1(_15820_),
    .Y(_17126_),
    .A1(_15835_),
    .A2(_17055_));
 sg13g2_nand2_1 _24090_ (.Y(_17127_),
    .A(_15840_),
    .B(_17126_));
 sg13g2_a21oi_1 _24091_ (.A1(_15809_),
    .A2(_17127_),
    .Y(_17128_),
    .B1(_15842_));
 sg13g2_nand2b_1 _24092_ (.Y(_17129_),
    .B(_15799_),
    .A_N(_17128_));
 sg13g2_xnor2_1 _24093_ (.Y(_17130_),
    .A(_15800_),
    .B(_17128_));
 sg13g2_o21ai_1 _24094_ (.B1(net5045),
    .Y(_17131_),
    .A1(\u_inv.f_next[206] ),
    .A2(net5756));
 sg13g2_a21oi_1 _24095_ (.A1(net5756),
    .A2(_17130_),
    .Y(_17132_),
    .B1(_17131_));
 sg13g2_a21oi_1 _24096_ (.A1(_16576_),
    .A2(_17062_),
    .Y(_17133_),
    .B1(_16557_));
 sg13g2_nor2b_2 _24097_ (.A(_17133_),
    .B_N(_16593_),
    .Y(_17134_));
 sg13g2_nor2_1 _24098_ (.A(_16555_),
    .B(_17134_),
    .Y(_17135_));
 sg13g2_o21ai_1 _24099_ (.B1(_16580_),
    .Y(_17136_),
    .A1(_16555_),
    .A2(_17134_));
 sg13g2_xnor2_1 _24100_ (.Y(_17137_),
    .A(_15799_),
    .B(_17136_));
 sg13g2_a21oi_1 _24101_ (.A1(net4954),
    .A2(_17137_),
    .Y(_17138_),
    .B1(_17132_));
 sg13g2_inv_2 _24102_ (.Y(_17139_),
    .A(_17138_));
 sg13g2_o21ai_1 _24103_ (.B1(_15837_),
    .Y(_17140_),
    .A1(_15813_),
    .A2(_17057_));
 sg13g2_xnor2_1 _24104_ (.Y(_17141_),
    .A(_15816_),
    .B(_17140_));
 sg13g2_nor2_1 _24105_ (.A(\u_inv.f_next[202] ),
    .B(net5755),
    .Y(_17142_));
 sg13g2_o21ai_1 _24106_ (.B1(net5045),
    .Y(_17143_),
    .A1(net5672),
    .A2(_17141_));
 sg13g2_nand3_1 _24107_ (.B(_16588_),
    .C(_17065_),
    .A(_15815_),
    .Y(_17144_));
 sg13g2_a21o_1 _24108_ (.A2(_17065_),
    .A1(_16588_),
    .B1(_15815_),
    .X(_17145_));
 sg13g2_nand3_1 _24109_ (.B(_17144_),
    .C(_17145_),
    .A(net4953),
    .Y(_17146_));
 sg13g2_o21ai_1 _24110_ (.B1(_17146_),
    .Y(_17147_),
    .A1(_17142_),
    .A2(_17143_));
 sg13g2_a21oi_1 _24111_ (.A1(_16561_),
    .A2(_16595_),
    .Y(_17148_),
    .B1(_14913_));
 sg13g2_o21ai_1 _24112_ (.B1(_14912_),
    .Y(_17149_),
    .A1(_16003_),
    .A2(_17148_));
 sg13g2_nand2_1 _24113_ (.Y(_17150_),
    .A(_16002_),
    .B(_17149_));
 sg13g2_xnor2_1 _24114_ (.Y(_17151_),
    .A(_14894_),
    .B(_17150_));
 sg13g2_nand3_1 _24115_ (.B(_14898_),
    .C(_16713_),
    .A(_14894_),
    .Y(_17152_));
 sg13g2_a21oi_1 _24116_ (.A1(_14898_),
    .A2(_16713_),
    .Y(_17153_),
    .B1(_14894_));
 sg13g2_nand3b_1 _24117_ (.B(net5755),
    .C(_17152_),
    .Y(_17154_),
    .A_N(_17153_));
 sg13g2_a21oi_1 _24118_ (.A1(\u_inv.f_next[210] ),
    .A2(net5673),
    .Y(_17155_),
    .B1(net4954));
 sg13g2_a22oi_1 _24119_ (.Y(_17156_),
    .B1(_17154_),
    .B2(_17155_),
    .A2(_17151_),
    .A1(net4953));
 sg13g2_a21oi_1 _24120_ (.A1(_15782_),
    .A2(_17042_),
    .Y(_17157_),
    .B1(_15833_));
 sg13g2_nand2b_1 _24121_ (.Y(_17158_),
    .B(_15775_),
    .A_N(_17157_));
 sg13g2_xor2_1 _24122_ (.B(_17157_),
    .A(_15775_),
    .X(_17159_));
 sg13g2_o21ai_1 _24123_ (.B1(net5052),
    .Y(_17160_),
    .A1(\u_inv.f_next[198] ),
    .A2(net5762));
 sg13g2_a21oi_1 _24124_ (.A1(net5762),
    .A2(_17159_),
    .Y(_17161_),
    .B1(_17160_));
 sg13g2_nand3_1 _24125_ (.B(_16562_),
    .C(_17051_),
    .A(_15775_),
    .Y(_17162_));
 sg13g2_a21oi_1 _24126_ (.A1(_16562_),
    .A2(_17051_),
    .Y(_17163_),
    .B1(_15775_));
 sg13g2_nor2_1 _24127_ (.A(net5052),
    .B(_17163_),
    .Y(_17164_));
 sg13g2_a21o_1 _24128_ (.A2(_17164_),
    .A1(_17162_),
    .B1(_17161_),
    .X(_17165_));
 sg13g2_nor2_1 _24129_ (.A(_16490_),
    .B(_16949_),
    .Y(_17166_));
 sg13g2_o21ai_1 _24130_ (.B1(_14971_),
    .Y(_17167_),
    .A1(_16490_),
    .A2(_16949_));
 sg13g2_a21oi_1 _24131_ (.A1(_16492_),
    .A2(_17167_),
    .Y(_17168_),
    .B1(_14972_));
 sg13g2_o21ai_1 _24132_ (.B1(_14968_),
    .Y(_17169_),
    .A1(_16491_),
    .A2(_17168_));
 sg13g2_nand2b_1 _24133_ (.Y(_17170_),
    .B(_17169_),
    .A_N(_16495_));
 sg13g2_o21ai_1 _24134_ (.B1(net4978),
    .Y(_17171_),
    .A1(_14966_),
    .A2(_17170_));
 sg13g2_a21oi_1 _24135_ (.A1(_14966_),
    .A2(_17170_),
    .Y(_17172_),
    .B1(_17171_));
 sg13g2_o21ai_1 _24136_ (.B1(_14980_),
    .Y(_17173_),
    .A1(_14964_),
    .A2(_16962_));
 sg13g2_and2_1 _24137_ (.A(_14988_),
    .B(_17173_),
    .X(_17174_));
 sg13g2_a21o_1 _24138_ (.A2(_17173_),
    .A1(_14988_),
    .B1(_14975_),
    .X(_17175_));
 sg13g2_a21o_1 _24139_ (.A2(_17175_),
    .A1(_14983_),
    .B1(_14968_),
    .X(_17176_));
 sg13g2_nand2_1 _24140_ (.Y(_17177_),
    .A(_14967_),
    .B(_17176_));
 sg13g2_xnor2_1 _24141_ (.Y(_17178_),
    .A(_14965_),
    .B(_17177_));
 sg13g2_o21ai_1 _24142_ (.B1(net5068),
    .Y(_17179_),
    .A1(\u_inv.f_next[167] ),
    .A2(net5782));
 sg13g2_a21oi_1 _24143_ (.A1(net5782),
    .A2(_17178_),
    .Y(_17180_),
    .B1(_17179_));
 sg13g2_or2_1 _24144_ (.X(_17181_),
    .B(_17180_),
    .A(_17172_));
 sg13g2_nand3_1 _24145_ (.B(_15906_),
    .C(_16734_),
    .A(_15872_),
    .Y(_17182_));
 sg13g2_a21oi_1 _24146_ (.A1(_16826_),
    .A2(_17182_),
    .Y(_17183_),
    .B1(net5665));
 sg13g2_a21oi_1 _24147_ (.A1(_13948_),
    .A2(net5666),
    .Y(_17184_),
    .B1(_17183_));
 sg13g2_or3_1 _24148_ (.A(_15872_),
    .B(_16617_),
    .C(_16725_),
    .X(_17185_));
 sg13g2_and2_1 _24149_ (.A(_16822_),
    .B(_17185_),
    .X(_17186_));
 sg13g2_mux2_1 _24150_ (.A0(_17184_),
    .A1(_17186_),
    .S(net4942),
    .X(_17187_));
 sg13g2_a21oi_1 _24151_ (.A1(_15915_),
    .A2(_16691_),
    .Y(_17188_),
    .B1(_15892_));
 sg13g2_and3_1 _24152_ (.X(_17189_),
    .A(_15892_),
    .B(_15915_),
    .C(_16691_));
 sg13g2_nor2_1 _24153_ (.A(_13942_),
    .B(net5741),
    .Y(_17190_));
 sg13g2_nor3_1 _24154_ (.A(net5665),
    .B(_17188_),
    .C(_17189_),
    .Y(_17191_));
 sg13g2_xnor2_1 _24155_ (.Y(_17192_),
    .A(_15893_),
    .B(_16683_));
 sg13g2_nor3_1 _24156_ (.A(net4942),
    .B(_17190_),
    .C(_17191_),
    .Y(_17193_));
 sg13g2_a21oi_2 _24157_ (.B1(_17193_),
    .Y(_17194_),
    .A2(_17192_),
    .A1(net4942));
 sg13g2_a21oi_1 _24158_ (.A1(_16033_),
    .A2(_17069_),
    .Y(_17195_),
    .B1(_15092_));
 sg13g2_o21ai_1 _24159_ (.B1(_15090_),
    .Y(_17196_),
    .A1(_16020_),
    .A2(_17195_));
 sg13g2_a21oi_1 _24160_ (.A1(_16019_),
    .A2(_17196_),
    .Y(_17197_),
    .B1(_15087_));
 sg13g2_nor2_1 _24161_ (.A(_16018_),
    .B(_17197_),
    .Y(_17198_));
 sg13g2_o21ai_1 _24162_ (.B1(net4988),
    .Y(_17199_),
    .A1(_15085_),
    .A2(_17198_));
 sg13g2_a21oi_1 _24163_ (.A1(_15085_),
    .A2(_17198_),
    .Y(_17200_),
    .B1(_17199_));
 sg13g2_o21ai_1 _24164_ (.B1(_15109_),
    .Y(_17201_),
    .A1(_15093_),
    .A2(_17078_));
 sg13g2_nand2_1 _24165_ (.Y(_17202_),
    .A(_15087_),
    .B(_17201_));
 sg13g2_nand2_1 _24166_ (.Y(_17203_),
    .A(_15086_),
    .B(_17202_));
 sg13g2_xnor2_1 _24167_ (.Y(_17204_),
    .A(_15085_),
    .B(_17203_));
 sg13g2_o21ai_1 _24168_ (.B1(net5074),
    .Y(_17205_),
    .A1(\u_inv.f_next[151] ),
    .A2(net5791));
 sg13g2_a21oi_1 _24169_ (.A1(net5791),
    .A2(_17204_),
    .Y(_17206_),
    .B1(_17205_));
 sg13g2_or2_1 _24170_ (.X(_17207_),
    .B(_17206_),
    .A(_17200_));
 sg13g2_o21ai_1 _24171_ (.B1(_15008_),
    .Y(_17208_),
    .A1(_16508_),
    .A2(_16952_));
 sg13g2_a21oi_1 _24172_ (.A1(_16509_),
    .A2(_17208_),
    .Y(_17209_),
    .B1(_15005_));
 sg13g2_nand3_1 _24173_ (.B(_16509_),
    .C(_17208_),
    .A(_15005_),
    .Y(_17210_));
 sg13g2_nand2_1 _24174_ (.Y(_17211_),
    .A(net4976),
    .B(_17210_));
 sg13g2_o21ai_1 _24175_ (.B1(_15007_),
    .Y(_17212_),
    .A1(_15008_),
    .A2(_16966_));
 sg13g2_xnor2_1 _24176_ (.Y(_17213_),
    .A(_15005_),
    .B(_17212_));
 sg13g2_a21oi_1 _24177_ (.A1(net5779),
    .A2(_17213_),
    .Y(_17214_),
    .B1(net4976));
 sg13g2_o21ai_1 _24178_ (.B1(_17214_),
    .Y(_17215_),
    .A1(\u_inv.f_next[171] ),
    .A2(net5779));
 sg13g2_o21ai_1 _24179_ (.B1(_17215_),
    .Y(_17216_),
    .A1(_17209_),
    .A2(_17211_));
 sg13g2_a21oi_2 _24180_ (.B1(_16441_),
    .Y(_17217_),
    .A2(_16417_),
    .A1(_16414_));
 sg13g2_o21ai_1 _24181_ (.B1(_16448_),
    .Y(_17218_),
    .A1(_16420_),
    .A2(_17217_));
 sg13g2_nand2_1 _24182_ (.Y(_17219_),
    .A(_15693_),
    .B(_17218_));
 sg13g2_a21oi_1 _24183_ (.A1(_16450_),
    .A2(_17219_),
    .Y(_17220_),
    .B1(_15690_));
 sg13g2_o21ai_1 _24184_ (.B1(_15688_),
    .Y(_17221_),
    .A1(_16449_),
    .A2(_17220_));
 sg13g2_nand3_1 _24185_ (.B(_16453_),
    .C(_17221_),
    .A(_15685_),
    .Y(_17222_));
 sg13g2_a21o_1 _24186_ (.A2(_17221_),
    .A1(_16453_),
    .B1(_15685_),
    .X(_17223_));
 sg13g2_nand3_1 _24187_ (.B(_17222_),
    .C(_17223_),
    .A(net4990),
    .Y(_17224_));
 sg13g2_a21oi_1 _24188_ (.A1(_15656_),
    .A2(_15680_),
    .Y(_17225_),
    .B1(_15734_));
 sg13g2_nor2_2 _24189_ (.A(_15740_),
    .B(_17225_),
    .Y(_17226_));
 sg13g2_a21oi_2 _24190_ (.B1(_15745_),
    .Y(_17227_),
    .A2(_17225_),
    .A1(_15721_));
 sg13g2_o21ai_1 _24191_ (.B1(_15753_),
    .Y(_17228_),
    .A1(_15703_),
    .A2(_17227_));
 sg13g2_a21oi_2 _24192_ (.B1(_15755_),
    .Y(_17229_),
    .A2(_17228_),
    .A1(_15708_));
 sg13g2_o21ai_1 _24193_ (.B1(_15748_),
    .Y(_17230_),
    .A1(_15694_),
    .A2(_17229_));
 sg13g2_a21oi_1 _24194_ (.A1(_15687_),
    .A2(_17230_),
    .Y(_17231_),
    .B1(_15686_));
 sg13g2_xnor2_1 _24195_ (.Y(_17232_),
    .A(_15685_),
    .B(_17231_));
 sg13g2_nor2_1 _24196_ (.A(\u_inv.f_next[143] ),
    .B(net5794),
    .Y(_17233_));
 sg13g2_o21ai_1 _24197_ (.B1(net5077),
    .Y(_17234_),
    .A1(net5697),
    .A2(_17232_));
 sg13g2_o21ai_1 _24198_ (.B1(_17224_),
    .Y(_17235_),
    .A1(_17233_),
    .A2(_17234_));
 sg13g2_a21oi_1 _24199_ (.A1(\u_inv.f_next[188] ),
    .A2(_14442_),
    .Y(_17236_),
    .B1(_14923_));
 sg13g2_o21ai_1 _24200_ (.B1(_17236_),
    .Y(_17237_),
    .A1(_14921_),
    .A2(_16863_));
 sg13g2_and4_1 _24201_ (.A(net4962),
    .B(_16522_),
    .C(_16864_),
    .D(_17237_),
    .X(_17238_));
 sg13g2_a21oi_1 _24202_ (.A1(_14921_),
    .A2(_16855_),
    .Y(_17239_),
    .B1(_14920_));
 sg13g2_xnor2_1 _24203_ (.Y(_17240_),
    .A(_14923_),
    .B(_17239_));
 sg13g2_o21ai_1 _24204_ (.B1(net5053),
    .Y(_17241_),
    .A1(\u_inv.f_next[189] ),
    .A2(net5764));
 sg13g2_a21oi_2 _24205_ (.B1(_17241_),
    .Y(_17242_),
    .A2(_17240_),
    .A1(net5763));
 sg13g2_nor2_1 _24206_ (.A(_17238_),
    .B(_17242_),
    .Y(_17243_));
 sg13g2_inv_1 _24207_ (.Y(_17244_),
    .A(_17243_));
 sg13g2_and2_1 _24208_ (.A(_16047_),
    .B(_17072_),
    .X(_17245_));
 sg13g2_o21ai_1 _24209_ (.B1(_16043_),
    .Y(_17246_),
    .A1(_15066_),
    .A2(_17245_));
 sg13g2_o21ai_1 _24210_ (.B1(net4988),
    .Y(_17247_),
    .A1(_15064_),
    .A2(_17246_));
 sg13g2_a21oi_1 _24211_ (.A1(_15064_),
    .A2(_17246_),
    .Y(_17248_),
    .B1(_17247_));
 sg13g2_a21o_1 _24212_ (.A2(_17082_),
    .A1(_15099_),
    .B1(_15067_),
    .X(_17249_));
 sg13g2_nand2_1 _24213_ (.Y(_17250_),
    .A(_15065_),
    .B(_17249_));
 sg13g2_xnor2_1 _24214_ (.Y(_17251_),
    .A(_15063_),
    .B(_17250_));
 sg13g2_o21ai_1 _24215_ (.B1(net5074),
    .Y(_17252_),
    .A1(\u_inv.f_next[155] ),
    .A2(net5791));
 sg13g2_a21oi_1 _24216_ (.A1(net5791),
    .A2(_17251_),
    .Y(_17253_),
    .B1(_17252_));
 sg13g2_or2_1 _24217_ (.X(_17254_),
    .B(_17253_),
    .A(_17248_));
 sg13g2_nand3_1 _24218_ (.B(_16621_),
    .C(_16727_),
    .A(_15856_),
    .Y(_17255_));
 sg13g2_nor3_1 _24219_ (.A(net5035),
    .B(_16622_),
    .C(_16728_),
    .Y(_17256_));
 sg13g2_a21oi_1 _24220_ (.A1(_15858_),
    .A2(_16735_),
    .Y(_17257_),
    .B1(_15857_));
 sg13g2_xor2_1 _24221_ (.B(_17257_),
    .A(_15856_),
    .X(_17258_));
 sg13g2_nand2_1 _24222_ (.Y(_17259_),
    .A(_13945_),
    .B(net5665));
 sg13g2_a21oi_1 _24223_ (.A1(net5739),
    .A2(_17258_),
    .Y(_17260_),
    .B1(net4941));
 sg13g2_a22oi_1 _24224_ (.Y(_17261_),
    .B1(_17259_),
    .B2(_17260_),
    .A2(_17256_),
    .A1(_17255_));
 sg13g2_inv_1 _24225_ (.Y(_17262_),
    .A(_17261_));
 sg13g2_xnor2_1 _24226_ (.Y(_17263_),
    .A(_15883_),
    .B(_16685_));
 sg13g2_a21oi_1 _24227_ (.A1(_15883_),
    .A2(_16693_),
    .Y(_17264_),
    .B1(net5665));
 sg13g2_o21ai_1 _24228_ (.B1(_17264_),
    .Y(_17265_),
    .A1(_15883_),
    .A2(_16693_));
 sg13g2_a21oi_1 _24229_ (.A1(\u_inv.f_next[236] ),
    .A2(net5665),
    .Y(_17266_),
    .B1(net4941));
 sg13g2_a22oi_1 _24230_ (.Y(_17267_),
    .B1(_17265_),
    .B2(_17266_),
    .A2(_17263_),
    .A1(net4941));
 sg13g2_inv_1 _24231_ (.Y(_17268_),
    .A(_17267_));
 sg13g2_xnor2_1 _24232_ (.Y(_17269_),
    .A(_14889_),
    .B(_17012_));
 sg13g2_o21ai_1 _24233_ (.B1(net5044),
    .Y(_17270_),
    .A1(\u_inv.f_next[212] ),
    .A2(net5754));
 sg13g2_a21oi_1 _24234_ (.A1(net5754),
    .A2(_17269_),
    .Y(_17271_),
    .B1(_17270_));
 sg13g2_xnor2_1 _24235_ (.Y(_17272_),
    .A(_14888_),
    .B(_17020_));
 sg13g2_a21oi_1 _24236_ (.A1(net4953),
    .A2(_17272_),
    .Y(_17273_),
    .B1(_17271_));
 sg13g2_inv_2 _24237_ (.Y(_17274_),
    .A(_17273_));
 sg13g2_a21oi_1 _24238_ (.A1(\u_inv.f_next[212] ),
    .A2(_14466_),
    .Y(_17275_),
    .B1(_14886_));
 sg13g2_o21ai_1 _24239_ (.B1(_17275_),
    .Y(_17276_),
    .A1(_14889_),
    .A2(_17020_));
 sg13g2_nor3_1 _24240_ (.A(net5044),
    .B(_16009_),
    .C(_17021_),
    .Y(_17277_));
 sg13g2_a21oi_1 _24241_ (.A1(_14889_),
    .A2(_17012_),
    .Y(_17278_),
    .B1(_14887_));
 sg13g2_xnor2_1 _24242_ (.Y(_17279_),
    .A(_14886_),
    .B(_17278_));
 sg13g2_nand2_1 _24243_ (.Y(_17280_),
    .A(_13961_),
    .B(net5672));
 sg13g2_a21oi_1 _24244_ (.A1(net5754),
    .A2(_17279_),
    .Y(_17281_),
    .B1(net4953));
 sg13g2_a22oi_1 _24245_ (.Y(_17282_),
    .B1(_17280_),
    .B2(_17281_),
    .A2(_17277_),
    .A1(_17276_));
 sg13g2_inv_1 _24246_ (.Y(_17283_),
    .A(_17282_));
 sg13g2_nor2b_1 _24247_ (.A(_15808_),
    .B_N(_16578_),
    .Y(_17284_));
 sg13g2_o21ai_1 _24248_ (.B1(_17284_),
    .Y(_17285_),
    .A1(_15805_),
    .A2(_17134_));
 sg13g2_nor3_1 _24249_ (.A(net5045),
    .B(_16579_),
    .C(_17135_),
    .Y(_17286_));
 sg13g2_a21oi_1 _24250_ (.A1(_15840_),
    .A2(_17126_),
    .Y(_17287_),
    .B1(_15804_));
 sg13g2_o21ai_1 _24251_ (.B1(_15808_),
    .Y(_17288_),
    .A1(_15803_),
    .A2(_17287_));
 sg13g2_or3_1 _24252_ (.A(_15803_),
    .B(_15808_),
    .C(_17287_),
    .X(_17289_));
 sg13g2_nand3_1 _24253_ (.B(_17288_),
    .C(_17289_),
    .A(net5764),
    .Y(_17290_));
 sg13g2_a21oi_1 _24254_ (.A1(_13969_),
    .A2(net5672),
    .Y(_17291_),
    .B1(net4954));
 sg13g2_a22oi_1 _24255_ (.Y(_17292_),
    .B1(_17290_),
    .B2(_17291_),
    .A2(_17286_),
    .A1(_17285_));
 sg13g2_inv_1 _24256_ (.Y(_17293_),
    .A(_17292_));
 sg13g2_or3_1 _24257_ (.A(_15786_),
    .B(_16566_),
    .C(_17027_),
    .X(_17294_));
 sg13g2_nand2_1 _24258_ (.Y(_17295_),
    .A(_17028_),
    .B(_17294_));
 sg13g2_xnor2_1 _24259_ (.Y(_17296_),
    .A(_15785_),
    .B(_17034_));
 sg13g2_o21ai_1 _24260_ (.B1(net5053),
    .Y(_17297_),
    .A1(_13980_),
    .A2(net5763));
 sg13g2_a21oi_1 _24261_ (.A1(net5763),
    .A2(_17296_),
    .Y(_17298_),
    .B1(_17297_));
 sg13g2_a21oi_1 _24262_ (.A1(net4961),
    .A2(_17295_),
    .Y(_17299_),
    .B1(_17298_));
 sg13g2_a21oi_1 _24263_ (.A1(_14988_),
    .A2(_17173_),
    .Y(_17300_),
    .B1(_14971_));
 sg13g2_o21ai_1 _24264_ (.B1(_14973_),
    .Y(_17301_),
    .A1(_14970_),
    .A2(_17300_));
 sg13g2_or3_1 _24265_ (.A(_14970_),
    .B(_14973_),
    .C(_17300_),
    .X(_17302_));
 sg13g2_nand3_1 _24266_ (.B(_17301_),
    .C(_17302_),
    .A(net5782),
    .Y(_17303_));
 sg13g2_a21oi_1 _24267_ (.A1(_14009_),
    .A2(net5691),
    .Y(_17304_),
    .B1(net4977));
 sg13g2_nand3_1 _24268_ (.B(_16492_),
    .C(_17167_),
    .A(_14972_),
    .Y(_17305_));
 sg13g2_nor2_1 _24269_ (.A(net5068),
    .B(_17168_),
    .Y(_17306_));
 sg13g2_a22oi_1 _24270_ (.Y(_17307_),
    .B1(_17305_),
    .B2(_17306_),
    .A2(_17304_),
    .A1(_17303_));
 sg13g2_a21oi_1 _24271_ (.A1(_16381_),
    .A2(_16413_),
    .Y(_17308_),
    .B1(_16415_));
 sg13g2_o21ai_1 _24272_ (.B1(_15720_),
    .Y(_17309_),
    .A1(_16430_),
    .A2(_17308_));
 sg13g2_nor2b_1 _24273_ (.A(_17309_),
    .B_N(_15718_),
    .Y(_17310_));
 sg13g2_o21ai_1 _24274_ (.B1(_15712_),
    .Y(_17311_),
    .A1(_16438_),
    .A2(_17310_));
 sg13g2_a21o_1 _24275_ (.A2(_17311_),
    .A1(_16433_),
    .B1(_15713_),
    .X(_17312_));
 sg13g2_nand3_1 _24276_ (.B(_16433_),
    .C(_17311_),
    .A(_15713_),
    .Y(_17313_));
 sg13g2_nand3_1 _24277_ (.B(_17312_),
    .C(_17313_),
    .A(net5001),
    .Y(_17314_));
 sg13g2_or3_1 _24278_ (.A(_15718_),
    .B(_15720_),
    .C(_17226_),
    .X(_17315_));
 sg13g2_a21o_1 _24279_ (.A2(_17315_),
    .A1(_15742_),
    .B1(_15712_),
    .X(_17316_));
 sg13g2_nand2_1 _24280_ (.Y(_17317_),
    .A(_15711_),
    .B(_17316_));
 sg13g2_xnor2_1 _24281_ (.Y(_17318_),
    .A(_15714_),
    .B(_17317_));
 sg13g2_nor2_1 _24282_ (.A(net5706),
    .B(_17318_),
    .Y(_17319_));
 sg13g2_o21ai_1 _24283_ (.B1(net5085),
    .Y(_17320_),
    .A1(\u_inv.f_next[135] ),
    .A2(net5805));
 sg13g2_o21ai_1 _24284_ (.B1(_17314_),
    .Y(_17321_),
    .A1(_17319_),
    .A2(_17320_));
 sg13g2_xnor2_1 _24285_ (.Y(_17322_),
    .A(_15812_),
    .B(_17056_));
 sg13g2_o21ai_1 _24286_ (.B1(net5052),
    .Y(_17323_),
    .A1(\u_inv.f_next[200] ),
    .A2(net5762));
 sg13g2_a21oi_1 _24287_ (.A1(net5762),
    .A2(_17322_),
    .Y(_17324_),
    .B1(_17323_));
 sg13g2_nand3_1 _24288_ (.B(_16576_),
    .C(_17062_),
    .A(_15811_),
    .Y(_17325_));
 sg13g2_nor2_1 _24289_ (.A(net5052),
    .B(_17063_),
    .Y(_17326_));
 sg13g2_a21o_2 _24290_ (.A2(_17326_),
    .A1(_17325_),
    .B1(_17324_),
    .X(_17327_));
 sg13g2_xor2_1 _24291_ (.B(_16994_),
    .A(_14943_),
    .X(_17328_));
 sg13g2_a21oi_1 _24292_ (.A1(net5767),
    .A2(_17328_),
    .Y(_17329_),
    .B1(net4963));
 sg13g2_o21ai_1 _24293_ (.B1(_17329_),
    .Y(_17330_),
    .A1(\u_inv.f_next[180] ),
    .A2(net5767));
 sg13g2_nand3_1 _24294_ (.B(_16538_),
    .C(_17001_),
    .A(_14943_),
    .Y(_17331_));
 sg13g2_nand2_1 _24295_ (.Y(_17332_),
    .A(net4963),
    .B(_17331_));
 sg13g2_o21ai_1 _24296_ (.B1(_17330_),
    .Y(_17333_),
    .A1(_17002_),
    .A2(_17332_));
 sg13g2_a21oi_1 _24297_ (.A1(_16542_),
    .A2(_16861_),
    .Y(_17334_),
    .B1(_14932_));
 sg13g2_nand3_1 _24298_ (.B(_16542_),
    .C(_16861_),
    .A(_14932_),
    .Y(_17335_));
 sg13g2_nand2b_1 _24299_ (.Y(_17336_),
    .B(_17335_),
    .A_N(_17334_));
 sg13g2_or3_1 _24300_ (.A(_14932_),
    .B(_15046_),
    .C(_16852_),
    .X(_17337_));
 sg13g2_nand3_1 _24301_ (.B(_16853_),
    .C(_17337_),
    .A(net5767),
    .Y(_17338_));
 sg13g2_a21oi_1 _24302_ (.A1(\u_inv.f_next[184] ),
    .A2(net5680),
    .Y(_17339_),
    .B1(net4962));
 sg13g2_a22oi_1 _24303_ (.Y(_17340_),
    .B1(_17338_),
    .B2(_17339_),
    .A2(_17336_),
    .A1(net4962));
 sg13g2_a21oi_1 _24304_ (.A1(\u_inv.f_next[192] ),
    .A2(\u_inv.f_reg[192] ),
    .Y(_17341_),
    .B1(_17032_));
 sg13g2_xnor2_1 _24305_ (.Y(_17342_),
    .A(_15792_),
    .B(_17341_));
 sg13g2_o21ai_1 _24306_ (.B1(net5053),
    .Y(_17343_),
    .A1(\u_inv.f_next[193] ),
    .A2(net5763));
 sg13g2_a21oi_1 _24307_ (.A1(net5763),
    .A2(_17342_),
    .Y(_17344_),
    .B1(_17343_));
 sg13g2_nand3_1 _24308_ (.B(_16567_),
    .C(_17026_),
    .A(_15791_),
    .Y(_17345_));
 sg13g2_nor2_1 _24309_ (.A(net5053),
    .B(_17027_),
    .Y(_17346_));
 sg13g2_a21oi_1 _24310_ (.A1(_17345_),
    .A2(_17346_),
    .Y(_17347_),
    .B1(_17344_));
 sg13g2_inv_4 _24311_ (.A(_17347_),
    .Y(_17348_));
 sg13g2_xnor2_1 _24312_ (.Y(_17349_),
    .A(_14913_),
    .B(_16712_));
 sg13g2_o21ai_1 _24313_ (.B1(net5044),
    .Y(_17350_),
    .A1(\u_inv.f_next[208] ),
    .A2(net5754));
 sg13g2_a21oi_1 _24314_ (.A1(net5754),
    .A2(_17349_),
    .Y(_17351_),
    .B1(_17350_));
 sg13g2_nand3_1 _24315_ (.B(_16561_),
    .C(_16595_),
    .A(_14913_),
    .Y(_17352_));
 sg13g2_nor2_1 _24316_ (.A(net5044),
    .B(_17148_),
    .Y(_17353_));
 sg13g2_a21o_2 _24317_ (.A2(_17353_),
    .A1(_17352_),
    .B1(_17351_),
    .X(_17354_));
 sg13g2_a21oi_1 _24318_ (.A1(_15058_),
    .A2(_17083_),
    .Y(_17355_),
    .B1(_15057_));
 sg13g2_xnor2_1 _24319_ (.Y(_17356_),
    .A(_15056_),
    .B(_17355_));
 sg13g2_o21ai_1 _24320_ (.B1(net5068),
    .Y(_17357_),
    .A1(\u_inv.f_next[157] ),
    .A2(net5783));
 sg13g2_a21oi_1 _24321_ (.A1(net5783),
    .A2(_17356_),
    .Y(_17358_),
    .B1(_17357_));
 sg13g2_nand3_1 _24322_ (.B(_16050_),
    .C(_17074_),
    .A(_15055_),
    .Y(_17359_));
 sg13g2_and4_1 _24323_ (.A(net4978),
    .B(_16052_),
    .C(_17114_),
    .D(_17359_),
    .X(_17360_));
 sg13g2_or2_1 _24324_ (.X(_17361_),
    .B(_17360_),
    .A(_17358_));
 sg13g2_nand3_1 _24325_ (.B(_15988_),
    .C(_16704_),
    .A(_14876_),
    .Y(_17362_));
 sg13g2_nor3_1 _24326_ (.A(net5042),
    .B(_15989_),
    .C(_16705_),
    .Y(_17363_));
 sg13g2_o21ai_1 _24327_ (.B1(_14863_),
    .Y(_17364_),
    .A1(_14875_),
    .A2(_16716_));
 sg13g2_xnor2_1 _24328_ (.Y(_17365_),
    .A(_14876_),
    .B(_17364_));
 sg13g2_o21ai_1 _24329_ (.B1(net5042),
    .Y(_17366_),
    .A1(\u_inv.f_next[217] ),
    .A2(net5752));
 sg13g2_a21oi_1 _24330_ (.A1(net5752),
    .A2(_17365_),
    .Y(_17367_),
    .B1(_17366_));
 sg13g2_a21o_2 _24331_ (.A2(_17363_),
    .A1(_17362_),
    .B1(_17367_),
    .X(_17368_));
 sg13g2_or3_1 _24332_ (.A(_14968_),
    .B(_16491_),
    .C(_17168_),
    .X(_17369_));
 sg13g2_a21oi_1 _24333_ (.A1(_17169_),
    .A2(_17369_),
    .Y(_17370_),
    .B1(net5069));
 sg13g2_nand3_1 _24334_ (.B(_14983_),
    .C(_17175_),
    .A(_14968_),
    .Y(_17371_));
 sg13g2_nand3_1 _24335_ (.B(_17176_),
    .C(_17371_),
    .A(net5782),
    .Y(_17372_));
 sg13g2_a21oi_1 _24336_ (.A1(net3323),
    .A2(net5691),
    .Y(_17373_),
    .B1(net4978));
 sg13g2_a21oi_2 _24337_ (.B1(_17370_),
    .Y(_17374_),
    .A2(_17373_),
    .A1(_17372_));
 sg13g2_xnor2_1 _24338_ (.Y(_17375_),
    .A(_14937_),
    .B(_16995_));
 sg13g2_a21oi_1 _24339_ (.A1(net5767),
    .A2(_17375_),
    .Y(_17376_),
    .B1(net4963));
 sg13g2_o21ai_1 _24340_ (.B1(_17376_),
    .Y(_17377_),
    .A1(\u_inv.f_next[182] ),
    .A2(net5767));
 sg13g2_xnor2_1 _24341_ (.Y(_17378_),
    .A(_14938_),
    .B(_17004_));
 sg13g2_o21ai_1 _24342_ (.B1(_17377_),
    .Y(_17379_),
    .A1(net5056),
    .A2(_17378_));
 sg13g2_xnor2_1 _24343_ (.Y(_17380_),
    .A(_14875_),
    .B(_16716_));
 sg13g2_nand2_1 _24344_ (.Y(_17381_),
    .A(net5755),
    .B(_17380_));
 sg13g2_a21oi_1 _24345_ (.A1(_13958_),
    .A2(net5672),
    .Y(_17382_),
    .B1(net4952));
 sg13g2_a21oi_1 _24346_ (.A1(_14874_),
    .A2(_16703_),
    .Y(_17383_),
    .B1(net5041));
 sg13g2_and2_1 _24347_ (.A(_16704_),
    .B(_17383_),
    .X(_17384_));
 sg13g2_a22oi_1 _24348_ (.Y(_17385_),
    .B1(_17383_),
    .B2(_16704_),
    .A2(_17382_),
    .A1(_17381_));
 sg13g2_a21o_1 _24349_ (.A2(_17382_),
    .A1(_17381_),
    .B1(_17384_),
    .X(_17386_));
 sg13g2_xnor2_1 _24350_ (.Y(_17387_),
    .A(_15001_),
    .B(_16955_));
 sg13g2_nand2_1 _24351_ (.Y(_17388_),
    .A(_15002_),
    .B(_16968_));
 sg13g2_a21oi_1 _24352_ (.A1(_15001_),
    .A2(_16969_),
    .Y(_17389_),
    .B1(net5689));
 sg13g2_a221oi_1 _24353_ (.B2(_17389_),
    .C1(net4975),
    .B1(_17388_),
    .A1(\u_inv.f_next[172] ),
    .Y(_17390_),
    .A2(net5692));
 sg13g2_a21oi_2 _24354_ (.B1(_17390_),
    .Y(_17391_),
    .A2(_17387_),
    .A1(net4975));
 sg13g2_xnor2_1 _24355_ (.Y(_17392_),
    .A(_14950_),
    .B(_16993_));
 sg13g2_a21oi_1 _24356_ (.A1(net5777),
    .A2(_17392_),
    .Y(_17393_),
    .B1(net4975));
 sg13g2_o21ai_1 _24357_ (.B1(_17393_),
    .Y(_17394_),
    .A1(\u_inv.f_next[178] ),
    .A2(net5777));
 sg13g2_nor3_1 _24358_ (.A(_14950_),
    .B(_16534_),
    .C(_17089_),
    .Y(_17395_));
 sg13g2_nand2_1 _24359_ (.Y(_17396_),
    .A(net4975),
    .B(_17090_));
 sg13g2_o21ai_1 _24360_ (.B1(_17394_),
    .Y(_17397_),
    .A1(_17395_),
    .A2(_17396_));
 sg13g2_xnor2_1 _24361_ (.Y(_17398_),
    .A(_15805_),
    .B(_17134_));
 sg13g2_and3_1 _24362_ (.X(_17399_),
    .A(_15804_),
    .B(_15840_),
    .C(_17126_));
 sg13g2_nor3_1 _24363_ (.A(net5681),
    .B(_17287_),
    .C(_17399_),
    .Y(_17400_));
 sg13g2_nor2_1 _24364_ (.A(_13970_),
    .B(net5764),
    .Y(_17401_));
 sg13g2_o21ai_1 _24365_ (.B1(net5045),
    .Y(_17402_),
    .A1(_17400_),
    .A2(_17401_));
 sg13g2_o21ai_1 _24366_ (.B1(_17402_),
    .Y(_17403_),
    .A1(net5045),
    .A2(_17398_));
 sg13g2_a21oi_1 _24367_ (.A1(_14913_),
    .A2(_16712_),
    .Y(_17404_),
    .B1(_14896_));
 sg13g2_xnor2_1 _24368_ (.Y(_17405_),
    .A(_14912_),
    .B(_17404_));
 sg13g2_o21ai_1 _24369_ (.B1(net5044),
    .Y(_17406_),
    .A1(\u_inv.f_next[209] ),
    .A2(net5754));
 sg13g2_a21o_1 _24370_ (.A2(_17405_),
    .A1(net5756),
    .B1(_17406_),
    .X(_17407_));
 sg13g2_nor3_1 _24371_ (.A(_14912_),
    .B(_16003_),
    .C(_17148_),
    .Y(_17408_));
 sg13g2_nand2_1 _24372_ (.Y(_17409_),
    .A(net4953),
    .B(_17149_));
 sg13g2_o21ai_1 _24373_ (.B1(_17407_),
    .Y(_17410_),
    .A1(_17408_),
    .A2(_17409_));
 sg13g2_and3_1 _24374_ (.X(_17411_),
    .A(net5622),
    .B(_15029_),
    .C(_16854_));
 sg13g2_o21ai_1 _24375_ (.B1(net5766),
    .Y(_17412_),
    .A1(_17104_),
    .A2(_17411_));
 sg13g2_a21oi_1 _24376_ (.A1(_13988_),
    .A2(net5682),
    .Y(_17413_),
    .B1(net4962));
 sg13g2_xnor2_1 _24377_ (.Y(_17414_),
    .A(net5622),
    .B(_17099_));
 sg13g2_a22oi_1 _24378_ (.Y(_17415_),
    .B1(_17414_),
    .B2(net4962),
    .A2(_17413_),
    .A1(_17412_));
 sg13g2_inv_1 _24379_ (.Y(_17416_),
    .A(_17415_));
 sg13g2_xnor2_1 _24380_ (.Y(_17417_),
    .A(_14921_),
    .B(_16863_));
 sg13g2_o21ai_1 _24381_ (.B1(net5766),
    .Y(_17418_),
    .A1(_14921_),
    .A2(_16855_));
 sg13g2_a21o_1 _24382_ (.A2(_16855_),
    .A1(_14921_),
    .B1(_17418_),
    .X(_17419_));
 sg13g2_a21oi_1 _24383_ (.A1(\u_inv.f_next[188] ),
    .A2(net5680),
    .Y(_17420_),
    .B1(net4962));
 sg13g2_a22oi_1 _24384_ (.Y(_17421_),
    .B1(_17419_),
    .B2(_17420_),
    .A2(_17417_),
    .A1(net4962));
 sg13g2_a21oi_1 _24385_ (.A1(\u_inv.f_next[232] ),
    .A2(_14486_),
    .Y(_17422_),
    .B1(_15891_));
 sg13g2_o21ai_1 _24386_ (.B1(_17422_),
    .Y(_17423_),
    .A1(_15893_),
    .A2(_16683_));
 sg13g2_nand4_1 _24387_ (.B(_16631_),
    .C(_16767_),
    .A(net4941),
    .Y(_17424_),
    .D(_17423_));
 sg13g2_a21o_1 _24388_ (.A2(\u_inv.f_reg[232] ),
    .A1(\u_inv.f_next[232] ),
    .B1(_17188_),
    .X(_17425_));
 sg13g2_o21ai_1 _24389_ (.B1(net5738),
    .Y(_17426_),
    .A1(_15891_),
    .A2(_17425_));
 sg13g2_a21oi_1 _24390_ (.A1(_15891_),
    .A2(_17425_),
    .Y(_17427_),
    .B1(_17426_));
 sg13g2_o21ai_1 _24391_ (.B1(net5034),
    .Y(_17428_),
    .A1(\u_inv.f_next[233] ),
    .A2(net5738));
 sg13g2_o21ai_1 _24392_ (.B1(_17424_),
    .Y(_17429_),
    .A1(_17427_),
    .A2(_17428_));
 sg13g2_a21oi_1 _24393_ (.A1(_15904_),
    .A2(_15927_),
    .Y(_17430_),
    .B1(_15929_));
 sg13g2_nand3_1 _24394_ (.B(_15927_),
    .C(_15929_),
    .A(_15904_),
    .Y(_17431_));
 sg13g2_nand2b_1 _24395_ (.Y(_17432_),
    .B(_17431_),
    .A_N(_17430_));
 sg13g2_nor2_1 _24396_ (.A(\u_inv.f_next[240] ),
    .B(net5735),
    .Y(_17433_));
 sg13g2_a21oi_1 _24397_ (.A1(net5735),
    .A2(_17432_),
    .Y(_17434_),
    .B1(_17433_));
 sg13g2_nand2_1 _24398_ (.Y(_17435_),
    .A(_15929_),
    .B(_16646_));
 sg13g2_nor2_1 _24399_ (.A(_15929_),
    .B(_16646_),
    .Y(_17436_));
 sg13g2_nor2_1 _24400_ (.A(net5032),
    .B(_17436_),
    .Y(_17437_));
 sg13g2_a22oi_1 _24401_ (.Y(_17438_),
    .B1(_17435_),
    .B2(_17437_),
    .A2(_17434_),
    .A1(net5032));
 sg13g2_inv_4 _24402_ (.A(_17438_),
    .Y(_17439_));
 sg13g2_nor2_1 _24403_ (.A(_15930_),
    .B(_16657_),
    .Y(_17440_));
 sg13g2_nand3_1 _24404_ (.B(_16658_),
    .C(_16778_),
    .A(net4939),
    .Y(_17441_));
 sg13g2_a21oi_1 _24405_ (.A1(_17435_),
    .A2(_17440_),
    .Y(_17442_),
    .B1(_17441_));
 sg13g2_o21ai_1 _24406_ (.B1(_15930_),
    .Y(_17443_),
    .A1(_15928_),
    .A2(_17430_));
 sg13g2_or3_1 _24407_ (.A(_15928_),
    .B(_15930_),
    .C(_17430_),
    .X(_17444_));
 sg13g2_nand3_1 _24408_ (.B(_17443_),
    .C(_17444_),
    .A(net5737),
    .Y(_17445_));
 sg13g2_a21oi_1 _24409_ (.A1(_13933_),
    .A2(net5664),
    .Y(_17446_),
    .B1(net4939));
 sg13g2_a21oi_1 _24410_ (.A1(_17445_),
    .A2(_17446_),
    .Y(_17447_),
    .B1(_17442_));
 sg13g2_inv_2 _24411_ (.Y(_17448_),
    .A(_17447_));
 sg13g2_and3_1 _24412_ (.X(_17449_),
    .A(_14992_),
    .B(_15013_),
    .C(_16964_));
 sg13g2_o21ai_1 _24413_ (.B1(net5779),
    .Y(_17450_),
    .A1(_16965_),
    .A2(_17449_));
 sg13g2_o21ai_1 _24414_ (.B1(_17450_),
    .Y(_17451_),
    .A1(\u_inv.f_next[168] ),
    .A2(net5778));
 sg13g2_a21oi_1 _24415_ (.A1(_15013_),
    .A2(_16951_),
    .Y(_17452_),
    .B1(net5065));
 sg13g2_o21ai_1 _24416_ (.B1(_17452_),
    .Y(_17453_),
    .A1(_15013_),
    .A2(_16951_));
 sg13g2_o21ai_1 _24417_ (.B1(_17453_),
    .Y(_17454_),
    .A1(net4976),
    .A2(_17451_));
 sg13g2_a21oi_1 _24418_ (.A1(\u_inv.f_next[168] ),
    .A2(_14422_),
    .Y(_17455_),
    .B1(_15011_));
 sg13g2_o21ai_1 _24419_ (.B1(_17455_),
    .Y(_17456_),
    .A1(_15012_),
    .A2(_16950_));
 sg13g2_nand4_1 _24420_ (.B(_16507_),
    .C(_16953_),
    .A(net4976),
    .Y(_17457_),
    .D(_17456_));
 sg13g2_a21o_1 _24421_ (.A2(\u_inv.f_reg[168] ),
    .A1(\u_inv.f_next[168] ),
    .B1(_16965_),
    .X(_17458_));
 sg13g2_o21ai_1 _24422_ (.B1(net5778),
    .Y(_17459_),
    .A1(_15011_),
    .A2(_17458_));
 sg13g2_a21oi_1 _24423_ (.A1(_15011_),
    .A2(_17458_),
    .Y(_17460_),
    .B1(_17459_));
 sg13g2_o21ai_1 _24424_ (.B1(net5066),
    .Y(_17461_),
    .A1(\u_inv.f_next[169] ),
    .A2(net5778));
 sg13g2_o21ai_1 _24425_ (.B1(_17457_),
    .Y(_17462_),
    .A1(_17460_),
    .A2(_17461_));
 sg13g2_o21ai_1 _24426_ (.B1(_15692_),
    .Y(_17463_),
    .A1(_15693_),
    .A2(_17229_));
 sg13g2_xnor2_1 _24427_ (.Y(_17464_),
    .A(_15690_),
    .B(_17463_));
 sg13g2_o21ai_1 _24428_ (.B1(net5077),
    .Y(_17465_),
    .A1(\u_inv.f_next[141] ),
    .A2(net5795));
 sg13g2_a21oi_1 _24429_ (.A1(net5795),
    .A2(_17464_),
    .Y(_17466_),
    .B1(_17465_));
 sg13g2_nand3_1 _24430_ (.B(_16450_),
    .C(_17219_),
    .A(_15690_),
    .Y(_17467_));
 sg13g2_nor2_1 _24431_ (.A(net5077),
    .B(_17220_),
    .Y(_17468_));
 sg13g2_a21oi_2 _24432_ (.B1(_17466_),
    .Y(_17469_),
    .A2(_17468_),
    .A1(_17467_));
 sg13g2_a21oi_1 _24433_ (.A1(_15092_),
    .A2(_17079_),
    .Y(_17470_),
    .B1(_15091_));
 sg13g2_xnor2_1 _24434_ (.Y(_17471_),
    .A(_15090_),
    .B(_17470_));
 sg13g2_o21ai_1 _24435_ (.B1(net5074),
    .Y(_17472_),
    .A1(\u_inv.f_next[149] ),
    .A2(net5792));
 sg13g2_a21oi_1 _24436_ (.A1(net5792),
    .A2(_17471_),
    .Y(_17473_),
    .B1(_17472_));
 sg13g2_nor3_1 _24437_ (.A(_15090_),
    .B(_16020_),
    .C(_17195_),
    .Y(_17474_));
 sg13g2_nor2_1 _24438_ (.A(net5075),
    .B(_17474_),
    .Y(_17475_));
 sg13g2_a21o_2 _24439_ (.A2(_17475_),
    .A1(_17196_),
    .B1(_17473_),
    .X(_17476_));
 sg13g2_a21oi_1 _24440_ (.A1(_15596_),
    .A2(_15609_),
    .Y(_17477_),
    .B1(_15650_));
 sg13g2_o21ai_1 _24441_ (.B1(_15649_),
    .Y(_17478_),
    .A1(_15595_),
    .A2(_15608_));
 sg13g2_a21oi_2 _24442_ (.B1(_15659_),
    .Y(_17479_),
    .A2(_17477_),
    .A1(_15651_));
 sg13g2_o21ai_1 _24443_ (.B1(_15658_),
    .Y(_17480_),
    .A1(_15652_),
    .A2(_17478_));
 sg13g2_a21oi_1 _24444_ (.A1(_15647_),
    .A2(_17480_),
    .Y(_17481_),
    .B1(_15661_));
 sg13g2_o21ai_1 _24445_ (.B1(_15662_),
    .Y(_17482_),
    .A1(_15646_),
    .A2(_17479_));
 sg13g2_a21oi_1 _24446_ (.A1(_15639_),
    .A2(_17482_),
    .Y(_17483_),
    .B1(_15666_));
 sg13g2_o21ai_1 _24447_ (.B1(_15632_),
    .Y(_17484_),
    .A1(_15633_),
    .A2(_17483_));
 sg13g2_o21ai_1 _24448_ (.B1(net5808),
    .Y(_17485_),
    .A1(_15631_),
    .A2(_17484_));
 sg13g2_a21oi_1 _24449_ (.A1(_15631_),
    .A2(_17484_),
    .Y(_17486_),
    .B1(_17485_));
 sg13g2_o21ai_1 _24450_ (.B1(net5086),
    .Y(_17487_),
    .A1(\u_inv.f_next[119] ),
    .A2(net5808));
 sg13g2_a21oi_1 _24451_ (.A1(_16352_),
    .A2(_16368_),
    .Y(_17488_),
    .B1(_16375_));
 sg13g2_o21ai_1 _24452_ (.B1(_15636_),
    .Y(_17489_),
    .A1(_16393_),
    .A2(_17488_));
 sg13g2_a21oi_1 _24453_ (.A1(_16384_),
    .A2(_17489_),
    .Y(_17490_),
    .B1(_15637_));
 sg13g2_o21ai_1 _24454_ (.B1(_15633_),
    .Y(_17491_),
    .A1(_16383_),
    .A2(_17490_));
 sg13g2_nand2b_1 _24455_ (.Y(_17492_),
    .B(_17491_),
    .A_N(_16382_));
 sg13g2_a21oi_1 _24456_ (.A1(_15631_),
    .A2(_17492_),
    .Y(_17493_),
    .B1(net5087));
 sg13g2_o21ai_1 _24457_ (.B1(_17493_),
    .Y(_17494_),
    .A1(_15631_),
    .A2(_17492_));
 sg13g2_o21ai_1 _24458_ (.B1(_17494_),
    .Y(_17495_),
    .A1(_17486_),
    .A2(_17487_));
 sg13g2_o21ai_1 _24459_ (.B1(_16396_),
    .Y(_17496_),
    .A1(_16369_),
    .A2(_16379_));
 sg13g2_a21oi_1 _24460_ (.A1(_15627_),
    .A2(_17496_),
    .Y(_17497_),
    .B1(_16406_));
 sg13g2_nor2_1 _24461_ (.A(_15628_),
    .B(_17497_),
    .Y(_17498_));
 sg13g2_o21ai_1 _24462_ (.B1(_16405_),
    .Y(_17499_),
    .A1(_15628_),
    .A2(_17497_));
 sg13g2_a21o_1 _24463_ (.A2(_17499_),
    .A1(_15624_),
    .B1(_16404_),
    .X(_17500_));
 sg13g2_and2_1 _24464_ (.A(_15622_),
    .B(_17500_),
    .X(_17501_));
 sg13g2_o21ai_1 _24465_ (.B1(net5002),
    .Y(_17502_),
    .A1(_15622_),
    .A2(_17500_));
 sg13g2_o21ai_1 _24466_ (.B1(_15653_),
    .Y(_17503_),
    .A1(_15595_),
    .A2(_15608_));
 sg13g2_and2_1 _24467_ (.A(_15669_),
    .B(_17503_),
    .X(_17504_));
 sg13g2_a21oi_1 _24468_ (.A1(_15669_),
    .A2(_17503_),
    .Y(_17505_),
    .B1(_15629_));
 sg13g2_nor2_1 _24469_ (.A(_15671_),
    .B(_17505_),
    .Y(_17506_));
 sg13g2_o21ai_1 _24470_ (.B1(_15623_),
    .Y(_17507_),
    .A1(_15624_),
    .A2(_17506_));
 sg13g2_xnor2_1 _24471_ (.Y(_17508_),
    .A(_15622_),
    .B(_17507_));
 sg13g2_a21oi_1 _24472_ (.A1(_14051_),
    .A2(net5707),
    .Y(_17509_),
    .B1(net5002));
 sg13g2_o21ai_1 _24473_ (.B1(_17509_),
    .Y(_17510_),
    .A1(net5707),
    .A2(_17508_));
 sg13g2_o21ai_1 _24474_ (.B1(_17510_),
    .Y(_17511_),
    .A1(_17501_),
    .A2(_17502_));
 sg13g2_xnor2_1 _24475_ (.Y(_17512_),
    .A(_15706_),
    .B(_17228_));
 sg13g2_a21oi_1 _24476_ (.A1(net5794),
    .A2(_17512_),
    .Y(_17513_),
    .B1(net4990));
 sg13g2_o21ai_1 _24477_ (.B1(_17513_),
    .Y(_17514_),
    .A1(\u_inv.f_next[138] ),
    .A2(net5794));
 sg13g2_or2_1 _24478_ (.X(_17515_),
    .B(_17217_),
    .A(_15698_));
 sg13g2_a21oi_1 _24479_ (.A1(_16444_),
    .A2(_17515_),
    .Y(_17516_),
    .B1(_15702_));
 sg13g2_nor3_1 _24480_ (.A(_15707_),
    .B(_16443_),
    .C(_17516_),
    .Y(_17517_));
 sg13g2_o21ai_1 _24481_ (.B1(_15707_),
    .Y(_17518_),
    .A1(_16443_),
    .A2(_17516_));
 sg13g2_nand2_1 _24482_ (.Y(_17519_),
    .A(net4991),
    .B(_17518_));
 sg13g2_o21ai_1 _24483_ (.B1(_17514_),
    .Y(_17520_),
    .A1(_17517_),
    .A2(_17519_));
 sg13g2_a21oi_1 _24484_ (.A1(_16060_),
    .A2(_17068_),
    .Y(_17521_),
    .B1(_16028_));
 sg13g2_o21ai_1 _24485_ (.B1(_16032_),
    .Y(_17522_),
    .A1(_15079_),
    .A2(_17521_));
 sg13g2_a21oi_1 _24486_ (.A1(_15077_),
    .A2(_17522_),
    .Y(_17523_),
    .B1(net5074));
 sg13g2_o21ai_1 _24487_ (.B1(_17523_),
    .Y(_17524_),
    .A1(_15077_),
    .A2(_17522_));
 sg13g2_o21ai_1 _24488_ (.B1(_17076_),
    .Y(_17525_),
    .A1(_14030_),
    .A2(_14398_));
 sg13g2_a21oi_1 _24489_ (.A1(_15113_),
    .A2(_17076_),
    .Y(_17526_),
    .B1(_15082_));
 sg13g2_a21oi_1 _24490_ (.A1(_15079_),
    .A2(_17526_),
    .Y(_17527_),
    .B1(_15078_));
 sg13g2_xnor2_1 _24491_ (.Y(_17528_),
    .A(_15076_),
    .B(_17527_));
 sg13g2_nor2_1 _24492_ (.A(\u_inv.f_next[147] ),
    .B(net5792),
    .Y(_17529_));
 sg13g2_o21ai_1 _24493_ (.B1(net5074),
    .Y(_17530_),
    .A1(net5697),
    .A2(_17528_));
 sg13g2_o21ai_1 _24494_ (.B1(_17524_),
    .Y(_17531_),
    .A1(_17529_),
    .A2(_17530_));
 sg13g2_xnor2_1 _24495_ (.Y(_17532_),
    .A(_15066_),
    .B(_17245_));
 sg13g2_nand3_1 _24496_ (.B(_15099_),
    .C(_17082_),
    .A(_15067_),
    .Y(_17533_));
 sg13g2_nand3_1 _24497_ (.B(_17249_),
    .C(_17533_),
    .A(net5791),
    .Y(_17534_));
 sg13g2_a21oi_1 _24498_ (.A1(\u_inv.f_next[154] ),
    .A2(net5698),
    .Y(_17535_),
    .B1(net4988));
 sg13g2_a22oi_1 _24499_ (.Y(_17536_),
    .B1(_17534_),
    .B2(_17535_),
    .A2(_17532_),
    .A1(net4988));
 sg13g2_a21oi_1 _24500_ (.A1(_16381_),
    .A2(_16413_),
    .Y(_17537_),
    .B1(_15730_));
 sg13g2_o21ai_1 _24501_ (.B1(_15728_),
    .Y(_17538_),
    .A1(_16424_),
    .A2(_17537_));
 sg13g2_a21oi_1 _24502_ (.A1(_16426_),
    .A2(_17538_),
    .Y(_17539_),
    .B1(_15723_));
 sg13g2_o21ai_1 _24503_ (.B1(_15726_),
    .Y(_17540_),
    .A1(_16425_),
    .A2(_17539_));
 sg13g2_nor3_1 _24504_ (.A(_15726_),
    .B(_16425_),
    .C(_17539_),
    .Y(_17541_));
 sg13g2_nand2_1 _24505_ (.Y(_17542_),
    .A(net5000),
    .B(_17540_));
 sg13g2_a21oi_1 _24506_ (.A1(_15682_),
    .A2(_15732_),
    .Y(_17543_),
    .B1(_15738_));
 sg13g2_o21ai_1 _24507_ (.B1(_15722_),
    .Y(_17544_),
    .A1(_15724_),
    .A2(_17543_));
 sg13g2_xor2_1 _24508_ (.B(_17544_),
    .A(_15726_),
    .X(_17545_));
 sg13g2_a21oi_1 _24509_ (.A1(net5806),
    .A2(_17545_),
    .Y(_17546_),
    .B1(net5000));
 sg13g2_o21ai_1 _24510_ (.B1(_17546_),
    .Y(_17547_),
    .A1(\u_inv.f_next[131] ),
    .A2(net5806));
 sg13g2_o21ai_1 _24511_ (.B1(_17547_),
    .Y(_17548_),
    .A1(_17541_),
    .A2(_17542_));
 sg13g2_nand3_1 _24512_ (.B(_16044_),
    .C(_17071_),
    .A(_15069_),
    .Y(_17549_));
 sg13g2_nand4_1 _24513_ (.B(_16046_),
    .C(_17072_),
    .A(net4988),
    .Y(_17550_),
    .D(_17549_));
 sg13g2_and3_1 _24514_ (.X(_17551_),
    .A(_15069_),
    .B(_15071_),
    .C(_17081_));
 sg13g2_a21oi_1 _24515_ (.A1(_15071_),
    .A2(_17081_),
    .Y(_17552_),
    .B1(_15069_));
 sg13g2_nor3_1 _24516_ (.A(net5698),
    .B(_17551_),
    .C(_17552_),
    .Y(_17553_));
 sg13g2_o21ai_1 _24517_ (.B1(net5074),
    .Y(_17554_),
    .A1(\u_inv.f_next[153] ),
    .A2(net5791));
 sg13g2_o21ai_1 _24518_ (.B1(_17550_),
    .Y(_17555_),
    .A1(_17553_),
    .A2(_17554_));
 sg13g2_or3_1 _24519_ (.A(_15072_),
    .B(_16024_),
    .C(_17070_),
    .X(_17556_));
 sg13g2_a21oi_1 _24520_ (.A1(_17071_),
    .A2(_17556_),
    .Y(_17557_),
    .B1(net5074));
 sg13g2_nand3_1 _24521_ (.B(_15112_),
    .C(_17080_),
    .A(_15072_),
    .Y(_17558_));
 sg13g2_nand3_1 _24522_ (.B(_17081_),
    .C(_17558_),
    .A(net5792),
    .Y(_17559_));
 sg13g2_a21oi_1 _24523_ (.A1(\u_inv.f_next[152] ),
    .A2(net5698),
    .Y(_17560_),
    .B1(net4988));
 sg13g2_a21oi_1 _24524_ (.A1(_17559_),
    .A2(_17560_),
    .Y(_17561_),
    .B1(_17557_));
 sg13g2_nor3_1 _24525_ (.A(_15780_),
    .B(_15828_),
    .C(_17040_),
    .Y(_17562_));
 sg13g2_o21ai_1 _24526_ (.B1(net5764),
    .Y(_17563_),
    .A1(_17043_),
    .A2(_17562_));
 sg13g2_a21oi_1 _24527_ (.A1(_13978_),
    .A2(net5681),
    .Y(_17564_),
    .B1(net4965));
 sg13g2_and3_1 _24528_ (.X(_17565_),
    .A(_15780_),
    .B(_16570_),
    .C(_17048_));
 sg13g2_nor3_1 _24529_ (.A(net5053),
    .B(_17049_),
    .C(_17565_),
    .Y(_17566_));
 sg13g2_a21o_1 _24530_ (.A2(_17564_),
    .A1(_17563_),
    .B1(_17566_),
    .X(_17567_));
 sg13g2_o21ai_1 _24531_ (.B1(_14930_),
    .Y(_17568_),
    .A1(_13990_),
    .A2(\u_inv.f_reg[184] ));
 sg13g2_nor3_1 _24532_ (.A(net5055),
    .B(_16518_),
    .C(_16862_),
    .Y(_17569_));
 sg13g2_o21ai_1 _24533_ (.B1(_17569_),
    .Y(_17570_),
    .A1(_17334_),
    .A2(_17568_));
 sg13g2_and3_1 _24534_ (.X(_17571_),
    .A(_14930_),
    .B(_14931_),
    .C(_16853_));
 sg13g2_a21oi_1 _24535_ (.A1(_14931_),
    .A2(_16853_),
    .Y(_17572_),
    .B1(_14930_));
 sg13g2_nor3_1 _24536_ (.A(net5681),
    .B(_17571_),
    .C(_17572_),
    .Y(_17573_));
 sg13g2_o21ai_1 _24537_ (.B1(net5055),
    .Y(_17574_),
    .A1(\u_inv.f_next[185] ),
    .A2(net5766));
 sg13g2_o21ai_1 _24538_ (.B1(_17570_),
    .Y(_17575_),
    .A1(_17573_),
    .A2(_17574_));
 sg13g2_or2_1 _24539_ (.X(_17576_),
    .B(_16478_),
    .A(_16459_));
 sg13g2_a21o_1 _24540_ (.A2(_17576_),
    .A1(_16487_),
    .B1(_14979_),
    .X(_17577_));
 sg13g2_a21oi_1 _24541_ (.A1(_16484_),
    .A2(_17577_),
    .Y(_17578_),
    .B1(_14977_));
 sg13g2_nand3_1 _24542_ (.B(_16484_),
    .C(_17577_),
    .A(_14977_),
    .Y(_17579_));
 sg13g2_nand2_1 _24543_ (.Y(_17580_),
    .A(net4977),
    .B(_17579_));
 sg13g2_a21oi_1 _24544_ (.A1(_14979_),
    .A2(_16963_),
    .Y(_17581_),
    .B1(_14978_));
 sg13g2_xor2_1 _24545_ (.B(_17581_),
    .A(_14977_),
    .X(_17582_));
 sg13g2_a21oi_1 _24546_ (.A1(net5782),
    .A2(_17582_),
    .Y(_17583_),
    .B1(net4977));
 sg13g2_o21ai_1 _24547_ (.B1(_17583_),
    .Y(_17584_),
    .A1(net2744),
    .A2(net5782));
 sg13g2_o21ai_1 _24548_ (.B1(_17584_),
    .Y(_17585_),
    .A1(_17578_),
    .A2(_17580_));
 sg13g2_nor3_1 _24549_ (.A(_14953_),
    .B(_14957_),
    .C(_16991_),
    .Y(_17586_));
 sg13g2_o21ai_1 _24550_ (.B1(_14957_),
    .Y(_17587_),
    .A1(_14953_),
    .A2(_16991_));
 sg13g2_nand2_1 _24551_ (.Y(_17588_),
    .A(net5777),
    .B(_17587_));
 sg13g2_a21oi_1 _24552_ (.A1(_13997_),
    .A2(net5680),
    .Y(_17589_),
    .B1(net4962));
 sg13g2_o21ai_1 _24553_ (.B1(_17589_),
    .Y(_17590_),
    .A1(_17586_),
    .A2(_17588_));
 sg13g2_nand3_1 _24554_ (.B(_16532_),
    .C(_17088_),
    .A(_14956_),
    .Y(_17591_));
 sg13g2_nand2_1 _24555_ (.Y(_17592_),
    .A(net4975),
    .B(_17591_));
 sg13g2_o21ai_1 _24556_ (.B1(_17590_),
    .Y(_17593_),
    .A1(_17089_),
    .A2(_17592_));
 sg13g2_xnor2_1 _24557_ (.Y(_17594_),
    .A(_15633_),
    .B(_17483_));
 sg13g2_o21ai_1 _24558_ (.B1(net5086),
    .Y(_17595_),
    .A1(\u_inv.f_next[118] ),
    .A2(net5807));
 sg13g2_a21oi_1 _24559_ (.A1(net5807),
    .A2(_17594_),
    .Y(_17596_),
    .B1(_17595_));
 sg13g2_nor3_1 _24560_ (.A(_15633_),
    .B(_16383_),
    .C(_17490_),
    .Y(_17597_));
 sg13g2_nor2_1 _24561_ (.A(net5086),
    .B(_17597_),
    .Y(_17598_));
 sg13g2_a21o_2 _24562_ (.A2(_17598_),
    .A1(_17491_),
    .B1(_17596_),
    .X(_17599_));
 sg13g2_xnor2_1 _24563_ (.Y(_17600_),
    .A(_15079_),
    .B(_17526_));
 sg13g2_o21ai_1 _24564_ (.B1(net5074),
    .Y(_17601_),
    .A1(\u_inv.f_next[146] ),
    .A2(net5796));
 sg13g2_a21oi_1 _24565_ (.A1(net5796),
    .A2(_17600_),
    .Y(_17602_),
    .B1(_17601_));
 sg13g2_o21ai_1 _24566_ (.B1(net4991),
    .Y(_17603_),
    .A1(_15079_),
    .A2(_17521_));
 sg13g2_a21oi_1 _24567_ (.A1(_15079_),
    .A2(_17521_),
    .Y(_17604_),
    .B1(_17603_));
 sg13g2_nor2_1 _24568_ (.A(_17602_),
    .B(_17604_),
    .Y(_17605_));
 sg13g2_inv_2 _24569_ (.Y(_17606_),
    .A(_17605_));
 sg13g2_a21oi_1 _24570_ (.A1(_15625_),
    .A2(_17505_),
    .Y(_17607_),
    .B1(_15673_));
 sg13g2_nand2b_1 _24571_ (.Y(_17608_),
    .B(_15618_),
    .A_N(_17607_));
 sg13g2_a21oi_1 _24572_ (.A1(_15617_),
    .A2(_17608_),
    .Y(_17609_),
    .B1(_15616_));
 sg13g2_nand3_1 _24573_ (.B(_15617_),
    .C(_17608_),
    .A(_15616_),
    .Y(_17610_));
 sg13g2_nand3b_1 _24574_ (.B(_17610_),
    .C(net5809),
    .Y(_17611_),
    .A_N(_17609_));
 sg13g2_o21ai_1 _24575_ (.B1(_17611_),
    .Y(_17612_),
    .A1(\u_inv.f_next[125] ),
    .A2(net5809));
 sg13g2_and2_1 _24576_ (.A(_16372_),
    .B(_17496_),
    .X(_17613_));
 sg13g2_o21ai_1 _24577_ (.B1(_15619_),
    .Y(_17614_),
    .A1(_16411_),
    .A2(_17613_));
 sg13g2_nand3_1 _24578_ (.B(_16399_),
    .C(_17614_),
    .A(_15616_),
    .Y(_17615_));
 sg13g2_a21oi_1 _24579_ (.A1(_16399_),
    .A2(_17614_),
    .Y(_17616_),
    .B1(_15616_));
 sg13g2_nor2_1 _24580_ (.A(net5088),
    .B(_17616_),
    .Y(_17617_));
 sg13g2_nand2_1 _24581_ (.Y(_17618_),
    .A(_17615_),
    .B(_17617_));
 sg13g2_o21ai_1 _24582_ (.B1(_17618_),
    .Y(_17619_),
    .A1(net5003),
    .A2(_17612_));
 sg13g2_a21oi_1 _24583_ (.A1(_16331_),
    .A2(_16345_),
    .Y(_17620_),
    .B1(_16347_));
 sg13g2_nor2_1 _24584_ (.A(_16359_),
    .B(_17620_),
    .Y(_17621_));
 sg13g2_o21ai_1 _24585_ (.B1(_15581_),
    .Y(_17622_),
    .A1(_16359_),
    .A2(_17620_));
 sg13g2_a21oi_1 _24586_ (.A1(_16361_),
    .A2(_17622_),
    .Y(_17623_),
    .B1(_15577_));
 sg13g2_a21oi_1 _24587_ (.A1(\u_inv.f_next[109] ),
    .A2(_14363_),
    .Y(_17624_),
    .B1(_17623_));
 sg13g2_nor2_1 _24588_ (.A(_15575_),
    .B(_17624_),
    .Y(_17625_));
 sg13g2_o21ai_1 _24589_ (.B1(_15572_),
    .Y(_17626_),
    .A1(_16365_),
    .A2(_17625_));
 sg13g2_nor3_1 _24590_ (.A(_15572_),
    .B(_16365_),
    .C(_17625_),
    .Y(_17627_));
 sg13g2_nor2_1 _24591_ (.A(net5096),
    .B(_17627_),
    .Y(_17628_));
 sg13g2_nand2_1 _24592_ (.Y(_17629_),
    .A(_17626_),
    .B(_17628_));
 sg13g2_a21oi_2 _24593_ (.B1(_15599_),
    .Y(_17630_),
    .A2(_15593_),
    .A1(_15570_));
 sg13g2_o21ai_1 _24594_ (.B1(_15601_),
    .Y(_17631_),
    .A1(_15589_),
    .A2(_17630_));
 sg13g2_a21oi_1 _24595_ (.A1(_15582_),
    .A2(_17631_),
    .Y(_17632_),
    .B1(_15606_));
 sg13g2_o21ai_1 _24596_ (.B1(_15573_),
    .Y(_17633_),
    .A1(_15574_),
    .A2(_17632_));
 sg13g2_a21oi_1 _24597_ (.A1(_15572_),
    .A2(_17633_),
    .Y(_17634_),
    .B1(net5715));
 sg13g2_o21ai_1 _24598_ (.B1(_17634_),
    .Y(_17635_),
    .A1(_15572_),
    .A2(_17633_));
 sg13g2_nor2_1 _24599_ (.A(\u_inv.f_next[111] ),
    .B(net5819),
    .Y(_17636_));
 sg13g2_nor2_1 _24600_ (.A(net5011),
    .B(_17636_),
    .Y(_17637_));
 sg13g2_nand2_1 _24601_ (.Y(_17638_),
    .A(net5096),
    .B(_17635_));
 sg13g2_a22oi_1 _24602_ (.Y(_17639_),
    .B1(_17635_),
    .B2(_17637_),
    .A2(_17628_),
    .A1(_17626_));
 sg13g2_o21ai_1 _24603_ (.B1(_17629_),
    .Y(_17640_),
    .A1(_17636_),
    .A2(_17638_));
 sg13g2_xnor2_1 _24604_ (.Y(_17641_),
    .A(_15624_),
    .B(_17506_));
 sg13g2_o21ai_1 _24605_ (.B1(net5088),
    .Y(_17642_),
    .A1(\u_inv.f_next[122] ),
    .A2(net5809));
 sg13g2_a21o_1 _24606_ (.A2(_17641_),
    .A1(net5807),
    .B1(_17642_),
    .X(_17643_));
 sg13g2_xnor2_1 _24607_ (.Y(_17644_),
    .A(_15624_),
    .B(_17499_));
 sg13g2_o21ai_1 _24608_ (.B1(_17643_),
    .Y(_17645_),
    .A1(net5088),
    .A2(_17644_));
 sg13g2_nand2b_1 _24609_ (.Y(_17646_),
    .B(_15698_),
    .A_N(_17227_));
 sg13g2_o21ai_1 _24610_ (.B1(_15696_),
    .Y(_17647_),
    .A1(_15699_),
    .A2(_17227_));
 sg13g2_xnor2_1 _24611_ (.Y(_17648_),
    .A(_15702_),
    .B(_17647_));
 sg13g2_o21ai_1 _24612_ (.B1(net5078),
    .Y(_17649_),
    .A1(\u_inv.f_next[137] ),
    .A2(net5795));
 sg13g2_a21oi_1 _24613_ (.A1(net5794),
    .A2(_17648_),
    .Y(_17650_),
    .B1(_17649_));
 sg13g2_nand3_1 _24614_ (.B(_16444_),
    .C(_17515_),
    .A(_15702_),
    .Y(_17651_));
 sg13g2_nor2_1 _24615_ (.A(net5077),
    .B(_17516_),
    .Y(_17652_));
 sg13g2_a21oi_2 _24616_ (.B1(_17650_),
    .Y(_17653_),
    .A2(_17652_),
    .A1(_17651_));
 sg13g2_nand2b_1 _24617_ (.Y(_17654_),
    .B(_17653_),
    .A_N(_17645_));
 sg13g2_o21ai_1 _24618_ (.B1(_15650_),
    .Y(_17655_),
    .A1(_16351_),
    .A2(_16367_));
 sg13g2_a21o_1 _24619_ (.A2(_17655_),
    .A1(_16390_),
    .B1(_15651_),
    .X(_17656_));
 sg13g2_a21oi_1 _24620_ (.A1(_16389_),
    .A2(_17656_),
    .Y(_17657_),
    .B1(_15644_));
 sg13g2_o21ai_1 _24621_ (.B1(_15642_),
    .Y(_17658_),
    .A1(_16388_),
    .A2(_17657_));
 sg13g2_nor3_1 _24622_ (.A(_15642_),
    .B(_16388_),
    .C(_17657_),
    .Y(_17659_));
 sg13g2_nor2_1 _24623_ (.A(net5096),
    .B(_17659_),
    .Y(_17660_));
 sg13g2_o21ai_1 _24624_ (.B1(_15643_),
    .Y(_17661_),
    .A1(_15645_),
    .A2(_17479_));
 sg13g2_xnor2_1 _24625_ (.Y(_17662_),
    .A(_15641_),
    .B(_17661_));
 sg13g2_o21ai_1 _24626_ (.B1(net5096),
    .Y(_17663_),
    .A1(\u_inv.f_next[115] ),
    .A2(net5820));
 sg13g2_a21oi_1 _24627_ (.A1(net5820),
    .A2(_17662_),
    .Y(_17664_),
    .B1(_17663_));
 sg13g2_a21o_2 _24628_ (.A2(_17660_),
    .A1(_17658_),
    .B1(_17664_),
    .X(_17665_));
 sg13g2_xnor2_1 _24629_ (.Y(_17666_),
    .A(_15693_),
    .B(_17229_));
 sg13g2_o21ai_1 _24630_ (.B1(net5077),
    .Y(_17667_),
    .A1(\u_inv.f_next[140] ),
    .A2(net5794));
 sg13g2_a21o_1 _24631_ (.A2(_17666_),
    .A1(net5795),
    .B1(_17667_),
    .X(_17668_));
 sg13g2_a21oi_1 _24632_ (.A1(_15693_),
    .A2(_17218_),
    .Y(_17669_),
    .B1(net5077));
 sg13g2_o21ai_1 _24633_ (.B1(_17669_),
    .Y(_17670_),
    .A1(_15693_),
    .A2(_17218_));
 sg13g2_nand2_1 _24634_ (.Y(_17671_),
    .A(_17668_),
    .B(_17670_));
 sg13g2_nand3b_1 _24635_ (.B(_15618_),
    .C(_15616_),
    .Y(_17672_),
    .A_N(_17607_));
 sg13g2_nor2b_1 _24636_ (.A(_15677_),
    .B_N(_17672_),
    .Y(_17673_));
 sg13g2_xnor2_1 _24637_ (.Y(_17674_),
    .A(_15614_),
    .B(_17673_));
 sg13g2_o21ai_1 _24638_ (.B1(net5088),
    .Y(_17675_),
    .A1(net5707),
    .A2(_17674_));
 sg13g2_a21oi_1 _24639_ (.A1(_14048_),
    .A2(net5708),
    .Y(_17676_),
    .B1(_17675_));
 sg13g2_nor3_1 _24640_ (.A(_15613_),
    .B(_16398_),
    .C(_17616_),
    .Y(_17677_));
 sg13g2_o21ai_1 _24641_ (.B1(_15613_),
    .Y(_17678_),
    .A1(_16398_),
    .A2(_17616_));
 sg13g2_nor2_1 _24642_ (.A(net5088),
    .B(_17677_),
    .Y(_17679_));
 sg13g2_nand2_1 _24643_ (.Y(_17680_),
    .A(_17678_),
    .B(_17679_));
 sg13g2_nor2b_1 _24644_ (.A(_17676_),
    .B_N(_17680_),
    .Y(_17681_));
 sg13g2_nand2b_1 _24645_ (.Y(_17682_),
    .B(_17680_),
    .A_N(_17676_));
 sg13g2_xnor2_1 _24646_ (.Y(_17683_),
    .A(_15724_),
    .B(_17543_));
 sg13g2_o21ai_1 _24647_ (.B1(net5085),
    .Y(_17684_),
    .A1(\u_inv.f_next[130] ),
    .A2(net5805));
 sg13g2_a21oi_1 _24648_ (.A1(net5805),
    .A2(_17683_),
    .Y(_17685_),
    .B1(_17684_));
 sg13g2_nand3_1 _24649_ (.B(_16426_),
    .C(_17538_),
    .A(_15723_),
    .Y(_17686_));
 sg13g2_nor2_1 _24650_ (.A(net5085),
    .B(_17539_),
    .Y(_17687_));
 sg13g2_a21o_1 _24651_ (.A2(_17687_),
    .A1(_17686_),
    .B1(_17685_),
    .X(_17688_));
 sg13g2_xnor2_1 _24652_ (.Y(_17689_),
    .A(_15092_),
    .B(_17079_));
 sg13g2_o21ai_1 _24653_ (.B1(net5075),
    .Y(_17690_),
    .A1(\u_inv.f_next[148] ),
    .A2(net5792));
 sg13g2_a21oi_1 _24654_ (.A1(net5792),
    .A2(_17689_),
    .Y(_17691_),
    .B1(_17690_));
 sg13g2_nand3_1 _24655_ (.B(_16033_),
    .C(_17069_),
    .A(_15092_),
    .Y(_17692_));
 sg13g2_nor2_1 _24656_ (.A(net5075),
    .B(_17195_),
    .Y(_17693_));
 sg13g2_a21o_2 _24657_ (.A2(_17693_),
    .A1(_17692_),
    .B1(_17691_),
    .X(_17694_));
 sg13g2_o21ai_1 _24658_ (.B1(_15565_),
    .Y(_17695_),
    .A1(_16308_),
    .A2(_16324_));
 sg13g2_o21ai_1 _24659_ (.B1(_16329_),
    .Y(_17696_),
    .A1(_16308_),
    .A2(_16324_));
 sg13g2_nand2_1 _24660_ (.Y(_17697_),
    .A(_16338_),
    .B(_17696_));
 sg13g2_a21oi_1 _24661_ (.A1(_16326_),
    .A2(_17697_),
    .Y(_17698_),
    .B1(_16334_));
 sg13g2_nor2_1 _24662_ (.A(_15130_),
    .B(_17698_),
    .Y(_17699_));
 sg13g2_or2_1 _24663_ (.X(_17700_),
    .B(_17699_),
    .A(_16332_));
 sg13g2_and2_1 _24664_ (.A(_15128_),
    .B(_17700_),
    .X(_17701_));
 sg13g2_o21ai_1 _24665_ (.B1(_15125_),
    .Y(_17702_),
    .A1(_16335_),
    .A2(_17701_));
 sg13g2_nand3_1 _24666_ (.B(_16343_),
    .C(_17702_),
    .A(_15123_),
    .Y(_17703_));
 sg13g2_a21oi_1 _24667_ (.A1(_16343_),
    .A2(_17702_),
    .Y(_17704_),
    .B1(_15123_));
 sg13g2_nand2_1 _24668_ (.Y(_17705_),
    .A(net5013),
    .B(_17703_));
 sg13g2_a21oi_2 _24669_ (.B1(_15139_),
    .Y(_17706_),
    .A2(_15566_),
    .A1(_15562_));
 sg13g2_o21ai_1 _24670_ (.B1(_15143_),
    .Y(_17707_),
    .A1(_15137_),
    .A2(_17706_));
 sg13g2_a21oi_1 _24671_ (.A1(_15131_),
    .A2(_17707_),
    .Y(_17708_),
    .B1(_15147_));
 sg13g2_o21ai_1 _24672_ (.B1(_15120_),
    .Y(_17709_),
    .A1(_15125_),
    .A2(_17708_));
 sg13g2_xnor2_1 _24673_ (.Y(_17710_),
    .A(_15123_),
    .B(_17709_));
 sg13g2_a21oi_1 _24674_ (.A1(net5826),
    .A2(_17710_),
    .Y(_17711_),
    .B1(net5013));
 sg13g2_o21ai_1 _24675_ (.B1(_17711_),
    .Y(_17712_),
    .A1(\u_inv.f_next[103] ),
    .A2(net5826));
 sg13g2_o21ai_1 _24676_ (.B1(_17712_),
    .Y(_17713_),
    .A1(_17704_),
    .A2(_17705_));
 sg13g2_xor2_1 _24677_ (.B(_16963_),
    .A(_14979_),
    .X(_17714_));
 sg13g2_nor2_1 _24678_ (.A(net5691),
    .B(_17714_),
    .Y(_17715_));
 sg13g2_o21ai_1 _24679_ (.B1(net5068),
    .Y(_17716_),
    .A1(\u_inv.f_next[162] ),
    .A2(net5782));
 sg13g2_nand3_1 _24680_ (.B(_16487_),
    .C(_17576_),
    .A(_14979_),
    .Y(_17717_));
 sg13g2_nand3_1 _24681_ (.B(_17577_),
    .C(_17717_),
    .A(net4977),
    .Y(_17718_));
 sg13g2_o21ai_1 _24682_ (.B1(_17718_),
    .Y(_17719_),
    .A1(_17715_),
    .A2(_17716_));
 sg13g2_nand3_1 _24683_ (.B(_15742_),
    .C(_17315_),
    .A(_15712_),
    .Y(_17720_));
 sg13g2_a21oi_1 _24684_ (.A1(_17316_),
    .A2(_17720_),
    .Y(_17721_),
    .B1(net5707));
 sg13g2_o21ai_1 _24685_ (.B1(net5085),
    .Y(_17722_),
    .A1(\u_inv.f_next[134] ),
    .A2(net5805));
 sg13g2_nor3_1 _24686_ (.A(_15712_),
    .B(_16438_),
    .C(_17310_),
    .Y(_17723_));
 sg13g2_nor2_1 _24687_ (.A(net5090),
    .B(_17723_),
    .Y(_17724_));
 sg13g2_nand2_1 _24688_ (.Y(_17725_),
    .A(_17311_),
    .B(_17724_));
 sg13g2_o21ai_1 _24689_ (.B1(_17725_),
    .Y(_17726_),
    .A1(_17721_),
    .A2(_17722_));
 sg13g2_nand3_1 _24690_ (.B(_15026_),
    .C(_16851_),
    .A(_14955_),
    .Y(_17727_));
 sg13g2_nand2b_1 _24691_ (.Y(_17728_),
    .B(_17727_),
    .A_N(_16991_));
 sg13g2_a21oi_1 _24692_ (.A1(net5777),
    .A2(_17728_),
    .Y(_17729_),
    .B1(net4975));
 sg13g2_o21ai_1 _24693_ (.B1(_17729_),
    .Y(_17730_),
    .A1(\u_inv.f_next[176] ),
    .A2(net5777));
 sg13g2_nor3_1 _24694_ (.A(_14955_),
    .B(_16514_),
    .C(_16860_),
    .Y(_17731_));
 sg13g2_nand2_1 _24695_ (.Y(_17732_),
    .A(net4975),
    .B(_17088_));
 sg13g2_o21ai_1 _24696_ (.B1(_17730_),
    .Y(_17733_),
    .A1(_17731_),
    .A2(_17732_));
 sg13g2_xnor2_1 _24697_ (.Y(_17734_),
    .A(_15793_),
    .B(_16548_));
 sg13g2_nand3_1 _24698_ (.B(_15773_),
    .C(_15794_),
    .A(_15049_),
    .Y(_17735_));
 sg13g2_nand3b_1 _24699_ (.B(_17735_),
    .C(net5763),
    .Y(_17736_),
    .A_N(_17032_));
 sg13g2_a21oi_1 _24700_ (.A1(\u_inv.f_next[192] ),
    .A2(net5681),
    .Y(_17737_),
    .B1(net4961));
 sg13g2_a22oi_1 _24701_ (.Y(_17738_),
    .B1(_17736_),
    .B2(_17737_),
    .A2(_17734_),
    .A1(net4961));
 sg13g2_xnor2_1 _24702_ (.Y(_17739_),
    .A(_15125_),
    .B(_17708_));
 sg13g2_nor2_1 _24703_ (.A(\u_inv.f_next[102] ),
    .B(net5825),
    .Y(_17740_));
 sg13g2_a21oi_1 _24704_ (.A1(net5824),
    .A2(_17739_),
    .Y(_17741_),
    .B1(_17740_));
 sg13g2_nor3_1 _24705_ (.A(_15125_),
    .B(_16335_),
    .C(_17701_),
    .Y(_17742_));
 sg13g2_nor2_1 _24706_ (.A(net5100),
    .B(_17742_),
    .Y(_17743_));
 sg13g2_a22oi_1 _24707_ (.Y(_17744_),
    .B1(_17743_),
    .B2(_17702_),
    .A2(_17741_),
    .A1(net5101));
 sg13g2_inv_1 _24708_ (.Y(_17745_),
    .A(_17744_));
 sg13g2_xnor2_1 _24709_ (.Y(_17746_),
    .A(_15575_),
    .B(_17632_));
 sg13g2_nor2_1 _24710_ (.A(\u_inv.f_next[110] ),
    .B(net5819),
    .Y(_17747_));
 sg13g2_o21ai_1 _24711_ (.B1(net5097),
    .Y(_17748_),
    .A1(net5715),
    .A2(_17746_));
 sg13g2_a21oi_1 _24712_ (.A1(_15575_),
    .A2(_17624_),
    .Y(_17749_),
    .B1(net5097));
 sg13g2_nand2b_1 _24713_ (.Y(_17750_),
    .B(_17749_),
    .A_N(_17625_));
 sg13g2_o21ai_1 _24714_ (.B1(_17750_),
    .Y(_17751_),
    .A1(_17747_),
    .A2(_17748_));
 sg13g2_nand2b_1 _24715_ (.Y(_17752_),
    .B(_16346_),
    .A_N(_15591_));
 sg13g2_a21o_1 _24716_ (.A2(_17752_),
    .A1(_16356_),
    .B1(_15592_),
    .X(_17753_));
 sg13g2_a21oi_1 _24717_ (.A1(_16355_),
    .A2(_17753_),
    .Y(_17754_),
    .B1(_15587_));
 sg13g2_nor3_1 _24718_ (.A(_15585_),
    .B(_16354_),
    .C(_17754_),
    .Y(_17755_));
 sg13g2_o21ai_1 _24719_ (.B1(_15585_),
    .Y(_17756_),
    .A1(_16354_),
    .A2(_17754_));
 sg13g2_nand2_1 _24720_ (.Y(_17757_),
    .A(net5011),
    .B(_17756_));
 sg13g2_o21ai_1 _24721_ (.B1(_15586_),
    .Y(_17758_),
    .A1(_15588_),
    .A2(_17630_));
 sg13g2_xnor2_1 _24722_ (.Y(_17759_),
    .A(_15584_),
    .B(_17758_));
 sg13g2_a21oi_1 _24723_ (.A1(net5826),
    .A2(_17759_),
    .Y(_17760_),
    .B1(net5011));
 sg13g2_o21ai_1 _24724_ (.B1(_17760_),
    .Y(_17761_),
    .A1(\u_inv.f_next[107] ),
    .A2(net5818));
 sg13g2_o21ai_1 _24725_ (.B1(_17761_),
    .Y(_17762_),
    .A1(_17755_),
    .A2(_17757_));
 sg13g2_a21oi_2 _24726_ (.B1(_16305_),
    .Y(_17763_),
    .A2(_16298_),
    .A1(_16291_));
 sg13g2_o21ai_1 _24727_ (.B1(_16303_),
    .Y(_17764_),
    .A1(_16314_),
    .A2(_17763_));
 sg13g2_a21o_1 _24728_ (.A2(_17764_),
    .A1(_16311_),
    .B1(_15533_),
    .X(_17765_));
 sg13g2_nand2_1 _24729_ (.Y(_17766_),
    .A(_16321_),
    .B(_17765_));
 sg13g2_nand2_1 _24730_ (.Y(_17767_),
    .A(_15535_),
    .B(_17766_));
 sg13g2_nand2_1 _24731_ (.Y(_17768_),
    .A(_16320_),
    .B(_17767_));
 sg13g2_and2_1 _24732_ (.A(_15532_),
    .B(_17768_),
    .X(_17769_));
 sg13g2_o21ai_1 _24733_ (.B1(_15530_),
    .Y(_17770_),
    .A1(_16318_),
    .A2(_17769_));
 sg13g2_nor3_1 _24734_ (.A(_15530_),
    .B(_16318_),
    .C(_17769_),
    .Y(_17771_));
 sg13g2_nand2_1 _24735_ (.Y(_17772_),
    .A(net5013),
    .B(_17770_));
 sg13g2_nand3_1 _24736_ (.B(_15527_),
    .C(_15549_),
    .A(_15168_),
    .Y(_17773_));
 sg13g2_a21oi_1 _24737_ (.A1(_15553_),
    .A2(_17773_),
    .Y(_17774_),
    .B1(_15541_));
 sg13g2_nor2_1 _24738_ (.A(_15560_),
    .B(_17774_),
    .Y(_17775_));
 sg13g2_or2_1 _24739_ (.X(_17776_),
    .B(_17775_),
    .A(_15536_));
 sg13g2_a21oi_1 _24740_ (.A1(_15555_),
    .A2(_17776_),
    .Y(_17777_),
    .B1(_15532_));
 sg13g2_nor2_1 _24741_ (.A(_15531_),
    .B(_17777_),
    .Y(_17778_));
 sg13g2_xnor2_1 _24742_ (.Y(_17779_),
    .A(_15530_),
    .B(_17778_));
 sg13g2_a21oi_1 _24743_ (.A1(net5821),
    .A2(_17779_),
    .Y(_17780_),
    .B1(net5013));
 sg13g2_o21ai_1 _24744_ (.B1(_17780_),
    .Y(_17781_),
    .A1(\u_inv.f_next[95] ),
    .A2(net5821));
 sg13g2_o21ai_1 _24745_ (.B1(_17781_),
    .Y(_17782_),
    .A1(_17771_),
    .A2(_17772_));
 sg13g2_xnor2_1 _24746_ (.Y(_17783_),
    .A(_15130_),
    .B(_17707_));
 sg13g2_o21ai_1 _24747_ (.B1(net5100),
    .Y(_17784_),
    .A1(\u_inv.f_next[100] ),
    .A2(net5825));
 sg13g2_a21o_1 _24748_ (.A2(_17783_),
    .A1(net5825),
    .B1(_17784_),
    .X(_17785_));
 sg13g2_xnor2_1 _24749_ (.Y(_17786_),
    .A(_15130_),
    .B(_17698_));
 sg13g2_o21ai_1 _24750_ (.B1(_17785_),
    .Y(_17787_),
    .A1(net5100),
    .A2(_17786_));
 sg13g2_a21oi_1 _24751_ (.A1(_15610_),
    .A2(_15650_),
    .Y(_17788_),
    .B1(net5715));
 sg13g2_xnor2_1 _24752_ (.Y(_17789_),
    .A(_15649_),
    .B(_16369_));
 sg13g2_a221oi_1 _24753_ (.B2(_17788_),
    .C1(net5011),
    .B1(_17478_),
    .A1(\u_inv.f_next[112] ),
    .Y(_17790_),
    .A2(net5715));
 sg13g2_a21oi_1 _24754_ (.A1(net5011),
    .A2(_17789_),
    .Y(_17791_),
    .B1(_17790_));
 sg13g2_xor2_1 _24755_ (.B(_17621_),
    .A(_15581_),
    .X(_17792_));
 sg13g2_xnor2_1 _24756_ (.Y(_17793_),
    .A(_15581_),
    .B(_17631_));
 sg13g2_o21ai_1 _24757_ (.B1(net5097),
    .Y(_17794_),
    .A1(_14066_),
    .A2(net5818));
 sg13g2_a21oi_1 _24758_ (.A1(net5818),
    .A2(_17793_),
    .Y(_17795_),
    .B1(_17794_));
 sg13g2_a21oi_1 _24759_ (.A1(net5011),
    .A2(_17792_),
    .Y(_17796_),
    .B1(_17795_));
 sg13g2_o21ai_1 _24760_ (.B1(_15533_),
    .Y(_17797_),
    .A1(_15560_),
    .A2(_17774_));
 sg13g2_o21ai_1 _24761_ (.B1(_17797_),
    .Y(_17798_),
    .A1(_14082_),
    .A2(_14346_));
 sg13g2_xnor2_1 _24762_ (.Y(_17799_),
    .A(_15534_),
    .B(_17798_));
 sg13g2_o21ai_1 _24763_ (.B1(net5098),
    .Y(_17800_),
    .A1(\u_inv.f_next[93] ),
    .A2(net5822));
 sg13g2_a21oi_1 _24764_ (.A1(net5822),
    .A2(_17799_),
    .Y(_17801_),
    .B1(_17800_));
 sg13g2_nor2_1 _24765_ (.A(_15535_),
    .B(_17766_),
    .Y(_17802_));
 sg13g2_nor2_1 _24766_ (.A(net5098),
    .B(_17802_),
    .Y(_17803_));
 sg13g2_a21oi_1 _24767_ (.A1(_17767_),
    .A2(_17803_),
    .Y(_17804_),
    .B1(_17801_));
 sg13g2_inv_4 _24768_ (.A(_17804_),
    .Y(_17805_));
 sg13g2_nand2_1 _24769_ (.Y(_17806_),
    .A(_15136_),
    .B(_17697_));
 sg13g2_a21o_1 _24770_ (.A2(_17806_),
    .A1(_16333_),
    .B1(_15133_),
    .X(_17807_));
 sg13g2_nand3_1 _24771_ (.B(_16333_),
    .C(_17806_),
    .A(_15133_),
    .Y(_17808_));
 sg13g2_nand3_1 _24772_ (.B(_17807_),
    .C(_17808_),
    .A(net5013),
    .Y(_17809_));
 sg13g2_o21ai_1 _24773_ (.B1(_15134_),
    .Y(_17810_),
    .A1(_15136_),
    .A2(_17706_));
 sg13g2_xor2_1 _24774_ (.B(_17810_),
    .A(_15133_),
    .X(_17811_));
 sg13g2_nor2_1 _24775_ (.A(net5715),
    .B(_17811_),
    .Y(_17812_));
 sg13g2_o21ai_1 _24776_ (.B1(net5100),
    .Y(_17813_),
    .A1(\u_inv.f_next[99] ),
    .A2(net5824));
 sg13g2_o21ai_1 _24777_ (.B1(_17809_),
    .Y(_17814_),
    .A1(_17812_),
    .A2(_17813_));
 sg13g2_a21oi_1 _24778_ (.A1(_15570_),
    .A2(_15591_),
    .Y(_17815_),
    .B1(_15590_));
 sg13g2_xor2_1 _24779_ (.B(_17815_),
    .A(_15592_),
    .X(_17816_));
 sg13g2_o21ai_1 _24780_ (.B1(net5097),
    .Y(_17817_),
    .A1(\u_inv.f_next[105] ),
    .A2(net5818));
 sg13g2_a21oi_1 _24781_ (.A1(net5818),
    .A2(_17816_),
    .Y(_17818_),
    .B1(_17817_));
 sg13g2_nand3_1 _24782_ (.B(_16356_),
    .C(_17752_),
    .A(_15592_),
    .Y(_17819_));
 sg13g2_nand3_1 _24783_ (.B(_17753_),
    .C(_17819_),
    .A(net5012),
    .Y(_17820_));
 sg13g2_nor2b_1 _24784_ (.A(_17818_),
    .B_N(_17820_),
    .Y(_17821_));
 sg13g2_inv_1 _24785_ (.Y(_17822_),
    .A(_17821_));
 sg13g2_xnor2_1 _24786_ (.Y(_17823_),
    .A(_15528_),
    .B(_15548_));
 sg13g2_o21ai_1 _24787_ (.B1(net5099),
    .Y(_17824_),
    .A1(\u_inv.f_next[88] ),
    .A2(net5821));
 sg13g2_a21o_1 _24788_ (.A2(_17823_),
    .A1(net5821),
    .B1(_17824_),
    .X(_17825_));
 sg13g2_nand2_1 _24789_ (.Y(_17826_),
    .A(_15548_),
    .B(_16299_));
 sg13g2_xnor2_1 _24790_ (.Y(_17827_),
    .A(_15548_),
    .B(_16299_));
 sg13g2_o21ai_1 _24791_ (.B1(_17825_),
    .Y(_17828_),
    .A1(net5099),
    .A2(_17827_));
 sg13g2_nor3_1 _24792_ (.A(_15509_),
    .B(_15517_),
    .C(_15519_),
    .Y(_17829_));
 sg13g2_or2_1 _24793_ (.X(_17830_),
    .B(_17829_),
    .A(_15522_));
 sg13g2_xnor2_1 _24794_ (.Y(_17831_),
    .A(_15513_),
    .B(_17830_));
 sg13g2_a21oi_1 _24795_ (.A1(net5806),
    .A2(_17831_),
    .Y(_17832_),
    .B1(net5000));
 sg13g2_o21ai_1 _24796_ (.B1(_17832_),
    .Y(_17833_),
    .A1(\u_inv.f_next[82] ),
    .A2(net5806));
 sg13g2_a21oi_1 _24797_ (.A1(_16263_),
    .A2(_16278_),
    .Y(_17834_),
    .B1(_15516_));
 sg13g2_o21ai_1 _24798_ (.B1(_15519_),
    .Y(_17835_),
    .A1(_16284_),
    .A2(_17834_));
 sg13g2_nand3_1 _24799_ (.B(_16283_),
    .C(_17835_),
    .A(_15513_),
    .Y(_17836_));
 sg13g2_a21oi_1 _24800_ (.A1(_16283_),
    .A2(_17835_),
    .Y(_17837_),
    .B1(_15513_));
 sg13g2_nand2_1 _24801_ (.Y(_17838_),
    .A(net5000),
    .B(_17836_));
 sg13g2_o21ai_1 _24802_ (.B1(_17833_),
    .Y(_17839_),
    .A1(_17837_),
    .A2(_17838_));
 sg13g2_nand3_1 _24803_ (.B(_16312_),
    .C(_17826_),
    .A(_15545_),
    .Y(_17840_));
 sg13g2_nor3_1 _24804_ (.A(net5099),
    .B(_16313_),
    .C(_17763_),
    .Y(_17841_));
 sg13g2_o21ai_1 _24805_ (.B1(_15546_),
    .Y(_17842_),
    .A1(_15528_),
    .A2(_15548_));
 sg13g2_xnor2_1 _24806_ (.Y(_17843_),
    .A(_15545_),
    .B(_17842_));
 sg13g2_o21ai_1 _24807_ (.B1(net5098),
    .Y(_17844_),
    .A1(\u_inv.f_next[89] ),
    .A2(net5821));
 sg13g2_a21oi_1 _24808_ (.A1(net5821),
    .A2(_17843_),
    .Y(_17845_),
    .B1(_17844_));
 sg13g2_a21oi_2 _24809_ (.B1(_17845_),
    .Y(_17846_),
    .A2(_17841_),
    .A1(_17840_));
 sg13g2_inv_1 _24810_ (.Y(_17847_),
    .A(_17846_));
 sg13g2_a21o_2 _24811_ (.A2(_16238_),
    .A1(_16222_),
    .B1(_15467_),
    .X(_17848_));
 sg13g2_a21o_1 _24812_ (.A2(_17848_),
    .A1(_16247_),
    .B1(_15469_),
    .X(_17849_));
 sg13g2_a21o_1 _24813_ (.A2(_17849_),
    .A1(_16246_),
    .B1(_15181_),
    .X(_17850_));
 sg13g2_a21oi_1 _24814_ (.A1(_16245_),
    .A2(_17850_),
    .Y(_17851_),
    .B1(_15180_));
 sg13g2_nand3_1 _24815_ (.B(_16245_),
    .C(_17850_),
    .A(_15180_),
    .Y(_17852_));
 sg13g2_nand2_1 _24816_ (.Y(_17853_),
    .A(net4979),
    .B(_17852_));
 sg13g2_a21oi_1 _24817_ (.A1(_15466_),
    .A2(_15470_),
    .Y(_17854_),
    .B1(_15187_));
 sg13g2_nor2b_1 _24818_ (.A(_17854_),
    .B_N(_15181_),
    .Y(_17855_));
 sg13g2_a21oi_1 _24819_ (.A1(\u_inv.f_next[66] ),
    .A2(\u_inv.f_reg[66] ),
    .Y(_17856_),
    .B1(_17855_));
 sg13g2_xor2_1 _24820_ (.B(_17856_),
    .A(_15180_),
    .X(_17857_));
 sg13g2_a21oi_1 _24821_ (.A1(net5781),
    .A2(_17857_),
    .Y(_17858_),
    .B1(net4979));
 sg13g2_o21ai_1 _24822_ (.B1(_17858_),
    .Y(_17859_),
    .A1(\u_inv.f_next[67] ),
    .A2(net5781));
 sg13g2_o21ai_1 _24823_ (.B1(_17859_),
    .Y(_17860_),
    .A1(_17851_),
    .A2(_17853_));
 sg13g2_o21ai_1 _24824_ (.B1(_15515_),
    .Y(_17861_),
    .A1(_15509_),
    .A2(_15517_));
 sg13g2_a21oi_1 _24825_ (.A1(_15519_),
    .A2(_17861_),
    .Y(_17862_),
    .B1(net5706));
 sg13g2_o21ai_1 _24826_ (.B1(_17862_),
    .Y(_17863_),
    .A1(_15519_),
    .A2(_17861_));
 sg13g2_a21oi_1 _24827_ (.A1(_14093_),
    .A2(net5706),
    .Y(_17864_),
    .B1(net5000));
 sg13g2_nor3_1 _24828_ (.A(_15519_),
    .B(_16284_),
    .C(_17834_),
    .Y(_17865_));
 sg13g2_nand2_1 _24829_ (.Y(_17866_),
    .A(net5000),
    .B(_17835_));
 sg13g2_nor2_1 _24830_ (.A(_17865_),
    .B(_17866_),
    .Y(_17867_));
 sg13g2_a21oi_1 _24831_ (.A1(_17863_),
    .A2(_17864_),
    .Y(_17868_),
    .B1(_17867_));
 sg13g2_inv_1 _24832_ (.Y(_17869_),
    .A(_17868_));
 sg13g2_a21oi_1 _24833_ (.A1(_15474_),
    .A2(_15497_),
    .Y(_17870_),
    .B1(_15500_));
 sg13g2_xnor2_1 _24834_ (.Y(_17871_),
    .A(_15488_),
    .B(_17870_));
 sg13g2_o21ai_1 _24835_ (.B1(net5076),
    .Y(_17872_),
    .A1(net5698),
    .A2(_17871_));
 sg13g2_a21o_1 _24836_ (.A2(net5698),
    .A1(_14100_),
    .B1(_17872_),
    .X(_17873_));
 sg13g2_o21ai_1 _24837_ (.B1(_15494_),
    .Y(_17874_),
    .A1(_16244_),
    .A2(_16257_));
 sg13g2_a21oi_1 _24838_ (.A1(_16272_),
    .A2(_17874_),
    .Y(_17875_),
    .B1(_15495_));
 sg13g2_nor3_1 _24839_ (.A(_15489_),
    .B(_16271_),
    .C(_17875_),
    .Y(_17876_));
 sg13g2_o21ai_1 _24840_ (.B1(_15489_),
    .Y(_17877_),
    .A1(_16271_),
    .A2(_17875_));
 sg13g2_nand2_1 _24841_ (.Y(_17878_),
    .A(net4989),
    .B(_17877_));
 sg13g2_o21ai_1 _24842_ (.B1(_17873_),
    .Y(_17879_),
    .A1(_17876_),
    .A2(_17878_));
 sg13g2_o21ai_1 _24843_ (.B1(_15525_),
    .Y(_17880_),
    .A1(_15509_),
    .A2(_15520_));
 sg13g2_nand2_1 _24844_ (.Y(_17881_),
    .A(_15164_),
    .B(_17880_));
 sg13g2_xnor2_1 _24845_ (.Y(_17882_),
    .A(_15164_),
    .B(_17880_));
 sg13g2_o21ai_1 _24846_ (.B1(net5089),
    .Y(_17883_),
    .A1(\u_inv.f_next[84] ),
    .A2(net5810));
 sg13g2_a21oi_1 _24847_ (.A1(net5810),
    .A2(_17882_),
    .Y(_17884_),
    .B1(_17883_));
 sg13g2_nor3_1 _24848_ (.A(_15165_),
    .B(_16281_),
    .C(_16288_),
    .Y(_17885_));
 sg13g2_o21ai_1 _24849_ (.B1(_15165_),
    .Y(_17886_),
    .A1(_16281_),
    .A2(_16288_));
 sg13g2_nor2_1 _24850_ (.A(net5089),
    .B(_17885_),
    .Y(_17887_));
 sg13g2_a21o_2 _24851_ (.A2(_17887_),
    .A1(_17886_),
    .B1(_17884_),
    .X(_17888_));
 sg13g2_o21ai_1 _24852_ (.B1(_15452_),
    .Y(_17889_),
    .A1(_15426_),
    .A2(_15446_));
 sg13g2_a21oi_2 _24853_ (.B1(_15455_),
    .Y(_17890_),
    .A2(_17889_),
    .A1(_15441_));
 sg13g2_nor3_1 _24854_ (.A(_15434_),
    .B(_15436_),
    .C(_17890_),
    .Y(_17891_));
 sg13g2_nor2_1 _24855_ (.A(_15450_),
    .B(_17891_),
    .Y(_17892_));
 sg13g2_xnor2_1 _24856_ (.Y(_17893_),
    .A(_15431_),
    .B(_17892_));
 sg13g2_nor2_1 _24857_ (.A(net5680),
    .B(_17893_),
    .Y(_17894_));
 sg13g2_o21ai_1 _24858_ (.B1(net5057),
    .Y(_17895_),
    .A1(\u_inv.f_next[54] ),
    .A2(net5768));
 sg13g2_o21ai_1 _24859_ (.B1(_15444_),
    .Y(_17896_),
    .A1(_16175_),
    .A2(_16191_));
 sg13g2_o21ai_1 _24860_ (.B1(_16195_),
    .Y(_17897_),
    .A1(_16175_),
    .A2(_16191_));
 sg13g2_nand2_1 _24861_ (.Y(_17898_),
    .A(_16203_),
    .B(_17897_));
 sg13g2_a21oi_1 _24862_ (.A1(_16203_),
    .A2(_17897_),
    .Y(_17899_),
    .B1(_16193_));
 sg13g2_o21ai_1 _24863_ (.B1(_15436_),
    .Y(_17900_),
    .A1(_16209_),
    .A2(_17899_));
 sg13g2_inv_1 _24864_ (.Y(_17901_),
    .A(_17900_));
 sg13g2_o21ai_1 _24865_ (.B1(_15434_),
    .Y(_17902_),
    .A1(_16206_),
    .A2(_17901_));
 sg13g2_nand3_1 _24866_ (.B(_16205_),
    .C(_17902_),
    .A(_15431_),
    .Y(_17903_));
 sg13g2_a21o_1 _24867_ (.A2(_17902_),
    .A1(_16205_),
    .B1(_15431_),
    .X(_17904_));
 sg13g2_nand3_1 _24868_ (.B(_17903_),
    .C(_17904_),
    .A(net4964),
    .Y(_17905_));
 sg13g2_o21ai_1 _24869_ (.B1(_17905_),
    .Y(_17906_),
    .A1(_17894_),
    .A2(_17895_));
 sg13g2_xnor2_1 _24870_ (.Y(_17907_),
    .A(_15181_),
    .B(_17854_));
 sg13g2_nor2_1 _24871_ (.A(\u_inv.f_next[66] ),
    .B(net5781),
    .Y(_17908_));
 sg13g2_o21ai_1 _24872_ (.B1(net5067),
    .Y(_17909_),
    .A1(net5690),
    .A2(_17907_));
 sg13g2_nand3_1 _24873_ (.B(_16246_),
    .C(_17849_),
    .A(_15181_),
    .Y(_17910_));
 sg13g2_nand3_1 _24874_ (.B(_17850_),
    .C(_17910_),
    .A(net4979),
    .Y(_17911_));
 sg13g2_o21ai_1 _24875_ (.B1(_17911_),
    .Y(_17912_),
    .A1(_17908_),
    .A2(_17909_));
 sg13g2_xnor2_1 _24876_ (.Y(_17913_),
    .A(_15509_),
    .B(_15516_));
 sg13g2_nor2_1 _24877_ (.A(\u_inv.f_next[80] ),
    .B(net5806),
    .Y(_17914_));
 sg13g2_o21ai_1 _24878_ (.B1(net5085),
    .Y(_17915_),
    .A1(net5706),
    .A2(_17913_));
 sg13g2_nand3_1 _24879_ (.B(_16263_),
    .C(_16278_),
    .A(_15516_),
    .Y(_17916_));
 sg13g2_nor2_1 _24880_ (.A(net5085),
    .B(_17834_),
    .Y(_17917_));
 sg13g2_nand2_1 _24881_ (.Y(_17918_),
    .A(_17916_),
    .B(_17917_));
 sg13g2_o21ai_1 _24882_ (.B1(_17918_),
    .Y(_17919_),
    .A1(_17914_),
    .A2(_17915_));
 sg13g2_nor2_1 _24883_ (.A(_17912_),
    .B(_17919_),
    .Y(_17920_));
 sg13g2_a21o_2 _24884_ (.A2(_16147_),
    .A1(_16138_),
    .B1(_15390_),
    .X(_17921_));
 sg13g2_a21o_1 _24885_ (.A2(_17921_),
    .A1(_16153_),
    .B1(_16149_),
    .X(_17922_));
 sg13g2_a21oi_1 _24886_ (.A1(_16158_),
    .A2(_17922_),
    .Y(_17923_),
    .B1(_15232_));
 sg13g2_o21ai_1 _24887_ (.B1(_15235_),
    .Y(_17924_),
    .A1(_16161_),
    .A2(_17923_));
 sg13g2_a21o_1 _24888_ (.A2(_17924_),
    .A1(_16160_),
    .B1(_15229_),
    .X(_17925_));
 sg13g2_nand3_1 _24889_ (.B(_16163_),
    .C(_17925_),
    .A(_15226_),
    .Y(_17926_));
 sg13g2_a21oi_1 _24890_ (.A1(_16163_),
    .A2(_17925_),
    .Y(_17927_),
    .B1(_15226_));
 sg13g2_nand2_1 _24891_ (.Y(_17928_),
    .A(net4951),
    .B(_17926_));
 sg13g2_a21oi_1 _24892_ (.A1(_15387_),
    .A2(_15391_),
    .Y(_17929_),
    .B1(_15245_));
 sg13g2_nor2b_1 _24893_ (.A(_17929_),
    .B_N(_15242_),
    .Y(_17930_));
 sg13g2_nor2_1 _24894_ (.A(_15247_),
    .B(_17930_),
    .Y(_17931_));
 sg13g2_nor2b_1 _24895_ (.A(_17931_),
    .B_N(_15236_),
    .Y(_17932_));
 sg13g2_nor2_1 _24896_ (.A(_15250_),
    .B(_17932_),
    .Y(_17933_));
 sg13g2_o21ai_1 _24897_ (.B1(_15227_),
    .Y(_17934_),
    .A1(_15228_),
    .A2(_17933_));
 sg13g2_xnor2_1 _24898_ (.Y(_17935_),
    .A(_15226_),
    .B(_17934_));
 sg13g2_a21oi_1 _24899_ (.A1(net5749),
    .A2(_17935_),
    .Y(_17936_),
    .B1(net4951));
 sg13g2_o21ai_1 _24900_ (.B1(_17936_),
    .Y(_17937_),
    .A1(\u_inv.f_next[39] ),
    .A2(net5750));
 sg13g2_o21ai_1 _24901_ (.B1(_17937_),
    .Y(_17938_),
    .A1(_17927_),
    .A2(_17928_));
 sg13g2_a21oi_2 _24902_ (.B1(_16219_),
    .Y(_17939_),
    .A2(_16214_),
    .A1(_16199_));
 sg13g2_o21ai_1 _24903_ (.B1(_15211_),
    .Y(_17940_),
    .A1(_16227_),
    .A2(_17939_));
 sg13g2_nor2b_1 _24904_ (.A(_16224_),
    .B_N(_17940_),
    .Y(_17941_));
 sg13g2_a21oi_1 _24905_ (.A1(_15208_),
    .A2(_17941_),
    .Y(_17942_),
    .B1(net5065));
 sg13g2_o21ai_1 _24906_ (.B1(_17942_),
    .Y(_17943_),
    .A1(_15208_),
    .A2(_17941_));
 sg13g2_a21oi_2 _24907_ (.B1(_15215_),
    .Y(_17944_),
    .A2(_15463_),
    .A1(_15459_));
 sg13g2_o21ai_1 _24908_ (.B1(_15209_),
    .Y(_17945_),
    .A1(_15211_),
    .A2(_17944_));
 sg13g2_xnor2_1 _24909_ (.Y(_17946_),
    .A(_15208_),
    .B(_17945_));
 sg13g2_a21oi_1 _24910_ (.A1(net5780),
    .A2(_17946_),
    .Y(_17947_),
    .B1(net4974));
 sg13g2_o21ai_1 _24911_ (.B1(_17947_),
    .Y(_17948_),
    .A1(net3109),
    .A2(net5780));
 sg13g2_nand2_1 _24912_ (.Y(_17949_),
    .A(_17943_),
    .B(_17948_));
 sg13g2_a21oi_1 _24913_ (.A1(_16167_),
    .A2(_16172_),
    .Y(_17950_),
    .B1(_16182_));
 sg13g2_a21o_1 _24914_ (.A2(_15400_),
    .A1(_15399_),
    .B1(_17950_),
    .X(_17951_));
 sg13g2_a21oi_1 _24915_ (.A1(_16185_),
    .A2(_17951_),
    .Y(_17952_),
    .B1(_15402_));
 sg13g2_o21ai_1 _24916_ (.B1(_15397_),
    .Y(_17953_),
    .A1(_16184_),
    .A2(_17952_));
 sg13g2_nand2b_1 _24917_ (.Y(_17954_),
    .B(_17953_),
    .A_N(_16188_));
 sg13g2_a21oi_1 _24918_ (.A1(_15395_),
    .A2(_17954_),
    .Y(_17955_),
    .B1(net5054));
 sg13g2_o21ai_1 _24919_ (.B1(_17955_),
    .Y(_17956_),
    .A1(_15395_),
    .A2(_17954_));
 sg13g2_a21oi_2 _24920_ (.B1(_15417_),
    .Y(_17957_),
    .A2(_15414_),
    .A1(_15394_));
 sg13g2_nor2b_1 _24921_ (.A(_17957_),
    .B_N(_15408_),
    .Y(_17958_));
 sg13g2_nor2_1 _24922_ (.A(_15419_),
    .B(_17958_),
    .Y(_17959_));
 sg13g2_or2_1 _24923_ (.X(_17960_),
    .B(_17958_),
    .A(_15419_));
 sg13g2_a21oi_1 _24924_ (.A1(_15403_),
    .A2(_17960_),
    .Y(_17961_),
    .B1(_15423_));
 sg13g2_o21ai_1 _24925_ (.B1(_15396_),
    .Y(_17962_),
    .A1(_15397_),
    .A2(_17961_));
 sg13g2_xor2_1 _24926_ (.B(_17962_),
    .A(_15395_),
    .X(_17963_));
 sg13g2_a21oi_1 _24927_ (.A1(net5765),
    .A2(_17963_),
    .Y(_17964_),
    .B1(net4961));
 sg13g2_o21ai_1 _24928_ (.B1(_17964_),
    .Y(_17965_),
    .A1(\u_inv.f_next[47] ),
    .A2(net5765));
 sg13g2_nand2_2 _24929_ (.Y(_17966_),
    .A(_17956_),
    .B(_17965_));
 sg13g2_xnor2_1 _24930_ (.Y(_17967_),
    .A(_15474_),
    .B(_15493_));
 sg13g2_nand2_1 _24931_ (.Y(_17968_),
    .A(net5793),
    .B(_17967_));
 sg13g2_o21ai_1 _24932_ (.B1(_17968_),
    .Y(_17969_),
    .A1(\u_inv.f_next[72] ),
    .A2(net5793));
 sg13g2_or3_1 _24933_ (.A(_15494_),
    .B(_16244_),
    .C(_16257_),
    .X(_17970_));
 sg13g2_nand3_1 _24934_ (.B(_17874_),
    .C(_17970_),
    .A(net4989),
    .Y(_17971_));
 sg13g2_o21ai_1 _24935_ (.B1(_17971_),
    .Y(_17972_),
    .A1(net4989),
    .A2(_17969_));
 sg13g2_nand2_1 _24936_ (.Y(_17973_),
    .A(_15466_),
    .B(_15467_));
 sg13g2_nand2_1 _24937_ (.Y(_17974_),
    .A(_15186_),
    .B(_17973_));
 sg13g2_xor2_1 _24938_ (.B(_17974_),
    .A(_15469_),
    .X(_17975_));
 sg13g2_nor2_1 _24939_ (.A(net5690),
    .B(_17975_),
    .Y(_17976_));
 sg13g2_o21ai_1 _24940_ (.B1(net5067),
    .Y(_17977_),
    .A1(\u_inv.f_next[65] ),
    .A2(net5781));
 sg13g2_nand3_1 _24941_ (.B(_16247_),
    .C(_17848_),
    .A(_15469_),
    .Y(_17978_));
 sg13g2_nand3_1 _24942_ (.B(_17849_),
    .C(_17978_),
    .A(net4979),
    .Y(_17979_));
 sg13g2_o21ai_1 _24943_ (.B1(_17979_),
    .Y(_17980_),
    .A1(_17976_),
    .A2(_17977_));
 sg13g2_o21ai_1 _24944_ (.B1(_15435_),
    .Y(_17981_),
    .A1(_15436_),
    .A2(_17890_));
 sg13g2_xor2_1 _24945_ (.B(_17981_),
    .A(_15434_),
    .X(_17982_));
 sg13g2_o21ai_1 _24946_ (.B1(net5057),
    .Y(_17983_),
    .A1(\u_inv.f_next[53] ),
    .A2(net5768));
 sg13g2_a21oi_1 _24947_ (.A1(net5768),
    .A2(_17982_),
    .Y(_17984_),
    .B1(_17983_));
 sg13g2_nor3_1 _24948_ (.A(_15434_),
    .B(_16206_),
    .C(_17901_),
    .Y(_17985_));
 sg13g2_nor2_1 _24949_ (.A(net5057),
    .B(_17985_),
    .Y(_17986_));
 sg13g2_a21o_2 _24950_ (.A2(_17986_),
    .A1(_17902_),
    .B1(_17984_),
    .X(_17987_));
 sg13g2_xnor2_1 _24951_ (.Y(_17988_),
    .A(_15211_),
    .B(_17944_));
 sg13g2_nor2_1 _24952_ (.A(\u_inv.f_next[58] ),
    .B(net5780),
    .Y(_17989_));
 sg13g2_a21oi_1 _24953_ (.A1(net5780),
    .A2(_17988_),
    .Y(_17990_),
    .B1(_17989_));
 sg13g2_nor3_1 _24954_ (.A(_15211_),
    .B(_16227_),
    .C(_17939_),
    .Y(_17991_));
 sg13g2_nor2_1 _24955_ (.A(net5065),
    .B(_17991_),
    .Y(_17992_));
 sg13g2_a22oi_1 _24956_ (.Y(_17993_),
    .B1(_17992_),
    .B2(_17940_),
    .A2(_17990_),
    .A1(net5065));
 sg13g2_inv_2 _24957_ (.Y(_17994_),
    .A(_17993_));
 sg13g2_nand2_1 _24958_ (.Y(_17995_),
    .A(_15410_),
    .B(_16167_));
 sg13g2_a21oi_1 _24959_ (.A1(_16178_),
    .A2(_17995_),
    .Y(_17996_),
    .B1(_15411_));
 sg13g2_o21ai_1 _24960_ (.B1(net5620),
    .Y(_17997_),
    .A1(_16177_),
    .A2(_17996_));
 sg13g2_nand2b_1 _24961_ (.Y(_17998_),
    .B(_17997_),
    .A_N(_16176_));
 sg13g2_a21oi_1 _24962_ (.A1(_15405_),
    .A2(_17998_),
    .Y(_17999_),
    .B1(net5046));
 sg13g2_o21ai_1 _24963_ (.B1(_17999_),
    .Y(_18000_),
    .A1(_15405_),
    .A2(_17998_));
 sg13g2_o21ai_1 _24964_ (.B1(_15406_),
    .Y(_18001_),
    .A1(net5620),
    .A2(_17957_));
 sg13g2_xor2_1 _24965_ (.B(_18001_),
    .A(_15405_),
    .X(_18002_));
 sg13g2_a21oi_1 _24966_ (.A1(net5753),
    .A2(_18002_),
    .Y(_18003_),
    .B1(net4955));
 sg13g2_o21ai_1 _24967_ (.B1(_18003_),
    .Y(_18004_),
    .A1(net2698),
    .A2(net5753));
 sg13g2_nand2_1 _24968_ (.Y(_18005_),
    .A(_18000_),
    .B(_18004_));
 sg13g2_xnor2_1 _24969_ (.Y(_18006_),
    .A(_15397_),
    .B(_17961_));
 sg13g2_o21ai_1 _24970_ (.B1(net5054),
    .Y(_18007_),
    .A1(\u_inv.f_next[46] ),
    .A2(net5765));
 sg13g2_a21oi_1 _24971_ (.A1(net5765),
    .A2(_18006_),
    .Y(_18008_),
    .B1(_18007_));
 sg13g2_nor3_1 _24972_ (.A(_15397_),
    .B(_16184_),
    .C(_17952_),
    .Y(_18009_));
 sg13g2_nor2_1 _24973_ (.A(net5054),
    .B(_18009_),
    .Y(_18010_));
 sg13g2_a21o_2 _24974_ (.A2(_18010_),
    .A1(_17953_),
    .B1(_18008_),
    .X(_18011_));
 sg13g2_o21ai_1 _24975_ (.B1(_16258_),
    .Y(_18012_),
    .A1(_16244_),
    .A2(_16257_));
 sg13g2_a21oi_1 _24976_ (.A1(_16276_),
    .A2(_18012_),
    .Y(_18013_),
    .B1(_15482_));
 sg13g2_nand3_1 _24977_ (.B(_16276_),
    .C(_18012_),
    .A(_15482_),
    .Y(_18014_));
 sg13g2_nand2b_1 _24978_ (.Y(_18015_),
    .B(_18014_),
    .A_N(_18013_));
 sg13g2_nor2_1 _24979_ (.A(_15491_),
    .B(_17870_),
    .Y(_18016_));
 sg13g2_nor2_1 _24980_ (.A(_15502_),
    .B(_18016_),
    .Y(_18017_));
 sg13g2_or2_1 _24981_ (.X(_18018_),
    .B(_18016_),
    .A(_15502_));
 sg13g2_a21oi_1 _24982_ (.A1(_15483_),
    .A2(_18017_),
    .Y(_18019_),
    .B1(net5697));
 sg13g2_o21ai_1 _24983_ (.B1(_18019_),
    .Y(_18020_),
    .A1(_15483_),
    .A2(_18017_));
 sg13g2_a21oi_1 _24984_ (.A1(\u_inv.f_next[76] ),
    .A2(net5697),
    .Y(_18021_),
    .B1(net4990));
 sg13g2_a22oi_1 _24985_ (.Y(_18022_),
    .B1(_18020_),
    .B2(_18021_),
    .A2(_18015_),
    .A1(net4990));
 sg13g2_o21ai_1 _24986_ (.B1(_15492_),
    .Y(_18023_),
    .A1(_15473_),
    .A2(_15494_));
 sg13g2_xnor2_1 _24987_ (.Y(_18024_),
    .A(_15495_),
    .B(_18023_));
 sg13g2_o21ai_1 _24988_ (.B1(net5076),
    .Y(_18025_),
    .A1(\u_inv.f_next[73] ),
    .A2(net5793));
 sg13g2_a21oi_1 _24989_ (.A1(net5793),
    .A2(_18024_),
    .Y(_18026_),
    .B1(_18025_));
 sg13g2_nand3_1 _24990_ (.B(_16272_),
    .C(_17874_),
    .A(_15495_),
    .Y(_18027_));
 sg13g2_nor2_1 _24991_ (.A(net5076),
    .B(_17875_),
    .Y(_18028_));
 sg13g2_a21oi_1 _24992_ (.A1(_18027_),
    .A2(_18028_),
    .Y(_18029_),
    .B1(_18026_));
 sg13g2_inv_1 _24993_ (.Y(_18030_),
    .A(_18029_));
 sg13g2_nand3_1 _24994_ (.B(_16212_),
    .C(_17904_),
    .A(_15428_),
    .Y(_18031_));
 sg13g2_a21oi_1 _24995_ (.A1(_16212_),
    .A2(_17904_),
    .Y(_18032_),
    .B1(_15428_));
 sg13g2_nand2_1 _24996_ (.Y(_18033_),
    .A(net4964),
    .B(_18031_));
 sg13g2_o21ai_1 _24997_ (.B1(_15430_),
    .Y(_18034_),
    .A1(_15432_),
    .A2(_17892_));
 sg13g2_xnor2_1 _24998_ (.Y(_18035_),
    .A(_15428_),
    .B(_18034_));
 sg13g2_a21oi_1 _24999_ (.A1(net5768),
    .A2(_18035_),
    .Y(_18036_),
    .B1(net4964));
 sg13g2_o21ai_1 _25000_ (.B1(_18036_),
    .Y(_18037_),
    .A1(\u_inv.f_next[55] ),
    .A2(net5768));
 sg13g2_o21ai_1 _25001_ (.B1(_18037_),
    .Y(_18038_),
    .A1(_18032_),
    .A2(_18033_));
 sg13g2_o21ai_1 _25002_ (.B1(_15481_),
    .Y(_18039_),
    .A1(_15483_),
    .A2(_18017_));
 sg13g2_xor2_1 _25003_ (.B(_18039_),
    .A(_15480_),
    .X(_18040_));
 sg13g2_o21ai_1 _25004_ (.B1(net5079),
    .Y(_18041_),
    .A1(\u_inv.f_next[77] ),
    .A2(net5797));
 sg13g2_a21o_1 _25005_ (.A2(_18040_),
    .A1(net5797),
    .B1(_18041_),
    .X(_18042_));
 sg13g2_nor3_1 _25006_ (.A(_15480_),
    .B(_16267_),
    .C(_18013_),
    .Y(_18043_));
 sg13g2_o21ai_1 _25007_ (.B1(_15480_),
    .Y(_18044_),
    .A1(_16267_),
    .A2(_18013_));
 sg13g2_nand2_1 _25008_ (.Y(_18045_),
    .A(net4990),
    .B(_18044_));
 sg13g2_o21ai_1 _25009_ (.B1(_18042_),
    .Y(_18046_),
    .A1(_18043_),
    .A2(_18045_));
 sg13g2_o21ai_1 _25010_ (.B1(_15487_),
    .Y(_18047_),
    .A1(_15489_),
    .A2(_17870_));
 sg13g2_xnor2_1 _25011_ (.Y(_18048_),
    .A(_15486_),
    .B(_18047_));
 sg13g2_o21ai_1 _25012_ (.B1(net5079),
    .Y(_18049_),
    .A1(\u_inv.f_next[75] ),
    .A2(net5797));
 sg13g2_a21oi_1 _25013_ (.A1(net5797),
    .A2(_18048_),
    .Y(_18050_),
    .B1(_18049_));
 sg13g2_a21oi_1 _25014_ (.A1(_16270_),
    .A2(_17877_),
    .Y(_18051_),
    .B1(_15486_));
 sg13g2_nand3_1 _25015_ (.B(_16270_),
    .C(_17877_),
    .A(_15486_),
    .Y(_18052_));
 sg13g2_nor2_1 _25016_ (.A(net5076),
    .B(_18051_),
    .Y(_18053_));
 sg13g2_a21o_1 _25017_ (.A2(_18053_),
    .A1(_18052_),
    .B1(_18050_),
    .X(_18054_));
 sg13g2_a21oi_1 _25018_ (.A1(_15484_),
    .A2(_18018_),
    .Y(_18055_),
    .B1(_15506_));
 sg13g2_xnor2_1 _25019_ (.Y(_18056_),
    .A(_15478_),
    .B(_18055_));
 sg13g2_nor2_1 _25020_ (.A(\u_inv.f_next[78] ),
    .B(net5797),
    .Y(_18057_));
 sg13g2_o21ai_1 _25021_ (.B1(net5079),
    .Y(_18058_),
    .A1(net5697),
    .A2(_18056_));
 sg13g2_a21o_1 _25022_ (.A2(_18044_),
    .A1(_16266_),
    .B1(_15478_),
    .X(_18059_));
 sg13g2_nand3_1 _25023_ (.B(_16266_),
    .C(_18044_),
    .A(_15478_),
    .Y(_18060_));
 sg13g2_nand3_1 _25024_ (.B(_18059_),
    .C(_18060_),
    .A(net4990),
    .Y(_18061_));
 sg13g2_o21ai_1 _25025_ (.B1(_18061_),
    .Y(_18062_),
    .A1(_18057_),
    .A2(_18058_));
 sg13g2_a21oi_1 _25026_ (.A1(_15553_),
    .A2(_17773_),
    .Y(_18063_),
    .B1(_15539_));
 sg13g2_nand3_1 _25027_ (.B(_15553_),
    .C(_17773_),
    .A(_15539_),
    .Y(_18064_));
 sg13g2_nand2b_1 _25028_ (.Y(_18065_),
    .B(_18064_),
    .A_N(_18063_));
 sg13g2_o21ai_1 _25029_ (.B1(net5098),
    .Y(_18066_),
    .A1(\u_inv.f_next[90] ),
    .A2(net5823));
 sg13g2_a21oi_1 _25030_ (.A1(net5823),
    .A2(_18065_),
    .Y(_18067_),
    .B1(_18066_));
 sg13g2_nor3_1 _25031_ (.A(_15539_),
    .B(_16314_),
    .C(_17763_),
    .Y(_18068_));
 sg13g2_o21ai_1 _25032_ (.B1(_15539_),
    .Y(_18069_),
    .A1(_16314_),
    .A2(_17763_));
 sg13g2_nor2b_1 _25033_ (.A(_18068_),
    .B_N(_18069_),
    .Y(_18070_));
 sg13g2_a21o_2 _25034_ (.A2(_18070_),
    .A1(net5013),
    .B1(_18067_),
    .X(_18071_));
 sg13g2_a21oi_1 _25035_ (.A1(\u_inv.f_next[90] ),
    .A2(_14344_),
    .Y(_18072_),
    .B1(_15538_));
 sg13g2_nor2b_1 _25036_ (.A(_16310_),
    .B_N(_17764_),
    .Y(_18073_));
 sg13g2_a21oi_1 _25037_ (.A1(_18069_),
    .A2(_18072_),
    .Y(_18074_),
    .B1(net5098));
 sg13g2_a21oi_1 _25038_ (.A1(\u_inv.f_next[90] ),
    .A2(\u_inv.f_reg[90] ),
    .Y(_18075_),
    .B1(_18063_));
 sg13g2_xnor2_1 _25039_ (.Y(_18076_),
    .A(_15538_),
    .B(_18075_));
 sg13g2_o21ai_1 _25040_ (.B1(net5098),
    .Y(_18077_),
    .A1(\u_inv.f_next[91] ),
    .A2(net5823));
 sg13g2_a21oi_1 _25041_ (.A1(net5823),
    .A2(_18076_),
    .Y(_18078_),
    .B1(_18077_));
 sg13g2_a21o_2 _25042_ (.A2(_18074_),
    .A1(_18073_),
    .B1(_18078_),
    .X(_18079_));
 sg13g2_inv_1 _25043_ (.Y(_18080_),
    .A(_18079_));
 sg13g2_nor2b_1 _25044_ (.A(_17886_),
    .B_N(_15163_),
    .Y(_18081_));
 sg13g2_nand2b_1 _25045_ (.Y(_18082_),
    .B(_15163_),
    .A_N(_17886_));
 sg13g2_nor2_1 _25046_ (.A(_16295_),
    .B(_18081_),
    .Y(_18083_));
 sg13g2_o21ai_1 _25047_ (.B1(_15153_),
    .Y(_18084_),
    .A1(_16295_),
    .A2(_18081_));
 sg13g2_and2_1 _25048_ (.A(_16292_),
    .B(_18084_),
    .X(_18085_));
 sg13g2_a21oi_1 _25049_ (.A1(_15150_),
    .A2(_18085_),
    .Y(_18086_),
    .B1(net5089));
 sg13g2_o21ai_1 _25050_ (.B1(_18086_),
    .Y(_18087_),
    .A1(_15150_),
    .A2(_18085_));
 sg13g2_a21oi_1 _25051_ (.A1(_15166_),
    .A2(_17880_),
    .Y(_18088_),
    .B1(_15159_));
 sg13g2_or2_1 _25052_ (.X(_18089_),
    .B(_18088_),
    .A(_15153_));
 sg13g2_nand3_1 _25053_ (.B(_15152_),
    .C(_18089_),
    .A(_15150_),
    .Y(_18090_));
 sg13g2_a21oi_1 _25054_ (.A1(_15152_),
    .A2(_18089_),
    .Y(_18091_),
    .B1(_15150_));
 sg13g2_nand2_1 _25055_ (.Y(_18092_),
    .A(net5810),
    .B(_18090_));
 sg13g2_nor2_1 _25056_ (.A(\u_inv.f_next[87] ),
    .B(net5810),
    .Y(_18093_));
 sg13g2_o21ai_1 _25057_ (.B1(net5089),
    .Y(_18094_),
    .A1(_18091_),
    .A2(_18092_));
 sg13g2_o21ai_1 _25058_ (.B1(_18087_),
    .Y(_18095_),
    .A1(_18093_),
    .A2(_18094_));
 sg13g2_xor2_1 _25059_ (.B(_18083_),
    .A(_15153_),
    .X(_18096_));
 sg13g2_xor2_1 _25060_ (.B(_18088_),
    .A(_15153_),
    .X(_18097_));
 sg13g2_nand2_1 _25061_ (.Y(_18098_),
    .A(net2951),
    .B(net5707));
 sg13g2_a21oi_1 _25062_ (.A1(net5810),
    .A2(_18097_),
    .Y(_18099_),
    .B1(net5002));
 sg13g2_a22oi_1 _25063_ (.Y(_18100_),
    .B1(_18098_),
    .B2(_18099_),
    .A2(_18096_),
    .A1(net5002));
 sg13g2_o21ai_1 _25064_ (.B1(_16250_),
    .Y(_18101_),
    .A1(_16242_),
    .A2(_17848_));
 sg13g2_and2_1 _25065_ (.A(_15176_),
    .B(_18101_),
    .X(_18102_));
 sg13g2_a21oi_1 _25066_ (.A1(\u_inv.f_next[68] ),
    .A2(_14322_),
    .Y(_18103_),
    .B1(_18102_));
 sg13g2_nor2_1 _25067_ (.A(_15177_),
    .B(_18103_),
    .Y(_18104_));
 sg13g2_o21ai_1 _25068_ (.B1(_15172_),
    .Y(_18105_),
    .A1(_16252_),
    .A2(_18104_));
 sg13g2_nand3_1 _25069_ (.B(_16251_),
    .C(_18105_),
    .A(_15169_),
    .Y(_18106_));
 sg13g2_a21oi_1 _25070_ (.A1(_16251_),
    .A2(_18105_),
    .Y(_18107_),
    .B1(_15169_));
 sg13g2_nand2_1 _25071_ (.Y(_18108_),
    .A(net4989),
    .B(_18106_));
 sg13g2_o21ai_1 _25072_ (.B1(_15190_),
    .Y(_18109_),
    .A1(_15183_),
    .A2(_17854_));
 sg13g2_a21oi_1 _25073_ (.A1(_15178_),
    .A2(_18109_),
    .Y(_18110_),
    .B1(_15195_));
 sg13g2_o21ai_1 _25074_ (.B1(_15171_),
    .Y(_18111_),
    .A1(_15172_),
    .A2(_18110_));
 sg13g2_xnor2_1 _25075_ (.Y(_18112_),
    .A(_15169_),
    .B(_18111_));
 sg13g2_a21oi_1 _25076_ (.A1(net5793),
    .A2(_18112_),
    .Y(_18113_),
    .B1(net4989));
 sg13g2_o21ai_1 _25077_ (.B1(_18113_),
    .Y(_18114_),
    .A1(\u_inv.f_next[71] ),
    .A2(net5793));
 sg13g2_o21ai_1 _25078_ (.B1(_18114_),
    .Y(_18115_),
    .A1(_18107_),
    .A2(_18108_));
 sg13g2_a21oi_1 _25079_ (.A1(_16218_),
    .A2(_17939_),
    .Y(_18116_),
    .B1(_16229_));
 sg13g2_o21ai_1 _25080_ (.B1(_16232_),
    .Y(_18117_),
    .A1(_15203_),
    .A2(_18116_));
 sg13g2_and2_1 _25081_ (.A(_15205_),
    .B(_18117_),
    .X(_18118_));
 sg13g2_o21ai_1 _25082_ (.B1(_15200_),
    .Y(_18119_),
    .A1(_16231_),
    .A2(_18118_));
 sg13g2_nand2b_1 _25083_ (.Y(_18120_),
    .B(_18119_),
    .A_N(_16235_));
 sg13g2_o21ai_1 _25084_ (.B1(net4980),
    .Y(_18121_),
    .A1(_15198_),
    .A2(_18120_));
 sg13g2_a21oi_1 _25085_ (.A1(_15198_),
    .A2(_18120_),
    .Y(_18122_),
    .B1(_18121_));
 sg13g2_o21ai_1 _25086_ (.B1(_15219_),
    .Y(_18123_),
    .A1(_15212_),
    .A2(_17944_));
 sg13g2_a21oi_1 _25087_ (.A1(_15206_),
    .A2(_18123_),
    .Y(_18124_),
    .B1(_15223_));
 sg13g2_o21ai_1 _25088_ (.B1(_15199_),
    .Y(_18125_),
    .A1(_15200_),
    .A2(_18124_));
 sg13g2_xnor2_1 _25089_ (.Y(_18126_),
    .A(_15198_),
    .B(_18125_));
 sg13g2_a21oi_1 _25090_ (.A1(_14111_),
    .A2(net5689),
    .Y(_18127_),
    .B1(net4974));
 sg13g2_o21ai_1 _25091_ (.B1(_18127_),
    .Y(_18128_),
    .A1(net5689),
    .A2(_18126_));
 sg13g2_nand2b_2 _25092_ (.Y(_18129_),
    .B(_18128_),
    .A_N(_18122_));
 sg13g2_xnor2_1 _25093_ (.Y(_18130_),
    .A(_15200_),
    .B(_18124_));
 sg13g2_o21ai_1 _25094_ (.B1(net5067),
    .Y(_18131_),
    .A1(\u_inv.f_next[62] ),
    .A2(net5781));
 sg13g2_a21o_1 _25095_ (.A2(_18130_),
    .A1(net5781),
    .B1(_18131_),
    .X(_18132_));
 sg13g2_nor3_1 _25096_ (.A(_15200_),
    .B(_16231_),
    .C(_18118_),
    .Y(_18133_));
 sg13g2_nand2_1 _25097_ (.Y(_18134_),
    .A(net4974),
    .B(_18119_));
 sg13g2_o21ai_1 _25098_ (.B1(_18132_),
    .Y(_18135_),
    .A1(_18133_),
    .A2(_18134_));
 sg13g2_a21o_1 _25099_ (.A2(_18109_),
    .A1(_15175_),
    .B1(_15174_),
    .X(_18136_));
 sg13g2_xnor2_1 _25100_ (.Y(_18137_),
    .A(_15177_),
    .B(_18136_));
 sg13g2_o21ai_1 _25101_ (.B1(net5067),
    .Y(_18138_),
    .A1(\u_inv.f_next[69] ),
    .A2(net5781));
 sg13g2_a21o_1 _25102_ (.A2(_18137_),
    .A1(net5784),
    .B1(_18138_),
    .X(_18139_));
 sg13g2_a21o_1 _25103_ (.A2(_18103_),
    .A1(_15177_),
    .B1(net5067),
    .X(_18140_));
 sg13g2_o21ai_1 _25104_ (.B1(_18139_),
    .Y(_18141_),
    .A1(_18104_),
    .A2(_18140_));
 sg13g2_xnor2_1 _25105_ (.Y(_18142_),
    .A(_15176_),
    .B(_18109_));
 sg13g2_nor2_1 _25106_ (.A(\u_inv.f_next[68] ),
    .B(net5781),
    .Y(_18143_));
 sg13g2_o21ai_1 _25107_ (.B1(net5067),
    .Y(_18144_),
    .A1(net5690),
    .A2(_18142_));
 sg13g2_nor2_1 _25108_ (.A(net5068),
    .B(_18102_),
    .Y(_18145_));
 sg13g2_o21ai_1 _25109_ (.B1(_18145_),
    .Y(_18146_),
    .A1(_15176_),
    .A2(_18101_));
 sg13g2_o21ai_1 _25110_ (.B1(_18146_),
    .Y(_18147_),
    .A1(_18143_),
    .A2(_18144_));
 sg13g2_a21oi_1 _25111_ (.A1(_15203_),
    .A2(_18123_),
    .Y(_18148_),
    .B1(_15202_));
 sg13g2_xnor2_1 _25112_ (.Y(_18149_),
    .A(_15205_),
    .B(_18148_));
 sg13g2_o21ai_1 _25113_ (.B1(net5065),
    .Y(_18150_),
    .A1(\u_inv.f_next[61] ),
    .A2(net5780));
 sg13g2_a21o_1 _25114_ (.A2(_18149_),
    .A1(net5780),
    .B1(_18150_),
    .X(_18151_));
 sg13g2_o21ai_1 _25115_ (.B1(net4974),
    .Y(_18152_),
    .A1(_15205_),
    .A2(_18117_));
 sg13g2_o21ai_1 _25116_ (.B1(_18151_),
    .Y(_18153_),
    .A1(_18118_),
    .A2(_18152_));
 sg13g2_xnor2_1 _25117_ (.Y(_18154_),
    .A(_15229_),
    .B(_17933_));
 sg13g2_nor2_1 _25118_ (.A(\u_inv.f_next[38] ),
    .B(net5750),
    .Y(_18155_));
 sg13g2_o21ai_1 _25119_ (.B1(net5043),
    .Y(_18156_),
    .A1(net5674),
    .A2(_18154_));
 sg13g2_nand3_1 _25120_ (.B(_16160_),
    .C(_17924_),
    .A(_15229_),
    .Y(_18157_));
 sg13g2_nand3_1 _25121_ (.B(_17925_),
    .C(_18157_),
    .A(net4951),
    .Y(_18158_));
 sg13g2_o21ai_1 _25122_ (.B1(_18158_),
    .Y(_18159_),
    .A1(_18155_),
    .A2(_18156_));
 sg13g2_nand2b_1 _25123_ (.Y(_18160_),
    .B(_17960_),
    .A_N(_15401_));
 sg13g2_nand2_1 _25124_ (.Y(_18161_),
    .A(_15399_),
    .B(_18160_));
 sg13g2_xor2_1 _25125_ (.B(_18161_),
    .A(_15402_),
    .X(_18162_));
 sg13g2_nor2_1 _25126_ (.A(net5673),
    .B(_18162_),
    .Y(_18163_));
 sg13g2_o21ai_1 _25127_ (.B1(net5046),
    .Y(_18164_),
    .A1(\u_inv.f_next[45] ),
    .A2(net5753));
 sg13g2_nand3_1 _25128_ (.B(_16185_),
    .C(_17951_),
    .A(_15402_),
    .Y(_18165_));
 sg13g2_nor2_1 _25129_ (.A(net5046),
    .B(_17952_),
    .Y(_18166_));
 sg13g2_nand2_1 _25130_ (.Y(_18167_),
    .A(_18165_),
    .B(_18166_));
 sg13g2_o21ai_1 _25131_ (.B1(_18167_),
    .Y(_18168_),
    .A1(_18163_),
    .A2(_18164_));
 sg13g2_xnor2_1 _25132_ (.Y(_18169_),
    .A(_15407_),
    .B(_17957_));
 sg13g2_o21ai_1 _25133_ (.B1(net5046),
    .Y(_18170_),
    .A1(\u_inv.f_next[42] ),
    .A2(net5753));
 sg13g2_a21o_1 _25134_ (.A2(_18169_),
    .A1(net5756),
    .B1(_18170_),
    .X(_18171_));
 sg13g2_nor3_1 _25135_ (.A(net5620),
    .B(_16177_),
    .C(_17996_),
    .Y(_18172_));
 sg13g2_nand2_1 _25136_ (.Y(_18173_),
    .A(net4955),
    .B(_17997_));
 sg13g2_o21ai_1 _25137_ (.B1(_18171_),
    .Y(_18174_),
    .A1(_18172_),
    .A2(_18173_));
 sg13g2_a21oi_1 _25138_ (.A1(_16199_),
    .A2(_16214_),
    .Y(_18175_),
    .B1(_15461_));
 sg13g2_xnor2_1 _25139_ (.Y(_18176_),
    .A(_15462_),
    .B(_16215_));
 sg13g2_a21oi_1 _25140_ (.A1(_15459_),
    .A2(_15461_),
    .Y(_18177_),
    .B1(net5689));
 sg13g2_o21ai_1 _25141_ (.B1(_18177_),
    .Y(_18178_),
    .A1(_15459_),
    .A2(_15461_));
 sg13g2_a21oi_1 _25142_ (.A1(net2546),
    .A2(net5689),
    .Y(_18179_),
    .B1(net4974));
 sg13g2_a22oi_1 _25143_ (.Y(_18180_),
    .B1(_18178_),
    .B2(_18179_),
    .A2(_18176_),
    .A1(net4974));
 sg13g2_xnor2_1 _25144_ (.Y(_18181_),
    .A(_15436_),
    .B(_17890_));
 sg13g2_a21oi_1 _25145_ (.A1(net5768),
    .A2(_18181_),
    .Y(_18182_),
    .B1(net4964));
 sg13g2_o21ai_1 _25146_ (.B1(_18182_),
    .Y(_18183_),
    .A1(\u_inv.f_next[52] ),
    .A2(net5768));
 sg13g2_nor3_1 _25147_ (.A(_15436_),
    .B(_16209_),
    .C(_17899_),
    .Y(_18184_));
 sg13g2_nand2_1 _25148_ (.Y(_18185_),
    .A(net4964),
    .B(_17900_));
 sg13g2_o21ai_1 _25149_ (.B1(_18183_),
    .Y(_18186_),
    .A1(_18184_),
    .A2(_18185_));
 sg13g2_nand3_1 _25150_ (.B(_16222_),
    .C(_16238_),
    .A(_15467_),
    .Y(_18187_));
 sg13g2_a21oi_1 _25151_ (.A1(_17848_),
    .A2(_18187_),
    .Y(_18188_),
    .B1(net5067));
 sg13g2_a21oi_1 _25152_ (.A1(_15465_),
    .A2(_15468_),
    .Y(_18189_),
    .B1(net5690));
 sg13g2_a22oi_1 _25153_ (.Y(_18190_),
    .B1(_17973_),
    .B2(_18189_),
    .A2(net5690),
    .A1(\u_inv.f_next[64] ));
 sg13g2_a21oi_2 _25154_ (.B1(_18188_),
    .Y(_18191_),
    .A2(_18190_),
    .A1(net5067));
 sg13g2_xnor2_1 _25155_ (.Y(_18192_),
    .A(_15203_),
    .B(_18116_));
 sg13g2_a21oi_1 _25156_ (.A1(_15203_),
    .A2(_18123_),
    .Y(_18193_),
    .B1(net5689));
 sg13g2_o21ai_1 _25157_ (.B1(_18193_),
    .Y(_18194_),
    .A1(_15203_),
    .A2(_18123_));
 sg13g2_a21oi_1 _25158_ (.A1(\u_inv.f_next[60] ),
    .A2(net5689),
    .Y(_18195_),
    .B1(net4974));
 sg13g2_a22oi_1 _25159_ (.Y(_18196_),
    .B1(_18194_),
    .B2(_18195_),
    .A2(_18192_),
    .A1(net4974));
 sg13g2_nor2b_1 _25160_ (.A(_15439_),
    .B_N(_17889_),
    .Y(_18197_));
 sg13g2_xnor2_1 _25161_ (.Y(_18198_),
    .A(_15439_),
    .B(_17889_));
 sg13g2_nor2_1 _25162_ (.A(\u_inv.f_next[50] ),
    .B(net5768),
    .Y(_18199_));
 sg13g2_o21ai_1 _25163_ (.B1(net5054),
    .Y(_18200_),
    .A1(net5681),
    .A2(_18198_));
 sg13g2_nand2_1 _25164_ (.Y(_18201_),
    .A(_15439_),
    .B(_17898_));
 sg13g2_o21ai_1 _25165_ (.B1(net4964),
    .Y(_18202_),
    .A1(_15439_),
    .A2(_17898_));
 sg13g2_nand2b_1 _25166_ (.Y(_18203_),
    .B(_18201_),
    .A_N(_18202_));
 sg13g2_o21ai_1 _25167_ (.B1(_18203_),
    .Y(_18204_),
    .A1(_18199_),
    .A2(_18200_));
 sg13g2_nor3_1 _25168_ (.A(_15460_),
    .B(_16225_),
    .C(_18175_),
    .Y(_18205_));
 sg13g2_nor4_1 _25169_ (.A(net5065),
    .B(_16226_),
    .C(_17939_),
    .D(_18205_),
    .Y(_18206_));
 sg13g2_a21oi_1 _25170_ (.A1(_15459_),
    .A2(_15461_),
    .Y(_18207_),
    .B1(_15213_));
 sg13g2_xnor2_1 _25171_ (.Y(_18208_),
    .A(_15460_),
    .B(_18207_));
 sg13g2_o21ai_1 _25172_ (.B1(net5065),
    .Y(_18209_),
    .A1(\u_inv.f_next[57] ),
    .A2(net5780));
 sg13g2_a21oi_1 _25173_ (.A1(net5780),
    .A2(_18208_),
    .Y(_18210_),
    .B1(_18209_));
 sg13g2_nor2_1 _25174_ (.A(_18206_),
    .B(_18210_),
    .Y(_18211_));
 sg13g2_inv_1 _25175_ (.Y(_18212_),
    .A(_18211_));
 sg13g2_o21ai_1 _25176_ (.B1(_15231_),
    .Y(_18213_),
    .A1(_15233_),
    .A2(_17931_));
 sg13g2_xnor2_1 _25177_ (.Y(_18214_),
    .A(_15234_),
    .B(_18213_));
 sg13g2_o21ai_1 _25178_ (.B1(net5043),
    .Y(_18215_),
    .A1(\u_inv.f_next[37] ),
    .A2(net5750));
 sg13g2_a21oi_1 _25179_ (.A1(net5750),
    .A2(_18214_),
    .Y(_18216_),
    .B1(_18215_));
 sg13g2_nor3_1 _25180_ (.A(_15235_),
    .B(_16161_),
    .C(_17923_),
    .Y(_18217_));
 sg13g2_nor2_1 _25181_ (.A(net5043),
    .B(_18217_),
    .Y(_18218_));
 sg13g2_a21o_1 _25182_ (.A2(_18218_),
    .A1(_17924_),
    .B1(_18216_),
    .X(_18219_));
 sg13g2_a21oi_1 _25183_ (.A1(_16153_),
    .A2(_17921_),
    .Y(_18220_),
    .B1(_15388_));
 sg13g2_o21ai_1 _25184_ (.B1(_15241_),
    .Y(_18221_),
    .A1(_16155_),
    .A2(_18220_));
 sg13g2_a21oi_1 _25185_ (.A1(_16154_),
    .A2(_18221_),
    .Y(_18222_),
    .B1(_15238_));
 sg13g2_nand3_1 _25186_ (.B(_16154_),
    .C(_18221_),
    .A(_15238_),
    .Y(_18223_));
 sg13g2_nand2_1 _25187_ (.Y(_18224_),
    .A(net4951),
    .B(_18223_));
 sg13g2_o21ai_1 _25188_ (.B1(_15240_),
    .Y(_18225_),
    .A1(_15241_),
    .A2(_17929_));
 sg13g2_xnor2_1 _25189_ (.Y(_18226_),
    .A(_15238_),
    .B(_18225_));
 sg13g2_a21oi_1 _25190_ (.A1(net5749),
    .A2(_18226_),
    .Y(_18227_),
    .B1(net4951));
 sg13g2_o21ai_1 _25191_ (.B1(_18227_),
    .Y(_18228_),
    .A1(\u_inv.f_next[35] ),
    .A2(net5749));
 sg13g2_o21ai_1 _25192_ (.B1(_18228_),
    .Y(_18229_),
    .A1(_18222_),
    .A2(_18224_));
 sg13g2_o21ai_1 _25193_ (.B1(_15377_),
    .Y(_18230_),
    .A1(_15371_),
    .A2(_15379_));
 sg13g2_xnor2_1 _25194_ (.Y(_18231_),
    .A(_15380_),
    .B(_18230_));
 sg13g2_a21oi_1 _25195_ (.A1(net5740),
    .A2(_18231_),
    .Y(_18232_),
    .B1(net4943));
 sg13g2_o21ai_1 _25196_ (.B1(_18232_),
    .Y(_18233_),
    .A1(\u_inv.f_next[29] ),
    .A2(net5740));
 sg13g2_nand2_1 _25197_ (.Y(_18234_),
    .A(_15379_),
    .B(_16135_));
 sg13g2_and2_1 _25198_ (.A(_16142_),
    .B(_18234_),
    .X(_18235_));
 sg13g2_xnor2_1 _25199_ (.Y(_18236_),
    .A(_15380_),
    .B(_18235_));
 sg13g2_o21ai_1 _25200_ (.B1(_18233_),
    .Y(_18237_),
    .A1(net5036),
    .A2(_18236_));
 sg13g2_xnor2_1 _25201_ (.Y(_18238_),
    .A(_15371_),
    .B(_15379_));
 sg13g2_o21ai_1 _25202_ (.B1(net5036),
    .Y(_18239_),
    .A1(\u_inv.f_next[28] ),
    .A2(net5740));
 sg13g2_a21o_1 _25203_ (.A2(_18238_),
    .A1(net5740),
    .B1(_18239_),
    .X(_18240_));
 sg13g2_xnor2_1 _25204_ (.Y(_18241_),
    .A(_15379_),
    .B(_16135_));
 sg13g2_o21ai_1 _25205_ (.B1(_18240_),
    .Y(_18242_),
    .A1(net5036),
    .A2(_18241_));
 sg13g2_a21oi_1 _25206_ (.A1(_15354_),
    .A2(_15364_),
    .Y(_18243_),
    .B1(_15363_));
 sg13g2_xor2_1 _25207_ (.B(_18243_),
    .A(_15365_),
    .X(_18244_));
 sg13g2_o21ai_1 _25208_ (.B1(net5033),
    .Y(_18245_),
    .A1(\u_inv.f_next[25] ),
    .A2(net5734));
 sg13g2_a21oi_1 _25209_ (.A1(net5734),
    .A2(_18244_),
    .Y(_18246_),
    .B1(_18245_));
 sg13g2_nor2_1 _25210_ (.A(_15364_),
    .B(_16125_),
    .Y(_18247_));
 sg13g2_a21oi_1 _25211_ (.A1(\u_inv.f_next[24] ),
    .A2(_14278_),
    .Y(_18248_),
    .B1(_18247_));
 sg13g2_or2_1 _25212_ (.X(_18249_),
    .B(_18248_),
    .A(_15365_));
 sg13g2_a21oi_1 _25213_ (.A1(_15365_),
    .A2(_18248_),
    .Y(_18250_),
    .B1(net5033));
 sg13g2_a21o_1 _25214_ (.A2(_18250_),
    .A1(_18249_),
    .B1(_18246_),
    .X(_18251_));
 sg13g2_xnor2_1 _25215_ (.Y(_18252_),
    .A(_15354_),
    .B(_15364_));
 sg13g2_o21ai_1 _25216_ (.B1(net5033),
    .Y(_18253_),
    .A1(\u_inv.f_next[24] ),
    .A2(net5734));
 sg13g2_a21o_1 _25217_ (.A2(_18252_),
    .A1(net5734),
    .B1(_18253_),
    .X(_18254_));
 sg13g2_xnor2_1 _25218_ (.Y(_18255_),
    .A(_15364_),
    .B(_16125_));
 sg13g2_o21ai_1 _25219_ (.B1(_18254_),
    .Y(_18256_),
    .A1(net5033),
    .A2(_18255_));
 sg13g2_a21oi_1 _25220_ (.A1(_15334_),
    .A2(_15347_),
    .Y(_18257_),
    .B1(_15351_));
 sg13g2_xnor2_1 _25221_ (.Y(_18258_),
    .A(_15340_),
    .B(_18257_));
 sg13g2_o21ai_1 _25222_ (.B1(net5030),
    .Y(_18259_),
    .A1(\u_inv.f_next[22] ),
    .A2(net5733));
 sg13g2_a21oi_1 _25223_ (.A1(net5733),
    .A2(_18258_),
    .Y(_18260_),
    .B1(_18259_));
 sg13g2_a21oi_1 _25224_ (.A1(_15344_),
    .A2(_16114_),
    .Y(_18261_),
    .B1(_16121_));
 sg13g2_nor2_1 _25225_ (.A(_15339_),
    .B(_18261_),
    .Y(_18262_));
 sg13g2_xnor2_1 _25226_ (.Y(_18263_),
    .A(_15340_),
    .B(_18261_));
 sg13g2_a21o_1 _25227_ (.A2(_18263_),
    .A1(net4940),
    .B1(_18260_),
    .X(_18264_));
 sg13g2_xnor2_1 _25228_ (.Y(_18265_),
    .A(_15334_),
    .B(_15346_));
 sg13g2_a21oi_1 _25229_ (.A1(net5727),
    .A2(_18265_),
    .Y(_18266_),
    .B1(net4928));
 sg13g2_o21ai_1 _25230_ (.B1(_18266_),
    .Y(_18267_),
    .A1(net3392),
    .A2(net5727));
 sg13g2_nand3_1 _25231_ (.B(_16111_),
    .C(_16113_),
    .A(_15346_),
    .Y(_18268_));
 sg13g2_nand2_1 _25232_ (.Y(_18269_),
    .A(net4928),
    .B(_18268_));
 sg13g2_o21ai_1 _25233_ (.B1(_18267_),
    .Y(_18270_),
    .A1(_16114_),
    .A2(_18269_));
 sg13g2_nor2_1 _25234_ (.A(_15318_),
    .B(_15327_),
    .Y(_18271_));
 sg13g2_a21oi_1 _25235_ (.A1(\u_inv.f_next[16] ),
    .A2(\u_inv.f_reg[16] ),
    .Y(_18272_),
    .B1(_18271_));
 sg13g2_o21ai_1 _25236_ (.B1(net5727),
    .Y(_18273_),
    .A1(net5621),
    .A2(_18272_));
 sg13g2_a21oi_1 _25237_ (.A1(net5621),
    .A2(_18272_),
    .Y(_18274_),
    .B1(_18273_));
 sg13g2_o21ai_1 _25238_ (.B1(net5025),
    .Y(_18275_),
    .A1(\u_inv.f_next[17] ),
    .A2(net5727));
 sg13g2_nand3_1 _25239_ (.B(_16104_),
    .C(_16105_),
    .A(_15325_),
    .Y(_18276_));
 sg13g2_nand3_1 _25240_ (.B(_16108_),
    .C(_18276_),
    .A(net4929),
    .Y(_18277_));
 sg13g2_o21ai_1 _25241_ (.B1(_18277_),
    .Y(_18278_),
    .A1(_18274_),
    .A2(_18275_));
 sg13g2_and2_1 _25242_ (.A(_15323_),
    .B(_16109_),
    .X(_18279_));
 sg13g2_nor2_1 _25243_ (.A(net5025),
    .B(_18279_),
    .Y(_18280_));
 sg13g2_o21ai_1 _25244_ (.B1(_18280_),
    .Y(_18281_),
    .A1(_15323_),
    .A2(_16109_));
 sg13g2_nor2_1 _25245_ (.A(_15318_),
    .B(_15328_),
    .Y(_18282_));
 sg13g2_nor2_1 _25246_ (.A(_15332_),
    .B(_18282_),
    .Y(_18283_));
 sg13g2_xnor2_1 _25247_ (.Y(_18284_),
    .A(_15323_),
    .B(_18283_));
 sg13g2_nand2_1 _25248_ (.Y(_18285_),
    .A(net5727),
    .B(_18284_));
 sg13g2_o21ai_1 _25249_ (.B1(_18285_),
    .Y(_18286_),
    .A1(\u_inv.f_next[18] ),
    .A2(net5727));
 sg13g2_o21ai_1 _25250_ (.B1(_18281_),
    .Y(_18287_),
    .A1(net4929),
    .A2(_18286_));
 sg13g2_a21oi_1 _25251_ (.A1(_15326_),
    .A2(_16103_),
    .Y(_18288_),
    .B1(net5025));
 sg13g2_xnor2_1 _25252_ (.Y(_18289_),
    .A(_15318_),
    .B(_15327_));
 sg13g2_o21ai_1 _25253_ (.B1(net5026),
    .Y(_18290_),
    .A1(\u_inv.f_next[16] ),
    .A2(net5728));
 sg13g2_a21oi_1 _25254_ (.A1(net5728),
    .A2(_18289_),
    .Y(_18291_),
    .B1(_18290_));
 sg13g2_a21o_1 _25255_ (.A2(_18288_),
    .A1(_16104_),
    .B1(_18291_),
    .X(_18292_));
 sg13g2_xnor2_1 _25256_ (.Y(_18293_),
    .A(_15313_),
    .B(_15315_));
 sg13g2_o21ai_1 _25257_ (.B1(net5026),
    .Y(_18294_),
    .A1(\u_inv.f_next[15] ),
    .A2(net5728));
 sg13g2_a21o_1 _25258_ (.A2(_18293_),
    .A1(net5728),
    .B1(_18294_),
    .X(_18295_));
 sg13g2_nor3_1 _25259_ (.A(_15315_),
    .B(_16097_),
    .C(_16098_),
    .Y(_18296_));
 sg13g2_nand2_1 _25260_ (.Y(_18297_),
    .A(net4929),
    .B(_16101_));
 sg13g2_or2_1 _25261_ (.X(_18298_),
    .B(_18297_),
    .A(_16100_));
 sg13g2_o21ai_1 _25262_ (.B1(_18295_),
    .Y(_18299_),
    .A1(_18296_),
    .A2(_18298_));
 sg13g2_a21oi_1 _25263_ (.A1(_15310_),
    .A2(_16096_),
    .Y(_18300_),
    .B1(net5026));
 sg13g2_nand2b_1 _25264_ (.Y(_18301_),
    .B(_18300_),
    .A_N(_16097_));
 sg13g2_nor3_1 _25265_ (.A(_15305_),
    .B(_15308_),
    .C(_15310_),
    .Y(_18302_));
 sg13g2_o21ai_1 _25266_ (.B1(net5728),
    .Y(_18303_),
    .A1(_15312_),
    .A2(_18302_));
 sg13g2_o21ai_1 _25267_ (.B1(_18303_),
    .Y(_18304_),
    .A1(\u_inv.f_next[14] ),
    .A2(net5728));
 sg13g2_o21ai_1 _25268_ (.B1(_18301_),
    .Y(_18305_),
    .A1(net4929),
    .A2(_18304_));
 sg13g2_nand3_1 _25269_ (.B(_16089_),
    .C(_16090_),
    .A(_15302_),
    .Y(_18306_));
 sg13g2_nor2_1 _25270_ (.A(net5024),
    .B(_16091_),
    .Y(_18307_));
 sg13g2_xnor2_1 _25271_ (.Y(_18308_),
    .A(_15301_),
    .B(_15302_));
 sg13g2_nor2_1 _25272_ (.A(\u_inv.f_next[12] ),
    .B(net5724),
    .Y(_18309_));
 sg13g2_a21oi_1 _25273_ (.A1(net5726),
    .A2(_18308_),
    .Y(_18310_),
    .B1(_18309_));
 sg13g2_a22oi_1 _25274_ (.Y(_18311_),
    .B1(_18310_),
    .B2(net5023),
    .A2(_18307_),
    .A1(_18306_));
 sg13g2_xor2_1 _25275_ (.B(_16067_),
    .A(_15299_),
    .X(_18312_));
 sg13g2_o21ai_1 _25276_ (.B1(net5024),
    .Y(_18313_),
    .A1(\u_inv.f_next[11] ),
    .A2(net5724));
 sg13g2_a21oi_1 _25277_ (.A1(net5724),
    .A2(_18312_),
    .Y(_18314_),
    .B1(_18313_));
 sg13g2_nand3_1 _25278_ (.B(_16068_),
    .C(_16088_),
    .A(_16067_),
    .Y(_18315_));
 sg13g2_nand3_1 _25279_ (.B(_16089_),
    .C(_18315_),
    .A(net4927),
    .Y(_18316_));
 sg13g2_nand2b_1 _25280_ (.Y(_18317_),
    .B(_18316_),
    .A_N(_18314_));
 sg13g2_nand3_1 _25281_ (.B(_16069_),
    .C(_16087_),
    .A(_15262_),
    .Y(_18318_));
 sg13g2_nand3_1 _25282_ (.B(_16088_),
    .C(_18318_),
    .A(net4927),
    .Y(_18319_));
 sg13g2_o21ai_1 _25283_ (.B1(_15263_),
    .Y(_18320_),
    .A1(_15264_),
    .A2(_15297_));
 sg13g2_nor2b_1 _25284_ (.A(_15298_),
    .B_N(_18320_),
    .Y(_18321_));
 sg13g2_nor2_1 _25285_ (.A(net5656),
    .B(_18321_),
    .Y(_18322_));
 sg13g2_o21ai_1 _25286_ (.B1(net5023),
    .Y(_18323_),
    .A1(net3207),
    .A2(net5724));
 sg13g2_o21ai_1 _25287_ (.B1(_18319_),
    .Y(_18324_),
    .A1(_18322_),
    .A2(_18323_));
 sg13g2_nand3_1 _25288_ (.B(_16072_),
    .C(_16085_),
    .A(_15266_),
    .Y(_18325_));
 sg13g2_nor2b_1 _25289_ (.A(_16086_),
    .B_N(_18325_),
    .Y(_18326_));
 sg13g2_xnor2_1 _25290_ (.Y(_18327_),
    .A(_15266_),
    .B(_15295_));
 sg13g2_a21oi_1 _25291_ (.A1(\u_inv.f_next[8] ),
    .A2(net5656),
    .Y(_18328_),
    .B1(net4927));
 sg13g2_o21ai_1 _25292_ (.B1(_18328_),
    .Y(_18329_),
    .A1(net5656),
    .A2(_18327_));
 sg13g2_o21ai_1 _25293_ (.B1(_18329_),
    .Y(_18330_),
    .A1(net5023),
    .A2(_18326_));
 sg13g2_nor3_1 _25294_ (.A(_15268_),
    .B(_16073_),
    .C(_16084_),
    .Y(_18331_));
 sg13g2_nor2_1 _25295_ (.A(net5023),
    .B(_18331_),
    .Y(_18332_));
 sg13g2_xnor2_1 _25296_ (.Y(_18333_),
    .A(_15268_),
    .B(_15294_));
 sg13g2_o21ai_1 _25297_ (.B1(net5023),
    .Y(_18334_),
    .A1(\u_inv.f_next[7] ),
    .A2(net5724));
 sg13g2_a21oi_1 _25298_ (.A1(net5724),
    .A2(_18333_),
    .Y(_18335_),
    .B1(_18334_));
 sg13g2_a21o_1 _25299_ (.A2(_18332_),
    .A1(_16085_),
    .B1(_18335_),
    .X(_18336_));
 sg13g2_inv_1 _25300_ (.Y(_18337_),
    .A(_18336_));
 sg13g2_or3_1 _25301_ (.A(_15272_),
    .B(_16075_),
    .C(_16082_),
    .X(_18338_));
 sg13g2_nand2_1 _25302_ (.Y(_18339_),
    .A(_16083_),
    .B(_18338_));
 sg13g2_nand2_1 _25303_ (.Y(_18340_),
    .A(_15272_),
    .B(_15290_));
 sg13g2_nand3_1 _25304_ (.B(_15291_),
    .C(_18340_),
    .A(net5725),
    .Y(_18341_));
 sg13g2_a21oi_1 _25305_ (.A1(net3352),
    .A2(net5656),
    .Y(_18342_),
    .B1(net4927));
 sg13g2_a22oi_1 _25306_ (.Y(_18343_),
    .B1(_18341_),
    .B2(_18342_),
    .A2(_18339_),
    .A1(net4927));
 sg13g2_nand3_1 _25307_ (.B(_16076_),
    .C(_16081_),
    .A(_15275_),
    .Y(_18344_));
 sg13g2_nand2b_1 _25308_ (.Y(_18345_),
    .B(_18344_),
    .A_N(_16082_));
 sg13g2_a21oi_1 _25309_ (.A1(_15275_),
    .A2(_15289_),
    .Y(_18346_),
    .B1(net5656));
 sg13g2_o21ai_1 _25310_ (.B1(_18346_),
    .Y(_18347_),
    .A1(_15275_),
    .A2(_15289_));
 sg13g2_a21oi_1 _25311_ (.A1(\u_inv.f_next[4] ),
    .A2(net5656),
    .Y(_18348_),
    .B1(net4927));
 sg13g2_a22oi_1 _25312_ (.Y(_18349_),
    .B1(_18347_),
    .B2(_18348_),
    .A2(_18345_),
    .A1(net4928));
 sg13g2_nand2_1 _25313_ (.Y(_18350_),
    .A(\u_inv.f_reg[0] ),
    .B(net4928));
 sg13g2_xnor2_1 _25314_ (.Y(_18351_),
    .A(_15285_),
    .B(_15286_));
 sg13g2_nand2_1 _25315_ (.Y(_18352_),
    .A(net5725),
    .B(_18351_));
 sg13g2_o21ai_1 _25316_ (.B1(_18352_),
    .Y(_18353_),
    .A1(\u_inv.f_next[1] ),
    .A2(net5726));
 sg13g2_xnor2_1 _25317_ (.Y(_18354_),
    .A(_18350_),
    .B(_18353_));
 sg13g2_xnor2_1 _25318_ (.Y(_18355_),
    .A(_15281_),
    .B(_15287_));
 sg13g2_nand2_1 _25319_ (.Y(_18356_),
    .A(net5725),
    .B(_18355_));
 sg13g2_o21ai_1 _25320_ (.B1(_18356_),
    .Y(_18357_),
    .A1(\u_inv.f_next[2] ),
    .A2(net5725));
 sg13g2_xnor2_1 _25321_ (.Y(_18358_),
    .A(_15281_),
    .B(_16079_));
 sg13g2_nand2_1 _25322_ (.Y(_18359_),
    .A(net5024),
    .B(_18357_));
 sg13g2_o21ai_1 _25323_ (.B1(_18359_),
    .Y(_18360_),
    .A1(net5024),
    .A2(_18358_));
 sg13g2_or3_1 _25324_ (.A(_15277_),
    .B(_16077_),
    .C(_16080_),
    .X(_18361_));
 sg13g2_nand2_1 _25325_ (.Y(_18362_),
    .A(_16081_),
    .B(_18361_));
 sg13g2_xor2_1 _25326_ (.B(_15288_),
    .A(_15277_),
    .X(_18363_));
 sg13g2_o21ai_1 _25327_ (.B1(net5024),
    .Y(_18364_),
    .A1(_14168_),
    .A2(net5725));
 sg13g2_a21oi_1 _25328_ (.A1(net5725),
    .A2(_18363_),
    .Y(_18365_),
    .B1(_18364_));
 sg13g2_a21o_1 _25329_ (.A2(_18362_),
    .A1(net4928),
    .B1(_18365_),
    .X(_18366_));
 sg13g2_inv_1 _25330_ (.Y(_18367_),
    .A(_18366_));
 sg13g2_nand3_1 _25331_ (.B(_18360_),
    .C(_18366_),
    .A(_18354_),
    .Y(_18368_));
 sg13g2_nor3_1 _25332_ (.A(_18343_),
    .B(_18349_),
    .C(_18368_),
    .Y(_18369_));
 sg13g2_and3_1 _25333_ (.X(_18370_),
    .A(_15270_),
    .B(_16074_),
    .C(_16083_));
 sg13g2_nor2_1 _25334_ (.A(_15270_),
    .B(_15292_),
    .Y(_18371_));
 sg13g2_nor3_1 _25335_ (.A(net5656),
    .B(_15293_),
    .C(_18371_),
    .Y(_18372_));
 sg13g2_a21o_1 _25336_ (.A2(net5656),
    .A1(\u_inv.f_next[6] ),
    .B1(_18372_),
    .X(_18373_));
 sg13g2_nor3_1 _25337_ (.A(net5023),
    .B(_16084_),
    .C(_18370_),
    .Y(_18374_));
 sg13g2_a21oi_1 _25338_ (.A1(net5023),
    .A2(_18373_),
    .Y(_18375_),
    .B1(_18374_));
 sg13g2_nand4_1 _25339_ (.B(_18337_),
    .C(_18369_),
    .A(_18330_),
    .Y(_18376_),
    .D(_18375_));
 sg13g2_xor2_1 _25340_ (.B(_16070_),
    .A(_15296_),
    .X(_18377_));
 sg13g2_o21ai_1 _25341_ (.B1(net5023),
    .Y(_18378_),
    .A1(\u_inv.f_next[9] ),
    .A2(net5724));
 sg13g2_a21o_1 _25342_ (.A2(_18377_),
    .A1(net5724),
    .B1(_18378_),
    .X(_18379_));
 sg13g2_nor3_1 _25343_ (.A(_16070_),
    .B(_16071_),
    .C(_16086_),
    .Y(_18380_));
 sg13g2_nand2_1 _25344_ (.Y(_18381_),
    .A(net4927),
    .B(_16087_));
 sg13g2_o21ai_1 _25345_ (.B1(_18379_),
    .Y(_18382_),
    .A1(_18380_),
    .A2(_18381_));
 sg13g2_nor4_1 _25346_ (.A(_18317_),
    .B(_18324_),
    .C(_18376_),
    .D(_18382_),
    .Y(_18383_));
 sg13g2_xnor2_1 _25347_ (.Y(_18384_),
    .A(_15304_),
    .B(_15306_));
 sg13g2_o21ai_1 _25348_ (.B1(net5025),
    .Y(_18385_),
    .A1(\u_inv.f_next[13] ),
    .A2(net5729));
 sg13g2_a21oi_1 _25349_ (.A1(net5729),
    .A2(_18384_),
    .Y(_18386_),
    .B1(_18385_));
 sg13g2_o21ai_1 _25350_ (.B1(net4927),
    .Y(_18387_),
    .A1(_15306_),
    .A2(_16093_));
 sg13g2_a21oi_1 _25351_ (.A1(_15306_),
    .A2(_16093_),
    .Y(_18388_),
    .B1(_18387_));
 sg13g2_nor2_1 _25352_ (.A(_18386_),
    .B(_18388_),
    .Y(_18389_));
 sg13g2_inv_1 _25353_ (.Y(_18390_),
    .A(_18389_));
 sg13g2_nand3_1 _25354_ (.B(_18383_),
    .C(_18389_),
    .A(_18311_),
    .Y(_18391_));
 sg13g2_or4_1 _25355_ (.A(_18292_),
    .B(_18299_),
    .C(_18305_),
    .D(_18391_),
    .X(_18392_));
 sg13g2_nor4_1 _25356_ (.A(_18270_),
    .B(_18278_),
    .C(_18287_),
    .D(_18392_),
    .Y(_18393_));
 sg13g2_a21oi_1 _25357_ (.A1(_15334_),
    .A2(_15346_),
    .Y(_18394_),
    .B1(_15345_));
 sg13g2_xnor2_1 _25358_ (.Y(_18395_),
    .A(_15344_),
    .B(_18394_));
 sg13g2_o21ai_1 _25359_ (.B1(net5020),
    .Y(_18396_),
    .A1(\u_inv.f_next[21] ),
    .A2(net5722));
 sg13g2_a21oi_1 _25360_ (.A1(net5722),
    .A2(_18395_),
    .Y(_18397_),
    .B1(_18396_));
 sg13g2_nor3_1 _25361_ (.A(_15344_),
    .B(_16114_),
    .C(_16119_),
    .Y(_18398_));
 sg13g2_nand3_1 _25362_ (.B(_16115_),
    .C(_16120_),
    .A(net4928),
    .Y(_18399_));
 sg13g2_nor2_1 _25363_ (.A(_18398_),
    .B(_18399_),
    .Y(_18400_));
 sg13g2_nor2_1 _25364_ (.A(_18397_),
    .B(_18400_),
    .Y(_18401_));
 sg13g2_o21ai_1 _25365_ (.B1(_15321_),
    .Y(_18402_),
    .A1(_15323_),
    .A2(_18283_));
 sg13g2_xnor2_1 _25366_ (.Y(_18403_),
    .A(_15319_),
    .B(_18402_));
 sg13g2_o21ai_1 _25367_ (.B1(net5025),
    .Y(_18404_),
    .A1(\u_inv.f_next[19] ),
    .A2(net5727));
 sg13g2_a21oi_1 _25368_ (.A1(net5727),
    .A2(_18403_),
    .Y(_18405_),
    .B1(_18404_));
 sg13g2_nor3_1 _25369_ (.A(_15320_),
    .B(_16065_),
    .C(_18279_),
    .Y(_18406_));
 sg13g2_o21ai_1 _25370_ (.B1(_15320_),
    .Y(_18407_),
    .A1(_16065_),
    .A2(_18279_));
 sg13g2_nor2_1 _25371_ (.A(net5025),
    .B(_18406_),
    .Y(_18408_));
 sg13g2_a21o_1 _25372_ (.A2(_18408_),
    .A1(_18407_),
    .B1(_18405_),
    .X(_18409_));
 sg13g2_nand2_1 _25373_ (.Y(_18410_),
    .A(_18393_),
    .B(_18401_));
 sg13g2_or4_1 _25374_ (.A(_18256_),
    .B(_18264_),
    .C(_18409_),
    .D(_18410_),
    .X(_18411_));
 sg13g2_nor2_1 _25375_ (.A(_16118_),
    .B(_18262_),
    .Y(_18412_));
 sg13g2_nor2_1 _25376_ (.A(_15337_),
    .B(_18412_),
    .Y(_18413_));
 sg13g2_nand2_1 _25377_ (.Y(_18414_),
    .A(_15337_),
    .B(_18412_));
 sg13g2_nor2_1 _25378_ (.A(net5033),
    .B(_18413_),
    .Y(_18415_));
 sg13g2_o21ai_1 _25379_ (.B1(_15338_),
    .Y(_18416_),
    .A1(_15340_),
    .A2(_18257_));
 sg13g2_xnor2_1 _25380_ (.Y(_18417_),
    .A(_15337_),
    .B(_18416_));
 sg13g2_nand2_1 _25381_ (.Y(_18418_),
    .A(_14151_),
    .B(net5664));
 sg13g2_a21oi_1 _25382_ (.A1(net5734),
    .A2(_18417_),
    .Y(_18419_),
    .B1(net4940));
 sg13g2_a22oi_1 _25383_ (.Y(_18420_),
    .B1(_18418_),
    .B2(_18419_),
    .A2(_18415_),
    .A1(_18414_));
 sg13g2_a21oi_1 _25384_ (.A1(_15354_),
    .A2(_15366_),
    .Y(_18421_),
    .B1(_15370_));
 sg13g2_xnor2_1 _25385_ (.Y(_18422_),
    .A(_15360_),
    .B(_18421_));
 sg13g2_nor2_1 _25386_ (.A(\u_inv.f_next[26] ),
    .B(net5734),
    .Y(_18423_));
 sg13g2_a21oi_1 _25387_ (.A1(net5734),
    .A2(_18422_),
    .Y(_18424_),
    .B1(_18423_));
 sg13g2_nand2_1 _25388_ (.Y(_18425_),
    .A(_16129_),
    .B(_18249_));
 sg13g2_nand3_1 _25389_ (.B(_16129_),
    .C(_18249_),
    .A(_15359_),
    .Y(_18426_));
 sg13g2_a21oi_1 _25390_ (.A1(_15360_),
    .A2(_18425_),
    .Y(_18427_),
    .B1(net5033));
 sg13g2_a22oi_1 _25391_ (.Y(_18428_),
    .B1(_18426_),
    .B2(_18427_),
    .A2(_18424_),
    .A1(net5033));
 sg13g2_nand3_1 _25392_ (.B(_16138_),
    .C(_16147_),
    .A(_15390_),
    .Y(_18429_));
 sg13g2_a21oi_1 _25393_ (.A1(_17921_),
    .A2(_18429_),
    .Y(_18430_),
    .B1(net5036));
 sg13g2_a21oi_1 _25394_ (.A1(_15387_),
    .A2(_15390_),
    .Y(_18431_),
    .B1(net5666));
 sg13g2_o21ai_1 _25395_ (.B1(_18431_),
    .Y(_18432_),
    .A1(_15387_),
    .A2(_15390_));
 sg13g2_a21oi_1 _25396_ (.A1(net3320),
    .A2(net5666),
    .Y(_18433_),
    .B1(net4943));
 sg13g2_a21oi_2 _25397_ (.B1(_18430_),
    .Y(_18434_),
    .A2(_18433_),
    .A1(_18432_));
 sg13g2_nor3_1 _25398_ (.A(_18242_),
    .B(_18251_),
    .C(_18411_),
    .Y(_18435_));
 sg13g2_nor2_1 _25399_ (.A(_18237_),
    .B(_18434_),
    .Y(_18436_));
 sg13g2_and4_1 _25400_ (.A(_18420_),
    .B(_18428_),
    .C(_18435_),
    .D(_18436_),
    .X(_18437_));
 sg13g2_o21ai_1 _25401_ (.B1(_15358_),
    .Y(_18438_),
    .A1(_15360_),
    .A2(_18421_));
 sg13g2_xnor2_1 _25402_ (.Y(_18439_),
    .A(_15357_),
    .B(_18438_));
 sg13g2_nand2_1 _25403_ (.Y(_18440_),
    .A(net5734),
    .B(_18439_));
 sg13g2_o21ai_1 _25404_ (.B1(_18440_),
    .Y(_18441_),
    .A1(\u_inv.f_next[27] ),
    .A2(net5737));
 sg13g2_a21oi_1 _25405_ (.A1(_15360_),
    .A2(_18425_),
    .Y(_18442_),
    .B1(_16128_));
 sg13g2_a21oi_1 _25406_ (.A1(_15357_),
    .A2(_18442_),
    .Y(_18443_),
    .B1(net5033));
 sg13g2_o21ai_1 _25407_ (.B1(_18443_),
    .Y(_18444_),
    .A1(_15357_),
    .A2(_18442_));
 sg13g2_o21ai_1 _25408_ (.B1(_18444_),
    .Y(_18445_),
    .A1(net4940),
    .A2(_18441_));
 sg13g2_xnor2_1 _25409_ (.Y(_18446_),
    .A(_15393_),
    .B(_15410_));
 sg13g2_a21oi_1 _25410_ (.A1(net5753),
    .A2(_18446_),
    .Y(_18447_),
    .B1(net4955));
 sg13g2_o21ai_1 _25411_ (.B1(_18447_),
    .Y(_18448_),
    .A1(\u_inv.f_next[40] ),
    .A2(net5753));
 sg13g2_nor2_1 _25412_ (.A(_15410_),
    .B(_16167_),
    .Y(_18449_));
 sg13g2_nand2_1 _25413_ (.Y(_18450_),
    .A(net4955),
    .B(_17995_));
 sg13g2_o21ai_1 _25414_ (.B1(_18448_),
    .Y(_18451_),
    .A1(_18449_),
    .A2(_18450_));
 sg13g2_a21oi_1 _25415_ (.A1(_15387_),
    .A2(_15390_),
    .Y(_18452_),
    .B1(_15243_));
 sg13g2_xnor2_1 _25416_ (.Y(_18453_),
    .A(_15389_),
    .B(_18452_));
 sg13g2_o21ai_1 _25417_ (.B1(net5043),
    .Y(_18454_),
    .A1(\u_inv.f_next[33] ),
    .A2(net5749));
 sg13g2_a21oi_1 _25418_ (.A1(net5749),
    .A2(_18453_),
    .Y(_18455_),
    .B1(_18454_));
 sg13g2_and3_1 _25419_ (.X(_18456_),
    .A(_15388_),
    .B(_16153_),
    .C(_17921_));
 sg13g2_nor3_1 _25420_ (.A(net5043),
    .B(_18220_),
    .C(_18456_),
    .Y(_18457_));
 sg13g2_nor2_1 _25421_ (.A(_18455_),
    .B(_18457_),
    .Y(_18458_));
 sg13g2_or2_1 _25422_ (.X(_18459_),
    .B(_18457_),
    .A(_18455_));
 sg13g2_nor2b_1 _25423_ (.A(_15371_),
    .B_N(_15381_),
    .Y(_18460_));
 sg13g2_nor2_1 _25424_ (.A(_15385_),
    .B(_18460_),
    .Y(_18461_));
 sg13g2_xnor2_1 _25425_ (.Y(_18462_),
    .A(_15375_),
    .B(_18461_));
 sg13g2_o21ai_1 _25426_ (.B1(net5036),
    .Y(_18463_),
    .A1(\u_inv.f_next[30] ),
    .A2(net5740));
 sg13g2_a21oi_1 _25427_ (.A1(net5740),
    .A2(_18462_),
    .Y(_18464_),
    .B1(_18463_));
 sg13g2_o21ai_1 _25428_ (.B1(_16141_),
    .Y(_18465_),
    .A1(_15380_),
    .A2(_18235_));
 sg13g2_nand2_1 _25429_ (.Y(_18466_),
    .A(_15375_),
    .B(_18465_));
 sg13g2_xnor2_1 _25430_ (.Y(_18467_),
    .A(_15374_),
    .B(_18465_));
 sg13g2_a21oi_2 _25431_ (.B1(_18464_),
    .Y(_18468_),
    .A2(_18467_),
    .A1(net4943));
 sg13g2_xnor2_1 _25432_ (.Y(_18469_),
    .A(_15426_),
    .B(_15444_));
 sg13g2_nor2_1 _25433_ (.A(\u_inv.f_next[48] ),
    .B(net5765),
    .Y(_18470_));
 sg13g2_a21oi_1 _25434_ (.A1(net5765),
    .A2(_18469_),
    .Y(_18471_),
    .B1(_18470_));
 sg13g2_or3_1 _25435_ (.A(_15444_),
    .B(_16175_),
    .C(_16191_),
    .X(_18472_));
 sg13g2_and2_1 _25436_ (.A(net4961),
    .B(_17896_),
    .X(_18473_));
 sg13g2_a22oi_1 _25437_ (.Y(_18474_),
    .B1(_18472_),
    .B2(_18473_),
    .A2(_18471_),
    .A1(net5054));
 sg13g2_inv_1 _25438_ (.Y(_18475_),
    .A(_18474_));
 sg13g2_nand3b_1 _25439_ (.B(_16200_),
    .C(_17896_),
    .Y(_18476_),
    .A_N(_15442_));
 sg13g2_nand4_1 _25440_ (.B(_16201_),
    .C(_17897_),
    .A(net4961),
    .Y(_18477_),
    .D(_18476_));
 sg13g2_o21ai_1 _25441_ (.B1(_15443_),
    .Y(_18478_),
    .A1(_15426_),
    .A2(_15444_));
 sg13g2_o21ai_1 _25442_ (.B1(net5765),
    .Y(_18479_),
    .A1(_15442_),
    .A2(_18478_));
 sg13g2_a21oi_1 _25443_ (.A1(_15442_),
    .A2(_18478_),
    .Y(_18480_),
    .B1(_18479_));
 sg13g2_o21ai_1 _25444_ (.B1(net5054),
    .Y(_18481_),
    .A1(\u_inv.f_next[49] ),
    .A2(net5765));
 sg13g2_o21ai_1 _25445_ (.B1(_18477_),
    .Y(_18482_),
    .A1(_18480_),
    .A2(_18481_));
 sg13g2_o21ai_1 _25446_ (.B1(_15409_),
    .Y(_18483_),
    .A1(_15393_),
    .A2(_15410_));
 sg13g2_xnor2_1 _25447_ (.Y(_18484_),
    .A(_15411_),
    .B(_18483_));
 sg13g2_o21ai_1 _25448_ (.B1(net5046),
    .Y(_18485_),
    .A1(\u_inv.f_next[41] ),
    .A2(net5753));
 sg13g2_a21oi_1 _25449_ (.A1(net5753),
    .A2(_18484_),
    .Y(_18486_),
    .B1(_18485_));
 sg13g2_nand3_1 _25450_ (.B(_16178_),
    .C(_17995_),
    .A(_15411_),
    .Y(_18487_));
 sg13g2_nor2_1 _25451_ (.A(net5046),
    .B(_17996_),
    .Y(_18488_));
 sg13g2_a21o_2 _25452_ (.A2(_18488_),
    .A1(_18487_),
    .B1(_18486_),
    .X(_18489_));
 sg13g2_o21ai_1 _25453_ (.B1(_15373_),
    .Y(_18490_),
    .A1(_15375_),
    .A2(_18461_));
 sg13g2_xnor2_1 _25454_ (.Y(_18491_),
    .A(_15372_),
    .B(_18490_));
 sg13g2_o21ai_1 _25455_ (.B1(net5036),
    .Y(_18492_),
    .A1(\u_inv.f_next[31] ),
    .A2(net5740));
 sg13g2_a21oi_1 _25456_ (.A1(net5740),
    .A2(_18491_),
    .Y(_18493_),
    .B1(_18492_));
 sg13g2_a21oi_1 _25457_ (.A1(_16140_),
    .A2(_18466_),
    .Y(_18494_),
    .B1(_15372_));
 sg13g2_nand3_1 _25458_ (.B(_16140_),
    .C(_18466_),
    .A(_15372_),
    .Y(_18495_));
 sg13g2_nor2_1 _25459_ (.A(net5036),
    .B(_18494_),
    .Y(_18496_));
 sg13g2_a21o_2 _25460_ (.A2(_18496_),
    .A1(_18495_),
    .B1(_18493_),
    .X(_18497_));
 sg13g2_o21ai_1 _25461_ (.B1(_18201_),
    .Y(_18498_),
    .A1(_14124_),
    .A2(\u_inv.f_reg[50] ));
 sg13g2_a21oi_1 _25462_ (.A1(_15440_),
    .A2(_18498_),
    .Y(_18499_),
    .B1(net5057));
 sg13g2_o21ai_1 _25463_ (.B1(_18499_),
    .Y(_18500_),
    .A1(_15440_),
    .A2(_18498_));
 sg13g2_nor2_1 _25464_ (.A(_15438_),
    .B(_18197_),
    .Y(_18501_));
 sg13g2_xor2_1 _25465_ (.B(_18501_),
    .A(_15440_),
    .X(_18502_));
 sg13g2_nand2_1 _25466_ (.Y(_18503_),
    .A(_14123_),
    .B(net5680));
 sg13g2_o21ai_1 _25467_ (.B1(_18503_),
    .Y(_18504_),
    .A1(net5680),
    .A2(_18502_));
 sg13g2_o21ai_1 _25468_ (.B1(_18500_),
    .Y(_18505_),
    .A1(net4964),
    .A2(_18504_));
 sg13g2_xor2_1 _25469_ (.B(_17950_),
    .A(_15401_),
    .X(_18506_));
 sg13g2_a21oi_1 _25470_ (.A1(_15401_),
    .A2(_17959_),
    .Y(_18507_),
    .B1(net5673));
 sg13g2_nand2_1 _25471_ (.Y(_18508_),
    .A(_18160_),
    .B(_18507_));
 sg13g2_a21oi_1 _25472_ (.A1(net2960),
    .A2(net5673),
    .Y(_18509_),
    .B1(net4955));
 sg13g2_a22oi_1 _25473_ (.Y(_18510_),
    .B1(_18508_),
    .B2(_18509_),
    .A2(_18506_),
    .A1(net4955));
 sg13g2_xnor2_1 _25474_ (.Y(_18511_),
    .A(_15241_),
    .B(_17929_));
 sg13g2_o21ai_1 _25475_ (.B1(net5043),
    .Y(_18512_),
    .A1(\u_inv.f_next[34] ),
    .A2(net5749));
 sg13g2_a21o_1 _25476_ (.A2(_18511_),
    .A1(net5749),
    .B1(_18512_),
    .X(_18513_));
 sg13g2_nor3_1 _25477_ (.A(_15241_),
    .B(_16155_),
    .C(_18220_),
    .Y(_18514_));
 sg13g2_nand2_1 _25478_ (.Y(_18515_),
    .A(net4951),
    .B(_18221_));
 sg13g2_o21ai_1 _25479_ (.B1(_18513_),
    .Y(_18516_),
    .A1(_18514_),
    .A2(_18515_));
 sg13g2_xnor2_1 _25480_ (.Y(_18517_),
    .A(_15233_),
    .B(_17931_));
 sg13g2_o21ai_1 _25481_ (.B1(net5043),
    .Y(_18518_),
    .A1(\u_inv.f_next[36] ),
    .A2(net5749));
 sg13g2_a21oi_1 _25482_ (.A1(net5750),
    .A2(_18517_),
    .Y(_18519_),
    .B1(_18518_));
 sg13g2_nand3_1 _25483_ (.B(_16158_),
    .C(_17922_),
    .A(_15232_),
    .Y(_18520_));
 sg13g2_nor2_1 _25484_ (.A(net5043),
    .B(_17923_),
    .Y(_18521_));
 sg13g2_a21o_1 _25485_ (.A2(_18521_),
    .A1(_18520_),
    .B1(_18519_),
    .X(_18522_));
 sg13g2_xnor2_1 _25486_ (.Y(_18523_),
    .A(_15172_),
    .B(_18110_));
 sg13g2_a21oi_1 _25487_ (.A1(net5793),
    .A2(_18523_),
    .Y(_18524_),
    .B1(net4979));
 sg13g2_o21ai_1 _25488_ (.B1(_18524_),
    .Y(_18525_),
    .A1(\u_inv.f_next[70] ),
    .A2(net5793));
 sg13g2_nor3_1 _25489_ (.A(_15172_),
    .B(_16252_),
    .C(_18104_),
    .Y(_18526_));
 sg13g2_nand2_1 _25490_ (.Y(_18527_),
    .A(net4979),
    .B(_18105_));
 sg13g2_o21ai_1 _25491_ (.B1(_18525_),
    .Y(_18528_),
    .A1(_18526_),
    .A2(_18527_));
 sg13g2_nand4_1 _25492_ (.B(_15157_),
    .C(_16293_),
    .A(_15156_),
    .Y(_18529_),
    .D(_17886_));
 sg13g2_nand4_1 _25493_ (.B(_16294_),
    .C(_18082_),
    .A(net5002),
    .Y(_18530_),
    .D(_18529_));
 sg13g2_nand2_1 _25494_ (.Y(_18531_),
    .A(_15158_),
    .B(_17881_));
 sg13g2_xor2_1 _25495_ (.B(_18531_),
    .A(_15163_),
    .X(_18532_));
 sg13g2_a21oi_1 _25496_ (.A1(net5810),
    .A2(_18532_),
    .Y(_18533_),
    .B1(net5002));
 sg13g2_o21ai_1 _25497_ (.B1(_18533_),
    .Y(_18534_),
    .A1(\u_inv.f_next[85] ),
    .A2(net5810));
 sg13g2_nand2_2 _25498_ (.Y(_18535_),
    .A(_18530_),
    .B(_18534_));
 sg13g2_xnor2_1 _25499_ (.Y(_18536_),
    .A(_15570_),
    .B(_15591_));
 sg13g2_o21ai_1 _25500_ (.B1(net5097),
    .Y(_18537_),
    .A1(\u_inv.f_next[104] ),
    .A2(net5818));
 sg13g2_a21oi_1 _25501_ (.A1(net5818),
    .A2(_18536_),
    .Y(_18538_),
    .B1(_18537_));
 sg13g2_xnor2_1 _25502_ (.Y(_18539_),
    .A(_15591_),
    .B(_16346_));
 sg13g2_a21oi_1 _25503_ (.A1(net5011),
    .A2(_18539_),
    .Y(_18540_),
    .B1(_18538_));
 sg13g2_inv_1 _25504_ (.Y(_18541_),
    .A(_18540_));
 sg13g2_a21oi_1 _25505_ (.A1(_16264_),
    .A2(_18059_),
    .Y(_18542_),
    .B1(_15475_));
 sg13g2_nand3_1 _25506_ (.B(_16264_),
    .C(_18059_),
    .A(_15475_),
    .Y(_18543_));
 sg13g2_nand2_1 _25507_ (.Y(_18544_),
    .A(net4990),
    .B(_18543_));
 sg13g2_o21ai_1 _25508_ (.B1(_15476_),
    .Y(_18545_),
    .A1(_15477_),
    .A2(_18055_));
 sg13g2_xnor2_1 _25509_ (.Y(_18546_),
    .A(_15475_),
    .B(_18545_));
 sg13g2_a21oi_1 _25510_ (.A1(net5797),
    .A2(_18546_),
    .Y(_18547_),
    .B1(net4990));
 sg13g2_o21ai_1 _25511_ (.B1(_18547_),
    .Y(_18548_),
    .A1(\u_inv.f_next[79] ),
    .A2(net5797));
 sg13g2_o21ai_1 _25512_ (.B1(_18548_),
    .Y(_18549_),
    .A1(_18542_),
    .A2(_18544_));
 sg13g2_nand3_1 _25513_ (.B(_16336_),
    .C(_17695_),
    .A(_15563_),
    .Y(_18550_));
 sg13g2_nand3_1 _25514_ (.B(_17696_),
    .C(_18550_),
    .A(net5014),
    .Y(_18551_));
 sg13g2_nand2_1 _25515_ (.Y(_18552_),
    .A(_15562_),
    .B(_15564_));
 sg13g2_o21ai_1 _25516_ (.B1(_18552_),
    .Y(_18553_),
    .A1(_14078_),
    .A2(_14350_));
 sg13g2_xnor2_1 _25517_ (.Y(_18554_),
    .A(_15563_),
    .B(_18553_));
 sg13g2_o21ai_1 _25518_ (.B1(net5100),
    .Y(_18555_),
    .A1(\u_inv.f_next[97] ),
    .A2(net5824));
 sg13g2_a21o_1 _25519_ (.A2(_18554_),
    .A1(net5824),
    .B1(_18555_),
    .X(_18556_));
 sg13g2_o21ai_1 _25520_ (.B1(_18556_),
    .Y(_18557_),
    .A1(_16337_),
    .A2(_18551_));
 sg13g2_nand3_1 _25521_ (.B(_16309_),
    .C(_16325_),
    .A(_15564_),
    .Y(_18558_));
 sg13g2_o21ai_1 _25522_ (.B1(net5824),
    .Y(_18559_),
    .A1(_15562_),
    .A2(_15564_));
 sg13g2_nor2b_1 _25523_ (.A(_18559_),
    .B_N(_18552_),
    .Y(_18560_));
 sg13g2_a21oi_1 _25524_ (.A1(\u_inv.f_next[96] ),
    .A2(net5716),
    .Y(_18561_),
    .B1(_18560_));
 sg13g2_nand3_1 _25525_ (.B(_17695_),
    .C(_18558_),
    .A(net5014),
    .Y(_18562_));
 sg13g2_o21ai_1 _25526_ (.B1(_18562_),
    .Y(_18563_),
    .A1(net5013),
    .A2(_18561_));
 sg13g2_a21oi_1 _25527_ (.A1(_15513_),
    .A2(_17830_),
    .Y(_18564_),
    .B1(_15512_));
 sg13g2_a21oi_1 _25528_ (.A1(_15510_),
    .A2(_18564_),
    .Y(_18565_),
    .B1(net5706));
 sg13g2_o21ai_1 _25529_ (.B1(_18565_),
    .Y(_18566_),
    .A1(_15510_),
    .A2(_18564_));
 sg13g2_o21ai_1 _25530_ (.B1(_18566_),
    .Y(_18567_),
    .A1(\u_inv.f_next[83] ),
    .A2(net5806));
 sg13g2_nor3_1 _25531_ (.A(_15511_),
    .B(_16282_),
    .C(_17837_),
    .Y(_18568_));
 sg13g2_o21ai_1 _25532_ (.B1(_15511_),
    .Y(_18569_),
    .A1(_16282_),
    .A2(_17837_));
 sg13g2_nor2_1 _25533_ (.A(net5085),
    .B(_18568_),
    .Y(_18570_));
 sg13g2_nand2_1 _25534_ (.Y(_18571_),
    .A(_18569_),
    .B(_18570_));
 sg13g2_o21ai_1 _25535_ (.B1(_18571_),
    .Y(_18572_),
    .A1(net5000),
    .A2(_18567_));
 sg13g2_xnor2_1 _25536_ (.Y(_18573_),
    .A(_15136_),
    .B(_17706_));
 sg13g2_nor2_1 _25537_ (.A(\u_inv.f_next[98] ),
    .B(net5824),
    .Y(_18574_));
 sg13g2_a21oi_1 _25538_ (.A1(net5824),
    .A2(_18573_),
    .Y(_18575_),
    .B1(_18574_));
 sg13g2_nor2_1 _25539_ (.A(_15136_),
    .B(_17697_),
    .Y(_18576_));
 sg13g2_nor2_1 _25540_ (.A(net5100),
    .B(_18576_),
    .Y(_18577_));
 sg13g2_a22oi_1 _25541_ (.Y(_18578_),
    .B1(_18577_),
    .B2(_17806_),
    .A2(_18575_),
    .A1(net5100));
 sg13g2_inv_1 _25542_ (.Y(_18579_),
    .A(_18578_));
 sg13g2_xor2_1 _25543_ (.B(_17775_),
    .A(_15533_),
    .X(_18580_));
 sg13g2_nor2_1 _25544_ (.A(\u_inv.f_next[92] ),
    .B(net5822),
    .Y(_18581_));
 sg13g2_a21oi_1 _25545_ (.A1(net5821),
    .A2(_18580_),
    .Y(_18582_),
    .B1(_18581_));
 sg13g2_nand3_1 _25546_ (.B(_16311_),
    .C(_17764_),
    .A(_15533_),
    .Y(_18583_));
 sg13g2_and2_1 _25547_ (.A(net5013),
    .B(_17765_),
    .X(_18584_));
 sg13g2_a22oi_1 _25548_ (.Y(_18585_),
    .B1(_18583_),
    .B2(_18584_),
    .A2(_18582_),
    .A1(net5098));
 sg13g2_inv_1 _25549_ (.Y(_18586_),
    .A(_18585_));
 sg13g2_or2_1 _25550_ (.X(_18587_),
    .B(_18011_),
    .A(_17994_));
 sg13g2_or2_1 _25551_ (.X(_18588_),
    .B(_18115_),
    .A(_18100_));
 sg13g2_xnor2_1 _25552_ (.Y(_18589_),
    .A(_15588_),
    .B(_17630_));
 sg13g2_a21oi_1 _25553_ (.A1(net5826),
    .A2(_18589_),
    .Y(_18590_),
    .B1(net5012));
 sg13g2_o21ai_1 _25554_ (.B1(_18590_),
    .Y(_18591_),
    .A1(\u_inv.f_next[106] ),
    .A2(net5819));
 sg13g2_nand3_1 _25555_ (.B(_16355_),
    .C(_17753_),
    .A(_15587_),
    .Y(_18592_));
 sg13g2_nand2_1 _25556_ (.Y(_18593_),
    .A(net5012),
    .B(_18592_));
 sg13g2_o21ai_1 _25557_ (.B1(_18591_),
    .Y(_18594_),
    .A1(_17754_),
    .A2(_18593_));
 sg13g2_a21oi_1 _25558_ (.A1(_15580_),
    .A2(_17631_),
    .Y(_18595_),
    .B1(_15579_));
 sg13g2_xnor2_1 _25559_ (.Y(_18596_),
    .A(_15578_),
    .B(_18595_));
 sg13g2_o21ai_1 _25560_ (.B1(net5097),
    .Y(_18597_),
    .A1(\u_inv.f_next[109] ),
    .A2(net5818));
 sg13g2_a21oi_1 _25561_ (.A1(net5819),
    .A2(_18596_),
    .Y(_18598_),
    .B1(_18597_));
 sg13g2_nand3_1 _25562_ (.B(_16361_),
    .C(_17622_),
    .A(_15577_),
    .Y(_18599_));
 sg13g2_nor2_1 _25563_ (.A(net5097),
    .B(_17623_),
    .Y(_18600_));
 sg13g2_a21o_2 _25564_ (.A2(_18600_),
    .A1(_18599_),
    .B1(_18598_),
    .X(_18601_));
 sg13g2_and3_1 _25565_ (.X(_18602_),
    .A(_15532_),
    .B(_15555_),
    .C(_17776_));
 sg13g2_o21ai_1 _25566_ (.B1(net5822),
    .Y(_18603_),
    .A1(_17777_),
    .A2(_18602_));
 sg13g2_o21ai_1 _25567_ (.B1(net5098),
    .Y(_18604_),
    .A1(\u_inv.f_next[94] ),
    .A2(net5821));
 sg13g2_nand2b_1 _25568_ (.Y(_18605_),
    .B(_18603_),
    .A_N(_18604_));
 sg13g2_xnor2_1 _25569_ (.Y(_18606_),
    .A(_15532_),
    .B(_17768_));
 sg13g2_o21ai_1 _25570_ (.B1(_18605_),
    .Y(_18607_),
    .A1(net5099),
    .A2(_18606_));
 sg13g2_xnor2_1 _25571_ (.Y(_18608_),
    .A(_15636_),
    .B(_17481_));
 sg13g2_o21ai_1 _25572_ (.B1(net5087),
    .Y(_18609_),
    .A1(\u_inv.f_next[116] ),
    .A2(net5820));
 sg13g2_a21oi_1 _25573_ (.A1(net5820),
    .A2(_18608_),
    .Y(_18610_),
    .B1(_18609_));
 sg13g2_nor3_1 _25574_ (.A(_15636_),
    .B(_16393_),
    .C(_17488_),
    .Y(_18611_));
 sg13g2_nor2_1 _25575_ (.A(net5096),
    .B(_18611_),
    .Y(_18612_));
 sg13g2_a21o_2 _25576_ (.A2(_18612_),
    .A1(_17489_),
    .B1(_18610_),
    .X(_18613_));
 sg13g2_or4_1 _25577_ (.A(_18594_),
    .B(_18601_),
    .C(_18607_),
    .D(_18613_),
    .X(_18614_));
 sg13g2_xnor2_1 _25578_ (.Y(_18615_),
    .A(_15645_),
    .B(_17479_));
 sg13g2_o21ai_1 _25579_ (.B1(net5096),
    .Y(_18616_),
    .A1(\u_inv.f_next[114] ),
    .A2(net5820));
 sg13g2_a21oi_1 _25580_ (.A1(net5820),
    .A2(_18615_),
    .Y(_18617_),
    .B1(_18616_));
 sg13g2_nand3_1 _25581_ (.B(_16389_),
    .C(_17656_),
    .A(_15644_),
    .Y(_18618_));
 sg13g2_nor2_1 _25582_ (.A(net5096),
    .B(_17657_),
    .Y(_18619_));
 sg13g2_a21o_1 _25583_ (.A2(_18619_),
    .A1(_18618_),
    .B1(_18617_),
    .X(_18620_));
 sg13g2_xnor2_1 _25584_ (.Y(_18621_),
    .A(_15627_),
    .B(_17504_));
 sg13g2_nor2_1 _25585_ (.A(\u_inv.f_next[120] ),
    .B(net5807),
    .Y(_18622_));
 sg13g2_a21oi_1 _25586_ (.A1(net5807),
    .A2(_18621_),
    .Y(_18623_),
    .B1(_18622_));
 sg13g2_or2_1 _25587_ (.X(_18624_),
    .B(_17496_),
    .A(_15627_));
 sg13g2_a21oi_1 _25588_ (.A1(_15627_),
    .A2(_17496_),
    .Y(_18625_),
    .B1(net5086));
 sg13g2_a22oi_1 _25589_ (.Y(_18626_),
    .B1(_18624_),
    .B2(_18625_),
    .A2(_18623_),
    .A1(net5086));
 sg13g2_inv_1 _25590_ (.Y(_18627_),
    .A(_18626_));
 sg13g2_xnor2_1 _25591_ (.Y(_18628_),
    .A(_15731_),
    .B(_16414_));
 sg13g2_a21oi_1 _25592_ (.A1(_15682_),
    .A2(_15730_),
    .Y(_18629_),
    .B1(net5706));
 sg13g2_o21ai_1 _25593_ (.B1(_18629_),
    .Y(_18630_),
    .A1(_15682_),
    .A2(_15730_));
 sg13g2_a21oi_1 _25594_ (.A1(\u_inv.f_next[128] ),
    .A2(net5706),
    .Y(_18631_),
    .B1(net5000));
 sg13g2_a22oi_1 _25595_ (.Y(_18632_),
    .B1(_18630_),
    .B2(_18631_),
    .A2(_18628_),
    .A1(net5001));
 sg13g2_nor2_2 _25596_ (.A(_18627_),
    .B(_18632_),
    .Y(_18633_));
 sg13g2_a21oi_1 _25597_ (.A1(_15130_),
    .A2(_17707_),
    .Y(_18634_),
    .B1(_15129_));
 sg13g2_xnor2_1 _25598_ (.Y(_18635_),
    .A(_15128_),
    .B(_18634_));
 sg13g2_o21ai_1 _25599_ (.B1(net5100),
    .Y(_18636_),
    .A1(\u_inv.f_next[101] ),
    .A2(net5825));
 sg13g2_a21oi_1 _25600_ (.A1(net5824),
    .A2(_18635_),
    .Y(_18637_),
    .B1(_18636_));
 sg13g2_nor2_1 _25601_ (.A(_15128_),
    .B(_17700_),
    .Y(_18638_));
 sg13g2_nor3_1 _25602_ (.A(net5101),
    .B(_17701_),
    .C(_18638_),
    .Y(_18639_));
 sg13g2_nor2_2 _25603_ (.A(_18637_),
    .B(_18639_),
    .Y(_18640_));
 sg13g2_inv_1 _25604_ (.Y(_18641_),
    .A(_18640_));
 sg13g2_nand3_1 _25605_ (.B(_16390_),
    .C(_17655_),
    .A(_15651_),
    .Y(_18642_));
 sg13g2_nand3_1 _25606_ (.B(_17656_),
    .C(_18642_),
    .A(net5011),
    .Y(_18643_));
 sg13g2_a21oi_1 _25607_ (.A1(_15648_),
    .A2(_17478_),
    .Y(_18644_),
    .B1(_15651_));
 sg13g2_nand3_1 _25608_ (.B(_15651_),
    .C(_17478_),
    .A(_15648_),
    .Y(_18645_));
 sg13g2_nand2_1 _25609_ (.Y(_18646_),
    .A(net5820),
    .B(_18645_));
 sg13g2_nor2_1 _25610_ (.A(\u_inv.f_next[113] ),
    .B(net5820),
    .Y(_18647_));
 sg13g2_o21ai_1 _25611_ (.B1(net5096),
    .Y(_18648_),
    .A1(_18644_),
    .A2(_18646_));
 sg13g2_o21ai_1 _25612_ (.B1(_18643_),
    .Y(_18649_),
    .A1(_18647_),
    .A2(_18648_));
 sg13g2_a21oi_1 _25613_ (.A1(_15619_),
    .A2(_17607_),
    .Y(_18650_),
    .B1(net5707));
 sg13g2_a22oi_1 _25614_ (.Y(_18651_),
    .B1(_17608_),
    .B2(_18650_),
    .A2(net5707),
    .A1(\u_inv.f_next[124] ));
 sg13g2_or3_1 _25615_ (.A(_15619_),
    .B(_16411_),
    .C(_17613_),
    .X(_18652_));
 sg13g2_nand3_1 _25616_ (.B(_17614_),
    .C(_18652_),
    .A(net5003),
    .Y(_18653_));
 sg13g2_o21ai_1 _25617_ (.B1(_18653_),
    .Y(_18654_),
    .A1(net5003),
    .A2(_18651_));
 sg13g2_a21oi_1 _25618_ (.A1(_15699_),
    .A2(_17227_),
    .Y(_18655_),
    .B1(net5697));
 sg13g2_a22oi_1 _25619_ (.Y(_18656_),
    .B1(_17646_),
    .B2(_18655_),
    .A2(net5697),
    .A1(\u_inv.f_next[136] ));
 sg13g2_nand2_1 _25620_ (.Y(_18657_),
    .A(_15698_),
    .B(_17217_));
 sg13g2_a21oi_1 _25621_ (.A1(_17515_),
    .A2(_18657_),
    .Y(_18658_),
    .B1(net5078));
 sg13g2_a21oi_2 _25622_ (.B1(_18658_),
    .Y(_18659_),
    .A2(_18656_),
    .A1(net5077));
 sg13g2_xnor2_1 _25623_ (.Y(_18660_),
    .A(_15720_),
    .B(_17226_));
 sg13g2_o21ai_1 _25624_ (.B1(net5090),
    .Y(_18661_),
    .A1(\u_inv.f_next[132] ),
    .A2(net5805));
 sg13g2_a21o_1 _25625_ (.A2(_18660_),
    .A1(net5805),
    .B1(_18661_),
    .X(_18662_));
 sg13g2_nor3_1 _25626_ (.A(_15720_),
    .B(_16430_),
    .C(_17308_),
    .Y(_18663_));
 sg13g2_nand2_1 _25627_ (.Y(_18664_),
    .A(net5001),
    .B(_17309_));
 sg13g2_o21ai_1 _25628_ (.B1(_18662_),
    .Y(_18665_),
    .A1(_18663_),
    .A2(_18664_));
 sg13g2_o21ai_1 _25629_ (.B1(_15635_),
    .Y(_18666_),
    .A1(_15636_),
    .A2(_17481_));
 sg13g2_xnor2_1 _25630_ (.Y(_18667_),
    .A(_15637_),
    .B(_18666_));
 sg13g2_o21ai_1 _25631_ (.B1(net5087),
    .Y(_18668_),
    .A1(\u_inv.f_next[117] ),
    .A2(net5808));
 sg13g2_a21oi_1 _25632_ (.A1(net5807),
    .A2(_18667_),
    .Y(_18669_),
    .B1(_18668_));
 sg13g2_nand3_1 _25633_ (.B(_16384_),
    .C(_17489_),
    .A(_15637_),
    .Y(_18670_));
 sg13g2_nor2_1 _25634_ (.A(net5086),
    .B(_17490_),
    .Y(_18671_));
 sg13g2_a21o_2 _25635_ (.A2(_18671_),
    .A1(_18670_),
    .B1(_18669_),
    .X(_18672_));
 sg13g2_o21ai_1 _25636_ (.B1(_15626_),
    .Y(_18673_),
    .A1(_15627_),
    .A2(_17504_));
 sg13g2_xnor2_1 _25637_ (.Y(_18674_),
    .A(_15628_),
    .B(_18673_));
 sg13g2_o21ai_1 _25638_ (.B1(net5086),
    .Y(_18675_),
    .A1(\u_inv.f_next[121] ),
    .A2(net5807));
 sg13g2_a21oi_1 _25639_ (.A1(net5807),
    .A2(_18674_),
    .Y(_18676_),
    .B1(_18675_));
 sg13g2_nand2_1 _25640_ (.Y(_18677_),
    .A(_15628_),
    .B(_17497_));
 sg13g2_nor2_1 _25641_ (.A(net5086),
    .B(_17498_),
    .Y(_18678_));
 sg13g2_a21oi_2 _25642_ (.B1(_18676_),
    .Y(_18679_),
    .A2(_18678_),
    .A1(_18677_));
 sg13g2_inv_1 _25643_ (.Y(_18680_),
    .A(_18679_));
 sg13g2_nand3_1 _25644_ (.B(_15736_),
    .C(_15758_),
    .A(_15095_),
    .Y(_18681_));
 sg13g2_a21oi_1 _25645_ (.A1(_17076_),
    .A2(_18681_),
    .Y(_18682_),
    .B1(net5699));
 sg13g2_o21ai_1 _25646_ (.B1(net5078),
    .Y(_18683_),
    .A1(\u_inv.f_next[144] ),
    .A2(net5796));
 sg13g2_nand2_1 _25647_ (.Y(_18684_),
    .A(_15095_),
    .B(_17068_));
 sg13g2_a21oi_1 _25648_ (.A1(_15095_),
    .A2(_17068_),
    .Y(_18685_),
    .B1(net5078));
 sg13g2_o21ai_1 _25649_ (.B1(_18685_),
    .Y(_18686_),
    .A1(_15095_),
    .A2(_17068_));
 sg13g2_o21ai_1 _25650_ (.B1(_18686_),
    .Y(_18687_),
    .A1(_18682_),
    .A2(_18683_));
 sg13g2_a21oi_1 _25651_ (.A1(_15682_),
    .A2(_15730_),
    .Y(_18688_),
    .B1(_15729_));
 sg13g2_xnor2_1 _25652_ (.Y(_18689_),
    .A(_15728_),
    .B(_18688_));
 sg13g2_nand2_1 _25653_ (.Y(_18690_),
    .A(net5806),
    .B(_18689_));
 sg13g2_a21oi_1 _25654_ (.A1(_14045_),
    .A2(net5706),
    .Y(_18691_),
    .B1(net5001));
 sg13g2_nor3_1 _25655_ (.A(_15728_),
    .B(_16424_),
    .C(_17537_),
    .Y(_18692_));
 sg13g2_nor2_1 _25656_ (.A(net5085),
    .B(_18692_),
    .Y(_18693_));
 sg13g2_a22oi_1 _25657_ (.Y(_18694_),
    .B1(_18693_),
    .B2(_17538_),
    .A2(_18691_),
    .A1(_18690_));
 sg13g2_a21oi_1 _25658_ (.A1(\u_inv.f_next[144] ),
    .A2(_14398_),
    .Y(_18695_),
    .B1(_15083_));
 sg13g2_nand2_1 _25659_ (.Y(_18696_),
    .A(net4991),
    .B(_16027_));
 sg13g2_a221oi_1 _25660_ (.B2(_18695_),
    .C1(_18696_),
    .B1(_18684_),
    .A1(_16060_),
    .Y(_18697_),
    .A2(_17068_));
 sg13g2_xnor2_1 _25661_ (.Y(_18698_),
    .A(_15083_),
    .B(_17525_));
 sg13g2_nor2_1 _25662_ (.A(net5699),
    .B(_18698_),
    .Y(_18699_));
 sg13g2_o21ai_1 _25663_ (.B1(net5078),
    .Y(_18700_),
    .A1(\u_inv.f_next[145] ),
    .A2(net5796));
 sg13g2_nor2_1 _25664_ (.A(_18699_),
    .B(_18700_),
    .Y(_18701_));
 sg13g2_nor2_1 _25665_ (.A(_18697_),
    .B(_18701_),
    .Y(_18702_));
 sg13g2_inv_1 _25666_ (.Y(_18703_),
    .A(_18702_));
 sg13g2_xor2_1 _25667_ (.B(_17166_),
    .A(_14971_),
    .X(_18704_));
 sg13g2_a21oi_1 _25668_ (.A1(_14971_),
    .A2(_17174_),
    .Y(_18705_),
    .B1(net5691));
 sg13g2_nand2b_1 _25669_ (.Y(_18706_),
    .B(_18705_),
    .A_N(_17300_));
 sg13g2_a21oi_1 _25670_ (.A1(\u_inv.f_next[164] ),
    .A2(net5691),
    .Y(_18707_),
    .B1(net4977));
 sg13g2_a22oi_1 _25671_ (.Y(_18708_),
    .B1(_18706_),
    .B2(_18707_),
    .A2(_18704_),
    .A1(net4977));
 sg13g2_xnor2_1 _25672_ (.Y(_18709_),
    .A(_15767_),
    .B(_16459_));
 sg13g2_a21oi_1 _25673_ (.A1(_15765_),
    .A2(_15766_),
    .Y(_18710_),
    .B1(net5690));
 sg13g2_o21ai_1 _25674_ (.B1(_18710_),
    .Y(_18711_),
    .A1(_15765_),
    .A2(_15766_));
 sg13g2_a21oi_1 _25675_ (.A1(\u_inv.f_next[160] ),
    .A2(net5690),
    .Y(_18712_),
    .B1(net4978));
 sg13g2_a22oi_1 _25676_ (.Y(_18713_),
    .B1(_18711_),
    .B2(_18712_),
    .A2(_18709_),
    .A1(net4978));
 sg13g2_a21oi_1 _25677_ (.A1(\u_inv.f_next[160] ),
    .A2(_14414_),
    .Y(_18714_),
    .B1(_15768_));
 sg13g2_o21ai_1 _25678_ (.B1(_18714_),
    .Y(_18715_),
    .A1(_15767_),
    .A2(_16459_));
 sg13g2_and3_1 _25679_ (.X(_18716_),
    .A(net4977),
    .B(_16485_),
    .C(_17576_));
 sg13g2_o21ai_1 _25680_ (.B1(_14962_),
    .Y(_18717_),
    .A1(_15765_),
    .A2(_15766_));
 sg13g2_xor2_1 _25681_ (.B(_18717_),
    .A(_15768_),
    .X(_18718_));
 sg13g2_nand2_1 _25682_ (.Y(_18719_),
    .A(_14013_),
    .B(net5690));
 sg13g2_a21oi_1 _25683_ (.A1(net5782),
    .A2(_18718_),
    .Y(_18720_),
    .B1(net4977));
 sg13g2_a22oi_1 _25684_ (.Y(_18721_),
    .B1(_18719_),
    .B2(_18720_),
    .A2(_18716_),
    .A1(_18715_));
 sg13g2_inv_1 _25685_ (.Y(_18722_),
    .A(_18721_));
 sg13g2_o21ai_1 _25686_ (.B1(_15719_),
    .Y(_18723_),
    .A1(_15720_),
    .A2(_17226_));
 sg13g2_xor2_1 _25687_ (.B(_18723_),
    .A(_15718_),
    .X(_18724_));
 sg13g2_o21ai_1 _25688_ (.B1(net5090),
    .Y(_18725_),
    .A1(\u_inv.f_next[133] ),
    .A2(net5805));
 sg13g2_a21o_1 _25689_ (.A2(_18724_),
    .A1(net5805),
    .B1(_18725_),
    .X(_18726_));
 sg13g2_nand4_1 _25690_ (.B(_15717_),
    .C(_16434_),
    .A(_15716_),
    .Y(_18727_),
    .D(_17309_));
 sg13g2_nand3_1 _25691_ (.B(_16435_),
    .C(_18727_),
    .A(net5001),
    .Y(_18728_));
 sg13g2_o21ai_1 _25692_ (.B1(_18726_),
    .Y(_18729_),
    .A1(_17310_),
    .A2(_18728_));
 sg13g2_xnor2_1 _25693_ (.Y(_18730_),
    .A(_15687_),
    .B(_17230_));
 sg13g2_a21oi_1 _25694_ (.A1(net5794),
    .A2(_18730_),
    .Y(_18731_),
    .B1(net4991));
 sg13g2_o21ai_1 _25695_ (.B1(_18731_),
    .Y(_18732_),
    .A1(\u_inv.f_next[142] ),
    .A2(net5794));
 sg13g2_nor3_1 _25696_ (.A(_15688_),
    .B(_16449_),
    .C(_17220_),
    .Y(_18733_));
 sg13g2_nand2_1 _25697_ (.Y(_18734_),
    .A(net4991),
    .B(_17221_));
 sg13g2_o21ai_1 _25698_ (.B1(_18732_),
    .Y(_18735_),
    .A1(_18733_),
    .A2(_18734_));
 sg13g2_a21oi_1 _25699_ (.A1(_16597_),
    .A2(_16599_),
    .Y(_18736_),
    .B1(_15876_));
 sg13g2_nor3_1 _25700_ (.A(_15874_),
    .B(_16615_),
    .C(_18736_),
    .Y(_18737_));
 sg13g2_nand2_1 _25701_ (.Y(_18738_),
    .A(net4952),
    .B(_16616_));
 sg13g2_nor3_1 _25702_ (.A(_16725_),
    .B(_18737_),
    .C(_18738_),
    .Y(_18739_));
 sg13g2_a21oi_1 _25703_ (.A1(_15875_),
    .A2(_16733_),
    .Y(_18740_),
    .B1(_15874_));
 sg13g2_and3_1 _25704_ (.X(_18741_),
    .A(_15874_),
    .B(_15875_),
    .C(_16733_));
 sg13g2_o21ai_1 _25705_ (.B1(net5751),
    .Y(_18742_),
    .A1(_18740_),
    .A2(_18741_));
 sg13g2_o21ai_1 _25706_ (.B1(net5041),
    .Y(_18743_),
    .A1(\u_inv.f_next[225] ),
    .A2(net5751));
 sg13g2_inv_1 _25707_ (.Y(_18744_),
    .A(_18743_));
 sg13g2_a21oi_2 _25708_ (.B1(_18739_),
    .Y(_18745_),
    .A2(_18744_),
    .A1(_18742_));
 sg13g2_inv_1 _25709_ (.Y(_18746_),
    .A(_18745_));
 sg13g2_nand3_1 _25710_ (.B(_16442_),
    .C(_17518_),
    .A(_15704_),
    .Y(_18747_));
 sg13g2_a21o_1 _25711_ (.A2(_17518_),
    .A1(_16442_),
    .B1(_15704_),
    .X(_18748_));
 sg13g2_nand3_1 _25712_ (.B(_18747_),
    .C(_18748_),
    .A(net4991),
    .Y(_18749_));
 sg13g2_a21oi_1 _25713_ (.A1(_15706_),
    .A2(_17228_),
    .Y(_18750_),
    .B1(_15705_));
 sg13g2_xnor2_1 _25714_ (.Y(_18751_),
    .A(_15704_),
    .B(_18750_));
 sg13g2_nor2_1 _25715_ (.A(\u_inv.f_next[139] ),
    .B(net5794),
    .Y(_18752_));
 sg13g2_o21ai_1 _25716_ (.B1(net5077),
    .Y(_18753_),
    .A1(net5697),
    .A2(_18751_));
 sg13g2_o21ai_1 _25717_ (.B1(_18749_),
    .Y(_18754_),
    .A1(_18752_),
    .A2(_18753_));
 sg13g2_nor3_1 _25718_ (.A(_15852_),
    .B(_15855_),
    .C(_15876_),
    .Y(_18755_));
 sg13g2_nor2_1 _25719_ (.A(_13950_),
    .B(net5751),
    .Y(_18756_));
 sg13g2_nor2_1 _25720_ (.A(net5674),
    .B(_18755_),
    .Y(_18757_));
 sg13g2_a21o_1 _25721_ (.A2(_18757_),
    .A1(_16733_),
    .B1(_18756_),
    .X(_18758_));
 sg13g2_and3_1 _25722_ (.X(_18759_),
    .A(_15876_),
    .B(_16597_),
    .C(_16599_));
 sg13g2_nor3_1 _25723_ (.A(net5041),
    .B(_18736_),
    .C(_18759_),
    .Y(_18760_));
 sg13g2_a21oi_2 _25724_ (.B1(_18760_),
    .Y(_18761_),
    .A2(_18758_),
    .A1(net5041));
 sg13g2_a21o_1 _25725_ (.A2(_18758_),
    .A1(net5041),
    .B1(_18760_),
    .X(_18762_));
 sg13g2_o21ai_1 _25726_ (.B1(_14941_),
    .Y(_18763_),
    .A1(_14942_),
    .A2(_16994_));
 sg13g2_xnor2_1 _25727_ (.Y(_18764_),
    .A(_14940_),
    .B(_18763_));
 sg13g2_o21ai_1 _25728_ (.B1(net5056),
    .Y(_18765_),
    .A1(\u_inv.f_next[181] ),
    .A2(net5767));
 sg13g2_a21oi_1 _25729_ (.A1(net5767),
    .A2(_18764_),
    .Y(_18766_),
    .B1(_18765_));
 sg13g2_nand3b_1 _25730_ (.B(_14940_),
    .C(_16528_),
    .Y(_18767_),
    .A_N(_17002_));
 sg13g2_nand4_1 _25731_ (.B(_16529_),
    .C(_17003_),
    .A(net4963),
    .Y(_18768_),
    .D(_18767_));
 sg13g2_nor2b_2 _25732_ (.A(_18766_),
    .B_N(_18768_),
    .Y(_18769_));
 sg13g2_inv_1 _25733_ (.Y(_18770_),
    .A(_18769_));
 sg13g2_xnor2_1 _25734_ (.Y(_18771_),
    .A(_15008_),
    .B(_16966_));
 sg13g2_o21ai_1 _25735_ (.B1(net5065),
    .Y(_18772_),
    .A1(\u_inv.f_next[170] ),
    .A2(net5779));
 sg13g2_a21oi_1 _25736_ (.A1(net5778),
    .A2(_18771_),
    .Y(_18773_),
    .B1(_18772_));
 sg13g2_or3_1 _25737_ (.A(_15008_),
    .B(_16508_),
    .C(_16952_),
    .X(_18774_));
 sg13g2_nand3_1 _25738_ (.B(_17208_),
    .C(_18774_),
    .A(net4976),
    .Y(_18775_));
 sg13g2_nor2b_1 _25739_ (.A(_18773_),
    .B_N(_18775_),
    .Y(_18776_));
 sg13g2_nand2b_1 _25740_ (.Y(_18777_),
    .B(_18775_),
    .A_N(_18773_));
 sg13g2_nand3_1 _25741_ (.B(_16401_),
    .C(_17678_),
    .A(_15611_),
    .Y(_18778_));
 sg13g2_a21o_1 _25742_ (.A2(_17678_),
    .A1(_16401_),
    .B1(_15611_),
    .X(_18779_));
 sg13g2_nand3_1 _25743_ (.B(_18778_),
    .C(_18779_),
    .A(net5003),
    .Y(_18780_));
 sg13g2_o21ai_1 _25744_ (.B1(_15612_),
    .Y(_18781_),
    .A1(_15613_),
    .A2(_17673_));
 sg13g2_xnor2_1 _25745_ (.Y(_18782_),
    .A(_15611_),
    .B(_18781_));
 sg13g2_a21oi_1 _25746_ (.A1(net5809),
    .A2(_18782_),
    .Y(_18783_),
    .B1(net5003));
 sg13g2_o21ai_1 _25747_ (.B1(_18783_),
    .Y(_18784_),
    .A1(net3175),
    .A2(net5809));
 sg13g2_nand2_1 _25748_ (.Y(_18785_),
    .A(_18780_),
    .B(_18784_));
 sg13g2_xnor2_1 _25749_ (.Y(_18786_),
    .A(_15087_),
    .B(_17201_));
 sg13g2_nand2_1 _25750_ (.Y(_18787_),
    .A(_14024_),
    .B(net5698));
 sg13g2_a21oi_1 _25751_ (.A1(net5792),
    .A2(_18786_),
    .Y(_18788_),
    .B1(net4989));
 sg13g2_nand2_1 _25752_ (.Y(_18789_),
    .A(_18787_),
    .B(_18788_));
 sg13g2_nand3_1 _25753_ (.B(_16019_),
    .C(_17196_),
    .A(_15087_),
    .Y(_18790_));
 sg13g2_nor2_1 _25754_ (.A(net5075),
    .B(_17197_),
    .Y(_18791_));
 sg13g2_nand2_1 _25755_ (.Y(_18792_),
    .A(_18790_),
    .B(_18791_));
 sg13g2_a22oi_1 _25756_ (.Y(_18793_),
    .B1(_18790_),
    .B2(_18791_),
    .A2(_18788_),
    .A1(_18787_));
 sg13g2_nand2_1 _25757_ (.Y(_18794_),
    .A(_18789_),
    .B(_18792_));
 sg13g2_a21oi_1 _25758_ (.A1(_16055_),
    .A2(_17116_),
    .Y(_18795_),
    .B1(_15050_));
 sg13g2_nand3_1 _25759_ (.B(_16055_),
    .C(_17116_),
    .A(_15050_),
    .Y(_18796_));
 sg13g2_nand2_1 _25760_ (.Y(_18797_),
    .A(net4988),
    .B(_18796_));
 sg13g2_o21ai_1 _25761_ (.B1(_15051_),
    .Y(_18798_),
    .A1(_15053_),
    .A2(_17110_));
 sg13g2_xnor2_1 _25762_ (.Y(_18799_),
    .A(_15050_),
    .B(_18798_));
 sg13g2_a21oi_1 _25763_ (.A1(net5791),
    .A2(_18799_),
    .Y(_18800_),
    .B1(net4988));
 sg13g2_o21ai_1 _25764_ (.B1(_18800_),
    .Y(_18801_),
    .A1(\u_inv.f_next[159] ),
    .A2(net5791));
 sg13g2_o21ai_1 _25765_ (.B1(_18801_),
    .Y(_18802_),
    .A1(_18795_),
    .A2(_18797_));
 sg13g2_a21o_1 _25766_ (.A2(_16981_),
    .A1(_15987_),
    .B1(_14858_),
    .X(_18803_));
 sg13g2_nand3_1 _25767_ (.B(_15987_),
    .C(_16981_),
    .A(_14858_),
    .Y(_18804_));
 sg13g2_nand3_1 _25768_ (.B(_18803_),
    .C(_18804_),
    .A(net4952),
    .Y(_18805_));
 sg13g2_and3_1 _25769_ (.X(_18806_),
    .A(_14858_),
    .B(_14859_),
    .C(_16976_));
 sg13g2_a21oi_1 _25770_ (.A1(_14859_),
    .A2(_16976_),
    .Y(_18807_),
    .B1(_14858_));
 sg13g2_nor3_1 _25771_ (.A(net5674),
    .B(_18806_),
    .C(_18807_),
    .Y(_18808_));
 sg13g2_o21ai_1 _25772_ (.B1(net5042),
    .Y(_18809_),
    .A1(\u_inv.f_next[219] ),
    .A2(net5752));
 sg13g2_o21ai_1 _25773_ (.B1(_18805_),
    .Y(_18810_),
    .A1(_18808_),
    .A2(_18809_));
 sg13g2_nand2_1 _25774_ (.Y(_18811_),
    .A(_16013_),
    .B(_17023_));
 sg13g2_a21oi_1 _25775_ (.A1(_14885_),
    .A2(_18811_),
    .Y(_18812_),
    .B1(net5044));
 sg13g2_o21ai_1 _25776_ (.B1(_18812_),
    .Y(_18813_),
    .A1(_14885_),
    .A2(_18811_));
 sg13g2_nor2_1 _25777_ (.A(_14880_),
    .B(_17014_),
    .Y(_18814_));
 sg13g2_o21ai_1 _25778_ (.B1(net5754),
    .Y(_18815_),
    .A1(_14884_),
    .A2(_18814_));
 sg13g2_a21oi_1 _25779_ (.A1(_14884_),
    .A2(_18814_),
    .Y(_18816_),
    .B1(_18815_));
 sg13g2_o21ai_1 _25780_ (.B1(net5044),
    .Y(_18817_),
    .A1(\u_inv.f_next[215] ),
    .A2(net5755));
 sg13g2_o21ai_1 _25781_ (.B1(_18813_),
    .Y(_18818_),
    .A1(_18816_),
    .A2(_18817_));
 sg13g2_a21oi_1 _25782_ (.A1(\u_inv.f_next[198] ),
    .A2(_14452_),
    .Y(_18819_),
    .B1(_17163_));
 sg13g2_a21oi_1 _25783_ (.A1(_15776_),
    .A2(_18819_),
    .Y(_18820_),
    .B1(net5052));
 sg13g2_o21ai_1 _25784_ (.B1(_18820_),
    .Y(_18821_),
    .A1(_15776_),
    .A2(_18819_));
 sg13g2_and3_1 _25785_ (.X(_18822_),
    .A(_15774_),
    .B(_15776_),
    .C(_17158_));
 sg13g2_a21oi_1 _25786_ (.A1(_15774_),
    .A2(_17158_),
    .Y(_18823_),
    .B1(_15776_));
 sg13g2_nor3_1 _25787_ (.A(net5681),
    .B(_18822_),
    .C(_18823_),
    .Y(_18824_));
 sg13g2_o21ai_1 _25788_ (.B1(net5052),
    .Y(_18825_),
    .A1(\u_inv.f_next[199] ),
    .A2(net5762));
 sg13g2_o21ai_1 _25789_ (.B1(_18821_),
    .Y(_18826_),
    .A1(_18824_),
    .A2(_18825_));
 sg13g2_a21o_1 _25790_ (.A2(_17150_),
    .A1(_14894_),
    .B1(_16001_),
    .X(_18827_));
 sg13g2_o21ai_1 _25791_ (.B1(net4953),
    .Y(_18828_),
    .A1(_14892_),
    .A2(_18827_));
 sg13g2_a21oi_1 _25792_ (.A1(_14892_),
    .A2(_18827_),
    .Y(_18829_),
    .B1(_18828_));
 sg13g2_o21ai_1 _25793_ (.B1(_14892_),
    .Y(_18830_),
    .A1(_14893_),
    .A2(_17153_));
 sg13g2_nor3_1 _25794_ (.A(_14892_),
    .B(_14893_),
    .C(_17153_),
    .Y(_18831_));
 sg13g2_nor2_1 _25795_ (.A(net5672),
    .B(_18831_),
    .Y(_18832_));
 sg13g2_a221oi_1 _25796_ (.B2(_18832_),
    .C1(net4953),
    .B1(_18830_),
    .A1(_13963_),
    .Y(_18833_),
    .A2(net5672));
 sg13g2_or2_1 _25797_ (.X(_18834_),
    .B(_18833_),
    .A(_18829_));
 sg13g2_xnor2_1 _25798_ (.Y(_18835_),
    .A(_14996_),
    .B(_16970_));
 sg13g2_nor2_1 _25799_ (.A(\u_inv.f_next[174] ),
    .B(net5777),
    .Y(_18836_));
 sg13g2_o21ai_1 _25800_ (.B1(net5066),
    .Y(_18837_),
    .A1(net5692),
    .A2(_18835_));
 sg13g2_nand3_1 _25801_ (.B(_16500_),
    .C(_16957_),
    .A(_14996_),
    .Y(_18838_));
 sg13g2_nand3_1 _25802_ (.B(_16958_),
    .C(_18838_),
    .A(net4976),
    .Y(_18839_));
 sg13g2_o21ai_1 _25803_ (.B1(_18839_),
    .Y(_18840_),
    .A1(_18836_),
    .A2(_18837_));
 sg13g2_nand2_1 _25804_ (.Y(_18841_),
    .A(_16587_),
    .B(_17145_));
 sg13g2_a21oi_1 _25805_ (.A1(_15818_),
    .A2(_18841_),
    .Y(_18842_),
    .B1(net5045));
 sg13g2_o21ai_1 _25806_ (.B1(_18842_),
    .Y(_18843_),
    .A1(_15818_),
    .A2(_18841_));
 sg13g2_a21oi_1 _25807_ (.A1(_15815_),
    .A2(_17140_),
    .Y(_18844_),
    .B1(_15814_));
 sg13g2_xnor2_1 _25808_ (.Y(_18845_),
    .A(_15818_),
    .B(_18844_));
 sg13g2_a21oi_1 _25809_ (.A1(net5755),
    .A2(_18845_),
    .Y(_18846_),
    .B1(net4954));
 sg13g2_o21ai_1 _25810_ (.B1(_18846_),
    .Y(_18847_),
    .A1(\u_inv.f_next[203] ),
    .A2(net5755));
 sg13g2_nand2_1 _25811_ (.Y(_18848_),
    .A(_18843_),
    .B(_18847_));
 sg13g2_a21oi_1 _25812_ (.A1(_15800_),
    .A2(_17136_),
    .Y(_18849_),
    .B1(_16581_));
 sg13g2_a21oi_1 _25813_ (.A1(_15801_),
    .A2(_18849_),
    .Y(_18850_),
    .B1(net5045));
 sg13g2_o21ai_1 _25814_ (.B1(_18850_),
    .Y(_18851_),
    .A1(_15801_),
    .A2(_18849_));
 sg13g2_a21oi_1 _25815_ (.A1(_15798_),
    .A2(_17129_),
    .Y(_18852_),
    .B1(_15801_));
 sg13g2_and3_1 _25816_ (.X(_18853_),
    .A(_15798_),
    .B(_15801_),
    .C(_17129_));
 sg13g2_nor3_1 _25817_ (.A(net5672),
    .B(_18852_),
    .C(_18853_),
    .Y(_18854_));
 sg13g2_o21ai_1 _25818_ (.B1(net5045),
    .Y(_18855_),
    .A1(\u_inv.f_next[207] ),
    .A2(net5755));
 sg13g2_o21ai_1 _25819_ (.B1(_18851_),
    .Y(_18856_),
    .A1(_18854_),
    .A2(_18855_));
 sg13g2_nor2_1 _25820_ (.A(\u_inv.f_next[255] ),
    .B(\u_inv.f_reg[255] ),
    .Y(_18857_));
 sg13g2_nand2_1 _25821_ (.Y(_18858_),
    .A(\u_inv.f_next[255] ),
    .B(\u_inv.f_reg[255] ));
 sg13g2_nor2b_2 _25822_ (.A(_18857_),
    .B_N(_18858_),
    .Y(_18859_));
 sg13g2_nor2_1 _25823_ (.A(_13920_),
    .B(\u_inv.f_reg[254] ),
    .Y(_18860_));
 sg13g2_nand2_1 _25824_ (.Y(_18861_),
    .A(\u_inv.f_next[254] ),
    .B(\u_inv.f_reg[254] ));
 sg13g2_nor2_1 _25825_ (.A(\u_inv.f_next[254] ),
    .B(\u_inv.f_reg[254] ),
    .Y(_18862_));
 sg13g2_xor2_1 _25826_ (.B(\u_inv.f_reg[254] ),
    .A(\u_inv.f_next[254] ),
    .X(_18863_));
 sg13g2_nor2_1 _25827_ (.A(_13921_),
    .B(\u_inv.f_reg[253] ),
    .Y(_18864_));
 sg13g2_a21oi_1 _25828_ (.A1(_16936_),
    .A2(_16937_),
    .Y(_18865_),
    .B1(_18864_));
 sg13g2_a21oi_1 _25829_ (.A1(_16941_),
    .A2(_18865_),
    .Y(_18866_),
    .B1(_18863_));
 sg13g2_nor2_1 _25830_ (.A(_18860_),
    .B(_18866_),
    .Y(_18867_));
 sg13g2_a21oi_1 _25831_ (.A1(_18859_),
    .A2(_18867_),
    .Y(_18868_),
    .B1(net5031));
 sg13g2_o21ai_1 _25832_ (.B1(_18868_),
    .Y(_18869_),
    .A1(_18859_),
    .A2(_18867_));
 sg13g2_a21oi_1 _25833_ (.A1(\u_inv.f_next[253] ),
    .A2(\u_inv.f_reg[253] ),
    .Y(_18870_),
    .B1(_16916_));
 sg13g2_a21oi_1 _25834_ (.A1(_13921_),
    .A2(_14507_),
    .Y(_18871_),
    .B1(_18870_));
 sg13g2_or2_1 _25835_ (.X(_18872_),
    .B(_16936_),
    .A(_16917_));
 sg13g2_a221oi_1 _25836_ (.B2(_16920_),
    .C1(_18872_),
    .B1(_16922_),
    .A1(_15953_),
    .Y(_18873_),
    .A2(_16921_));
 sg13g2_o21ai_1 _25837_ (.B1(_18863_),
    .Y(_18874_),
    .A1(_18871_),
    .A2(_18873_));
 sg13g2_nand2_1 _25838_ (.Y(_18875_),
    .A(_18861_),
    .B(_18874_));
 sg13g2_xor2_1 _25839_ (.B(_18875_),
    .A(_18859_),
    .X(_18876_));
 sg13g2_nor2_1 _25840_ (.A(\u_inv.f_next[255] ),
    .B(net5736),
    .Y(_18877_));
 sg13g2_o21ai_1 _25841_ (.B1(net5031),
    .Y(_18878_),
    .A1(net5663),
    .A2(_18876_));
 sg13g2_o21ai_1 _25842_ (.B1(_18869_),
    .Y(_18879_),
    .A1(_18877_),
    .A2(_18878_));
 sg13g2_or3_1 _25843_ (.A(_18863_),
    .B(_18871_),
    .C(_18873_),
    .X(_18880_));
 sg13g2_a21o_1 _25844_ (.A2(_18880_),
    .A1(_18874_),
    .B1(net5663),
    .X(_18881_));
 sg13g2_a21oi_1 _25845_ (.A1(_13920_),
    .A2(net5663),
    .Y(_18882_),
    .B1(net4938));
 sg13g2_nand3_1 _25846_ (.B(_18863_),
    .C(_18865_),
    .A(_16941_),
    .Y(_18883_));
 sg13g2_nor2_1 _25847_ (.A(net5031),
    .B(_18866_),
    .Y(_18884_));
 sg13g2_a22oi_1 _25848_ (.Y(_18885_),
    .B1(_18883_),
    .B2(_18884_),
    .A2(_18882_),
    .A1(_18881_));
 sg13g2_inv_1 _25849_ (.Y(_18886_),
    .A(_18885_));
 sg13g2_nor2_1 _25850_ (.A(\u_inv.f_next[256] ),
    .B(net5839),
    .Y(_18887_));
 sg13g2_xnor2_1 _25851_ (.Y(_18888_),
    .A(\u_inv.f_next[256] ),
    .B(net5839));
 sg13g2_nor3_1 _25852_ (.A(_16940_),
    .B(_18859_),
    .C(_18863_),
    .Y(_18889_));
 sg13g2_nand2_1 _25853_ (.Y(_18890_),
    .A(\u_inv.f_next[255] ),
    .B(_14509_));
 sg13g2_nor2_1 _25854_ (.A(_18863_),
    .B(_18865_),
    .Y(_18891_));
 sg13g2_nor2_1 _25855_ (.A(_18860_),
    .B(_18891_),
    .Y(_18892_));
 sg13g2_o21ai_1 _25856_ (.B1(_18890_),
    .Y(_18893_),
    .A1(_18859_),
    .A2(_18892_));
 sg13g2_a21o_1 _25857_ (.A2(_18889_),
    .A1(_16932_),
    .B1(_18893_),
    .X(_18894_));
 sg13g2_a21oi_1 _25858_ (.A1(_18888_),
    .A2(_18894_),
    .Y(_18895_),
    .B1(net5031));
 sg13g2_or2_1 _25859_ (.X(_18896_),
    .B(_18894_),
    .A(_18888_));
 sg13g2_nand2_1 _25860_ (.Y(_18897_),
    .A(\u_inv.f_next[256] ),
    .B(net5663));
 sg13g2_o21ai_1 _25861_ (.B1(_18858_),
    .Y(_18898_),
    .A1(_18857_),
    .A2(_18861_));
 sg13g2_or2_1 _25862_ (.X(_18899_),
    .B(_18898_),
    .A(_18871_));
 sg13g2_a21oi_1 _25863_ (.A1(_18858_),
    .A2(_18862_),
    .Y(_18900_),
    .B1(_18857_));
 sg13g2_o21ai_1 _25864_ (.B1(_18900_),
    .Y(_18901_),
    .A1(_18873_),
    .A2(_18899_));
 sg13g2_o21ai_1 _25865_ (.B1(net5736),
    .Y(_18902_),
    .A1(_18888_),
    .A2(_18901_));
 sg13g2_and2_1 _25866_ (.A(_18888_),
    .B(_18901_),
    .X(_18903_));
 sg13g2_o21ai_1 _25867_ (.B1(_18897_),
    .Y(_18904_),
    .A1(_18902_),
    .A2(_18903_));
 sg13g2_a22oi_1 _25868_ (.Y(_18905_),
    .B1(_18904_),
    .B2(net5031),
    .A2(_18896_),
    .A1(_18895_));
 sg13g2_nand2b_1 _25869_ (.Y(_18906_),
    .B(net5839),
    .A_N(\u_inv.f_next[256] ));
 sg13g2_o21ai_1 _25870_ (.B1(_18897_),
    .Y(_18907_),
    .A1(_18887_),
    .A2(_18902_));
 sg13g2_a22oi_1 _25871_ (.Y(_18908_),
    .B1(_18907_),
    .B2(net5031),
    .A2(_18906_),
    .A1(_18895_));
 sg13g2_inv_1 _25872_ (.Y(_18909_),
    .A(_18908_));
 sg13g2_nor2_1 _25873_ (.A(_16783_),
    .B(_18810_),
    .Y(_18910_));
 sg13g2_nand3_1 _25874_ (.B(_16914_),
    .C(_18910_),
    .A(_16760_),
    .Y(_18911_));
 sg13g2_or4_1 _25875_ (.A(_16772_),
    .B(_16844_),
    .C(_16904_),
    .D(_16909_),
    .X(_18912_));
 sg13g2_or4_1 _25876_ (.A(_16681_),
    .B(_16896_),
    .C(_18911_),
    .D(_18912_),
    .X(_18913_));
 sg13g2_nand4_1 _25877_ (.B(_16812_),
    .C(_16869_),
    .A(_16798_),
    .Y(_18914_),
    .D(_17010_));
 sg13g2_nor4_1 _25878_ (.A(_16790_),
    .B(_16836_),
    .C(_16984_),
    .D(_17118_),
    .Y(_18915_));
 sg13g2_nand2b_1 _25879_ (.Y(_18916_),
    .B(_18915_),
    .A_N(_16748_));
 sg13g2_or4_1 _25880_ (.A(_16741_),
    .B(_18802_),
    .C(_18914_),
    .D(_18916_),
    .X(_18917_));
 sg13g2_nand3b_1 _25881_ (.B(_18885_),
    .C(_18908_),
    .Y(_18918_),
    .A_N(_16948_));
 sg13g2_nor4_2 _25882_ (.A(_16701_),
    .B(_18913_),
    .C(_18917_),
    .Y(_18919_),
    .D(_18918_));
 sg13g2_nor3_1 _25883_ (.A(_16850_),
    .B(_16887_),
    .C(_16975_),
    .Y(_18920_));
 sg13g2_or4_1 _25884_ (.A(_17039_),
    .B(_17147_),
    .C(_17156_),
    .D(_17165_),
    .X(_18921_));
 sg13g2_nand2_1 _25885_ (.Y(_18922_),
    .A(_17067_),
    .B(_17385_));
 sg13g2_or4_1 _25886_ (.A(_17125_),
    .B(_17274_),
    .C(_17391_),
    .D(_18922_),
    .X(_18923_));
 sg13g2_nand4_1 _25887_ (.B(_18761_),
    .C(_18776_),
    .A(_18745_),
    .Y(_18924_),
    .D(_18793_));
 sg13g2_nor3_1 _25888_ (.A(_17358_),
    .B(_17360_),
    .C(_18924_),
    .Y(_18925_));
 sg13g2_nor3_1 _25889_ (.A(_17327_),
    .B(_17567_),
    .C(_17575_),
    .Y(_18926_));
 sg13g2_and2_1 _25890_ (.A(_17292_),
    .B(_18926_),
    .X(_18927_));
 sg13g2_nor4_1 _25891_ (.A(_17713_),
    .B(_17726_),
    .C(_17733_),
    .D(_17738_),
    .Y(_18928_));
 sg13g2_or4_1 _25892_ (.A(_17751_),
    .B(_17782_),
    .C(_18620_),
    .D(_18672_),
    .X(_18929_));
 sg13g2_or4_1 _25893_ (.A(_17762_),
    .B(_18665_),
    .C(_18697_),
    .D(_18701_),
    .X(_18930_));
 sg13g2_nor4_1 _25894_ (.A(_17619_),
    .B(_17694_),
    .C(_18929_),
    .D(_18930_),
    .Y(_18931_));
 sg13g2_or2_1 _25895_ (.X(_18932_),
    .B(_18654_),
    .A(_18614_));
 sg13g2_nand2b_1 _25896_ (.Y(_18933_),
    .B(_17821_),
    .A_N(_17791_));
 sg13g2_nor4_1 _25897_ (.A(_17796_),
    .B(_17805_),
    .C(_18649_),
    .D(_18933_),
    .Y(_18934_));
 sg13g2_nor4_1 _25898_ (.A(_18071_),
    .B(_18549_),
    .C(_18563_),
    .D(_18572_),
    .Y(_18935_));
 sg13g2_nand4_1 _25899_ (.B(_18540_),
    .C(_18585_),
    .A(_18080_),
    .Y(_18936_),
    .D(_18935_));
 sg13g2_nand2b_1 _25900_ (.Y(_18937_),
    .B(_17846_),
    .A_N(_17839_));
 sg13g2_nor4_2 _25901_ (.A(_17906_),
    .B(_18038_),
    .C(_18135_),
    .Y(_18938_),
    .D(_18141_));
 sg13g2_nor3_1 _25902_ (.A(_17869_),
    .B(_17888_),
    .C(_18046_),
    .Y(_18939_));
 sg13g2_nand2_2 _25903_ (.Y(_18940_),
    .A(_18938_),
    .B(_18939_));
 sg13g2_nor4_1 _25904_ (.A(_18557_),
    .B(_18588_),
    .C(_18937_),
    .D(_18940_),
    .Y(_18941_));
 sg13g2_or3_1 _25905_ (.A(_18129_),
    .B(_18528_),
    .C(_18535_),
    .X(_18942_));
 sg13g2_or2_1 _25906_ (.X(_18943_),
    .B(_18062_),
    .A(_17828_));
 sg13g2_nor2_1 _25907_ (.A(_17987_),
    .B(_18153_),
    .Y(_18944_));
 sg13g2_nor2_1 _25908_ (.A(_18159_),
    .B(_18191_),
    .Y(_18945_));
 sg13g2_or3_1 _25909_ (.A(_18445_),
    .B(_18451_),
    .C(_18510_),
    .X(_18946_));
 sg13g2_nand4_1 _25910_ (.B(_18458_),
    .C(_18468_),
    .A(_18437_),
    .Y(_18947_),
    .D(_18474_));
 sg13g2_nor4_2 _25911_ (.A(_18204_),
    .B(_18482_),
    .C(_18946_),
    .Y(_18948_),
    .D(_18947_));
 sg13g2_nor3_1 _25912_ (.A(_18168_),
    .B(_18180_),
    .C(_18212_),
    .Y(_18949_));
 sg13g2_nand3_1 _25913_ (.B(_18948_),
    .C(_18949_),
    .A(_18945_),
    .Y(_18950_));
 sg13g2_nor4_1 _25914_ (.A(_17949_),
    .B(_17966_),
    .C(_17972_),
    .D(_18950_),
    .Y(_18951_));
 sg13g2_nand3_1 _25915_ (.B(_18944_),
    .C(_18951_),
    .A(_17920_),
    .Y(_18952_));
 sg13g2_nor4_1 _25916_ (.A(_18147_),
    .B(_18186_),
    .C(_18196_),
    .D(_18505_),
    .Y(_18953_));
 sg13g2_or4_1 _25917_ (.A(_18489_),
    .B(_18497_),
    .C(_18516_),
    .D(_18522_),
    .X(_18954_));
 sg13g2_nor4_1 _25918_ (.A(_18174_),
    .B(_18219_),
    .C(_18229_),
    .D(_18954_),
    .Y(_18955_));
 sg13g2_nand2b_2 _25919_ (.Y(_18956_),
    .B(_18955_),
    .A_N(_18005_));
 sg13g2_nor4_1 _25920_ (.A(_17938_),
    .B(_17980_),
    .C(_18587_),
    .D(_18956_),
    .Y(_18957_));
 sg13g2_nand2_2 _25921_ (.Y(_18958_),
    .A(_18953_),
    .B(_18957_));
 sg13g2_or4_1 _25922_ (.A(_17860_),
    .B(_18022_),
    .C(_18030_),
    .D(_18958_),
    .X(_18959_));
 sg13g2_or4_1 _25923_ (.A(_17879_),
    .B(_18054_),
    .C(_18952_),
    .D(_18959_),
    .X(_18960_));
 sg13g2_nor4_2 _25924_ (.A(_18095_),
    .B(_18942_),
    .C(_18943_),
    .Y(_18961_),
    .D(_18960_));
 sg13g2_nand3_1 _25925_ (.B(_18941_),
    .C(_18961_),
    .A(_18578_),
    .Y(_18962_));
 sg13g2_nor4_1 _25926_ (.A(_17787_),
    .B(_17814_),
    .C(_18936_),
    .D(_18962_),
    .Y(_18963_));
 sg13g2_nand4_1 _25927_ (.B(_18640_),
    .C(_18934_),
    .A(_18633_),
    .Y(_18964_),
    .D(_18963_));
 sg13g2_or2_1 _25928_ (.X(_18965_),
    .B(_18729_),
    .A(_18713_));
 sg13g2_nor4_1 _25929_ (.A(_18708_),
    .B(_18932_),
    .C(_18964_),
    .D(_18965_),
    .Y(_18966_));
 sg13g2_nor2_1 _25930_ (.A(_17665_),
    .B(_17688_),
    .Y(_18967_));
 sg13g2_nand4_1 _25931_ (.B(_17668_),
    .C(_17670_),
    .A(_17639_),
    .Y(_18968_),
    .D(_18967_));
 sg13g2_nor2_1 _25932_ (.A(_18659_),
    .B(_18687_),
    .Y(_18969_));
 sg13g2_and2_1 _25933_ (.A(_18679_),
    .B(_18694_),
    .X(_18970_));
 sg13g2_nand4_1 _25934_ (.B(_18721_),
    .C(_18969_),
    .A(_17744_),
    .Y(_18971_),
    .D(_18970_));
 sg13g2_nor4_1 _25935_ (.A(_17555_),
    .B(_17719_),
    .C(_18968_),
    .D(_18971_),
    .Y(_18972_));
 sg13g2_and4_1 _25936_ (.A(_18928_),
    .B(_18931_),
    .C(_18966_),
    .D(_18972_),
    .X(_18973_));
 sg13g2_nor4_1 _25937_ (.A(_17548_),
    .B(_17599_),
    .C(_17606_),
    .D(_17654_),
    .Y(_18974_));
 sg13g2_nor3_1 _25938_ (.A(_17495_),
    .B(_17511_),
    .C(_17531_),
    .Y(_18975_));
 sg13g2_and4_1 _25939_ (.A(_17469_),
    .B(_17681_),
    .C(_18974_),
    .D(_18975_),
    .X(_18976_));
 sg13g2_nand4_1 _25940_ (.B(_18927_),
    .C(_18973_),
    .A(_18925_),
    .Y(_18977_),
    .D(_18976_));
 sg13g2_a221oi_1 _25941_ (.B2(_17260_),
    .C1(_16831_),
    .B1(_17259_),
    .A1(_17255_),
    .Y(_18978_),
    .A2(_17256_));
 sg13g2_nor2_1 _25942_ (.A(_17087_),
    .B(_17194_),
    .Y(_18979_));
 sg13g2_nor3_1 _25943_ (.A(_17187_),
    .B(_17238_),
    .C(_17242_),
    .Y(_18980_));
 sg13g2_nand4_1 _25944_ (.B(_18978_),
    .C(_18979_),
    .A(_16879_),
    .Y(_18981_),
    .D(_18980_));
 sg13g2_nor4_2 _25945_ (.A(_18921_),
    .B(_18923_),
    .C(_18977_),
    .Y(_18982_),
    .D(_18981_));
 sg13g2_nor4_2 _25946_ (.A(_17139_),
    .B(_18818_),
    .C(_18826_),
    .Y(_18983_),
    .D(_18856_));
 sg13g2_nand4_1 _25947_ (.B(_18920_),
    .C(_18982_),
    .A(_18905_),
    .Y(_18984_),
    .D(_18983_));
 sg13g2_nor4_1 _25948_ (.A(_16990_),
    .B(_17098_),
    .C(_17181_),
    .D(_17254_),
    .Y(_18985_));
 sg13g2_nor2b_1 _25949_ (.A(_17536_),
    .B_N(_17053_),
    .Y(_18986_));
 sg13g2_nor4_1 _25950_ (.A(_17299_),
    .B(_17397_),
    .C(_17403_),
    .D(_17410_),
    .Y(_18987_));
 sg13g2_and4_1 _25951_ (.A(_17282_),
    .B(_17415_),
    .C(_18986_),
    .D(_18987_),
    .X(_18988_));
 sg13g2_nand3_1 _25952_ (.B(_18780_),
    .C(_18784_),
    .A(_18769_),
    .Y(_18989_));
 sg13g2_nor4_1 _25953_ (.A(_17421_),
    .B(_17462_),
    .C(_18754_),
    .D(_18989_),
    .Y(_18990_));
 sg13g2_nand2b_1 _25954_ (.Y(_18991_),
    .B(_17307_),
    .A_N(_17340_));
 sg13g2_or4_1 _25955_ (.A(_17333_),
    .B(_17374_),
    .C(_17593_),
    .D(_18991_),
    .X(_18992_));
 sg13g2_or4_1 _25956_ (.A(_17321_),
    .B(_17348_),
    .C(_17354_),
    .D(_17585_),
    .X(_18993_));
 sg13g2_or4_1 _25957_ (.A(_17454_),
    .B(_17476_),
    .C(_17520_),
    .D(_17561_),
    .X(_18994_));
 sg13g2_nor4_1 _25958_ (.A(_18735_),
    .B(_18992_),
    .C(_18993_),
    .D(_18994_),
    .Y(_18995_));
 sg13g2_nand4_1 _25959_ (.B(_18988_),
    .C(_18990_),
    .A(_18985_),
    .Y(_18996_),
    .D(_18995_));
 sg13g2_nor4_1 _25960_ (.A(_17216_),
    .B(_17235_),
    .C(_17429_),
    .D(_17448_),
    .Y(_18997_));
 sg13g2_nor4_2 _25961_ (.A(_17207_),
    .B(_17368_),
    .C(_17379_),
    .Y(_18998_),
    .D(_17439_));
 sg13g2_nand4_1 _25962_ (.B(_17268_),
    .C(_18997_),
    .A(_16820_),
    .Y(_18999_),
    .D(_18998_));
 sg13g2_or3_1 _25963_ (.A(_16804_),
    .B(_17025_),
    .C(_17109_),
    .X(_19000_));
 sg13g2_or4_1 _25964_ (.A(_18834_),
    .B(_18840_),
    .C(_18848_),
    .D(_19000_),
    .X(_19001_));
 sg13g2_or4_1 _25965_ (.A(_16935_),
    .B(_18996_),
    .C(_18999_),
    .D(_19001_),
    .X(_19002_));
 sg13g2_nor4_2 _25966_ (.A(_16724_),
    .B(_18879_),
    .C(_18984_),
    .Y(_19003_),
    .D(_19002_));
 sg13g2_and2_1 _25967_ (.A(_18919_),
    .B(_19003_),
    .X(_19004_));
 sg13g2_nor4_1 _25968_ (.A(net5829),
    .B(\u_inv.counter[3] ),
    .C(\u_inv.counter[4] ),
    .D(\u_inv.counter[8] ),
    .Y(_19005_));
 sg13g2_a21oi_1 _25969_ (.A1(_14249_),
    .A2(_19005_),
    .Y(_19006_),
    .B1(_14826_));
 sg13g2_nor2b_2 _25970_ (.A(_19006_),
    .B_N(_18354_),
    .Y(_19007_));
 sg13g2_inv_4 _25971_ (.A(_19007_),
    .Y(_19008_));
 sg13g2_a21oi_2 _25972_ (.B1(_19008_),
    .Y(_19009_),
    .A2(_19003_),
    .A1(_18919_));
 sg13g2_nand2b_2 _25973_ (.Y(_19010_),
    .B(_19007_),
    .A_N(net4451));
 sg13g2_nor2_1 _25974_ (.A(net5624),
    .B(net4353),
    .Y(_19011_));
 sg13g2_nand2_2 _25975_ (.Y(_19012_),
    .A(net5634),
    .B(net4389));
 sg13g2_and3_1 _25976_ (.X(_19013_),
    .A(_14826_),
    .B(net5633),
    .C(net4389));
 sg13g2_nand2_1 _25977_ (.Y(_19014_),
    .A(inv_done),
    .B(_14811_));
 sg13g2_nor2b_1 _25978_ (.A(net3378),
    .B_N(net3331),
    .Y(_19015_));
 sg13g2_nand2b_1 _25979_ (.Y(_19016_),
    .B(net3331),
    .A_N(\u_inv.state[0] ));
 sg13g2_nand3_1 _25980_ (.B(_14811_),
    .C(_19015_),
    .A(net3417),
    .Y(_19017_));
 sg13g2_nand4_1 _25981_ (.B(net5881),
    .C(\u_inv.counter[9] ),
    .A(\u_inv.counter[0] ),
    .Y(_19018_),
    .D(_14254_));
 sg13g2_nor4_1 _25982_ (.A(\u_inv.counter[1] ),
    .B(\u_inv.counter[3] ),
    .C(\u_inv.counter[4] ),
    .D(_19018_),
    .Y(_19019_));
 sg13g2_nand2b_1 _25983_ (.Y(_19020_),
    .B(_19019_),
    .A_N(_14823_));
 sg13g2_nand3_1 _25984_ (.B(_19008_),
    .C(_19020_),
    .A(net5633),
    .Y(_19021_));
 sg13g2_nor2_1 _25985_ (.A(net4451),
    .B(_19021_),
    .Y(_19022_));
 sg13g2_o21ai_1 _25986_ (.B1(_19017_),
    .Y(_19023_),
    .A1(net4451),
    .A2(_19021_));
 sg13g2_or2_1 _25987_ (.X(_19024_),
    .B(_19022_),
    .A(_19013_));
 sg13g2_or4_1 _25988_ (.A(net3378),
    .B(_14246_),
    .C(_19013_),
    .D(_19023_),
    .X(_19025_));
 sg13g2_inv_2 _25989_ (.Y(_20877_[0]),
    .A(_19025_));
 sg13g2_nand2_1 _25990_ (.Y(_00000_),
    .A(_19014_),
    .B(net3332));
 sg13g2_and2_1 _25991_ (.A(net5885),
    .B(net5634),
    .X(_19026_));
 sg13g2_nand2_1 _25992_ (.Y(_19027_),
    .A(net5885),
    .B(net5634));
 sg13g2_nand2_2 _25993_ (.Y(_19028_),
    .A(net5627),
    .B(_19025_));
 sg13g2_o21ai_1 _25994_ (.B1(net5903),
    .Y(_19029_),
    .A1(net5632),
    .A2(_20877_[0]));
 sg13g2_o21ai_1 _25995_ (.B1(net5535),
    .Y(_19030_),
    .A1(net1745),
    .A2(net4146));
 sg13g2_nor2_1 _25996_ (.A(net5626),
    .B(net4389),
    .Y(_19031_));
 sg13g2_nand2_2 _25997_ (.Y(_19032_),
    .A(net5634),
    .B(net4353));
 sg13g2_a22oi_1 _25998_ (.Y(_19033_),
    .B1(net4312),
    .B2(_18497_),
    .A2(net4268),
    .A1(_18434_));
 sg13g2_a22oi_1 _25999_ (.Y(_00001_),
    .B1(_19030_),
    .B2(_19033_),
    .A2(net4146),
    .A1(_14144_));
 sg13g2_o21ai_1 _26000_ (.B1(net5535),
    .Y(_19034_),
    .A1(net1838),
    .A2(net4146));
 sg13g2_a22oi_1 _26001_ (.Y(_19035_),
    .B1(net4312),
    .B2(_18434_),
    .A2(net4268),
    .A1(_18459_));
 sg13g2_a22oi_1 _26002_ (.Y(_00002_),
    .B1(_19034_),
    .B2(_19035_),
    .A2(net4146),
    .A1(_14143_));
 sg13g2_o21ai_1 _26003_ (.B1(net5535),
    .Y(_19036_),
    .A1(net1792),
    .A2(net4146));
 sg13g2_a22oi_1 _26004_ (.Y(_19037_),
    .B1(net4312),
    .B2(_18459_),
    .A2(net4268),
    .A1(_18516_));
 sg13g2_a22oi_1 _26005_ (.Y(_00003_),
    .B1(_19036_),
    .B2(_19037_),
    .A2(net4146),
    .A1(_14142_));
 sg13g2_o21ai_1 _26006_ (.B1(net5542),
    .Y(_19038_),
    .A1(net2286),
    .A2(net4158));
 sg13g2_a22oi_1 _26007_ (.Y(_19039_),
    .B1(net4316),
    .B2(_18516_),
    .A2(net4273),
    .A1(_18229_));
 sg13g2_a22oi_1 _26008_ (.Y(_00004_),
    .B1(_19038_),
    .B2(_19039_),
    .A2(net4158),
    .A1(_14141_));
 sg13g2_o21ai_1 _26009_ (.B1(net5542),
    .Y(_19040_),
    .A1(net1741),
    .A2(net4158));
 sg13g2_a22oi_1 _26010_ (.Y(_19041_),
    .B1(net4316),
    .B2(_18229_),
    .A2(net4273),
    .A1(_18522_));
 sg13g2_a22oi_1 _26011_ (.Y(_00005_),
    .B1(_19040_),
    .B2(_19041_),
    .A2(net4158),
    .A1(_14140_));
 sg13g2_o21ai_1 _26012_ (.B1(net5542),
    .Y(_19042_),
    .A1(net1753),
    .A2(net4157));
 sg13g2_a22oi_1 _26013_ (.Y(_19043_),
    .B1(net4316),
    .B2(_18522_),
    .A2(net4273),
    .A1(_18219_));
 sg13g2_a22oi_1 _26014_ (.Y(_00006_),
    .B1(_19042_),
    .B2(_19043_),
    .A2(net4157),
    .A1(_14139_));
 sg13g2_o21ai_1 _26015_ (.B1(net5542),
    .Y(_19044_),
    .A1(net1529),
    .A2(net4157));
 sg13g2_a22oi_1 _26016_ (.Y(_19045_),
    .B1(net4316),
    .B2(_18219_),
    .A2(net4273),
    .A1(_18159_));
 sg13g2_a22oi_1 _26017_ (.Y(_00007_),
    .B1(_19044_),
    .B2(_19045_),
    .A2(net4158),
    .A1(_14138_));
 sg13g2_o21ai_1 _26018_ (.B1(net5542),
    .Y(_19046_),
    .A1(net1755),
    .A2(net4157));
 sg13g2_a22oi_1 _26019_ (.Y(_19047_),
    .B1(net4316),
    .B2(_18159_),
    .A2(net4273),
    .A1(_17938_));
 sg13g2_a22oi_1 _26020_ (.Y(_00008_),
    .B1(_19046_),
    .B2(_19047_),
    .A2(net4158),
    .A1(_14137_));
 sg13g2_o21ai_1 _26021_ (.B1(net5542),
    .Y(_19048_),
    .A1(net1677),
    .A2(net4157));
 sg13g2_a22oi_1 _26022_ (.Y(_19049_),
    .B1(net4316),
    .B2(_17938_),
    .A2(net4273),
    .A1(_18451_));
 sg13g2_a22oi_1 _26023_ (.Y(_00009_),
    .B1(_19048_),
    .B2(_19049_),
    .A2(net4157),
    .A1(_14136_));
 sg13g2_o21ai_1 _26024_ (.B1(net5542),
    .Y(_19050_),
    .A1(net1928),
    .A2(net4157));
 sg13g2_a22oi_1 _26025_ (.Y(_19051_),
    .B1(net4316),
    .B2(_18451_),
    .A2(net4273),
    .A1(_18489_));
 sg13g2_a22oi_1 _26026_ (.Y(_00010_),
    .B1(_19050_),
    .B2(_19051_),
    .A2(net4157),
    .A1(_14135_));
 sg13g2_o21ai_1 _26027_ (.B1(net5545),
    .Y(_19052_),
    .A1(net1778),
    .A2(net4164));
 sg13g2_a22oi_1 _26028_ (.Y(_19053_),
    .B1(net4316),
    .B2(_18489_),
    .A2(net4276),
    .A1(_18174_));
 sg13g2_a22oi_1 _26029_ (.Y(_00011_),
    .B1(_19052_),
    .B2(_19053_),
    .A2(net4164),
    .A1(_14134_));
 sg13g2_o21ai_1 _26030_ (.B1(net5545),
    .Y(_19054_),
    .A1(net2048),
    .A2(net4164));
 sg13g2_a22oi_1 _26031_ (.Y(_19055_),
    .B1(net4319),
    .B2(_18174_),
    .A2(net4276),
    .A1(_18005_));
 sg13g2_a22oi_1 _26032_ (.Y(_00012_),
    .B1(_19054_),
    .B2(_19055_),
    .A2(net4164),
    .A1(_14133_));
 sg13g2_o21ai_1 _26033_ (.B1(net5545),
    .Y(_19056_),
    .A1(net1742),
    .A2(net4164));
 sg13g2_a22oi_1 _26034_ (.Y(_19057_),
    .B1(net4319),
    .B2(_18005_),
    .A2(net4276),
    .A1(_18510_));
 sg13g2_a22oi_1 _26035_ (.Y(_00013_),
    .B1(_19056_),
    .B2(_19057_),
    .A2(net4164),
    .A1(_14132_));
 sg13g2_o21ai_1 _26036_ (.B1(net5545),
    .Y(_19058_),
    .A1(net1690),
    .A2(net4169));
 sg13g2_a22oi_1 _26037_ (.Y(_19059_),
    .B1(net4319),
    .B2(_18510_),
    .A2(net4276),
    .A1(_18168_));
 sg13g2_a22oi_1 _26038_ (.Y(_00014_),
    .B1(_19058_),
    .B2(_19059_),
    .A2(net4169),
    .A1(_14131_));
 sg13g2_o21ai_1 _26039_ (.B1(net5552),
    .Y(_19060_),
    .A1(net1739),
    .A2(net4174));
 sg13g2_a22oi_1 _26040_ (.Y(_19061_),
    .B1(net4323),
    .B2(_18168_),
    .A2(net4278),
    .A1(_18011_));
 sg13g2_a22oi_1 _26041_ (.Y(_00015_),
    .B1(_19060_),
    .B2(_19061_),
    .A2(net4174),
    .A1(_14130_));
 sg13g2_o21ai_1 _26042_ (.B1(net5545),
    .Y(_19062_),
    .A1(net1797),
    .A2(net4169));
 sg13g2_a22oi_1 _26043_ (.Y(_19063_),
    .B1(net4323),
    .B2(_18011_),
    .A2(net4278),
    .A1(_17966_));
 sg13g2_a22oi_1 _26044_ (.Y(_00016_),
    .B1(_19062_),
    .B2(_19063_),
    .A2(net4164),
    .A1(_14129_));
 sg13g2_o21ai_1 _26045_ (.B1(net5552),
    .Y(_19064_),
    .A1(net1813),
    .A2(net4174));
 sg13g2_a22oi_1 _26046_ (.Y(_19065_),
    .B1(net4323),
    .B2(_17966_),
    .A2(net4278),
    .A1(_18475_));
 sg13g2_a22oi_1 _26047_ (.Y(_00017_),
    .B1(_19064_),
    .B2(_19065_),
    .A2(net4174),
    .A1(_14128_));
 sg13g2_o21ai_1 _26048_ (.B1(net5552),
    .Y(_19066_),
    .A1(net1672),
    .A2(net4174));
 sg13g2_a22oi_1 _26049_ (.Y(_19067_),
    .B1(net4323),
    .B2(_18475_),
    .A2(net4278),
    .A1(_18482_));
 sg13g2_a22oi_1 _26050_ (.Y(_00018_),
    .B1(_19066_),
    .B2(_19067_),
    .A2(net4174),
    .A1(_14127_));
 sg13g2_o21ai_1 _26051_ (.B1(net5552),
    .Y(_19068_),
    .A1(net1573),
    .A2(net4179));
 sg13g2_a22oi_1 _26052_ (.Y(_19069_),
    .B1(net4323),
    .B2(_18482_),
    .A2(net4278),
    .A1(_18204_));
 sg13g2_a22oi_1 _26053_ (.Y(_00019_),
    .B1(_19068_),
    .B2(_19069_),
    .A2(net4174),
    .A1(_14126_));
 sg13g2_o21ai_1 _26054_ (.B1(net5552),
    .Y(_19070_),
    .A1(net2187),
    .A2(net4174));
 sg13g2_a22oi_1 _26055_ (.Y(_19071_),
    .B1(net4323),
    .B2(_18204_),
    .A2(net4278),
    .A1(_18505_));
 sg13g2_a22oi_1 _26056_ (.Y(_00020_),
    .B1(_19070_),
    .B2(_19071_),
    .A2(net4179),
    .A1(_14125_));
 sg13g2_o21ai_1 _26057_ (.B1(net5552),
    .Y(_19072_),
    .A1(net1807),
    .A2(net4179));
 sg13g2_a22oi_1 _26058_ (.Y(_19073_),
    .B1(net4325),
    .B2(_18505_),
    .A2(net4280),
    .A1(_18186_));
 sg13g2_a22oi_1 _26059_ (.Y(_00021_),
    .B1(_19072_),
    .B2(_19073_),
    .A2(net4180),
    .A1(_14124_));
 sg13g2_o21ai_1 _26060_ (.B1(net5555),
    .Y(_19074_),
    .A1(net1750),
    .A2(net4180));
 sg13g2_a22oi_1 _26061_ (.Y(_19075_),
    .B1(net4325),
    .B2(_18186_),
    .A2(net4280),
    .A1(_17987_));
 sg13g2_a22oi_1 _26062_ (.Y(_00022_),
    .B1(_19074_),
    .B2(_19075_),
    .A2(net4180),
    .A1(_14123_));
 sg13g2_o21ai_1 _26063_ (.B1(net5555),
    .Y(_19076_),
    .A1(net1455),
    .A2(net4180));
 sg13g2_a22oi_1 _26064_ (.Y(_19077_),
    .B1(net4325),
    .B2(_17987_),
    .A2(net4280),
    .A1(_17906_));
 sg13g2_a22oi_1 _26065_ (.Y(_00023_),
    .B1(_19076_),
    .B2(_19077_),
    .A2(net4180),
    .A1(_14122_));
 sg13g2_o21ai_1 _26066_ (.B1(net5555),
    .Y(_19078_),
    .A1(net1663),
    .A2(net4180));
 sg13g2_a22oi_1 _26067_ (.Y(_19079_),
    .B1(net4325),
    .B2(_17906_),
    .A2(net4280),
    .A1(_18038_));
 sg13g2_a22oi_1 _26068_ (.Y(_00024_),
    .B1(_19078_),
    .B2(_19079_),
    .A2(net4181),
    .A1(_14121_));
 sg13g2_o21ai_1 _26069_ (.B1(net5555),
    .Y(_19080_),
    .A1(net1508),
    .A2(net4180));
 sg13g2_a22oi_1 _26070_ (.Y(_19081_),
    .B1(net4325),
    .B2(_18038_),
    .A2(net4280),
    .A1(_18180_));
 sg13g2_a22oi_1 _26071_ (.Y(_00025_),
    .B1(_19080_),
    .B2(_19081_),
    .A2(net4181),
    .A1(_14120_));
 sg13g2_o21ai_1 _26072_ (.B1(net5555),
    .Y(_19082_),
    .A1(net1483),
    .A2(net4180));
 sg13g2_a22oi_1 _26073_ (.Y(_19083_),
    .B1(net4325),
    .B2(_18180_),
    .A2(net4280),
    .A1(_18212_));
 sg13g2_a22oi_1 _26074_ (.Y(_00026_),
    .B1(_19082_),
    .B2(_19083_),
    .A2(net4181),
    .A1(_14119_));
 sg13g2_o21ai_1 _26075_ (.B1(net5555),
    .Y(_19084_),
    .A1(net2331),
    .A2(net4181));
 sg13g2_a22oi_1 _26076_ (.Y(_19085_),
    .B1(net4325),
    .B2(_18212_),
    .A2(net4280),
    .A1(_17994_));
 sg13g2_a22oi_1 _26077_ (.Y(_00027_),
    .B1(_19084_),
    .B2(_19085_),
    .A2(net4181),
    .A1(_14118_));
 sg13g2_o21ai_1 _26078_ (.B1(net5561),
    .Y(_19086_),
    .A1(net1699),
    .A2(net4196));
 sg13g2_a22oi_1 _26079_ (.Y(_19087_),
    .B1(net4329),
    .B2(_17994_),
    .A2(net4285),
    .A1(_17949_));
 sg13g2_a22oi_1 _26080_ (.Y(_00028_),
    .B1(_19086_),
    .B2(_19087_),
    .A2(net4196),
    .A1(_14117_));
 sg13g2_o21ai_1 _26081_ (.B1(net5561),
    .Y(_19088_),
    .A1(net1654),
    .A2(net4196));
 sg13g2_a22oi_1 _26082_ (.Y(_19089_),
    .B1(net4329),
    .B2(_17949_),
    .A2(net4285),
    .A1(_18196_));
 sg13g2_a22oi_1 _26083_ (.Y(_00029_),
    .B1(_19088_),
    .B2(_19089_),
    .A2(net4196),
    .A1(_14116_));
 sg13g2_o21ai_1 _26084_ (.B1(net5561),
    .Y(_19090_),
    .A1(net2240),
    .A2(net4195));
 sg13g2_a22oi_1 _26085_ (.Y(_19091_),
    .B1(net4329),
    .B2(_18196_),
    .A2(net4285),
    .A1(_18153_));
 sg13g2_a22oi_1 _26086_ (.Y(_00030_),
    .B1(_19090_),
    .B2(_19091_),
    .A2(net4195),
    .A1(_14115_));
 sg13g2_o21ai_1 _26087_ (.B1(net5561),
    .Y(_19092_),
    .A1(net1436),
    .A2(net4195));
 sg13g2_a22oi_1 _26088_ (.Y(_19093_),
    .B1(net4329),
    .B2(_18153_),
    .A2(net4285),
    .A1(_18135_));
 sg13g2_a22oi_1 _26089_ (.Y(_00031_),
    .B1(_19092_),
    .B2(_19093_),
    .A2(net4195),
    .A1(_14114_));
 sg13g2_o21ai_1 _26090_ (.B1(net5561),
    .Y(_19094_),
    .A1(net1538),
    .A2(net4195));
 sg13g2_a22oi_1 _26091_ (.Y(_19095_),
    .B1(net4329),
    .B2(_18135_),
    .A2(net4285),
    .A1(_18129_));
 sg13g2_a22oi_1 _26092_ (.Y(_00032_),
    .B1(_19094_),
    .B2(_19095_),
    .A2(net4195),
    .A1(_14113_));
 sg13g2_o21ai_1 _26093_ (.B1(net5563),
    .Y(_19096_),
    .A1(net1488),
    .A2(net4195));
 sg13g2_a22oi_1 _26094_ (.Y(_19097_),
    .B1(net4331),
    .B2(_18129_),
    .A2(net4286),
    .A1(_18191_));
 sg13g2_a22oi_1 _26095_ (.Y(_00033_),
    .B1(_19096_),
    .B2(_19097_),
    .A2(net4203),
    .A1(_14112_));
 sg13g2_o21ai_1 _26096_ (.B1(net5561),
    .Y(_19098_),
    .A1(net1457),
    .A2(net4195));
 sg13g2_a22oi_1 _26097_ (.Y(_19099_),
    .B1(net4329),
    .B2(_18191_),
    .A2(net4285),
    .A1(_17980_));
 sg13g2_a22oi_1 _26098_ (.Y(_00034_),
    .B1(_19098_),
    .B2(_19099_),
    .A2(net4196),
    .A1(_14111_));
 sg13g2_o21ai_1 _26099_ (.B1(net5563),
    .Y(_19100_),
    .A1(net1667),
    .A2(net4202));
 sg13g2_a22oi_1 _26100_ (.Y(_19101_),
    .B1(net4331),
    .B2(_17980_),
    .A2(net4286),
    .A1(_17912_));
 sg13g2_a22oi_1 _26101_ (.Y(_00035_),
    .B1(_19100_),
    .B2(_19101_),
    .A2(net4202),
    .A1(_14110_));
 sg13g2_o21ai_1 _26102_ (.B1(net5566),
    .Y(_19102_),
    .A1(net1542),
    .A2(net4202));
 sg13g2_a22oi_1 _26103_ (.Y(_19103_),
    .B1(net4331),
    .B2(_17912_),
    .A2(net4286),
    .A1(_17860_));
 sg13g2_a22oi_1 _26104_ (.Y(_00036_),
    .B1(_19102_),
    .B2(_19103_),
    .A2(net4202),
    .A1(_14109_));
 sg13g2_o21ai_1 _26105_ (.B1(net5566),
    .Y(_19104_),
    .A1(net1769),
    .A2(net4214));
 sg13g2_a22oi_1 _26106_ (.Y(_19105_),
    .B1(net4331),
    .B2(_17860_),
    .A2(net4286),
    .A1(_18147_));
 sg13g2_a22oi_1 _26107_ (.Y(_00037_),
    .B1(_19104_),
    .B2(_19105_),
    .A2(net4214),
    .A1(_14108_));
 sg13g2_o21ai_1 _26108_ (.B1(net5563),
    .Y(_19106_),
    .A1(net1802),
    .A2(net4202));
 sg13g2_a22oi_1 _26109_ (.Y(_19107_),
    .B1(net4331),
    .B2(_18147_),
    .A2(net4286),
    .A1(_18141_));
 sg13g2_a22oi_1 _26110_ (.Y(_00038_),
    .B1(_19106_),
    .B2(_19107_),
    .A2(net4202),
    .A1(_14107_));
 sg13g2_o21ai_1 _26111_ (.B1(net5563),
    .Y(_19108_),
    .A1(net2435),
    .A2(net4203));
 sg13g2_a22oi_1 _26112_ (.Y(_19109_),
    .B1(net4331),
    .B2(_18141_),
    .A2(net4286),
    .A1(_18528_));
 sg13g2_a22oi_1 _26113_ (.Y(_00039_),
    .B1(_19108_),
    .B2(_19109_),
    .A2(net4203),
    .A1(_14106_));
 sg13g2_o21ai_1 _26114_ (.B1(net5563),
    .Y(_19110_),
    .A1(net1547),
    .A2(net4202));
 sg13g2_a22oi_1 _26115_ (.Y(_19111_),
    .B1(net4333),
    .B2(_18528_),
    .A2(net4289),
    .A1(_18115_));
 sg13g2_a22oi_1 _26116_ (.Y(_00040_),
    .B1(_19110_),
    .B2(_19111_),
    .A2(net4202),
    .A1(_14105_));
 sg13g2_o21ai_1 _26117_ (.B1(net5565),
    .Y(_19112_),
    .A1(net1958),
    .A2(net4214));
 sg13g2_a22oi_1 _26118_ (.Y(_19113_),
    .B1(net4333),
    .B2(_18115_),
    .A2(net4289),
    .A1(_17972_));
 sg13g2_a22oi_1 _26119_ (.Y(_00041_),
    .B1(_19112_),
    .B2(_19113_),
    .A2(net4214),
    .A1(_14104_));
 sg13g2_o21ai_1 _26120_ (.B1(net5566),
    .Y(_19114_),
    .A1(net1514),
    .A2(net4214));
 sg13g2_a22oi_1 _26121_ (.Y(_19115_),
    .B1(net4333),
    .B2(_17972_),
    .A2(net4289),
    .A1(_18030_));
 sg13g2_a22oi_1 _26122_ (.Y(_00042_),
    .B1(_19114_),
    .B2(_19115_),
    .A2(net4214),
    .A1(_14103_));
 sg13g2_o21ai_1 _26123_ (.B1(net5566),
    .Y(_19116_),
    .A1(net1626),
    .A2(net4215));
 sg13g2_a22oi_1 _26124_ (.Y(_19117_),
    .B1(net4333),
    .B2(_18030_),
    .A2(net4289),
    .A1(_17879_));
 sg13g2_a22oi_1 _26125_ (.Y(_00043_),
    .B1(_19116_),
    .B2(_19117_),
    .A2(net4215),
    .A1(_14102_));
 sg13g2_o21ai_1 _26126_ (.B1(net5566),
    .Y(_19118_),
    .A1(net2079),
    .A2(net4215));
 sg13g2_a22oi_1 _26127_ (.Y(_19119_),
    .B1(net4333),
    .B2(_17879_),
    .A2(net4289),
    .A1(_18054_));
 sg13g2_a22oi_1 _26128_ (.Y(_00044_),
    .B1(_19118_),
    .B2(_19119_),
    .A2(net4214),
    .A1(_14101_));
 sg13g2_o21ai_1 _26129_ (.B1(net5566),
    .Y(_19120_),
    .A1(net1650),
    .A2(net4215));
 sg13g2_a22oi_1 _26130_ (.Y(_19121_),
    .B1(net4333),
    .B2(_18054_),
    .A2(net4289),
    .A1(_18022_));
 sg13g2_a22oi_1 _26131_ (.Y(_00045_),
    .B1(_19120_),
    .B2(_19121_),
    .A2(net4214),
    .A1(_14100_));
 sg13g2_o21ai_1 _26132_ (.B1(net5568),
    .Y(_19122_),
    .A1(net1591),
    .A2(net4223));
 sg13g2_a22oi_1 _26133_ (.Y(_19123_),
    .B1(net4335),
    .B2(_18022_),
    .A2(net4291),
    .A1(_18046_));
 sg13g2_a22oi_1 _26134_ (.Y(_00046_),
    .B1(_19122_),
    .B2(_19123_),
    .A2(net4219),
    .A1(_14099_));
 sg13g2_o21ai_1 _26135_ (.B1(net5568),
    .Y(_19124_),
    .A1(net1569),
    .A2(net4219));
 sg13g2_a22oi_1 _26136_ (.Y(_19125_),
    .B1(net4335),
    .B2(_18046_),
    .A2(net4291),
    .A1(_18062_));
 sg13g2_a22oi_1 _26137_ (.Y(_00047_),
    .B1(_19124_),
    .B2(_19125_),
    .A2(net4219),
    .A1(_14098_));
 sg13g2_o21ai_1 _26138_ (.B1(net5568),
    .Y(_19126_),
    .A1(net1562),
    .A2(net4219));
 sg13g2_a22oi_1 _26139_ (.Y(_19127_),
    .B1(net4335),
    .B2(_18062_),
    .A2(net4291),
    .A1(_18549_));
 sg13g2_a22oi_1 _26140_ (.Y(_00048_),
    .B1(_19126_),
    .B2(_19127_),
    .A2(net4219),
    .A1(_14097_));
 sg13g2_o21ai_1 _26141_ (.B1(net5568),
    .Y(_19128_),
    .A1(net1888),
    .A2(net4219));
 sg13g2_a22oi_1 _26142_ (.Y(_19129_),
    .B1(net4335),
    .B2(_18549_),
    .A2(net4291),
    .A1(_17919_));
 sg13g2_a22oi_1 _26143_ (.Y(_00049_),
    .B1(_19128_),
    .B2(_19129_),
    .A2(net4219),
    .A1(_14096_));
 sg13g2_o21ai_1 _26144_ (.B1(net5573),
    .Y(_19130_),
    .A1(net1461),
    .A2(net4219));
 sg13g2_a22oi_1 _26145_ (.Y(_19131_),
    .B1(net4337),
    .B2(_17919_),
    .A2(net4293),
    .A1(_17869_));
 sg13g2_a22oi_1 _26146_ (.Y(_00050_),
    .B1(_19130_),
    .B2(_19131_),
    .A2(net4223),
    .A1(_14095_));
 sg13g2_o21ai_1 _26147_ (.B1(net5574),
    .Y(_19132_),
    .A1(net1589),
    .A2(net4233));
 sg13g2_a22oi_1 _26148_ (.Y(_19133_),
    .B1(net4337),
    .B2(_17869_),
    .A2(net4293),
    .A1(_17839_));
 sg13g2_a22oi_1 _26149_ (.Y(_00051_),
    .B1(_19132_),
    .B2(_19133_),
    .A2(net4233),
    .A1(_14094_));
 sg13g2_o21ai_1 _26150_ (.B1(net5574),
    .Y(_19134_),
    .A1(net1578),
    .A2(net4233));
 sg13g2_a22oi_1 _26151_ (.Y(_19135_),
    .B1(net4337),
    .B2(_17839_),
    .A2(net4293),
    .A1(_18572_));
 sg13g2_a22oi_1 _26152_ (.Y(_00052_),
    .B1(_19134_),
    .B2(_19135_),
    .A2(net4233),
    .A1(_14093_));
 sg13g2_o21ai_1 _26153_ (.B1(net5574),
    .Y(_19136_),
    .A1(net1856),
    .A2(net4233));
 sg13g2_a22oi_1 _26154_ (.Y(_19137_),
    .B1(net4337),
    .B2(_18572_),
    .A2(net4293),
    .A1(_17888_));
 sg13g2_a22oi_1 _26155_ (.Y(_00053_),
    .B1(_19136_),
    .B2(_19137_),
    .A2(net4233),
    .A1(_14092_));
 sg13g2_o21ai_1 _26156_ (.B1(net5574),
    .Y(_19138_),
    .A1(net1522),
    .A2(net4233));
 sg13g2_a22oi_1 _26157_ (.Y(_19139_),
    .B1(net4337),
    .B2(_17888_),
    .A2(net4293),
    .A1(_18535_));
 sg13g2_a22oi_1 _26158_ (.Y(_00054_),
    .B1(_19138_),
    .B2(_19139_),
    .A2(net4233),
    .A1(_14091_));
 sg13g2_o21ai_1 _26159_ (.B1(net5577),
    .Y(_19140_),
    .A1(net2182),
    .A2(net4235));
 sg13g2_a22oi_1 _26160_ (.Y(_19141_),
    .B1(net4340),
    .B2(_18535_),
    .A2(net4296),
    .A1(_18100_));
 sg13g2_a22oi_1 _26161_ (.Y(_00055_),
    .B1(_19140_),
    .B2(_19141_),
    .A2(net4234),
    .A1(_14090_));
 sg13g2_o21ai_1 _26162_ (.B1(net5577),
    .Y(_19142_),
    .A1(net1907),
    .A2(net4235));
 sg13g2_a22oi_1 _26163_ (.Y(_19143_),
    .B1(net4340),
    .B2(_18100_),
    .A2(net4296),
    .A1(_18095_));
 sg13g2_a22oi_1 _26164_ (.Y(_00056_),
    .B1(_19142_),
    .B2(_19143_),
    .A2(net4234),
    .A1(_14089_));
 sg13g2_o21ai_1 _26165_ (.B1(net5577),
    .Y(_19144_),
    .A1(net1782),
    .A2(net4234));
 sg13g2_a22oi_1 _26166_ (.Y(_19145_),
    .B1(net4340),
    .B2(_18095_),
    .A2(net4296),
    .A1(_17828_));
 sg13g2_a22oi_1 _26167_ (.Y(_00057_),
    .B1(_19144_),
    .B2(_19145_),
    .A2(net4234),
    .A1(_14088_));
 sg13g2_o21ai_1 _26168_ (.B1(net5576),
    .Y(_19146_),
    .A1(net1575),
    .A2(net4234));
 sg13g2_a22oi_1 _26169_ (.Y(_19147_),
    .B1(net4345),
    .B2(_17828_),
    .A2(net4301),
    .A1(_17847_));
 sg13g2_a22oi_1 _26170_ (.Y(_00058_),
    .B1(_19146_),
    .B2(_19147_),
    .A2(net4234),
    .A1(_14087_));
 sg13g2_o21ai_1 _26171_ (.B1(net5582),
    .Y(_19148_),
    .A1(net1822),
    .A2(net4253));
 sg13g2_a22oi_1 _26172_ (.Y(_19149_),
    .B1(net4345),
    .B2(_17847_),
    .A2(net4301),
    .A1(_18071_));
 sg13g2_a22oi_1 _26173_ (.Y(_00059_),
    .B1(_19148_),
    .B2(_19149_),
    .A2(net4253),
    .A1(_14086_));
 sg13g2_o21ai_1 _26174_ (.B1(net5582),
    .Y(_19150_),
    .A1(net2077),
    .A2(net4253));
 sg13g2_a22oi_1 _26175_ (.Y(_19151_),
    .B1(net4345),
    .B2(_18071_),
    .A2(net4301),
    .A1(_18079_));
 sg13g2_a22oi_1 _26176_ (.Y(_00060_),
    .B1(_19150_),
    .B2(_19151_),
    .A2(net4253),
    .A1(_14085_));
 sg13g2_o21ai_1 _26177_ (.B1(net5582),
    .Y(_19152_),
    .A1(net1702),
    .A2(net4252));
 sg13g2_a22oi_1 _26178_ (.Y(_19153_),
    .B1(net4345),
    .B2(_18079_),
    .A2(net4301),
    .A1(_18586_));
 sg13g2_a22oi_1 _26179_ (.Y(_00061_),
    .B1(_19152_),
    .B2(_19153_),
    .A2(net4252),
    .A1(_14084_));
 sg13g2_o21ai_1 _26180_ (.B1(net5582),
    .Y(_19154_),
    .A1(net1599),
    .A2(net4253));
 sg13g2_a22oi_1 _26181_ (.Y(_19155_),
    .B1(net4345),
    .B2(_18586_),
    .A2(net4301),
    .A1(_17805_));
 sg13g2_a22oi_1 _26182_ (.Y(_00062_),
    .B1(_19154_),
    .B2(_19155_),
    .A2(net4257),
    .A1(_14083_));
 sg13g2_o21ai_1 _26183_ (.B1(net5582),
    .Y(_19156_),
    .A1(net1576),
    .A2(net4253));
 sg13g2_a22oi_1 _26184_ (.Y(_19157_),
    .B1(net4345),
    .B2(_17805_),
    .A2(net4301),
    .A1(_18607_));
 sg13g2_a22oi_1 _26185_ (.Y(_00063_),
    .B1(_19156_),
    .B2(_19157_),
    .A2(net4252),
    .A1(_14082_));
 sg13g2_o21ai_1 _26186_ (.B1(net5583),
    .Y(_19158_),
    .A1(net2314),
    .A2(net4253));
 sg13g2_a22oi_1 _26187_ (.Y(_19159_),
    .B1(net4345),
    .B2(_18607_),
    .A2(net4301),
    .A1(_17782_));
 sg13g2_a22oi_1 _26188_ (.Y(_00064_),
    .B1(_19158_),
    .B2(_19159_),
    .A2(net4252),
    .A1(_14081_));
 sg13g2_o21ai_1 _26189_ (.B1(net5584),
    .Y(_19160_),
    .A1(net1707),
    .A2(net4256));
 sg13g2_a22oi_1 _26190_ (.Y(_19161_),
    .B1(net4343),
    .B2(_17782_),
    .A2(net4299),
    .A1(_18563_));
 sg13g2_a22oi_1 _26191_ (.Y(_00065_),
    .B1(_19160_),
    .B2(_19161_),
    .A2(net4255),
    .A1(_14080_));
 sg13g2_o21ai_1 _26192_ (.B1(net5583),
    .Y(_19162_),
    .A1(net1494),
    .A2(net4254));
 sg13g2_a22oi_1 _26193_ (.Y(_19163_),
    .B1(net4344),
    .B2(_18563_),
    .A2(net4300),
    .A1(_18557_));
 sg13g2_a22oi_1 _26194_ (.Y(_00066_),
    .B1(_19162_),
    .B2(_19163_),
    .A2(net4256),
    .A1(_14079_));
 sg13g2_o21ai_1 _26195_ (.B1(net5584),
    .Y(_19164_),
    .A1(net1756),
    .A2(net4256));
 sg13g2_a22oi_1 _26196_ (.Y(_19165_),
    .B1(net4344),
    .B2(_18557_),
    .A2(net4300),
    .A1(_18579_));
 sg13g2_a22oi_1 _26197_ (.Y(_00067_),
    .B1(_19164_),
    .B2(_19165_),
    .A2(net4256),
    .A1(_14078_));
 sg13g2_o21ai_1 _26198_ (.B1(net5582),
    .Y(_19166_),
    .A1(net1728),
    .A2(net4252));
 sg13g2_a22oi_1 _26199_ (.Y(_19167_),
    .B1(net4344),
    .B2(_18579_),
    .A2(net4300),
    .A1(_17814_));
 sg13g2_a22oi_1 _26200_ (.Y(_00068_),
    .B1(_19166_),
    .B2(_19167_),
    .A2(net4255),
    .A1(_14077_));
 sg13g2_o21ai_1 _26201_ (.B1(net5583),
    .Y(_19168_),
    .A1(net2436),
    .A2(net4254));
 sg13g2_a22oi_1 _26202_ (.Y(_19169_),
    .B1(net4344),
    .B2(_17814_),
    .A2(net4300),
    .A1(_17787_));
 sg13g2_a22oi_1 _26203_ (.Y(_00069_),
    .B1(_19168_),
    .B2(_19169_),
    .A2(net4254),
    .A1(_14076_));
 sg13g2_o21ai_1 _26204_ (.B1(net5583),
    .Y(_19170_),
    .A1(net1512),
    .A2(net4254));
 sg13g2_a22oi_1 _26205_ (.Y(_19171_),
    .B1(net4343),
    .B2(_17787_),
    .A2(net4299),
    .A1(_18641_));
 sg13g2_a22oi_1 _26206_ (.Y(_00070_),
    .B1(_19170_),
    .B2(_19171_),
    .A2(net4255),
    .A1(_14075_));
 sg13g2_o21ai_1 _26207_ (.B1(net5584),
    .Y(_19172_),
    .A1(net2387),
    .A2(net4255));
 sg13g2_a22oi_1 _26208_ (.Y(_19173_),
    .B1(net4343),
    .B2(_18641_),
    .A2(net4299),
    .A1(_17745_));
 sg13g2_a22oi_1 _26209_ (.Y(_00071_),
    .B1(_19172_),
    .B2(_19173_),
    .A2(net4255),
    .A1(_14074_));
 sg13g2_o21ai_1 _26210_ (.B1(net5583),
    .Y(_19174_),
    .A1(net1879),
    .A2(net4254));
 sg13g2_a22oi_1 _26211_ (.Y(_19175_),
    .B1(net4343),
    .B2(_17745_),
    .A2(net4299),
    .A1(_17713_));
 sg13g2_a22oi_1 _26212_ (.Y(_00072_),
    .B1(_19174_),
    .B2(_19175_),
    .A2(net4254),
    .A1(_14073_));
 sg13g2_o21ai_1 _26213_ (.B1(net5583),
    .Y(_19176_),
    .A1(net1984),
    .A2(net4255));
 sg13g2_a22oi_1 _26214_ (.Y(_19177_),
    .B1(net4343),
    .B2(_17713_),
    .A2(net4299),
    .A1(_18541_));
 sg13g2_a22oi_1 _26215_ (.Y(_00073_),
    .B1(_19176_),
    .B2(_19177_),
    .A2(net4254),
    .A1(_14072_));
 sg13g2_o21ai_1 _26216_ (.B1(net5583),
    .Y(_19178_),
    .A1(net1485),
    .A2(net4255));
 sg13g2_a22oi_1 _26217_ (.Y(_19179_),
    .B1(net4343),
    .B2(_18541_),
    .A2(net4299),
    .A1(_17822_));
 sg13g2_a22oi_1 _26218_ (.Y(_00074_),
    .B1(_19178_),
    .B2(_19179_),
    .A2(net4254),
    .A1(_14071_));
 sg13g2_o21ai_1 _26219_ (.B1(net5580),
    .Y(_19180_),
    .A1(net1930),
    .A2(net4250));
 sg13g2_a22oi_1 _26220_ (.Y(_19181_),
    .B1(net4341),
    .B2(_17822_),
    .A2(net4297),
    .A1(_18594_));
 sg13g2_a22oi_1 _26221_ (.Y(_00075_),
    .B1(_19180_),
    .B2(_19181_),
    .A2(net4250),
    .A1(_14070_));
 sg13g2_o21ai_1 _26222_ (.B1(net5580),
    .Y(_19182_),
    .A1(net2015),
    .A2(net4250));
 sg13g2_a22oi_1 _26223_ (.Y(_19183_),
    .B1(net4342),
    .B2(_18594_),
    .A2(net4298),
    .A1(_17762_));
 sg13g2_a22oi_1 _26224_ (.Y(_00076_),
    .B1(_19182_),
    .B2(_19183_),
    .A2(net4250),
    .A1(_14069_));
 sg13g2_o21ai_1 _26225_ (.B1(net5583),
    .Y(_19184_),
    .A1(net1633),
    .A2(net4250));
 sg13g2_a22oi_1 _26226_ (.Y(_19185_),
    .B1(net4343),
    .B2(_17762_),
    .A2(net4299),
    .A1(_17796_));
 sg13g2_a22oi_1 _26227_ (.Y(_00077_),
    .B1(_19184_),
    .B2(_19185_),
    .A2(net4250),
    .A1(_14068_));
 sg13g2_o21ai_1 _26228_ (.B1(net5581),
    .Y(_19186_),
    .A1(net1447),
    .A2(net4250));
 sg13g2_a22oi_1 _26229_ (.Y(_19187_),
    .B1(net4343),
    .B2(_17796_),
    .A2(net4299),
    .A1(_18601_));
 sg13g2_a22oi_1 _26230_ (.Y(_00078_),
    .B1(_19186_),
    .B2(_19187_),
    .A2(net4251),
    .A1(_14067_));
 sg13g2_o21ai_1 _26231_ (.B1(net5581),
    .Y(_19188_),
    .A1(net1805),
    .A2(net4250));
 sg13g2_a22oi_1 _26232_ (.Y(_19189_),
    .B1(net4341),
    .B2(_18601_),
    .A2(net4297),
    .A1(_17751_));
 sg13g2_a22oi_1 _26233_ (.Y(_00079_),
    .B1(_19188_),
    .B2(_19189_),
    .A2(net4251),
    .A1(_14066_));
 sg13g2_o21ai_1 _26234_ (.B1(net5580),
    .Y(_19190_),
    .A1(net1717),
    .A2(net4248));
 sg13g2_a22oi_1 _26235_ (.Y(_19191_),
    .B1(net4341),
    .B2(_17751_),
    .A2(net4297),
    .A1(_17640_));
 sg13g2_a22oi_1 _26236_ (.Y(_00080_),
    .B1(_19190_),
    .B2(_19191_),
    .A2(net4249),
    .A1(_14065_));
 sg13g2_o21ai_1 _26237_ (.B1(net5580),
    .Y(_19192_),
    .A1(net1917),
    .A2(net4248));
 sg13g2_a22oi_1 _26238_ (.Y(_19193_),
    .B1(net4342),
    .B2(_17640_),
    .A2(net4298),
    .A1(_17791_));
 sg13g2_a22oi_1 _26239_ (.Y(_00081_),
    .B1(_19192_),
    .B2(_19193_),
    .A2(net4249),
    .A1(_14064_));
 sg13g2_o21ai_1 _26240_ (.B1(net5581),
    .Y(_19194_),
    .A1(net1549),
    .A2(net4248));
 sg13g2_a22oi_1 _26241_ (.Y(_19195_),
    .B1(net4342),
    .B2(_17791_),
    .A2(net4298),
    .A1(_18649_));
 sg13g2_a22oi_1 _26242_ (.Y(_00082_),
    .B1(_19194_),
    .B2(_19195_),
    .A2(net4249),
    .A1(_14063_));
 sg13g2_o21ai_1 _26243_ (.B1(net5580),
    .Y(_19196_),
    .A1(net1913),
    .A2(net4248));
 sg13g2_a22oi_1 _26244_ (.Y(_19197_),
    .B1(net4341),
    .B2(_18649_),
    .A2(net4297),
    .A1(_18620_));
 sg13g2_a22oi_1 _26245_ (.Y(_00083_),
    .B1(_19196_),
    .B2(_19197_),
    .A2(net4248),
    .A1(_14062_));
 sg13g2_o21ai_1 _26246_ (.B1(net5580),
    .Y(_19198_),
    .A1(net1892),
    .A2(net4248));
 sg13g2_a22oi_1 _26247_ (.Y(_19199_),
    .B1(net4341),
    .B2(_18620_),
    .A2(net4297),
    .A1(_17665_));
 sg13g2_a22oi_1 _26248_ (.Y(_00084_),
    .B1(_19198_),
    .B2(_19199_),
    .A2(net4248),
    .A1(_14061_));
 sg13g2_o21ai_1 _26249_ (.B1(net5580),
    .Y(_19200_),
    .A1(net1531),
    .A2(net4248));
 sg13g2_a22oi_1 _26250_ (.Y(_19201_),
    .B1(net4341),
    .B2(_17665_),
    .A2(net4297),
    .A1(_18613_));
 sg13g2_a22oi_1 _26251_ (.Y(_00085_),
    .B1(_19200_),
    .B2(_19201_),
    .A2(net4249),
    .A1(_14060_));
 sg13g2_o21ai_1 _26252_ (.B1(net5580),
    .Y(_19202_),
    .A1(net1527),
    .A2(net4238));
 sg13g2_a22oi_1 _26253_ (.Y(_19203_),
    .B1(net4341),
    .B2(_18613_),
    .A2(net4297),
    .A1(_18672_));
 sg13g2_a22oi_1 _26254_ (.Y(_00086_),
    .B1(_19202_),
    .B2(_19203_),
    .A2(net4238),
    .A1(_14059_));
 sg13g2_o21ai_1 _26255_ (.B1(net5576),
    .Y(_19204_),
    .A1(net1632),
    .A2(net4238));
 sg13g2_a22oi_1 _26256_ (.Y(_19205_),
    .B1(net4341),
    .B2(_18672_),
    .A2(net4297),
    .A1(_17599_));
 sg13g2_a22oi_1 _26257_ (.Y(_00087_),
    .B1(_19204_),
    .B2(_19205_),
    .A2(net4238),
    .A1(_14058_));
 sg13g2_o21ai_1 _26258_ (.B1(net5575),
    .Y(_19206_),
    .A1(net2157),
    .A2(net4238));
 sg13g2_a22oi_1 _26259_ (.Y(_19207_),
    .B1(net4340),
    .B2(_17599_),
    .A2(net4295),
    .A1(_17495_));
 sg13g2_a22oi_1 _26260_ (.Y(_00088_),
    .B1(_19206_),
    .B2(_19207_),
    .A2(net4238),
    .A1(_14057_));
 sg13g2_o21ai_1 _26261_ (.B1(net5575),
    .Y(_19208_),
    .A1(net2283),
    .A2(net4238));
 sg13g2_a22oi_1 _26262_ (.Y(_19209_),
    .B1(net4339),
    .B2(_17495_),
    .A2(net4296),
    .A1(_18627_));
 sg13g2_a22oi_1 _26263_ (.Y(_00089_),
    .B1(_19208_),
    .B2(_19209_),
    .A2(net4239),
    .A1(_14056_));
 sg13g2_o21ai_1 _26264_ (.B1(net5576),
    .Y(_19210_),
    .A1(net1646),
    .A2(net4238));
 sg13g2_a22oi_1 _26265_ (.Y(_19211_),
    .B1(net4340),
    .B2(_18627_),
    .A2(net4296),
    .A1(_18680_));
 sg13g2_a22oi_1 _26266_ (.Y(_00090_),
    .B1(_19210_),
    .B2(_19211_),
    .A2(net4239),
    .A1(_14055_));
 sg13g2_o21ai_1 _26267_ (.B1(net5576),
    .Y(_19212_),
    .A1(net1855),
    .A2(net4236));
 sg13g2_a22oi_1 _26268_ (.Y(_19213_),
    .B1(net4339),
    .B2(_18680_),
    .A2(net4295),
    .A1(_17645_));
 sg13g2_a22oi_1 _26269_ (.Y(_00091_),
    .B1(_19212_),
    .B2(_19213_),
    .A2(net4239),
    .A1(_14054_));
 sg13g2_o21ai_1 _26270_ (.B1(net5575),
    .Y(_19214_),
    .A1(net1681),
    .A2(net4236));
 sg13g2_a22oi_1 _26271_ (.Y(_19215_),
    .B1(net4339),
    .B2(_17645_),
    .A2(net4295),
    .A1(_17511_));
 sg13g2_a22oi_1 _26272_ (.Y(_00092_),
    .B1(_19214_),
    .B2(_19215_),
    .A2(net4236),
    .A1(_14053_));
 sg13g2_o21ai_1 _26273_ (.B1(net5575),
    .Y(_19216_),
    .A1(net1974),
    .A2(net4236));
 sg13g2_a22oi_1 _26274_ (.Y(_19217_),
    .B1(net4339),
    .B2(_17511_),
    .A2(net4295),
    .A1(_18654_));
 sg13g2_a22oi_1 _26275_ (.Y(_00093_),
    .B1(_19216_),
    .B2(_19217_),
    .A2(net4237),
    .A1(_14052_));
 sg13g2_o21ai_1 _26276_ (.B1(net5575),
    .Y(_19218_),
    .A1(net1912),
    .A2(net4236));
 sg13g2_a22oi_1 _26277_ (.Y(_19219_),
    .B1(net4339),
    .B2(_18654_),
    .A2(net4295),
    .A1(_17619_));
 sg13g2_a22oi_1 _26278_ (.Y(_00094_),
    .B1(_19218_),
    .B2(_19219_),
    .A2(net4237),
    .A1(_14051_));
 sg13g2_o21ai_1 _26279_ (.B1(net5575),
    .Y(_19220_),
    .A1(net2085),
    .A2(net4236));
 sg13g2_a22oi_1 _26280_ (.Y(_19221_),
    .B1(net4339),
    .B2(_17619_),
    .A2(net4295),
    .A1(_17682_));
 sg13g2_a22oi_1 _26281_ (.Y(_00095_),
    .B1(_19220_),
    .B2(_19221_),
    .A2(net4236),
    .A1(_14050_));
 sg13g2_o21ai_1 _26282_ (.B1(net5575),
    .Y(_19222_),
    .A1(net2064),
    .A2(net4236));
 sg13g2_a22oi_1 _26283_ (.Y(_19223_),
    .B1(net4339),
    .B2(_17682_),
    .A2(net4295),
    .A1(_18785_));
 sg13g2_a22oi_1 _26284_ (.Y(_00096_),
    .B1(_19222_),
    .B2(_19223_),
    .A2(net4237),
    .A1(_14049_));
 sg13g2_o21ai_1 _26285_ (.B1(net5575),
    .Y(_19224_),
    .A1(net2191),
    .A2(net4231));
 sg13g2_a22oi_1 _26286_ (.Y(_19225_),
    .B1(net4339),
    .B2(_18785_),
    .A2(net4295),
    .A1(_18632_));
 sg13g2_a22oi_1 _26287_ (.Y(_00097_),
    .B1(_19224_),
    .B2(_19225_),
    .A2(net4237),
    .A1(_14048_));
 sg13g2_o21ai_1 _26288_ (.B1(net5573),
    .Y(_19226_),
    .A1(net1884),
    .A2(net4231));
 sg13g2_nor2_1 _26289_ (.A(_18694_),
    .B(net4349),
    .Y(_19227_));
 sg13g2_a21oi_1 _26290_ (.A1(_18632_),
    .A2(net4337),
    .Y(_19228_),
    .B1(_19227_));
 sg13g2_a22oi_1 _26291_ (.Y(_00098_),
    .B1(_19226_),
    .B2(_19228_),
    .A2(net4231),
    .A1(_14047_));
 sg13g2_o21ai_1 _26292_ (.B1(net5573),
    .Y(_19229_),
    .A1(net1686),
    .A2(net4231));
 sg13g2_nor2_1 _26293_ (.A(_18694_),
    .B(net4260),
    .Y(_19230_));
 sg13g2_a21oi_1 _26294_ (.A1(_17688_),
    .A2(net4293),
    .Y(_19231_),
    .B1(_19230_));
 sg13g2_a22oi_1 _26295_ (.Y(_00099_),
    .B1(_19229_),
    .B2(_19231_),
    .A2(net4231),
    .A1(_14046_));
 sg13g2_o21ai_1 _26296_ (.B1(net5574),
    .Y(_19232_),
    .A1(net1715),
    .A2(net4231));
 sg13g2_a22oi_1 _26297_ (.Y(_19233_),
    .B1(net4337),
    .B2(_17688_),
    .A2(net4293),
    .A1(_17548_));
 sg13g2_a22oi_1 _26298_ (.Y(_00100_),
    .B1(_19232_),
    .B2(_19233_),
    .A2(net4231),
    .A1(_14045_));
 sg13g2_o21ai_1 _26299_ (.B1(net5574),
    .Y(_19234_),
    .A1(net1622),
    .A2(net4231));
 sg13g2_a22oi_1 _26300_ (.Y(_19235_),
    .B1(net4337),
    .B2(_17548_),
    .A2(net4293),
    .A1(_18665_));
 sg13g2_a22oi_1 _26301_ (.Y(_00101_),
    .B1(_19234_),
    .B2(_19235_),
    .A2(net4232),
    .A1(_14044_));
 sg13g2_o21ai_1 _26302_ (.B1(net5573),
    .Y(_19236_),
    .A1(net2067),
    .A2(net4230));
 sg13g2_a22oi_1 _26303_ (.Y(_19237_),
    .B1(net4338),
    .B2(_18665_),
    .A2(net4294),
    .A1(_18729_));
 sg13g2_a22oi_1 _26304_ (.Y(_00102_),
    .B1(_19236_),
    .B2(_19237_),
    .A2(net4230),
    .A1(_14043_));
 sg13g2_o21ai_1 _26305_ (.B1(net5573),
    .Y(_19238_),
    .A1(net1587),
    .A2(net4230));
 sg13g2_a22oi_1 _26306_ (.Y(_19239_),
    .B1(net4338),
    .B2(_18729_),
    .A2(net4294),
    .A1(_17726_));
 sg13g2_a22oi_1 _26307_ (.Y(_00103_),
    .B1(_19238_),
    .B2(_19239_),
    .A2(net4232),
    .A1(_14042_));
 sg13g2_o21ai_1 _26308_ (.B1(net5573),
    .Y(_19240_),
    .A1(net1693),
    .A2(net4230));
 sg13g2_a22oi_1 _26309_ (.Y(_19241_),
    .B1(net4338),
    .B2(_17726_),
    .A2(net4294),
    .A1(_17321_));
 sg13g2_a22oi_1 _26310_ (.Y(_00104_),
    .B1(_19240_),
    .B2(_19241_),
    .A2(net4230),
    .A1(_14041_));
 sg13g2_o21ai_1 _26311_ (.B1(net5573),
    .Y(_19242_),
    .A1(net1475),
    .A2(net4230));
 sg13g2_a22oi_1 _26312_ (.Y(_19243_),
    .B1(net4338),
    .B2(_17321_),
    .A2(net4294),
    .A1(_18659_));
 sg13g2_a22oi_1 _26313_ (.Y(_00105_),
    .B1(_19242_),
    .B2(_19243_),
    .A2(net4230),
    .A1(_14040_));
 sg13g2_o21ai_1 _26314_ (.B1(net5573),
    .Y(_19244_),
    .A1(net1665),
    .A2(net4230));
 sg13g2_nor2_1 _26315_ (.A(_17653_),
    .B(net4349),
    .Y(_19245_));
 sg13g2_a21oi_1 _26316_ (.A1(_18659_),
    .A2(net4338),
    .Y(_19246_),
    .B1(_19245_));
 sg13g2_a22oi_1 _26317_ (.Y(_00106_),
    .B1(_19244_),
    .B2(_19246_),
    .A2(net4232),
    .A1(_14039_));
 sg13g2_o21ai_1 _26318_ (.B1(net5567),
    .Y(_19247_),
    .A1(net2135),
    .A2(net4221));
 sg13g2_nor2_1 _26319_ (.A(_17653_),
    .B(net4260),
    .Y(_19248_));
 sg13g2_a21oi_1 _26320_ (.A1(_17520_),
    .A2(net4290),
    .Y(_19249_),
    .B1(_19248_));
 sg13g2_a22oi_1 _26321_ (.Y(_00107_),
    .B1(_19247_),
    .B2(_19249_),
    .A2(net4221),
    .A1(_14038_));
 sg13g2_o21ai_1 _26322_ (.B1(net5567),
    .Y(_19250_),
    .A1(net1556),
    .A2(net4221));
 sg13g2_a22oi_1 _26323_ (.Y(_19251_),
    .B1(net4334),
    .B2(_17520_),
    .A2(net4291),
    .A1(_18754_));
 sg13g2_a22oi_1 _26324_ (.Y(_00108_),
    .B1(_19250_),
    .B2(_19251_),
    .A2(net4221),
    .A1(_14037_));
 sg13g2_o21ai_1 _26325_ (.B1(net5567),
    .Y(_19252_),
    .A1(net1803),
    .A2(net4220));
 sg13g2_a22oi_1 _26326_ (.Y(_19253_),
    .B1(net4335),
    .B2(_18754_),
    .A2(net4291),
    .A1(_17671_));
 sg13g2_a22oi_1 _26327_ (.Y(_00109_),
    .B1(_19252_),
    .B2(_19253_),
    .A2(net4220),
    .A1(_14036_));
 sg13g2_o21ai_1 _26328_ (.B1(net5568),
    .Y(_19254_),
    .A1(net1506),
    .A2(net4221));
 sg13g2_nor2_1 _26329_ (.A(_17469_),
    .B(net4349),
    .Y(_19255_));
 sg13g2_a21oi_1 _26330_ (.A1(_17671_),
    .A2(net4334),
    .Y(_19256_),
    .B1(_19255_));
 sg13g2_a22oi_1 _26331_ (.Y(_00110_),
    .B1(_19254_),
    .B2(_19256_),
    .A2(net4221),
    .A1(_14035_));
 sg13g2_o21ai_1 _26332_ (.B1(net5567),
    .Y(_19257_),
    .A1(net2025),
    .A2(net4222));
 sg13g2_nor2_1 _26333_ (.A(_17469_),
    .B(_19032_),
    .Y(_19258_));
 sg13g2_a21oi_1 _26334_ (.A1(_18735_),
    .A2(net4290),
    .Y(_19259_),
    .B1(_19258_));
 sg13g2_a22oi_1 _26335_ (.Y(_00111_),
    .B1(_19257_),
    .B2(_19259_),
    .A2(net4222),
    .A1(_14034_));
 sg13g2_o21ai_1 _26336_ (.B1(net5568),
    .Y(_19260_),
    .A1(net2090),
    .A2(net4221));
 sg13g2_a22oi_1 _26337_ (.Y(_19261_),
    .B1(net4334),
    .B2(_18735_),
    .A2(net4290),
    .A1(_17235_));
 sg13g2_a22oi_1 _26338_ (.Y(_00112_),
    .B1(_19260_),
    .B2(_19261_),
    .A2(net4222),
    .A1(_14033_));
 sg13g2_o21ai_1 _26339_ (.B1(net5567),
    .Y(_19262_),
    .A1(net2263),
    .A2(net4220));
 sg13g2_a22oi_1 _26340_ (.Y(_19263_),
    .B1(net4334),
    .B2(_17235_),
    .A2(net4290),
    .A1(_18687_));
 sg13g2_a22oi_1 _26341_ (.Y(_00113_),
    .B1(_19262_),
    .B2(_19263_),
    .A2(net4220),
    .A1(_14032_));
 sg13g2_o21ai_1 _26342_ (.B1(net5567),
    .Y(_19264_),
    .A1(net1652),
    .A2(net4220));
 sg13g2_a22oi_1 _26343_ (.Y(_19265_),
    .B1(net4334),
    .B2(_18687_),
    .A2(net4290),
    .A1(_18703_));
 sg13g2_a22oi_1 _26344_ (.Y(_00114_),
    .B1(_19264_),
    .B2(_19265_),
    .A2(net4220),
    .A1(_14031_));
 sg13g2_o21ai_1 _26345_ (.B1(net5568),
    .Y(_19266_),
    .A1(net1883),
    .A2(net4221));
 sg13g2_a22oi_1 _26346_ (.Y(_19267_),
    .B1(net4334),
    .B2(_18703_),
    .A2(net4290),
    .A1(_17606_));
 sg13g2_a22oi_1 _26347_ (.Y(_00115_),
    .B1(_19266_),
    .B2(_19267_),
    .A2(net4220),
    .A1(_14030_));
 sg13g2_o21ai_1 _26348_ (.B1(net5565),
    .Y(_19268_),
    .A1(net1861),
    .A2(net4216));
 sg13g2_a22oi_1 _26349_ (.Y(_19269_),
    .B1(net4334),
    .B2(_17606_),
    .A2(net4290),
    .A1(_17531_));
 sg13g2_a22oi_1 _26350_ (.Y(_00116_),
    .B1(_19268_),
    .B2(_19269_),
    .A2(net4216),
    .A1(_14029_));
 sg13g2_o21ai_1 _26351_ (.B1(net5565),
    .Y(_19270_),
    .A1(net2014),
    .A2(net4216));
 sg13g2_a22oi_1 _26352_ (.Y(_19271_),
    .B1(net4334),
    .B2(_17531_),
    .A2(net4290),
    .A1(_17694_));
 sg13g2_a22oi_1 _26353_ (.Y(_00117_),
    .B1(_19270_),
    .B2(_19271_),
    .A2(net4218),
    .A1(_14028_));
 sg13g2_o21ai_1 _26354_ (.B1(net5567),
    .Y(_19272_),
    .A1(net1776),
    .A2(net4222));
 sg13g2_a22oi_1 _26355_ (.Y(_19273_),
    .B1(net4332),
    .B2(_17694_),
    .A2(net4288),
    .A1(_17476_));
 sg13g2_a22oi_1 _26356_ (.Y(_00118_),
    .B1(_19272_),
    .B2(_19273_),
    .A2(net4218),
    .A1(_14027_));
 sg13g2_o21ai_1 _26357_ (.B1(net5567),
    .Y(_19274_),
    .A1(net1759),
    .A2(net4220));
 sg13g2_a22oi_1 _26358_ (.Y(_19275_),
    .B1(net4332),
    .B2(_17476_),
    .A2(net4288),
    .A1(_18794_));
 sg13g2_a22oi_1 _26359_ (.Y(_00119_),
    .B1(_19274_),
    .B2(_19275_),
    .A2(net4216),
    .A1(_14026_));
 sg13g2_o21ai_1 _26360_ (.B1(net5565),
    .Y(_19276_),
    .A1(net2046),
    .A2(net4216));
 sg13g2_a22oi_1 _26361_ (.Y(_19277_),
    .B1(net4332),
    .B2(_18794_),
    .A2(net4288),
    .A1(_17207_));
 sg13g2_a22oi_1 _26362_ (.Y(_00120_),
    .B1(_19276_),
    .B2(_19277_),
    .A2(net4216),
    .A1(_14025_));
 sg13g2_o21ai_1 _26363_ (.B1(net5565),
    .Y(_19278_),
    .A1(net1851),
    .A2(net4217));
 sg13g2_a22oi_1 _26364_ (.Y(_19279_),
    .B1(net4332),
    .B2(_17207_),
    .A2(net4289),
    .A1(_17561_));
 sg13g2_a22oi_1 _26365_ (.Y(_00121_),
    .B1(_19278_),
    .B2(_19279_),
    .A2(net4217),
    .A1(_14024_));
 sg13g2_o21ai_1 _26366_ (.B1(net5565),
    .Y(_19280_),
    .A1(net1932),
    .A2(net4216));
 sg13g2_a22oi_1 _26367_ (.Y(_19281_),
    .B1(net4332),
    .B2(_17561_),
    .A2(net4288),
    .A1(_17555_));
 sg13g2_a22oi_1 _26368_ (.Y(_00122_),
    .B1(_19280_),
    .B2(_19281_),
    .A2(net4217),
    .A1(_14023_));
 sg13g2_o21ai_1 _26369_ (.B1(net5565),
    .Y(_19282_),
    .A1(net2376),
    .A2(net4216));
 sg13g2_a22oi_1 _26370_ (.Y(_19283_),
    .B1(net4333),
    .B2(_17555_),
    .A2(net4288),
    .A1(_17536_));
 sg13g2_a22oi_1 _26371_ (.Y(_00123_),
    .B1(_19282_),
    .B2(_19283_),
    .A2(net4218),
    .A1(_14022_));
 sg13g2_o21ai_1 _26372_ (.B1(net5566),
    .Y(_19284_),
    .A1(net1859),
    .A2(net4217));
 sg13g2_a22oi_1 _26373_ (.Y(_19285_),
    .B1(net4332),
    .B2(_17536_),
    .A2(net4288),
    .A1(_17254_));
 sg13g2_a22oi_1 _26374_ (.Y(_00124_),
    .B1(_19284_),
    .B2(_19285_),
    .A2(net4217),
    .A1(_14021_));
 sg13g2_o21ai_1 _26375_ (.B1(net5563),
    .Y(_19286_),
    .A1(net1886),
    .A2(net4205));
 sg13g2_a22oi_1 _26376_ (.Y(_19287_),
    .B1(net4330),
    .B2(_17254_),
    .A2(net4287),
    .A1(_17087_));
 sg13g2_a22oi_1 _26377_ (.Y(_00125_),
    .B1(_19286_),
    .B2(_19287_),
    .A2(net4204),
    .A1(_14020_));
 sg13g2_o21ai_1 _26378_ (.B1(net5565),
    .Y(_19288_),
    .A1(net1459),
    .A2(net4217));
 sg13g2_a22oi_1 _26379_ (.Y(_19289_),
    .B1(net4330),
    .B2(_17087_),
    .A2(net4287),
    .A1(_17361_));
 sg13g2_a22oi_1 _26380_ (.Y(_00126_),
    .B1(_19288_),
    .B2(_19289_),
    .A2(net4204),
    .A1(_14019_));
 sg13g2_o21ai_1 _26381_ (.B1(net5562),
    .Y(_19290_),
    .A1(net1816),
    .A2(net4205));
 sg13g2_a22oi_1 _26382_ (.Y(_19291_),
    .B1(net4330),
    .B2(_17361_),
    .A2(net4287),
    .A1(_17118_));
 sg13g2_a22oi_1 _26383_ (.Y(_00127_),
    .B1(_19290_),
    .B2(_19291_),
    .A2(net4205),
    .A1(_14018_));
 sg13g2_o21ai_1 _26384_ (.B1(net5562),
    .Y(_19292_),
    .A1(net2166),
    .A2(net4204));
 sg13g2_a22oi_1 _26385_ (.Y(_19293_),
    .B1(net4331),
    .B2(_17118_),
    .A2(net4286),
    .A1(_18802_));
 sg13g2_a22oi_1 _26386_ (.Y(_00128_),
    .B1(_19292_),
    .B2(_19293_),
    .A2(net4204),
    .A1(_14017_));
 sg13g2_o21ai_1 _26387_ (.B1(net5563),
    .Y(_19294_),
    .A1(net1940),
    .A2(net4204));
 sg13g2_a22oi_1 _26388_ (.Y(_19295_),
    .B1(net4330),
    .B2(_18802_),
    .A2(net4286),
    .A1(_18713_));
 sg13g2_a22oi_1 _26389_ (.Y(_00129_),
    .B1(_19294_),
    .B2(_19295_),
    .A2(net4204),
    .A1(_14016_));
 sg13g2_o21ai_1 _26390_ (.B1(net5562),
    .Y(_19296_),
    .A1(net1689),
    .A2(net4205));
 sg13g2_a22oi_1 _26391_ (.Y(_19297_),
    .B1(net4332),
    .B2(_18713_),
    .A2(net4288),
    .A1(_18722_));
 sg13g2_a22oi_1 _26392_ (.Y(_00130_),
    .B1(_19296_),
    .B2(_19297_),
    .A2(net4217),
    .A1(_14015_));
 sg13g2_o21ai_1 _26393_ (.B1(net5562),
    .Y(_19298_),
    .A1(net1595),
    .A2(net4204));
 sg13g2_a22oi_1 _26394_ (.Y(_19299_),
    .B1(net4332),
    .B2(_18722_),
    .A2(net4288),
    .A1(_17719_));
 sg13g2_a22oi_1 _26395_ (.Y(_00131_),
    .B1(_19298_),
    .B2(_19299_),
    .A2(net4204),
    .A1(_14014_));
 sg13g2_o21ai_1 _26396_ (.B1(net5562),
    .Y(_19300_),
    .A1(net1620),
    .A2(net4206));
 sg13g2_a22oi_1 _26397_ (.Y(_19301_),
    .B1(net4330),
    .B2(_17719_),
    .A2(net4287),
    .A1(_17585_));
 sg13g2_a22oi_1 _26398_ (.Y(_00132_),
    .B1(_19300_),
    .B2(_19301_),
    .A2(net4206),
    .A1(_14013_));
 sg13g2_o21ai_1 _26399_ (.B1(net5562),
    .Y(_19302_),
    .A1(net1935),
    .A2(net4206));
 sg13g2_a22oi_1 _26400_ (.Y(_19303_),
    .B1(net4330),
    .B2(_17585_),
    .A2(net4287),
    .A1(_18708_));
 sg13g2_a22oi_1 _26401_ (.Y(_00133_),
    .B1(_19302_),
    .B2(_19303_),
    .A2(net4206),
    .A1(_14012_));
 sg13g2_o21ai_1 _26402_ (.B1(net5562),
    .Y(_19304_),
    .A1(net1897),
    .A2(net4206));
 sg13g2_nor2_1 _26403_ (.A(_17307_),
    .B(net4349),
    .Y(_19305_));
 sg13g2_a21oi_1 _26404_ (.A1(_18708_),
    .A2(net4330),
    .Y(_19306_),
    .B1(_19305_));
 sg13g2_a22oi_1 _26405_ (.Y(_00134_),
    .B1(_19304_),
    .B2(_19306_),
    .A2(net4206),
    .A1(_14011_));
 sg13g2_o21ai_1 _26406_ (.B1(net5560),
    .Y(_19307_),
    .A1(net1607),
    .A2(net4199));
 sg13g2_nor2_1 _26407_ (.A(_17307_),
    .B(_19032_),
    .Y(_19308_));
 sg13g2_a21oi_1 _26408_ (.A1(_17374_),
    .A2(net4284),
    .Y(_19309_),
    .B1(_19308_));
 sg13g2_a22oi_1 _26409_ (.Y(_00135_),
    .B1(_19307_),
    .B2(_19309_),
    .A2(net4199),
    .A1(_14010_));
 sg13g2_o21ai_1 _26410_ (.B1(net5560),
    .Y(_19310_),
    .A1(net2156),
    .A2(net4199));
 sg13g2_a22oi_1 _26411_ (.Y(_19311_),
    .B1(net4328),
    .B2(_17374_),
    .A2(net4284),
    .A1(_17181_));
 sg13g2_a22oi_1 _26412_ (.Y(_00136_),
    .B1(_19310_),
    .B2(_19311_),
    .A2(net4200),
    .A1(_14009_));
 sg13g2_o21ai_1 _26413_ (.B1(net5562),
    .Y(_19312_),
    .A1(net1749),
    .A2(net4199));
 sg13g2_a22oi_1 _26414_ (.Y(_19313_),
    .B1(net4330),
    .B2(_17181_),
    .A2(net4287),
    .A1(_17454_));
 sg13g2_a22oi_1 _26415_ (.Y(_00137_),
    .B1(_19312_),
    .B2(_19313_),
    .A2(net4206),
    .A1(_14008_));
 sg13g2_o21ai_1 _26416_ (.B1(net5560),
    .Y(_19314_),
    .A1(net1704),
    .A2(net4199));
 sg13g2_a22oi_1 _26417_ (.Y(_19315_),
    .B1(net4328),
    .B2(_17454_),
    .A2(net4284),
    .A1(_17462_));
 sg13g2_a22oi_1 _26418_ (.Y(_00138_),
    .B1(_19314_),
    .B2(_19315_),
    .A2(net4200),
    .A1(_14007_));
 sg13g2_o21ai_1 _26419_ (.B1(net5559),
    .Y(_19316_),
    .A1(net1723),
    .A2(net4199));
 sg13g2_a22oi_1 _26420_ (.Y(_19317_),
    .B1(net4328),
    .B2(_17462_),
    .A2(net4284),
    .A1(_18777_));
 sg13g2_a22oi_1 _26421_ (.Y(_00139_),
    .B1(_19316_),
    .B2(_19317_),
    .A2(net4200),
    .A1(_14006_));
 sg13g2_o21ai_1 _26422_ (.B1(net5559),
    .Y(_19318_),
    .A1(net2109),
    .A2(net4199));
 sg13g2_a22oi_1 _26423_ (.Y(_19319_),
    .B1(net4328),
    .B2(_18777_),
    .A2(net4284),
    .A1(_17216_));
 sg13g2_a22oi_1 _26424_ (.Y(_00140_),
    .B1(_19318_),
    .B2(_19319_),
    .A2(net4200),
    .A1(_14005_));
 sg13g2_o21ai_1 _26425_ (.B1(net5560),
    .Y(_19320_),
    .A1(net1735),
    .A2(net4197));
 sg13g2_a22oi_1 _26426_ (.Y(_19321_),
    .B1(net4327),
    .B2(_17216_),
    .A2(net4283),
    .A1(_17391_));
 sg13g2_a22oi_1 _26427_ (.Y(_00141_),
    .B1(_19320_),
    .B2(_19321_),
    .A2(net4200),
    .A1(_14004_));
 sg13g2_o21ai_1 _26428_ (.B1(net5560),
    .Y(_19322_),
    .A1(net2088),
    .A2(net4199));
 sg13g2_a22oi_1 _26429_ (.Y(_19323_),
    .B1(net4327),
    .B2(_17391_),
    .A2(net4284),
    .A1(_17125_));
 sg13g2_a22oi_1 _26430_ (.Y(_00142_),
    .B1(_19322_),
    .B2(_19323_),
    .A2(net4200),
    .A1(_14003_));
 sg13g2_o21ai_1 _26431_ (.B1(net5559),
    .Y(_19324_),
    .A1(net2208),
    .A2(net4197));
 sg13g2_a22oi_1 _26432_ (.Y(_19325_),
    .B1(net4327),
    .B2(_17125_),
    .A2(net4283),
    .A1(_18840_));
 sg13g2_a22oi_1 _26433_ (.Y(_00143_),
    .B1(_19324_),
    .B2(_19325_),
    .A2(net4198),
    .A1(_14002_));
 sg13g2_o21ai_1 _26434_ (.B1(net5559),
    .Y(_19326_),
    .A1(net2086),
    .A2(net4197));
 sg13g2_a22oi_1 _26435_ (.Y(_19327_),
    .B1(net4327),
    .B2(_18840_),
    .A2(net4283),
    .A1(_16975_));
 sg13g2_a22oi_1 _26436_ (.Y(_00144_),
    .B1(_19326_),
    .B2(_19327_),
    .A2(net4198),
    .A1(_14001_));
 sg13g2_o21ai_1 _26437_ (.B1(net5559),
    .Y(_19328_),
    .A1(net1440),
    .A2(net4197));
 sg13g2_a22oi_1 _26438_ (.Y(_19329_),
    .B1(net4327),
    .B2(_16975_),
    .A2(net4283),
    .A1(_17733_));
 sg13g2_a22oi_1 _26439_ (.Y(_00145_),
    .B1(_19328_),
    .B2(_19329_),
    .A2(net4198),
    .A1(_14000_));
 sg13g2_o21ai_1 _26440_ (.B1(net5559),
    .Y(_19330_),
    .A1(net1695),
    .A2(net4197));
 sg13g2_a22oi_1 _26441_ (.Y(_19331_),
    .B1(net4327),
    .B2(_17733_),
    .A2(net4283),
    .A1(_17593_));
 sg13g2_a22oi_1 _26442_ (.Y(_00146_),
    .B1(_19330_),
    .B2(_19331_),
    .A2(net4198),
    .A1(_13999_));
 sg13g2_o21ai_1 _26443_ (.B1(net5553),
    .Y(_19332_),
    .A1(net1894),
    .A2(net4184));
 sg13g2_a22oi_1 _26444_ (.Y(_19333_),
    .B1(net4327),
    .B2(_17593_),
    .A2(net4283),
    .A1(_17397_));
 sg13g2_a22oi_1 _26445_ (.Y(_00147_),
    .B1(_19332_),
    .B2(_19333_),
    .A2(net4185),
    .A1(_13998_));
 sg13g2_o21ai_1 _26446_ (.B1(net5554),
    .Y(_19334_),
    .A1(net1571),
    .A2(net4184));
 sg13g2_a22oi_1 _26447_ (.Y(_19335_),
    .B1(net4324),
    .B2(_17397_),
    .A2(net4283),
    .A1(_17098_));
 sg13g2_a22oi_1 _26448_ (.Y(_00148_),
    .B1(_19334_),
    .B2(_19335_),
    .A2(net4185),
    .A1(_13997_));
 sg13g2_o21ai_1 _26449_ (.B1(net5559),
    .Y(_19336_),
    .A1(net1858),
    .A2(net4197));
 sg13g2_a22oi_1 _26450_ (.Y(_19337_),
    .B1(net4327),
    .B2(_17098_),
    .A2(net4283),
    .A1(_17333_));
 sg13g2_a22oi_1 _26451_ (.Y(_00149_),
    .B1(_19336_),
    .B2(_19337_),
    .A2(net4197),
    .A1(_13996_));
 sg13g2_o21ai_1 _26452_ (.B1(net5559),
    .Y(_19338_),
    .A1(net2098),
    .A2(net4197));
 sg13g2_a22oi_1 _26453_ (.Y(_19339_),
    .B1(net4324),
    .B2(_17333_),
    .A2(net4279),
    .A1(_18770_));
 sg13g2_a22oi_1 _26454_ (.Y(_00150_),
    .B1(_19338_),
    .B2(_19339_),
    .A2(net4185),
    .A1(_13995_));
 sg13g2_o21ai_1 _26455_ (.B1(net5554),
    .Y(_19340_),
    .A1(net1680),
    .A2(net4184));
 sg13g2_a22oi_1 _26456_ (.Y(_19341_),
    .B1(net4326),
    .B2(_18770_),
    .A2(net4279),
    .A1(_17379_));
 sg13g2_a22oi_1 _26457_ (.Y(_00151_),
    .B1(_19340_),
    .B2(_19341_),
    .A2(net4184),
    .A1(_13994_));
 sg13g2_o21ai_1 _26458_ (.B1(net5554),
    .Y(_19342_),
    .A1(net1536),
    .A2(net4184));
 sg13g2_a22oi_1 _26459_ (.Y(_19343_),
    .B1(net4326),
    .B2(_17379_),
    .A2(net4281),
    .A1(_17011_));
 sg13g2_a22oi_1 _26460_ (.Y(_00152_),
    .B1(_19342_),
    .B2(_19343_),
    .A2(net4184),
    .A1(_13993_));
 sg13g2_o21ai_1 _26461_ (.B1(net5554),
    .Y(_19344_),
    .A1(net1895),
    .A2(net4184));
 sg13g2_a22oi_1 _26462_ (.Y(_19345_),
    .B1(net4324),
    .B2(_17011_),
    .A2(net4279),
    .A1(_17340_));
 sg13g2_a22oi_1 _26463_ (.Y(_00153_),
    .B1(_19344_),
    .B2(_19345_),
    .A2(net4185),
    .A1(_13992_));
 sg13g2_o21ai_1 _26464_ (.B1(net5553),
    .Y(_19346_),
    .A1(net1688),
    .A2(net4182));
 sg13g2_a22oi_1 _26465_ (.Y(_19347_),
    .B1(net4324),
    .B2(_17340_),
    .A2(net4281),
    .A1(_17575_));
 sg13g2_a22oi_1 _26466_ (.Y(_00154_),
    .B1(_19346_),
    .B2(_19347_),
    .A2(net4184),
    .A1(_13991_));
 sg13g2_o21ai_1 _26467_ (.B1(net5553),
    .Y(_19348_),
    .A1(net1714),
    .A2(net4182));
 sg13g2_a22oi_1 _26468_ (.Y(_19349_),
    .B1(net4324),
    .B2(_17575_),
    .A2(net4279),
    .A1(_17416_));
 sg13g2_a22oi_1 _26469_ (.Y(_00155_),
    .B1(_19348_),
    .B2(_19349_),
    .A2(net4182),
    .A1(_13990_));
 sg13g2_o21ai_1 _26470_ (.B1(net5553),
    .Y(_19350_),
    .A1(net1826),
    .A2(net4182));
 sg13g2_a22oi_1 _26471_ (.Y(_19351_),
    .B1(net4324),
    .B2(_17416_),
    .A2(net4279),
    .A1(_17109_));
 sg13g2_a22oi_1 _26472_ (.Y(_00156_),
    .B1(_19350_),
    .B2(_19351_),
    .A2(net4182),
    .A1(_13989_));
 sg13g2_o21ai_1 _26473_ (.B1(net5553),
    .Y(_19352_),
    .A1(net1943),
    .A2(net4182));
 sg13g2_a22oi_1 _26474_ (.Y(_19353_),
    .B1(net4324),
    .B2(_17109_),
    .A2(net4279),
    .A1(_17421_));
 sg13g2_a22oi_1 _26475_ (.Y(_00157_),
    .B1(_19352_),
    .B2(_19353_),
    .A2(net4183),
    .A1(_13988_));
 sg13g2_o21ai_1 _26476_ (.B1(net5553),
    .Y(_19354_),
    .A1(net1875),
    .A2(net4182));
 sg13g2_a22oi_1 _26477_ (.Y(_19355_),
    .B1(net4324),
    .B2(_17421_),
    .A2(net4279),
    .A1(_17244_));
 sg13g2_a22oi_1 _26478_ (.Y(_00158_),
    .B1(_19354_),
    .B2(_19355_),
    .A2(net4183),
    .A1(_13987_));
 sg13g2_o21ai_1 _26479_ (.B1(net5550),
    .Y(_19356_),
    .A1(net1970),
    .A2(net4177));
 sg13g2_a22oi_1 _26480_ (.Y(_19357_),
    .B1(net4322),
    .B2(_17244_),
    .A2(net4277),
    .A1(_16870_));
 sg13g2_a22oi_1 _26481_ (.Y(_00159_),
    .B1(_19356_),
    .B2(_19357_),
    .A2(net4178),
    .A1(_13986_));
 sg13g2_o21ai_1 _26482_ (.B1(net5550),
    .Y(_19358_),
    .A1(net1780),
    .A2(net4178));
 sg13g2_a22oi_1 _26483_ (.Y(_19359_),
    .B1(net4322),
    .B2(_16870_),
    .A2(net4281),
    .A1(_16904_));
 sg13g2_a22oi_1 _26484_ (.Y(_00160_),
    .B1(_19358_),
    .B2(_19359_),
    .A2(net4178),
    .A1(_13985_));
 sg13g2_o21ai_1 _26485_ (.B1(net5553),
    .Y(_19360_),
    .A1(net1944),
    .A2(net4177));
 sg13g2_a22oi_1 _26486_ (.Y(_19361_),
    .B1(net4321),
    .B2(_16904_),
    .A2(net4277),
    .A1(_17738_));
 sg13g2_a22oi_1 _26487_ (.Y(_00161_),
    .B1(_19360_),
    .B2(_19361_),
    .A2(net4183),
    .A1(_13984_));
 sg13g2_o21ai_1 _26488_ (.B1(net5553),
    .Y(_19362_),
    .A1(net1683),
    .A2(net4182));
 sg13g2_a22oi_1 _26489_ (.Y(_19363_),
    .B1(net4321),
    .B2(_17738_),
    .A2(net4279),
    .A1(_17348_));
 sg13g2_a22oi_1 _26490_ (.Y(_00162_),
    .B1(_19362_),
    .B2(_19363_),
    .A2(net4183),
    .A1(_13983_));
 sg13g2_o21ai_1 _26491_ (.B1(net5551),
    .Y(_19364_),
    .A1(net1481),
    .A2(net4177));
 sg13g2_a22oi_1 _26492_ (.Y(_19365_),
    .B1(net4322),
    .B2(_17348_),
    .A2(net4281),
    .A1(_17299_));
 sg13g2_a22oi_1 _26493_ (.Y(_00163_),
    .B1(_19364_),
    .B2(_19365_),
    .A2(net4177),
    .A1(_13982_));
 sg13g2_o21ai_1 _26494_ (.B1(net5551),
    .Y(_19366_),
    .A1(net1564),
    .A2(net4177));
 sg13g2_a22oi_1 _26495_ (.Y(_19367_),
    .B1(net4321),
    .B2(_17299_),
    .A2(net4277),
    .A1(_17039_));
 sg13g2_a22oi_1 _26496_ (.Y(_00164_),
    .B1(_19366_),
    .B2(_19367_),
    .A2(net4177),
    .A1(_13981_));
 sg13g2_o21ai_1 _26497_ (.B1(net5551),
    .Y(_19368_),
    .A1(net1758),
    .A2(net4177));
 sg13g2_a22oi_1 _26498_ (.Y(_19369_),
    .B1(net4322),
    .B2(_17039_),
    .A2(net4278),
    .A1(_17567_));
 sg13g2_a22oi_1 _26499_ (.Y(_00165_),
    .B1(_19368_),
    .B2(_19369_),
    .A2(net4178),
    .A1(_13980_));
 sg13g2_o21ai_1 _26500_ (.B1(net5551),
    .Y(_19370_),
    .A1(net2006),
    .A2(net4177));
 sg13g2_a22oi_1 _26501_ (.Y(_19371_),
    .B1(net4321),
    .B2(_17567_),
    .A2(net4277),
    .A1(_17054_));
 sg13g2_a22oi_1 _26502_ (.Y(_00166_),
    .B1(_19370_),
    .B2(_19371_),
    .A2(net4178),
    .A1(_13979_));
 sg13g2_o21ai_1 _26503_ (.B1(net5550),
    .Y(_19372_),
    .A1(net1960),
    .A2(net4175));
 sg13g2_a22oi_1 _26504_ (.Y(_19373_),
    .B1(net4321),
    .B2(_17054_),
    .A2(net4277),
    .A1(_17165_));
 sg13g2_a22oi_1 _26505_ (.Y(_00167_),
    .B1(_19372_),
    .B2(_19373_),
    .A2(net4176),
    .A1(_13978_));
 sg13g2_o21ai_1 _26506_ (.B1(net5550),
    .Y(_19374_),
    .A1(net1978),
    .A2(net4176));
 sg13g2_a22oi_1 _26507_ (.Y(_19375_),
    .B1(net4321),
    .B2(_17165_),
    .A2(net4277),
    .A1(_18826_));
 sg13g2_a22oi_1 _26508_ (.Y(_00168_),
    .B1(_19374_),
    .B2(_19375_),
    .A2(net4176),
    .A1(_13977_));
 sg13g2_o21ai_1 _26509_ (.B1(net5550),
    .Y(_19376_),
    .A1(net1789),
    .A2(net4175));
 sg13g2_a22oi_1 _26510_ (.Y(_19377_),
    .B1(net4321),
    .B2(_18826_),
    .A2(net4277),
    .A1(_17327_));
 sg13g2_a22oi_1 _26511_ (.Y(_00169_),
    .B1(_19376_),
    .B2(_19377_),
    .A2(net4175),
    .A1(_13976_));
 sg13g2_o21ai_1 _26512_ (.B1(net5550),
    .Y(_19378_),
    .A1(net1764),
    .A2(net4176));
 sg13g2_nor2_1 _26513_ (.A(_17067_),
    .B(net4348),
    .Y(_19379_));
 sg13g2_a21oi_1 _26514_ (.A1(_17327_),
    .A2(net4321),
    .Y(_19380_),
    .B1(_19379_));
 sg13g2_a22oi_1 _26515_ (.Y(_00170_),
    .B1(_19378_),
    .B2(_19380_),
    .A2(net4175),
    .A1(_13975_));
 sg13g2_o21ai_1 _26516_ (.B1(net5550),
    .Y(_19381_),
    .A1(net1992),
    .A2(net4175));
 sg13g2_nor2_1 _26517_ (.A(_17067_),
    .B(net4260),
    .Y(_19382_));
 sg13g2_a21oi_1 _26518_ (.A1(_17147_),
    .A2(net4277),
    .Y(_19383_),
    .B1(_19382_));
 sg13g2_a22oi_1 _26519_ (.Y(_00171_),
    .B1(_19381_),
    .B2(_19383_),
    .A2(net4175),
    .A1(_13974_));
 sg13g2_o21ai_1 _26520_ (.B1(net5550),
    .Y(_19384_),
    .A1(net2065),
    .A2(net4175));
 sg13g2_a22oi_1 _26521_ (.Y(_19385_),
    .B1(net4318),
    .B2(_17147_),
    .A2(net4274),
    .A1(_18848_));
 sg13g2_a22oi_1 _26522_ (.Y(_00172_),
    .B1(_19384_),
    .B2(_19385_),
    .A2(net4175),
    .A1(_13973_));
 sg13g2_o21ai_1 _26523_ (.B1(net5543),
    .Y(_19386_),
    .A1(net1771),
    .A2(net4166));
 sg13g2_a22oi_1 _26524_ (.Y(_19387_),
    .B1(net4317),
    .B2(_18848_),
    .A2(net4274),
    .A1(_17403_));
 sg13g2_a22oi_1 _26525_ (.Y(_00173_),
    .B1(_19386_),
    .B2(_19387_),
    .A2(net4166),
    .A1(_13972_));
 sg13g2_o21ai_1 _26526_ (.B1(net5544),
    .Y(_19388_),
    .A1(net2001),
    .A2(net4166));
 sg13g2_a22oi_1 _26527_ (.Y(_19389_),
    .B1(net4318),
    .B2(_17403_),
    .A2(net4275),
    .A1(_17293_));
 sg13g2_a22oi_1 _26528_ (.Y(_00174_),
    .B1(_19388_),
    .B2(_19389_),
    .A2(net4167),
    .A1(_13971_));
 sg13g2_o21ai_1 _26529_ (.B1(net5543),
    .Y(_19390_),
    .A1(net1675),
    .A2(net4167));
 sg13g2_a22oi_1 _26530_ (.Y(_19391_),
    .B1(net4317),
    .B2(_17293_),
    .A2(net4274),
    .A1(_17139_));
 sg13g2_a22oi_1 _26531_ (.Y(_00175_),
    .B1(_19390_),
    .B2(_19391_),
    .A2(net4167),
    .A1(_13970_));
 sg13g2_o21ai_1 _26532_ (.B1(net5543),
    .Y(_19392_),
    .A1(net1927),
    .A2(net4167));
 sg13g2_a22oi_1 _26533_ (.Y(_19393_),
    .B1(net4317),
    .B2(_17139_),
    .A2(net4275),
    .A1(_18856_));
 sg13g2_a22oi_1 _26534_ (.Y(_00176_),
    .B1(_19392_),
    .B2(_19393_),
    .A2(net4167),
    .A1(_13969_));
 sg13g2_o21ai_1 _26535_ (.B1(net5543),
    .Y(_19394_),
    .A1(net1873),
    .A2(net4164));
 sg13g2_a22oi_1 _26536_ (.Y(_19395_),
    .B1(net4318),
    .B2(_18856_),
    .A2(net4275),
    .A1(_17354_));
 sg13g2_a22oi_1 _26537_ (.Y(_00177_),
    .B1(_19394_),
    .B2(_19395_),
    .A2(net4167),
    .A1(_13968_));
 sg13g2_o21ai_1 _26538_ (.B1(net5543),
    .Y(_19396_),
    .A1(net2133),
    .A2(net4166));
 sg13g2_a22oi_1 _26539_ (.Y(_19397_),
    .B1(net4318),
    .B2(_17354_),
    .A2(net4275),
    .A1(_17410_));
 sg13g2_a22oi_1 _26540_ (.Y(_00178_),
    .B1(_19396_),
    .B2(_19397_),
    .A2(net4167),
    .A1(_13967_));
 sg13g2_o21ai_1 _26541_ (.B1(net5543),
    .Y(_19398_),
    .A1(net1603),
    .A2(net4166));
 sg13g2_a22oi_1 _26542_ (.Y(_19399_),
    .B1(net4317),
    .B2(_17410_),
    .A2(net4274),
    .A1(_17156_));
 sg13g2_a22oi_1 _26543_ (.Y(_00179_),
    .B1(_19398_),
    .B2(_19399_),
    .A2(net4168),
    .A1(_13966_));
 sg13g2_o21ai_1 _26544_ (.B1(net5543),
    .Y(_19400_),
    .A1(net1747),
    .A2(net4166));
 sg13g2_a22oi_1 _26545_ (.Y(_19401_),
    .B1(net4317),
    .B2(_17156_),
    .A2(net4274),
    .A1(_18834_));
 sg13g2_a22oi_1 _26546_ (.Y(_00180_),
    .B1(_19400_),
    .B2(_19401_),
    .A2(net4168),
    .A1(_13965_));
 sg13g2_o21ai_1 _26547_ (.B1(net5543),
    .Y(_19402_),
    .A1(net1885),
    .A2(net4166));
 sg13g2_a22oi_1 _26548_ (.Y(_19403_),
    .B1(net4317),
    .B2(_18834_),
    .A2(net4274),
    .A1(_17274_));
 sg13g2_a22oi_1 _26549_ (.Y(_00181_),
    .B1(_19402_),
    .B2(_19403_),
    .A2(net4166),
    .A1(_13964_));
 sg13g2_o21ai_1 _26550_ (.B1(net5544),
    .Y(_19404_),
    .A1(net1783),
    .A2(net4165));
 sg13g2_a22oi_1 _26551_ (.Y(_19405_),
    .B1(net4317),
    .B2(_17274_),
    .A2(net4274),
    .A1(_17283_));
 sg13g2_a22oi_1 _26552_ (.Y(_00182_),
    .B1(_19404_),
    .B2(_19405_),
    .A2(net4165),
    .A1(_13963_));
 sg13g2_o21ai_1 _26553_ (.B1(net5544),
    .Y(_19406_),
    .A1(net2183),
    .A2(net4165));
 sg13g2_a22oi_1 _26554_ (.Y(_19407_),
    .B1(net4317),
    .B2(_17283_),
    .A2(net4274),
    .A1(_17025_));
 sg13g2_a22oi_1 _26555_ (.Y(_00183_),
    .B1(_19406_),
    .B2(_19407_),
    .A2(net4165),
    .A1(_13962_));
 sg13g2_o21ai_1 _26556_ (.B1(net5544),
    .Y(_19408_),
    .A1(net2152),
    .A2(net4165));
 sg13g2_a22oi_1 _26557_ (.Y(_19409_),
    .B1(net4314),
    .B2(_17025_),
    .A2(net4271),
    .A1(_18818_));
 sg13g2_a22oi_1 _26558_ (.Y(_00184_),
    .B1(_19408_),
    .B2(_19409_),
    .A2(net4165),
    .A1(_13961_));
 sg13g2_o21ai_1 _26559_ (.B1(net5540),
    .Y(_19410_),
    .A1(net1986),
    .A2(net4161));
 sg13g2_a22oi_1 _26560_ (.Y(_19411_),
    .B1(net4314),
    .B2(_18818_),
    .A2(net4271),
    .A1(_17386_));
 sg13g2_a22oi_1 _26561_ (.Y(_00185_),
    .B1(_19410_),
    .B2(_19411_),
    .A2(net4165),
    .A1(_13960_));
 sg13g2_o21ai_1 _26562_ (.B1(net5544),
    .Y(_19412_),
    .A1(net1844),
    .A2(net4161));
 sg13g2_a22oi_1 _26563_ (.Y(_19413_),
    .B1(net4315),
    .B2(_17386_),
    .A2(net4271),
    .A1(_17368_));
 sg13g2_a22oi_1 _26564_ (.Y(_00186_),
    .B1(_19412_),
    .B2(_19413_),
    .A2(net4165),
    .A1(_13959_));
 sg13g2_o21ai_1 _26565_ (.B1(net5541),
    .Y(_19414_),
    .A1(net1618),
    .A2(net4161));
 sg13g2_a22oi_1 _26566_ (.Y(_19415_),
    .B1(net4315),
    .B2(_17368_),
    .A2(net4272),
    .A1(_16984_));
 sg13g2_a22oi_1 _26567_ (.Y(_00187_),
    .B1(_19414_),
    .B2(_19415_),
    .A2(net4168),
    .A1(_13958_));
 sg13g2_o21ai_1 _26568_ (.B1(net5541),
    .Y(_19416_),
    .A1(net1560),
    .A2(net4162));
 sg13g2_a22oi_1 _26569_ (.Y(_19417_),
    .B1(net4315),
    .B2(_16984_),
    .A2(net4272),
    .A1(_18810_));
 sg13g2_a22oi_1 _26570_ (.Y(_00188_),
    .B1(_19416_),
    .B2(_19417_),
    .A2(net4162),
    .A1(_13957_));
 sg13g2_o21ai_1 _26571_ (.B1(net5540),
    .Y(_19418_),
    .A1(net1520),
    .A2(net4159));
 sg13g2_a22oi_1 _26572_ (.Y(_19419_),
    .B1(net4314),
    .B2(_18810_),
    .A2(net4271),
    .A1(_16804_));
 sg13g2_a22oi_1 _26573_ (.Y(_00189_),
    .B1(_19418_),
    .B2(_19419_),
    .A2(net4162),
    .A1(_13956_));
 sg13g2_o21ai_1 _26574_ (.B1(net5541),
    .Y(_19420_),
    .A1(net1540),
    .A2(net4161));
 sg13g2_a22oi_1 _26575_ (.Y(_19421_),
    .B1(net4315),
    .B2(_16804_),
    .A2(net4272),
    .A1(_16887_));
 sg13g2_a22oi_1 _26576_ (.Y(_00190_),
    .B1(_19420_),
    .B2(_19421_),
    .A2(net4162),
    .A1(_13955_));
 sg13g2_o21ai_1 _26577_ (.B1(net5540),
    .Y(_19422_),
    .A1(net1824),
    .A2(net4161));
 sg13g2_a22oi_1 _26578_ (.Y(_19423_),
    .B1(net4314),
    .B2(_16887_),
    .A2(net4272),
    .A1(_16850_));
 sg13g2_a22oi_1 _26579_ (.Y(_00191_),
    .B1(_19422_),
    .B2(_19423_),
    .A2(net4161),
    .A1(_13954_));
 sg13g2_o21ai_1 _26580_ (.B1(net5541),
    .Y(_19424_),
    .A1(net1662),
    .A2(net4161));
 sg13g2_a22oi_1 _26581_ (.Y(_19425_),
    .B1(net4314),
    .B2(_16850_),
    .A2(net4271),
    .A1(_16724_));
 sg13g2_a22oi_1 _26582_ (.Y(_00192_),
    .B1(_19424_),
    .B2(_19425_),
    .A2(net4161),
    .A1(_13953_));
 sg13g2_o21ai_1 _26583_ (.B1(net5540),
    .Y(_19426_),
    .A1(net1639),
    .A2(net4159));
 sg13g2_a22oi_1 _26584_ (.Y(_19427_),
    .B1(net4314),
    .B2(_16724_),
    .A2(net4271),
    .A1(_18762_));
 sg13g2_a22oi_1 _26585_ (.Y(_00193_),
    .B1(_19426_),
    .B2(_19427_),
    .A2(net4159),
    .A1(_13952_));
 sg13g2_o21ai_1 _26586_ (.B1(net5540),
    .Y(_19428_),
    .A1(net1909),
    .A2(net4159));
 sg13g2_a22oi_1 _26587_ (.Y(_19429_),
    .B1(net4314),
    .B2(_18762_),
    .A2(net4271),
    .A1(_18746_));
 sg13g2_a22oi_1 _26588_ (.Y(_00194_),
    .B1(_19428_),
    .B2(_19429_),
    .A2(net4160),
    .A1(_13951_));
 sg13g2_o21ai_1 _26589_ (.B1(net5540),
    .Y(_19430_),
    .A1(net1467),
    .A2(net4159));
 sg13g2_a22oi_1 _26590_ (.Y(_19431_),
    .B1(net4314),
    .B2(_18746_),
    .A2(net4271),
    .A1(_17187_));
 sg13g2_a22oi_1 _26591_ (.Y(_00195_),
    .B1(_19430_),
    .B2(_19431_),
    .A2(net4160),
    .A1(_13950_));
 sg13g2_o21ai_1 _26592_ (.B1(net5540),
    .Y(_19432_),
    .A1(net1985),
    .A2(net4159));
 sg13g2_a22oi_1 _26593_ (.Y(_19433_),
    .B1(net4310),
    .B2(_17187_),
    .A2(net4266),
    .A1(_16831_));
 sg13g2_a22oi_1 _26594_ (.Y(_00196_),
    .B1(_19432_),
    .B2(_19433_),
    .A2(net4160),
    .A1(_13949_));
 sg13g2_o21ai_1 _26595_ (.B1(net5533),
    .Y(_19434_),
    .A1(net1685),
    .A2(net4149));
 sg13g2_a22oi_1 _26596_ (.Y(_19435_),
    .B1(net4311),
    .B2(_16831_),
    .A2(net4267),
    .A1(_16990_));
 sg13g2_a22oi_1 _26597_ (.Y(_00197_),
    .B1(_19434_),
    .B2(_19435_),
    .A2(net4160),
    .A1(_13948_));
 sg13g2_o21ai_1 _26598_ (.B1(net5534),
    .Y(_19436_),
    .A1(net1905),
    .A2(net4149));
 sg13g2_a22oi_1 _26599_ (.Y(_19437_),
    .B1(net4311),
    .B2(_16990_),
    .A2(net4267),
    .A1(_17262_));
 sg13g2_a22oi_1 _26600_ (.Y(_00198_),
    .B1(_19436_),
    .B2(_19437_),
    .A2(net4150),
    .A1(_13947_));
 sg13g2_o21ai_1 _26601_ (.B1(net5540),
    .Y(_19438_),
    .A1(net1469),
    .A2(net4159));
 sg13g2_a22oi_1 _26602_ (.Y(_19439_),
    .B1(net4310),
    .B2(_17262_),
    .A2(net4266),
    .A1(_16909_));
 sg13g2_a22oi_1 _26603_ (.Y(_00199_),
    .B1(_19438_),
    .B2(_19439_),
    .A2(net4159),
    .A1(_13946_));
 sg13g2_o21ai_1 _26604_ (.B1(net5534),
    .Y(_19440_),
    .A1(net1586),
    .A2(net4149));
 sg13g2_a22oi_1 _26605_ (.Y(_19441_),
    .B1(net4311),
    .B2(_16909_),
    .A2(net4267),
    .A1(_16741_));
 sg13g2_a22oi_1 _26606_ (.Y(_00200_),
    .B1(_19440_),
    .B2(_19441_),
    .A2(net4149),
    .A1(_13945_));
 sg13g2_o21ai_1 _26607_ (.B1(net5534),
    .Y(_19442_),
    .A1(net2059),
    .A2(net4149));
 sg13g2_a22oi_1 _26608_ (.Y(_19443_),
    .B1(net4311),
    .B2(_16741_),
    .A2(net4267),
    .A1(_17194_));
 sg13g2_a22oi_1 _26609_ (.Y(_00201_),
    .B1(_19442_),
    .B2(_19443_),
    .A2(net4149),
    .A1(_13944_));
 sg13g2_o21ai_1 _26610_ (.B1(net5534),
    .Y(_19444_),
    .A1(net1551),
    .A2(net4149));
 sg13g2_a22oi_1 _26611_ (.Y(_19445_),
    .B1(net4311),
    .B2(_17194_),
    .A2(net4267),
    .A1(_17429_));
 sg13g2_a22oi_1 _26612_ (.Y(_00202_),
    .B1(_19444_),
    .B2(_19445_),
    .A2(net4150),
    .A1(_13943_));
 sg13g2_o21ai_1 _26613_ (.B1(net5534),
    .Y(_19446_),
    .A1(net1919),
    .A2(net4149));
 sg13g2_a22oi_1 _26614_ (.Y(_19447_),
    .B1(net4310),
    .B2(_17429_),
    .A2(net4266),
    .A1(_16880_));
 sg13g2_a22oi_1 _26615_ (.Y(_00203_),
    .B1(_19446_),
    .B2(_19447_),
    .A2(net4150),
    .A1(_13942_));
 sg13g2_o21ai_1 _26616_ (.B1(net5533),
    .Y(_19448_),
    .A1(net1814),
    .A2(net4147));
 sg13g2_a22oi_1 _26617_ (.Y(_19449_),
    .B1(net4310),
    .B2(_16880_),
    .A2(net4266),
    .A1(_16772_));
 sg13g2_a22oi_1 _26618_ (.Y(_00204_),
    .B1(_19448_),
    .B2(_19449_),
    .A2(net4148),
    .A1(_13941_));
 sg13g2_o21ai_1 _26619_ (.B1(net5533),
    .Y(_19450_),
    .A1(net1593),
    .A2(net4147));
 sg13g2_a22oi_1 _26620_ (.Y(_19451_),
    .B1(net4310),
    .B2(_16772_),
    .A2(net4266),
    .A1(_17267_));
 sg13g2_a22oi_1 _26621_ (.Y(_00205_),
    .B1(_19450_),
    .B2(_19451_),
    .A2(net4148),
    .A1(_13940_));
 sg13g2_o21ai_1 _26622_ (.B1(net5533),
    .Y(_19452_),
    .A1(net2179),
    .A2(net4148));
 sg13g2_a22oi_1 _26623_ (.Y(_19453_),
    .B1(net4310),
    .B2(_17267_),
    .A2(net4266),
    .A1(_16813_));
 sg13g2_a22oi_1 _26624_ (.Y(_00206_),
    .B1(_19452_),
    .B2(_19453_),
    .A2(net4148),
    .A1(_13939_));
 sg13g2_o21ai_1 _26625_ (.B1(net5533),
    .Y(_19454_),
    .A1(net1637),
    .A2(net4148));
 sg13g2_a22oi_1 _26626_ (.Y(_19455_),
    .B1(net4310),
    .B2(_16813_),
    .A2(net4266),
    .A1(_16915_));
 sg13g2_a22oi_1 _26627_ (.Y(_00207_),
    .B1(_19454_),
    .B2(_19455_),
    .A2(net4148),
    .A1(_13938_));
 sg13g2_o21ai_1 _26628_ (.B1(net5533),
    .Y(_19456_),
    .A1(net2089),
    .A2(net4147));
 sg13g2_a22oi_1 _26629_ (.Y(_19457_),
    .B1(net4310),
    .B2(_16915_),
    .A2(net4266),
    .A1(_16701_));
 sg13g2_a22oi_1 _26630_ (.Y(_00208_),
    .B1(_19456_),
    .B2(_19457_),
    .A2(net4147),
    .A1(_13937_));
 sg13g2_o21ai_1 _26631_ (.B1(net5533),
    .Y(_19458_),
    .A1(net2192),
    .A2(net4147));
 sg13g2_a22oi_1 _26632_ (.Y(_19459_),
    .B1(net4308),
    .B2(_16701_),
    .A2(net4264),
    .A1(_17439_));
 sg13g2_a22oi_1 _26633_ (.Y(_00209_),
    .B1(_19458_),
    .B2(_19459_),
    .A2(net4147),
    .A1(_13936_));
 sg13g2_o21ai_1 _26634_ (.B1(net5533),
    .Y(_19460_),
    .A1(net1706),
    .A2(net4147));
 sg13g2_a22oi_1 _26635_ (.Y(_19461_),
    .B1(net4308),
    .B2(_17439_),
    .A2(net4264),
    .A1(_17448_));
 sg13g2_a22oi_1 _26636_ (.Y(_00210_),
    .B1(_19460_),
    .B2(_19461_),
    .A2(net4147),
    .A1(_13935_));
 sg13g2_o21ai_1 _26637_ (.B1(net5531),
    .Y(_19462_),
    .A1(net1473),
    .A2(net4143));
 sg13g2_a22oi_1 _26638_ (.Y(_19463_),
    .B1(net4308),
    .B2(_17448_),
    .A2(net4264),
    .A1(_16821_));
 sg13g2_a22oi_1 _26639_ (.Y(_00211_),
    .B1(_19462_),
    .B2(_19463_),
    .A2(net4148),
    .A1(_13934_));
 sg13g2_o21ai_1 _26640_ (.B1(net5531),
    .Y(_19464_),
    .A1(net1498),
    .A2(net4140));
 sg13g2_a22oi_1 _26641_ (.Y(_19465_),
    .B1(net4308),
    .B2(_16821_),
    .A2(net4269),
    .A1(_16783_));
 sg13g2_a22oi_1 _26642_ (.Y(_00212_),
    .B1(_19464_),
    .B2(_19465_),
    .A2(net4144),
    .A1(_13933_));
 sg13g2_o21ai_1 _26643_ (.B1(net5531),
    .Y(_19466_),
    .A1(net1568),
    .A2(net4143));
 sg13g2_a22oi_1 _26644_ (.Y(_19467_),
    .B1(net4309),
    .B2(_16783_),
    .A2(net4269),
    .A1(_16790_));
 sg13g2_a22oi_1 _26645_ (.Y(_00213_),
    .B1(_19466_),
    .B2(_19467_),
    .A2(net4143),
    .A1(_13932_));
 sg13g2_o21ai_1 _26646_ (.B1(net5531),
    .Y(_19468_),
    .A1(net1553),
    .A2(net4143));
 sg13g2_a22oi_1 _26647_ (.Y(_19469_),
    .B1(net4308),
    .B2(_16790_),
    .A2(net4264),
    .A1(_16799_));
 sg13g2_a22oi_1 _26648_ (.Y(_00214_),
    .B1(_19468_),
    .B2(_19469_),
    .A2(net4143),
    .A1(_13931_));
 sg13g2_o21ai_1 _26649_ (.B1(net5532),
    .Y(_19470_),
    .A1(net1580),
    .A2(net4143));
 sg13g2_a22oi_1 _26650_ (.Y(_19471_),
    .B1(net4309),
    .B2(_16799_),
    .A2(net4265),
    .A1(_16761_));
 sg13g2_a22oi_1 _26651_ (.Y(_00215_),
    .B1(_19470_),
    .B2(_19471_),
    .A2(net4144),
    .A1(_13930_));
 sg13g2_o21ai_1 _26652_ (.B1(net5532),
    .Y(_19472_),
    .A1(net1833),
    .A2(net4143));
 sg13g2_a22oi_1 _26653_ (.Y(_19473_),
    .B1(net4308),
    .B2(_16761_),
    .A2(net4264),
    .A1(_16896_));
 sg13g2_a22oi_1 _26654_ (.Y(_00216_),
    .B1(_19472_),
    .B2(_19473_),
    .A2(net4144),
    .A1(_13929_));
 sg13g2_o21ai_1 _26655_ (.B1(net5531),
    .Y(_19474_),
    .A1(net1794),
    .A2(net4142));
 sg13g2_a22oi_1 _26656_ (.Y(_19475_),
    .B1(net4308),
    .B2(_16896_),
    .A2(net4264),
    .A1(_16836_));
 sg13g2_a22oi_1 _26657_ (.Y(_00217_),
    .B1(_19474_),
    .B2(_19475_),
    .A2(net4144),
    .A1(_13928_));
 sg13g2_o21ai_1 _26658_ (.B1(net5531),
    .Y(_19476_),
    .A1(net2215),
    .A2(net4142));
 sg13g2_a22oi_1 _26659_ (.Y(_19477_),
    .B1(net4308),
    .B2(_16836_),
    .A2(net4264),
    .A1(_16844_));
 sg13g2_a22oi_1 _26660_ (.Y(_00218_),
    .B1(_19476_),
    .B2(_19477_),
    .A2(net4144),
    .A1(_13927_));
 sg13g2_o21ai_1 _26661_ (.B1(net5528),
    .Y(_19478_),
    .A1(net1642),
    .A2(net4133));
 sg13g2_a22oi_1 _26662_ (.Y(_19479_),
    .B1(net4307),
    .B2(_16844_),
    .A2(net4262),
    .A1(_16748_));
 sg13g2_a22oi_1 _26663_ (.Y(_00219_),
    .B1(_19478_),
    .B2(_19479_),
    .A2(net4142),
    .A1(_13926_));
 sg13g2_o21ai_1 _26664_ (.B1(net5528),
    .Y(_19480_),
    .A1(net2780),
    .A2(net4133));
 sg13g2_a22oi_1 _26665_ (.Y(_19481_),
    .B1(net4306),
    .B2(_16748_),
    .A2(net4261),
    .A1(_16681_));
 sg13g2_a22oi_1 _26666_ (.Y(_00220_),
    .B1(_19480_),
    .B2(_19481_),
    .A2(net4132),
    .A1(_13925_));
 sg13g2_o21ai_1 _26667_ (.B1(net5528),
    .Y(_19482_),
    .A1(net1648),
    .A2(net4132));
 sg13g2_a22oi_1 _26668_ (.Y(_19483_),
    .B1(net4307),
    .B2(_16681_),
    .A2(net4261),
    .A1(_16935_));
 sg13g2_a22oi_1 _26669_ (.Y(_00221_),
    .B1(_19482_),
    .B2(_19483_),
    .A2(net4133),
    .A1(_13924_));
 sg13g2_o21ai_1 _26670_ (.B1(net5528),
    .Y(_19484_),
    .A1(net1490),
    .A2(net4132));
 sg13g2_a22oi_1 _26671_ (.Y(_19485_),
    .B1(net4307),
    .B2(_16935_),
    .A2(net4262),
    .A1(_16948_));
 sg13g2_a22oi_1 _26672_ (.Y(_00222_),
    .B1(_19484_),
    .B2(_19485_),
    .A2(net4132),
    .A1(_13923_));
 sg13g2_o21ai_1 _26673_ (.B1(net5531),
    .Y(_19486_),
    .A1(net1635),
    .A2(net4142));
 sg13g2_a22oi_1 _26674_ (.Y(_19487_),
    .B1(net4307),
    .B2(_16948_),
    .A2(net4261),
    .A1(_18886_));
 sg13g2_a22oi_1 _26675_ (.Y(_00223_),
    .B1(_19486_),
    .B2(_19487_),
    .A2(net4142),
    .A1(_13922_));
 sg13g2_o21ai_1 _26676_ (.B1(net5537),
    .Y(_19488_),
    .A1(net2288),
    .A2(net4132));
 sg13g2_a22oi_1 _26677_ (.Y(_19489_),
    .B1(net4307),
    .B2(_18886_),
    .A2(net4262),
    .A1(_18879_));
 sg13g2_a22oi_1 _26678_ (.Y(_00224_),
    .B1(_19488_),
    .B2(_19489_),
    .A2(net4142),
    .A1(_13921_));
 sg13g2_nand2_1 _26679_ (.Y(_19490_),
    .A(net1842),
    .B(net5627));
 sg13g2_nand2b_1 _26680_ (.Y(_19491_),
    .B(_19008_),
    .A_N(_18879_));
 sg13g2_a21oi_1 _26681_ (.A1(_18905_),
    .A2(_19007_),
    .Y(_19492_),
    .B1(net5537));
 sg13g2_a22oi_1 _26682_ (.Y(_19493_),
    .B1(_19491_),
    .B2(_19492_),
    .A2(net4132),
    .A1(\u_inv.f_next[254] ));
 sg13g2_o21ai_1 _26683_ (.B1(_19493_),
    .Y(_00225_),
    .A1(net4132),
    .A2(_19490_));
 sg13g2_o21ai_1 _26684_ (.B1(net5531),
    .Y(_19494_),
    .A1(net1605),
    .A2(net4142));
 sg13g2_nor2_1 _26685_ (.A(_18905_),
    .B(net4260),
    .Y(_19495_));
 sg13g2_a21oi_1 _26686_ (.A1(_18909_),
    .A2(net4264),
    .Y(_19496_),
    .B1(_19495_));
 sg13g2_a22oi_1 _26687_ (.Y(_00226_),
    .B1(_19494_),
    .B2(_19496_),
    .A2(net4142),
    .A1(_13919_));
 sg13g2_a21oi_1 _26688_ (.A1(_14246_),
    .A2(_14511_),
    .Y(_00227_),
    .B1(net1074));
 sg13g2_and2_1 _26689_ (.A(_14243_),
    .B(_14814_),
    .X(_19497_));
 sg13g2_nor2_1 _26690_ (.A(net5882),
    .B(_14815_),
    .Y(_19498_));
 sg13g2_a21oi_1 _26691_ (.A1(pipe_pending),
    .A2(_14815_),
    .Y(_19499_),
    .B1(net5882));
 sg13g2_a21oi_1 _26692_ (.A1(net1965),
    .A2(_14815_),
    .Y(_19500_),
    .B1(_14809_));
 sg13g2_nor4_1 _26693_ (.A(net5882),
    .B(_14816_),
    .C(_19497_),
    .D(_19500_),
    .Y(_19501_));
 sg13g2_or2_1 _26694_ (.X(_00228_),
    .B(_19501_),
    .A(_14812_));
 sg13g2_and2_1 _26695_ (.A(inv_done),
    .B(_14810_),
    .X(_19502_));
 sg13g2_nand2_2 _26696_ (.Y(_19503_),
    .A(inv_done),
    .B(_14810_));
 sg13g2_a21oi_1 _26697_ (.A1(uio_out[1]),
    .A2(_14816_),
    .Y(_19504_),
    .B1(net5482));
 sg13g2_inv_1 _26698_ (.Y(_00229_),
    .A(_19504_));
 sg13g2_nand2_2 _26699_ (.Y(_19505_),
    .A(_14809_),
    .B(net5442));
 sg13g2_nor2_1 _26700_ (.A(net2548),
    .B(_19505_),
    .Y(_19506_));
 sg13g2_a221oi_1 _26701_ (.B2(_14817_),
    .C1(_19498_),
    .B1(_14812_),
    .A1(\state[1] ),
    .Y(_19507_),
    .A2(\state[0] ));
 sg13g2_nor2_1 _26702_ (.A(_19500_),
    .B(_19506_),
    .Y(_19508_));
 sg13g2_nor2_1 _26703_ (.A(net2548),
    .B(net5230),
    .Y(_19509_));
 sg13g2_a21oi_1 _26704_ (.A1(net5230),
    .A2(_19508_),
    .Y(_00230_),
    .B1(_19509_));
 sg13g2_a21oi_1 _26705_ (.A1(\byte_cnt[0] ),
    .A2(net5230),
    .Y(_19510_),
    .B1(net1181));
 sg13g2_a21o_1 _26706_ (.A2(\byte_cnt[0] ),
    .A1(net1181),
    .B1(_19505_),
    .X(_19511_));
 sg13g2_a21oi_1 _26707_ (.A1(net5230),
    .A2(_19511_),
    .Y(_00231_),
    .B1(net1182));
 sg13g2_o21ai_1 _26708_ (.B1(net5230),
    .Y(_19512_),
    .A1(_14813_),
    .A2(_19505_));
 sg13g2_nand3_1 _26709_ (.B(net2548),
    .C(net5230),
    .A(net1181),
    .Y(_19513_));
 sg13g2_nand2b_1 _26710_ (.Y(_19514_),
    .B(_19513_),
    .A_N(net3313));
 sg13g2_and2_1 _26711_ (.A(_19512_),
    .B(_19514_),
    .X(_00232_));
 sg13g2_nand2b_1 _26712_ (.Y(_19515_),
    .B(_14813_),
    .A_N(net2831));
 sg13g2_nor2_1 _26713_ (.A(_19505_),
    .B(_19515_),
    .Y(_19516_));
 sg13g2_a22oi_1 _26714_ (.Y(_19517_),
    .B1(_19516_),
    .B2(net5230),
    .A2(_19512_),
    .A1(net2831));
 sg13g2_inv_1 _26715_ (.Y(_00233_),
    .A(net2832));
 sg13g2_nand3_1 _26716_ (.B(_14813_),
    .C(_19507_),
    .A(\byte_cnt[3] ),
    .Y(_19518_));
 sg13g2_nand3_1 _26717_ (.B(_14814_),
    .C(net5435),
    .A(_14809_),
    .Y(_19519_));
 sg13g2_a22oi_1 _26718_ (.Y(_00234_),
    .B1(_19519_),
    .B2(net5230),
    .A2(_19518_),
    .A1(_14247_));
 sg13g2_nor2_1 _26719_ (.A(_14243_),
    .B(_19499_),
    .Y(_19520_));
 sg13g2_nand3b_1 _26720_ (.B(net10),
    .C(\state[1] ),
    .Y(_19521_),
    .A_N(rd_prev));
 sg13g2_a221oi_1 _26721_ (.B2(_19521_),
    .C1(_19520_),
    .B1(_19498_),
    .A1(_14812_),
    .Y(_19522_),
    .A2(_14817_));
 sg13g2_a22oi_1 _26722_ (.Y(_19523_),
    .B1(net5296),
    .B2(net1),
    .A2(net5481),
    .A1(net1172));
 sg13g2_nor2_1 _26723_ (.A(net1397),
    .B(net5138),
    .Y(_19524_));
 sg13g2_a21oi_1 _26724_ (.A1(net5138),
    .A2(_19523_),
    .Y(_00235_),
    .B1(_19524_));
 sg13g2_a22oi_1 _26725_ (.Y(_19525_),
    .B1(net5296),
    .B2(net2),
    .A2(net5481),
    .A1(net1273));
 sg13g2_nor2_1 _26726_ (.A(net2066),
    .B(net5140),
    .Y(_19526_));
 sg13g2_a21oi_1 _26727_ (.A1(net5140),
    .A2(_19525_),
    .Y(_00236_),
    .B1(_19526_));
 sg13g2_a22oi_1 _26728_ (.Y(_19527_),
    .B1(net5296),
    .B2(net3),
    .A2(net5481),
    .A1(net1656));
 sg13g2_nor2_1 _26729_ (.A(net1312),
    .B(net5139),
    .Y(_19528_));
 sg13g2_a21oi_1 _26730_ (.A1(net5139),
    .A2(_19527_),
    .Y(_00237_),
    .B1(_19528_));
 sg13g2_a22oi_1 _26731_ (.Y(_19529_),
    .B1(net5296),
    .B2(net4),
    .A2(net5481),
    .A1(net1124));
 sg13g2_nor2_1 _26732_ (.A(net1287),
    .B(net5145),
    .Y(_19530_));
 sg13g2_a21oi_1 _26733_ (.A1(net5145),
    .A2(_19529_),
    .Y(_00238_),
    .B1(_19530_));
 sg13g2_a22oi_1 _26734_ (.Y(_19531_),
    .B1(net5296),
    .B2(net5),
    .A2(net5481),
    .A1(net1411));
 sg13g2_nor2_1 _26735_ (.A(net1326),
    .B(net5143),
    .Y(_19532_));
 sg13g2_a21oi_1 _26736_ (.A1(net5143),
    .A2(_19531_),
    .Y(_00239_),
    .B1(_19532_));
 sg13g2_a22oi_1 _26737_ (.Y(_19533_),
    .B1(net5296),
    .B2(net6),
    .A2(net5481),
    .A1(net1270));
 sg13g2_nor2_1 _26738_ (.A(net1629),
    .B(net5143),
    .Y(_19534_));
 sg13g2_a21oi_1 _26739_ (.A1(net5144),
    .A2(_19533_),
    .Y(_00240_),
    .B1(_19534_));
 sg13g2_a22oi_1 _26740_ (.Y(_19535_),
    .B1(net5296),
    .B2(net7),
    .A2(net5481),
    .A1(net1364));
 sg13g2_nor2_1 _26741_ (.A(net2319),
    .B(net5140),
    .Y(_19536_));
 sg13g2_a21oi_1 _26742_ (.A1(net5140),
    .A2(_19535_),
    .Y(_00241_),
    .B1(_19536_));
 sg13g2_a22oi_1 _26743_ (.Y(_19537_),
    .B1(net5296),
    .B2(net8),
    .A2(net5481),
    .A1(net1237));
 sg13g2_nor2_1 _26744_ (.A(net1644),
    .B(net5145),
    .Y(_19538_));
 sg13g2_a21oi_1 _26745_ (.A1(net5145),
    .A2(_19537_),
    .Y(_00242_),
    .B1(_19538_));
 sg13g2_and2_1 _26746_ (.A(net1397),
    .B(net5434),
    .X(_19539_));
 sg13g2_a21oi_1 _26747_ (.A1(net1132),
    .A2(net5482),
    .Y(_19540_),
    .B1(_19539_));
 sg13g2_nor2_1 _26748_ (.A(net2545),
    .B(net5142),
    .Y(_19541_));
 sg13g2_a21oi_1 _26749_ (.A1(net5139),
    .A2(_19540_),
    .Y(_00243_),
    .B1(_19541_));
 sg13g2_and2_1 _26750_ (.A(net2066),
    .B(net5434),
    .X(_19542_));
 sg13g2_a21oi_1 _26751_ (.A1(net1442),
    .A2(net5482),
    .Y(_19543_),
    .B1(_19542_));
 sg13g2_nor2_1 _26752_ (.A(net2453),
    .B(net5142),
    .Y(_19544_));
 sg13g2_a21oi_1 _26753_ (.A1(net5142),
    .A2(_19543_),
    .Y(_00244_),
    .B1(_19544_));
 sg13g2_nand3_1 _26754_ (.B(net5434),
    .C(net5142),
    .A(net1312),
    .Y(_19545_));
 sg13g2_o21ai_1 _26755_ (.B1(_19545_),
    .Y(_00245_),
    .A1(_14512_),
    .A2(net5142));
 sg13g2_nand3_1 _26756_ (.B(net5434),
    .C(net5143),
    .A(net1287),
    .Y(_19546_));
 sg13g2_o21ai_1 _26757_ (.B1(_19546_),
    .Y(_00246_),
    .A1(_14513_),
    .A2(net5143));
 sg13g2_nand3_1 _26758_ (.B(net5442),
    .C(net5150),
    .A(net1326),
    .Y(_19547_));
 sg13g2_o21ai_1 _26759_ (.B1(_19547_),
    .Y(_00247_),
    .A1(_14515_),
    .A2(net5150));
 sg13g2_nand3_1 _26760_ (.B(net5435),
    .C(net5143),
    .A(net1629),
    .Y(_19548_));
 sg13g2_o21ai_1 _26761_ (.B1(_19548_),
    .Y(_00248_),
    .A1(_14516_),
    .A2(net5144));
 sg13g2_nand3_1 _26762_ (.B(net5435),
    .C(net5142),
    .A(net2319),
    .Y(_19549_));
 sg13g2_o21ai_1 _26763_ (.B1(_19549_),
    .Y(_00249_),
    .A1(_14517_),
    .A2(net5143));
 sg13g2_nand3_1 _26764_ (.B(net5434),
    .C(net5142),
    .A(net1644),
    .Y(_19550_));
 sg13g2_o21ai_1 _26765_ (.B1(_19550_),
    .Y(_00250_),
    .A1(_14518_),
    .A2(net5143));
 sg13g2_and2_1 _26766_ (.A(\shift_reg[8] ),
    .B(net5434),
    .X(_19551_));
 sg13g2_a21oi_1 _26767_ (.A1(net1249),
    .A2(net5480),
    .Y(_19552_),
    .B1(_19551_));
 sg13g2_nor2_1 _26768_ (.A(net2460),
    .B(net5147),
    .Y(_19553_));
 sg13g2_a21oi_1 _26769_ (.A1(net5147),
    .A2(_19552_),
    .Y(_00251_),
    .B1(_19553_));
 sg13g2_and2_1 _26770_ (.A(\shift_reg[9] ),
    .B(net5433),
    .X(_19554_));
 sg13g2_a21oi_1 _26771_ (.A1(\inv_result[1] ),
    .A2(net5483),
    .Y(_19555_),
    .B1(_19554_));
 sg13g2_nor2_1 _26772_ (.A(net2228),
    .B(net5147),
    .Y(_19556_));
 sg13g2_a21oi_1 _26773_ (.A1(net5147),
    .A2(_19555_),
    .Y(_00252_),
    .B1(_19556_));
 sg13g2_nor2_1 _26774_ (.A(_14512_),
    .B(net5483),
    .Y(_19557_));
 sg13g2_a21oi_1 _26775_ (.A1(\inv_result[2] ),
    .A2(net5483),
    .Y(_19558_),
    .B1(_19557_));
 sg13g2_nor2_1 _26776_ (.A(net2211),
    .B(net5147),
    .Y(_19559_));
 sg13g2_a21oi_1 _26777_ (.A1(net5147),
    .A2(_19558_),
    .Y(_00253_),
    .B1(_19559_));
 sg13g2_nor2_1 _26778_ (.A(_14513_),
    .B(net5483),
    .Y(_19560_));
 sg13g2_a21oi_1 _26779_ (.A1(net1837),
    .A2(net5483),
    .Y(_19561_),
    .B1(_19560_));
 sg13g2_nor2_1 _26780_ (.A(net1910),
    .B(net5149),
    .Y(_19562_));
 sg13g2_a21oi_1 _26781_ (.A1(net5149),
    .A2(_19561_),
    .Y(_00254_),
    .B1(_19562_));
 sg13g2_nor2_1 _26782_ (.A(_14515_),
    .B(net5484),
    .Y(_19563_));
 sg13g2_a21oi_1 _26783_ (.A1(\inv_result[4] ),
    .A2(net5484),
    .Y(_19564_),
    .B1(_19563_));
 sg13g2_nor2_1 _26784_ (.A(net1962),
    .B(net5149),
    .Y(_19565_));
 sg13g2_a21oi_1 _26785_ (.A1(net5149),
    .A2(_19564_),
    .Y(_00255_),
    .B1(_19565_));
 sg13g2_nor2_1 _26786_ (.A(_14516_),
    .B(net5484),
    .Y(_19566_));
 sg13g2_a21oi_1 _26787_ (.A1(net1325),
    .A2(net5484),
    .Y(_19567_),
    .B1(_19566_));
 sg13g2_nor2_1 _26788_ (.A(net2126),
    .B(net5151),
    .Y(_19568_));
 sg13g2_a21oi_1 _26789_ (.A1(net5151),
    .A2(_19567_),
    .Y(_00256_),
    .B1(_19568_));
 sg13g2_nor2_1 _26790_ (.A(_14517_),
    .B(net5484),
    .Y(_19569_));
 sg13g2_a21oi_1 _26791_ (.A1(net1206),
    .A2(net5485),
    .Y(_19570_),
    .B1(_19569_));
 sg13g2_nor2_1 _26792_ (.A(net2028),
    .B(net5151),
    .Y(_19571_));
 sg13g2_a21oi_1 _26793_ (.A1(net5151),
    .A2(_19570_),
    .Y(_00257_),
    .B1(_19571_));
 sg13g2_nor2_1 _26794_ (.A(_14518_),
    .B(net5486),
    .Y(_19572_));
 sg13g2_a21oi_1 _26795_ (.A1(net1111),
    .A2(net5485),
    .Y(_19573_),
    .B1(_19572_));
 sg13g2_nor2_1 _26796_ (.A(net1465),
    .B(net5152),
    .Y(_19574_));
 sg13g2_a21oi_1 _26797_ (.A1(net5151),
    .A2(_19573_),
    .Y(_00258_),
    .B1(_19574_));
 sg13g2_and2_1 _26798_ (.A(\shift_reg[16] ),
    .B(net5436),
    .X(_19575_));
 sg13g2_a21oi_1 _26799_ (.A1(net1257),
    .A2(net5485),
    .Y(_19576_),
    .B1(_19575_));
 sg13g2_nor2_1 _26800_ (.A(net1731),
    .B(net5151),
    .Y(_19577_));
 sg13g2_a21oi_1 _26801_ (.A1(net5152),
    .A2(_19576_),
    .Y(_00259_),
    .B1(_19577_));
 sg13g2_and2_1 _26802_ (.A(\shift_reg[17] ),
    .B(net5437),
    .X(_19578_));
 sg13g2_a21oi_1 _26803_ (.A1(net1264),
    .A2(net5485),
    .Y(_19579_),
    .B1(_19578_));
 sg13g2_nor2_1 _26804_ (.A(net2161),
    .B(net5154),
    .Y(_19580_));
 sg13g2_a21oi_1 _26805_ (.A1(net5151),
    .A2(_19579_),
    .Y(_00260_),
    .B1(_19580_));
 sg13g2_and2_1 _26806_ (.A(\shift_reg[18] ),
    .B(net5436),
    .X(_19581_));
 sg13g2_a21oi_1 _26807_ (.A1(net1085),
    .A2(net5485),
    .Y(_19582_),
    .B1(_19581_));
 sg13g2_nor2_1 _26808_ (.A(net1500),
    .B(net5154),
    .Y(_19583_));
 sg13g2_a21oi_1 _26809_ (.A1(net5153),
    .A2(_19582_),
    .Y(_00261_),
    .B1(_19583_));
 sg13g2_and2_1 _26810_ (.A(\shift_reg[19] ),
    .B(net5436),
    .X(_19584_));
 sg13g2_a21oi_1 _26811_ (.A1(net1380),
    .A2(net5485),
    .Y(_19585_),
    .B1(_19584_));
 sg13g2_nor2_1 _26812_ (.A(net1900),
    .B(net5153),
    .Y(_19586_));
 sg13g2_a21oi_1 _26813_ (.A1(net5154),
    .A2(_19585_),
    .Y(_00262_),
    .B1(_19586_));
 sg13g2_and2_1 _26814_ (.A(net1962),
    .B(net5436),
    .X(_19587_));
 sg13g2_a21oi_1 _26815_ (.A1(net1080),
    .A2(net5485),
    .Y(_19588_),
    .B1(_19587_));
 sg13g2_nor2_1 _26816_ (.A(net2169),
    .B(net5153),
    .Y(_19589_));
 sg13g2_a21oi_1 _26817_ (.A1(net5151),
    .A2(_19588_),
    .Y(_00263_),
    .B1(_19589_));
 sg13g2_and2_1 _26818_ (.A(net2126),
    .B(net5436),
    .X(_19590_));
 sg13g2_a21oi_1 _26819_ (.A1(net1353),
    .A2(net5487),
    .Y(_19591_),
    .B1(_19590_));
 sg13g2_nor2_1 _26820_ (.A(net2631),
    .B(net5154),
    .Y(_19592_));
 sg13g2_a21oi_1 _26821_ (.A1(net5153),
    .A2(_19591_),
    .Y(_00264_),
    .B1(_19592_));
 sg13g2_and2_1 _26822_ (.A(net2028),
    .B(net5436),
    .X(_19593_));
 sg13g2_a21oi_1 _26823_ (.A1(net1372),
    .A2(net5485),
    .Y(_19594_),
    .B1(_19593_));
 sg13g2_nor2_1 _26824_ (.A(net2534),
    .B(net5153),
    .Y(_19595_));
 sg13g2_a21oi_1 _26825_ (.A1(net5153),
    .A2(_19594_),
    .Y(_00265_),
    .B1(_19595_));
 sg13g2_and2_1 _26826_ (.A(net1465),
    .B(net5436),
    .X(_19596_));
 sg13g2_a21oi_1 _26827_ (.A1(net1177),
    .A2(net5487),
    .Y(_19597_),
    .B1(_19596_));
 sg13g2_nor2_1 _26828_ (.A(net2350),
    .B(net5153),
    .Y(_19598_));
 sg13g2_a21oi_1 _26829_ (.A1(net5153),
    .A2(_19597_),
    .Y(_00266_),
    .B1(_19598_));
 sg13g2_and2_1 _26830_ (.A(net1731),
    .B(net5436),
    .X(_19599_));
 sg13g2_a21oi_1 _26831_ (.A1(net1087),
    .A2(net5487),
    .Y(_19600_),
    .B1(_19599_));
 sg13g2_nor2_1 _26832_ (.A(net2445),
    .B(net5159),
    .Y(_19601_));
 sg13g2_a21oi_1 _26833_ (.A1(net5159),
    .A2(_19600_),
    .Y(_00267_),
    .B1(_19601_));
 sg13g2_and2_1 _26834_ (.A(\shift_reg[25] ),
    .B(net5438),
    .X(_19602_));
 sg13g2_a21oi_1 _26835_ (.A1(\inv_result[17] ),
    .A2(net5490),
    .Y(_19603_),
    .B1(_19602_));
 sg13g2_nor2_1 _26836_ (.A(net1558),
    .B(net5159),
    .Y(_19604_));
 sg13g2_a21oi_1 _26837_ (.A1(net5162),
    .A2(_19603_),
    .Y(_00268_),
    .B1(_19604_));
 sg13g2_and2_1 _26838_ (.A(\shift_reg[26] ),
    .B(net5438),
    .X(_19605_));
 sg13g2_a21oi_1 _26839_ (.A1(net1076),
    .A2(net5493),
    .Y(_19606_),
    .B1(_19605_));
 sg13g2_nor2_1 _26840_ (.A(net1378),
    .B(net5164),
    .Y(_19607_));
 sg13g2_a21oi_1 _26841_ (.A1(net5164),
    .A2(_19606_),
    .Y(_00269_),
    .B1(_19607_));
 sg13g2_and2_1 _26842_ (.A(net1900),
    .B(net5441),
    .X(_19608_));
 sg13g2_a21oi_1 _26843_ (.A1(net1768),
    .A2(net5493),
    .Y(_19609_),
    .B1(_19608_));
 sg13g2_nor2_1 _26844_ (.A(net2103),
    .B(net5164),
    .Y(_19610_));
 sg13g2_a21oi_1 _26845_ (.A1(net5164),
    .A2(_19609_),
    .Y(_00270_),
    .B1(_19610_));
 sg13g2_and2_1 _26846_ (.A(\shift_reg[28] ),
    .B(net5441),
    .X(_19611_));
 sg13g2_a21oi_1 _26847_ (.A1(\inv_result[20] ),
    .A2(net5490),
    .Y(_19612_),
    .B1(_19611_));
 sg13g2_nor2_1 _26848_ (.A(net2075),
    .B(net5164),
    .Y(_19613_));
 sg13g2_a21oi_1 _26849_ (.A1(net5164),
    .A2(_19612_),
    .Y(_00271_),
    .B1(_19613_));
 sg13g2_and2_1 _26850_ (.A(\shift_reg[29] ),
    .B(net5443),
    .X(_19614_));
 sg13g2_a21oi_1 _26851_ (.A1(net1155),
    .A2(net5493),
    .Y(_19615_),
    .B1(_19614_));
 sg13g2_nor2_1 _26852_ (.A(net1449),
    .B(net5164),
    .Y(_19616_));
 sg13g2_a21oi_1 _26853_ (.A1(net5164),
    .A2(_19615_),
    .Y(_00272_),
    .B1(_19616_));
 sg13g2_and2_1 _26854_ (.A(\shift_reg[30] ),
    .B(net5443),
    .X(_19617_));
 sg13g2_a21oi_1 _26855_ (.A1(\inv_result[22] ),
    .A2(net5494),
    .Y(_19618_),
    .B1(_19617_));
 sg13g2_nor2_1 _26856_ (.A(net1354),
    .B(net5165),
    .Y(_19619_));
 sg13g2_a21oi_1 _26857_ (.A1(net5166),
    .A2(_19618_),
    .Y(_00273_),
    .B1(_19619_));
 sg13g2_and2_1 _26858_ (.A(net2350),
    .B(net5441),
    .X(_19620_));
 sg13g2_a21oi_1 _26859_ (.A1(net1228),
    .A2(net5493),
    .Y(_19621_),
    .B1(_19620_));
 sg13g2_nor2_1 _26860_ (.A(net2434),
    .B(net5165),
    .Y(_19622_));
 sg13g2_a21oi_1 _26861_ (.A1(net5166),
    .A2(_19621_),
    .Y(_00274_),
    .B1(_19622_));
 sg13g2_and2_1 _26862_ (.A(\shift_reg[32] ),
    .B(net5444),
    .X(_19623_));
 sg13g2_a21oi_1 _26863_ (.A1(net1262),
    .A2(net5493),
    .Y(_19624_),
    .B1(_19623_));
 sg13g2_nor2_1 _26864_ (.A(net2404),
    .B(net5166),
    .Y(_19625_));
 sg13g2_a21oi_1 _26865_ (.A1(net5166),
    .A2(_19624_),
    .Y(_00275_),
    .B1(_19625_));
 sg13g2_and2_1 _26866_ (.A(net1558),
    .B(net5443),
    .X(_19626_));
 sg13g2_a21oi_1 _26867_ (.A1(net1259),
    .A2(net5494),
    .Y(_19627_),
    .B1(_19626_));
 sg13g2_nor2_1 _26868_ (.A(net2721),
    .B(net5172),
    .Y(_19628_));
 sg13g2_a21oi_1 _26869_ (.A1(net5172),
    .A2(_19627_),
    .Y(_00276_),
    .B1(_19628_));
 sg13g2_and2_1 _26870_ (.A(net1378),
    .B(net5443),
    .X(_19629_));
 sg13g2_a21oi_1 _26871_ (.A1(net1175),
    .A2(net5494),
    .Y(_19630_),
    .B1(_19629_));
 sg13g2_nor2_1 _26872_ (.A(net1722),
    .B(net5172),
    .Y(_19631_));
 sg13g2_a21oi_1 _26873_ (.A1(net5172),
    .A2(_19630_),
    .Y(_00277_),
    .B1(_19631_));
 sg13g2_and2_1 _26874_ (.A(net2103),
    .B(net5443),
    .X(_19632_));
 sg13g2_a21oi_2 _26875_ (.B1(_19632_),
    .Y(_19633_),
    .A2(net5493),
    .A1(net2027));
 sg13g2_nor2_1 _26876_ (.A(net2144),
    .B(net5170),
    .Y(_19634_));
 sg13g2_a21oi_1 _26877_ (.A1(net5170),
    .A2(_19633_),
    .Y(_00278_),
    .B1(_19634_));
 sg13g2_and2_1 _26878_ (.A(\shift_reg[36] ),
    .B(net5443),
    .X(_19635_));
 sg13g2_a21oi_2 _26879_ (.B1(_19635_),
    .Y(_19636_),
    .A2(net5493),
    .A1(net1388));
 sg13g2_nor2_1 _26880_ (.A(net1865),
    .B(net5174),
    .Y(_19637_));
 sg13g2_a21oi_1 _26881_ (.A1(net5174),
    .A2(_19636_),
    .Y(_00279_),
    .B1(_19637_));
 sg13g2_and2_1 _26882_ (.A(net1449),
    .B(net5443),
    .X(_19638_));
 sg13g2_a21oi_1 _26883_ (.A1(net1339),
    .A2(net5493),
    .Y(_19639_),
    .B1(_19638_));
 sg13g2_nor2_1 _26884_ (.A(net2440),
    .B(net5172),
    .Y(_19640_));
 sg13g2_a21oi_1 _26885_ (.A1(net5172),
    .A2(_19639_),
    .Y(_00280_),
    .B1(_19640_));
 sg13g2_and2_1 _26886_ (.A(net1354),
    .B(net5444),
    .X(_19641_));
 sg13g2_a21oi_1 _26887_ (.A1(net1078),
    .A2(net5495),
    .Y(_19642_),
    .B1(_19641_));
 sg13g2_nor2_1 _26888_ (.A(net1721),
    .B(net5170),
    .Y(_19643_));
 sg13g2_a21oi_1 _26889_ (.A1(net5170),
    .A2(_19642_),
    .Y(_00281_),
    .B1(_19643_));
 sg13g2_and2_1 _26890_ (.A(\shift_reg[39] ),
    .B(net5445),
    .X(_19644_));
 sg13g2_a21oi_1 _26891_ (.A1(net1356),
    .A2(net5496),
    .Y(_19645_),
    .B1(_19644_));
 sg13g2_nor2_1 _26892_ (.A(net2312),
    .B(net5170),
    .Y(_19646_));
 sg13g2_a21oi_1 _26893_ (.A1(net5170),
    .A2(_19645_),
    .Y(_00282_),
    .B1(_19646_));
 sg13g2_and2_1 _26894_ (.A(\shift_reg[40] ),
    .B(net5446),
    .X(_19647_));
 sg13g2_a21oi_1 _26895_ (.A1(net1079),
    .A2(net5498),
    .Y(_19648_),
    .B1(_19647_));
 sg13g2_nor2_1 _26896_ (.A(net1967),
    .B(net5175),
    .Y(_19649_));
 sg13g2_a21oi_1 _26897_ (.A1(net5174),
    .A2(_19648_),
    .Y(_00283_),
    .B1(_19649_));
 sg13g2_and2_1 _26898_ (.A(\shift_reg[41] ),
    .B(net5448),
    .X(_19650_));
 sg13g2_a21oi_1 _26899_ (.A1(net1265),
    .A2(net5497),
    .Y(_19651_),
    .B1(_19650_));
 sg13g2_nor2_1 _26900_ (.A(net1310),
    .B(net5175),
    .Y(_19652_));
 sg13g2_a21oi_1 _26901_ (.A1(net5175),
    .A2(_19651_),
    .Y(_00284_),
    .B1(_19652_));
 sg13g2_and2_1 _26902_ (.A(\shift_reg[42] ),
    .B(net5445),
    .X(_19653_));
 sg13g2_a21oi_1 _26903_ (.A1(net1077),
    .A2(net5497),
    .Y(_19654_),
    .B1(_19653_));
 sg13g2_nor2_1 _26904_ (.A(net1516),
    .B(net5176),
    .Y(_19655_));
 sg13g2_a21oi_1 _26905_ (.A1(net5175),
    .A2(_19654_),
    .Y(_00285_),
    .B1(_19655_));
 sg13g2_and2_1 _26906_ (.A(\shift_reg[43] ),
    .B(net5448),
    .X(_19656_));
 sg13g2_a21oi_1 _26907_ (.A1(net1144),
    .A2(net5497),
    .Y(_19657_),
    .B1(_19656_));
 sg13g2_nor2_1 _26908_ (.A(net1416),
    .B(net5180),
    .Y(_19658_));
 sg13g2_a21oi_1 _26909_ (.A1(net5180),
    .A2(_19657_),
    .Y(_00286_),
    .B1(_19658_));
 sg13g2_and2_1 _26910_ (.A(net1865),
    .B(net5448),
    .X(_19659_));
 sg13g2_a21oi_1 _26911_ (.A1(net1171),
    .A2(net5497),
    .Y(_19660_),
    .B1(_19659_));
 sg13g2_nor2_1 _26912_ (.A(net2896),
    .B(net5175),
    .Y(_19661_));
 sg13g2_a21oi_1 _26913_ (.A1(net5175),
    .A2(_19660_),
    .Y(_00287_),
    .B1(_19661_));
 sg13g2_and2_1 _26914_ (.A(\shift_reg[45] ),
    .B(net5448),
    .X(_19662_));
 sg13g2_a21oi_1 _26915_ (.A1(net1352),
    .A2(net5500),
    .Y(_19663_),
    .B1(_19662_));
 sg13g2_nor2_1 _26916_ (.A(net2218),
    .B(net5180),
    .Y(_19664_));
 sg13g2_a21oi_1 _26917_ (.A1(net5180),
    .A2(_19663_),
    .Y(_00288_),
    .B1(_19664_));
 sg13g2_and2_1 _26918_ (.A(net1721),
    .B(net5448),
    .X(_19665_));
 sg13g2_a21oi_1 _26919_ (.A1(net1176),
    .A2(net5497),
    .Y(_19666_),
    .B1(_19665_));
 sg13g2_nor2_1 _26920_ (.A(net2245),
    .B(net5181),
    .Y(_19667_));
 sg13g2_a21oi_1 _26921_ (.A1(net5181),
    .A2(_19666_),
    .Y(_00289_),
    .B1(_19667_));
 sg13g2_and2_1 _26922_ (.A(net2312),
    .B(net5448),
    .X(_19668_));
 sg13g2_a21oi_1 _26923_ (.A1(net1188),
    .A2(net5497),
    .Y(_19669_),
    .B1(_19668_));
 sg13g2_nor2_1 _26924_ (.A(net2731),
    .B(net5175),
    .Y(_19670_));
 sg13g2_a21oi_1 _26925_ (.A1(net5175),
    .A2(_19669_),
    .Y(_00290_),
    .B1(_19670_));
 sg13g2_and2_1 _26926_ (.A(net1967),
    .B(net5448),
    .X(_19671_));
 sg13g2_a21oi_1 _26927_ (.A1(net1197),
    .A2(net5497),
    .Y(_19672_),
    .B1(_19671_));
 sg13g2_nor2_1 _26928_ (.A(net2819),
    .B(net5180),
    .Y(_19673_));
 sg13g2_a21oi_1 _26929_ (.A1(net5180),
    .A2(_19672_),
    .Y(_00291_),
    .B1(_19673_));
 sg13g2_and2_1 _26930_ (.A(net1310),
    .B(net5448),
    .X(_19674_));
 sg13g2_a21oi_1 _26931_ (.A1(net1246),
    .A2(net5500),
    .Y(_19675_),
    .B1(_19674_));
 sg13g2_nor2_1 _26932_ (.A(net2941),
    .B(net5180),
    .Y(_19676_));
 sg13g2_a21oi_1 _26933_ (.A1(net5180),
    .A2(_19675_),
    .Y(_00292_),
    .B1(_19676_));
 sg13g2_and2_1 _26934_ (.A(net1516),
    .B(net5451),
    .X(_19677_));
 sg13g2_a21oi_1 _26935_ (.A1(net1358),
    .A2(net5500),
    .Y(_19678_),
    .B1(_19677_));
 sg13g2_nor2_1 _26936_ (.A(net1660),
    .B(net5191),
    .Y(_19679_));
 sg13g2_a21oi_1 _26937_ (.A1(net5191),
    .A2(_19678_),
    .Y(_00293_),
    .B1(_19679_));
 sg13g2_and2_1 _26938_ (.A(net1416),
    .B(net5451),
    .X(_19680_));
 sg13g2_a21oi_1 _26939_ (.A1(net1306),
    .A2(net5500),
    .Y(_19681_),
    .B1(_19680_));
 sg13g2_nor2_1 _26940_ (.A(net1533),
    .B(net5191),
    .Y(_19682_));
 sg13g2_a21oi_1 _26941_ (.A1(net5191),
    .A2(_19681_),
    .Y(_00294_),
    .B1(_19682_));
 sg13g2_and2_1 _26942_ (.A(\shift_reg[52] ),
    .B(net5458),
    .X(_19683_));
 sg13g2_a21oi_1 _26943_ (.A1(net1290),
    .A2(net5503),
    .Y(_19684_),
    .B1(_19683_));
 sg13g2_nor2_1 _26944_ (.A(net1737),
    .B(net5192),
    .Y(_19685_));
 sg13g2_a21oi_1 _26945_ (.A1(net5191),
    .A2(_19684_),
    .Y(_00295_),
    .B1(_19685_));
 sg13g2_and2_1 _26946_ (.A(\shift_reg[53] ),
    .B(net5455),
    .X(_19686_));
 sg13g2_a21oi_1 _26947_ (.A1(net1178),
    .A2(net5507),
    .Y(_19687_),
    .B1(_19686_));
 sg13g2_nor2_1 _26948_ (.A(net1915),
    .B(net5192),
    .Y(_19688_));
 sg13g2_a21oi_1 _26949_ (.A1(net5192),
    .A2(_19687_),
    .Y(_00296_),
    .B1(_19688_));
 sg13g2_and2_1 _26950_ (.A(net2245),
    .B(net5458),
    .X(_19689_));
 sg13g2_a21oi_1 _26951_ (.A1(net1186),
    .A2(net5507),
    .Y(_19690_),
    .B1(_19689_));
 sg13g2_nor2_1 _26952_ (.A(net2556),
    .B(net5192),
    .Y(_19691_));
 sg13g2_a21oi_1 _26953_ (.A1(net5192),
    .A2(_19690_),
    .Y(_00297_),
    .B1(_19691_));
 sg13g2_and2_1 _26954_ (.A(\shift_reg[55] ),
    .B(net5455),
    .X(_19692_));
 sg13g2_a21oi_1 _26955_ (.A1(net1216),
    .A2(net5503),
    .Y(_19693_),
    .B1(_19692_));
 sg13g2_nor2_1 _26956_ (.A(net1952),
    .B(net5192),
    .Y(_19694_));
 sg13g2_a21oi_1 _26957_ (.A1(net5192),
    .A2(_19693_),
    .Y(_00298_),
    .B1(_19694_));
 sg13g2_and2_1 _26958_ (.A(\shift_reg[56] ),
    .B(net5458),
    .X(_19695_));
 sg13g2_a21oi_1 _26959_ (.A1(net1279),
    .A2(net5508),
    .Y(_19696_),
    .B1(_19695_));
 sg13g2_nor2_1 _26960_ (.A(net1479),
    .B(net5198),
    .Y(_19697_));
 sg13g2_a21oi_1 _26961_ (.A1(net5198),
    .A2(_19696_),
    .Y(_00299_),
    .B1(_19697_));
 sg13g2_and2_1 _26962_ (.A(\shift_reg[57] ),
    .B(net5460),
    .X(_19698_));
 sg13g2_a21oi_1 _26963_ (.A1(net1166),
    .A2(net5508),
    .Y(_19699_),
    .B1(_19698_));
 sg13g2_nor2_1 _26964_ (.A(net1463),
    .B(net5198),
    .Y(_19700_));
 sg13g2_a21oi_1 _26965_ (.A1(net5198),
    .A2(_19699_),
    .Y(_00300_),
    .B1(_19700_));
 sg13g2_and2_1 _26966_ (.A(net1660),
    .B(net5458),
    .X(_19701_));
 sg13g2_a21oi_1 _26967_ (.A1(net1299),
    .A2(net5509),
    .Y(_19702_),
    .B1(_19701_));
 sg13g2_nor2_1 _26968_ (.A(net2138),
    .B(net5197),
    .Y(_19703_));
 sg13g2_a21oi_1 _26969_ (.A1(net5197),
    .A2(_19702_),
    .Y(_00301_),
    .B1(_19703_));
 sg13g2_and2_1 _26970_ (.A(\shift_reg[59] ),
    .B(net5458),
    .X(_19704_));
 sg13g2_a21oi_1 _26971_ (.A1(net1147),
    .A2(net5508),
    .Y(_19705_),
    .B1(_19704_));
 sg13g2_nor2_1 _26972_ (.A(net1329),
    .B(net5198),
    .Y(_19706_));
 sg13g2_a21oi_1 _26973_ (.A1(net5198),
    .A2(_19705_),
    .Y(_00302_),
    .B1(_19706_));
 sg13g2_and2_1 _26974_ (.A(net1737),
    .B(net5458),
    .X(_19707_));
 sg13g2_a21oi_1 _26975_ (.A1(\inv_result[52] ),
    .A2(net5508),
    .Y(_19708_),
    .B1(_19707_));
 sg13g2_nor2_1 _26976_ (.A(net2073),
    .B(net5198),
    .Y(_19709_));
 sg13g2_a21oi_1 _26977_ (.A1(net5198),
    .A2(_19708_),
    .Y(_00303_),
    .B1(_19709_));
 sg13g2_and2_1 _26978_ (.A(\shift_reg[61] ),
    .B(net5458),
    .X(_19710_));
 sg13g2_a21oi_1 _26979_ (.A1(\inv_result[53] ),
    .A2(net5507),
    .Y(_19711_),
    .B1(_19710_));
 sg13g2_nor2_1 _26980_ (.A(net1853),
    .B(net5192),
    .Y(_19712_));
 sg13g2_a21oi_1 _26981_ (.A1(net5196),
    .A2(_19711_),
    .Y(_00304_),
    .B1(_19712_));
 sg13g2_and2_1 _26982_ (.A(\shift_reg[62] ),
    .B(net5460),
    .X(_19713_));
 sg13g2_a21oi_1 _26983_ (.A1(net1167),
    .A2(net5508),
    .Y(_19714_),
    .B1(_19713_));
 sg13g2_nor2_1 _26984_ (.A(net1510),
    .B(net5201),
    .Y(_19715_));
 sg13g2_a21oi_1 _26985_ (.A1(net5201),
    .A2(_19714_),
    .Y(_00305_),
    .B1(_19715_));
 sg13g2_and2_1 _26986_ (.A(\shift_reg[63] ),
    .B(net5458),
    .X(_19716_));
 sg13g2_a21oi_1 _26987_ (.A1(net1179),
    .A2(net5508),
    .Y(_19717_),
    .B1(_19716_));
 sg13g2_nor2_1 _26988_ (.A(net1810),
    .B(net5197),
    .Y(_19718_));
 sg13g2_a21oi_1 _26989_ (.A1(net5197),
    .A2(_19717_),
    .Y(_00306_),
    .B1(_19718_));
 sg13g2_and2_1 _26990_ (.A(net1479),
    .B(net5460),
    .X(_19719_));
 sg13g2_a21oi_1 _26991_ (.A1(net1090),
    .A2(net5508),
    .Y(_19720_),
    .B1(_19719_));
 sg13g2_nor2_1 _26992_ (.A(net2859),
    .B(net5197),
    .Y(_19721_));
 sg13g2_a21oi_1 _26993_ (.A1(net5197),
    .A2(_19720_),
    .Y(_00307_),
    .B1(_19721_));
 sg13g2_and2_1 _26994_ (.A(net1463),
    .B(net5460),
    .X(_19722_));
 sg13g2_a21oi_1 _26995_ (.A1(net1091),
    .A2(net5508),
    .Y(_19723_),
    .B1(_19722_));
 sg13g2_nor2_1 _26996_ (.A(net2897),
    .B(net5197),
    .Y(_19724_));
 sg13g2_a21oi_1 _26997_ (.A1(net5197),
    .A2(_19723_),
    .Y(_00308_),
    .B1(_19724_));
 sg13g2_and2_1 _26998_ (.A(net2138),
    .B(net5462),
    .X(_19725_));
 sg13g2_a21oi_1 _26999_ (.A1(net1084),
    .A2(net5510),
    .Y(_19726_),
    .B1(_19725_));
 sg13g2_nor2_1 _27000_ (.A(net2651),
    .B(net5205),
    .Y(_19727_));
 sg13g2_a21oi_1 _27001_ (.A1(net5205),
    .A2(_19726_),
    .Y(_00309_),
    .B1(_19727_));
 sg13g2_and2_1 _27002_ (.A(net1329),
    .B(net5460),
    .X(_19728_));
 sg13g2_a21oi_1 _27003_ (.A1(net1096),
    .A2(net5510),
    .Y(_19729_),
    .B1(_19728_));
 sg13g2_nor2_1 _27004_ (.A(net2168),
    .B(net5206),
    .Y(_19730_));
 sg13g2_a21oi_1 _27005_ (.A1(net5206),
    .A2(_19729_),
    .Y(_00310_),
    .B1(_19730_));
 sg13g2_and2_1 _27006_ (.A(net2073),
    .B(net5460),
    .X(_19731_));
 sg13g2_a21oi_1 _27007_ (.A1(net1086),
    .A2(net5510),
    .Y(_19732_),
    .B1(_19731_));
 sg13g2_nor2_1 _27008_ (.A(net2207),
    .B(net5205),
    .Y(_19733_));
 sg13g2_a21oi_1 _27009_ (.A1(net5205),
    .A2(_19732_),
    .Y(_00311_),
    .B1(_19733_));
 sg13g2_and2_1 _27010_ (.A(net1853),
    .B(net5460),
    .X(_19734_));
 sg13g2_a21oi_1 _27011_ (.A1(net1093),
    .A2(net5515),
    .Y(_19735_),
    .B1(_19734_));
 sg13g2_nor2_1 _27012_ (.A(net1923),
    .B(net5206),
    .Y(_19736_));
 sg13g2_a21oi_1 _27013_ (.A1(net5206),
    .A2(_19735_),
    .Y(_00312_),
    .B1(_19736_));
 sg13g2_and2_1 _27014_ (.A(net1510),
    .B(net5462),
    .X(_19737_));
 sg13g2_a21oi_1 _27015_ (.A1(net1219),
    .A2(net5510),
    .Y(_19738_),
    .B1(_19737_));
 sg13g2_nor2_1 _27016_ (.A(net2136),
    .B(net5205),
    .Y(_19739_));
 sg13g2_a21oi_1 _27017_ (.A1(net5205),
    .A2(_19738_),
    .Y(_00313_),
    .B1(_19739_));
 sg13g2_and2_1 _27018_ (.A(net1810),
    .B(net5462),
    .X(_19740_));
 sg13g2_a21oi_1 _27019_ (.A1(net1303),
    .A2(net5515),
    .Y(_19741_),
    .B1(_19740_));
 sg13g2_nor2_1 _27020_ (.A(net2551),
    .B(net5206),
    .Y(_19742_));
 sg13g2_a21oi_1 _27021_ (.A1(net5206),
    .A2(_19741_),
    .Y(_00314_),
    .B1(_19742_));
 sg13g2_and2_1 _27022_ (.A(\shift_reg[72] ),
    .B(net5466),
    .X(_19743_));
 sg13g2_a21oi_1 _27023_ (.A1(net1263),
    .A2(net5515),
    .Y(_19744_),
    .B1(_19743_));
 sg13g2_nor2_1 _27024_ (.A(net1903),
    .B(net5206),
    .Y(_19745_));
 sg13g2_a21oi_1 _27025_ (.A1(net5210),
    .A2(_19744_),
    .Y(_00315_),
    .B1(_19745_));
 sg13g2_and2_1 _27026_ (.A(\shift_reg[73] ),
    .B(net5468),
    .X(_19746_));
 sg13g2_a21oi_1 _27027_ (.A1(net1083),
    .A2(net5516),
    .Y(_19747_),
    .B1(_19746_));
 sg13g2_nor2_1 _27028_ (.A(net2742),
    .B(net5214),
    .Y(_19748_));
 sg13g2_a21oi_1 _27029_ (.A1(net5214),
    .A2(_19747_),
    .Y(_00316_),
    .B1(_19748_));
 sg13g2_and2_1 _27030_ (.A(\shift_reg[74] ),
    .B(net5468),
    .X(_19749_));
 sg13g2_a21oi_1 _27031_ (.A1(net1105),
    .A2(net5516),
    .Y(_19750_),
    .B1(_19749_));
 sg13g2_nor2_1 _27032_ (.A(net2310),
    .B(net5214),
    .Y(_19751_));
 sg13g2_a21oi_1 _27033_ (.A1(net5214),
    .A2(_19750_),
    .Y(_00317_),
    .B1(_19751_));
 sg13g2_and2_1 _27034_ (.A(net2168),
    .B(net5466),
    .X(_19752_));
 sg13g2_a21oi_1 _27035_ (.A1(net1081),
    .A2(net5515),
    .Y(_19753_),
    .B1(_19752_));
 sg13g2_nor2_1 _27036_ (.A(net2623),
    .B(net5206),
    .Y(_19754_));
 sg13g2_a21oi_1 _27037_ (.A1(net5210),
    .A2(_19753_),
    .Y(_00318_),
    .B1(_19754_));
 sg13g2_and2_1 _27038_ (.A(\shift_reg[76] ),
    .B(net5466),
    .X(_19755_));
 sg13g2_a21oi_1 _27039_ (.A1(net1128),
    .A2(net5516),
    .Y(_19756_),
    .B1(_19755_));
 sg13g2_nor2_1 _27040_ (.A(net1376),
    .B(net5215),
    .Y(_19757_));
 sg13g2_a21oi_1 _27041_ (.A1(net5215),
    .A2(_19756_),
    .Y(_00319_),
    .B1(_19757_));
 sg13g2_and2_1 _27042_ (.A(net1923),
    .B(net5466),
    .X(_19758_));
 sg13g2_a21oi_1 _27043_ (.A1(net1309),
    .A2(net5516),
    .Y(_19759_),
    .B1(_19758_));
 sg13g2_nor2_1 _27044_ (.A(net2037),
    .B(net5214),
    .Y(_19760_));
 sg13g2_a21oi_1 _27045_ (.A1(net5214),
    .A2(_19759_),
    .Y(_00320_),
    .B1(_19760_));
 sg13g2_and2_1 _27046_ (.A(\shift_reg[78] ),
    .B(net5466),
    .X(_19761_));
 sg13g2_a21oi_1 _27047_ (.A1(net1092),
    .A2(net5516),
    .Y(_19762_),
    .B1(_19761_));
 sg13g2_nor2_1 _27048_ (.A(net1492),
    .B(net5215),
    .Y(_19763_));
 sg13g2_a21oi_1 _27049_ (.A1(net5215),
    .A2(_19762_),
    .Y(_00321_),
    .B1(_19763_));
 sg13g2_and2_1 _27050_ (.A(\shift_reg[79] ),
    .B(net5468),
    .X(_19764_));
 sg13g2_a21oi_1 _27051_ (.A1(net1168),
    .A2(net5516),
    .Y(_19765_),
    .B1(_19764_));
 sg13g2_nor2_1 _27052_ (.A(net1395),
    .B(net5215),
    .Y(_19766_));
 sg13g2_a21oi_1 _27053_ (.A1(net5215),
    .A2(_19765_),
    .Y(_00322_),
    .B1(_19766_));
 sg13g2_and2_1 _27054_ (.A(net1903),
    .B(net5468),
    .X(_19767_));
 sg13g2_a21oi_1 _27055_ (.A1(net1126),
    .A2(net5516),
    .Y(_19768_),
    .B1(_19767_));
 sg13g2_nor2_1 _27056_ (.A(net2475),
    .B(net5215),
    .Y(_19769_));
 sg13g2_a21oi_1 _27057_ (.A1(net5218),
    .A2(_19768_),
    .Y(_00323_),
    .B1(_19769_));
 sg13g2_and2_1 _27058_ (.A(\shift_reg[81] ),
    .B(net5469),
    .X(_19770_));
 sg13g2_a21oi_1 _27059_ (.A1(net1526),
    .A2(net5522),
    .Y(_19771_),
    .B1(_19770_));
 sg13g2_nor2_1 _27060_ (.A(net2115),
    .B(net5220),
    .Y(_19772_));
 sg13g2_a21oi_1 _27061_ (.A1(net5220),
    .A2(_19771_),
    .Y(_00324_),
    .B1(_19772_));
 sg13g2_and2_1 _27062_ (.A(net2310),
    .B(net5469),
    .X(_19773_));
 sg13g2_a21oi_1 _27063_ (.A1(net1996),
    .A2(net5518),
    .Y(_19774_),
    .B1(_19773_));
 sg13g2_nor2_1 _27064_ (.A(net2454),
    .B(net5219),
    .Y(_19775_));
 sg13g2_a21oi_1 _27065_ (.A1(net5219),
    .A2(_19774_),
    .Y(_00325_),
    .B1(_19775_));
 sg13g2_and2_1 _27066_ (.A(\shift_reg[83] ),
    .B(net5469),
    .X(_19776_));
 sg13g2_a21oi_1 _27067_ (.A1(net1253),
    .A2(net5518),
    .Y(_19777_),
    .B1(_19776_));
 sg13g2_nor2_1 _27068_ (.A(net2374),
    .B(net5220),
    .Y(_19778_));
 sg13g2_a21oi_1 _27069_ (.A1(net5219),
    .A2(_19777_),
    .Y(_00326_),
    .B1(_19778_));
 sg13g2_and2_1 _27070_ (.A(net1376),
    .B(net5469),
    .X(_19779_));
 sg13g2_a21oi_1 _27071_ (.A1(net1143),
    .A2(net5518),
    .Y(_19780_),
    .B1(_19779_));
 sg13g2_nor2_1 _27072_ (.A(net2675),
    .B(net5220),
    .Y(_19781_));
 sg13g2_a21oi_1 _27073_ (.A1(net5219),
    .A2(_19780_),
    .Y(_00327_),
    .B1(_19781_));
 sg13g2_and2_1 _27074_ (.A(net2037),
    .B(net5469),
    .X(_19782_));
 sg13g2_a21oi_1 _27075_ (.A1(\inv_result[77] ),
    .A2(net5518),
    .Y(_19783_),
    .B1(_19782_));
 sg13g2_nor2_1 _27076_ (.A(net2400),
    .B(net5219),
    .Y(_19784_));
 sg13g2_a21oi_1 _27077_ (.A1(net5218),
    .A2(_19783_),
    .Y(_00328_),
    .B1(_19784_));
 sg13g2_and2_1 _27078_ (.A(net1492),
    .B(net5469),
    .X(_19785_));
 sg13g2_a21oi_1 _27079_ (.A1(net1207),
    .A2(net5518),
    .Y(_19786_),
    .B1(_19785_));
 sg13g2_nor2_1 _27080_ (.A(net2686),
    .B(net5216),
    .Y(_19787_));
 sg13g2_a21oi_1 _27081_ (.A1(net5215),
    .A2(_19786_),
    .Y(_00329_),
    .B1(_19787_));
 sg13g2_and2_1 _27082_ (.A(net1395),
    .B(net5469),
    .X(_19788_));
 sg13g2_a21oi_1 _27083_ (.A1(net1203),
    .A2(net5518),
    .Y(_19789_),
    .B1(_19788_));
 sg13g2_nor2_1 _27084_ (.A(net1775),
    .B(net5222),
    .Y(_19790_));
 sg13g2_a21oi_1 _27085_ (.A1(net5222),
    .A2(_19789_),
    .Y(_00330_),
    .B1(_19790_));
 sg13g2_and2_1 _27086_ (.A(\shift_reg[88] ),
    .B(net5471),
    .X(_19791_));
 sg13g2_a21oi_1 _27087_ (.A1(net1097),
    .A2(net5520),
    .Y(_19792_),
    .B1(_19791_));
 sg13g2_nor2_1 _27088_ (.A(net2230),
    .B(net5222),
    .Y(_19793_));
 sg13g2_a21oi_1 _27089_ (.A1(net5222),
    .A2(_19792_),
    .Y(_00331_),
    .B1(_19793_));
 sg13g2_and2_1 _27090_ (.A(net2115),
    .B(net5473),
    .X(_19794_));
 sg13g2_a21oi_1 _27091_ (.A1(net1832),
    .A2(net5521),
    .Y(_19795_),
    .B1(_19794_));
 sg13g2_nor2_1 _27092_ (.A(net2539),
    .B(net5223),
    .Y(_19796_));
 sg13g2_a21oi_1 _27093_ (.A1(net5223),
    .A2(_19795_),
    .Y(_00332_),
    .B1(_19796_));
 sg13g2_and2_1 _27094_ (.A(\shift_reg[90] ),
    .B(net5471),
    .X(_19797_));
 sg13g2_a21oi_1 _27095_ (.A1(net1282),
    .A2(net5520),
    .Y(_19798_),
    .B1(_19797_));
 sg13g2_nor2_1 _27096_ (.A(net1994),
    .B(net5221),
    .Y(_19799_));
 sg13g2_a21oi_1 _27097_ (.A1(net5221),
    .A2(_19798_),
    .Y(_00333_),
    .B1(_19799_));
 sg13g2_and2_1 _27098_ (.A(\shift_reg[91] ),
    .B(net5471),
    .X(_19800_));
 sg13g2_a21oi_1 _27099_ (.A1(\inv_result[83] ),
    .A2(net5520),
    .Y(_19801_),
    .B1(_19800_));
 sg13g2_nor2_1 _27100_ (.A(net1709),
    .B(net5221),
    .Y(_19802_));
 sg13g2_a21oi_1 _27101_ (.A1(net5221),
    .A2(_19801_),
    .Y(_00334_),
    .B1(_19802_));
 sg13g2_and2_1 _27102_ (.A(\shift_reg[92] ),
    .B(net5472),
    .X(_19803_));
 sg13g2_a21oi_1 _27103_ (.A1(net1152),
    .A2(net5521),
    .Y(_19804_),
    .B1(_19803_));
 sg13g2_nor2_1 _27104_ (.A(net2259),
    .B(net5221),
    .Y(_19805_));
 sg13g2_a21oi_1 _27105_ (.A1(net5221),
    .A2(_19804_),
    .Y(_00335_),
    .B1(_19805_));
 sg13g2_and2_1 _27106_ (.A(\shift_reg[93] ),
    .B(net5471),
    .X(_19806_));
 sg13g2_a21oi_1 _27107_ (.A1(net1387),
    .A2(net5521),
    .Y(_19807_),
    .B1(_19806_));
 sg13g2_nor2_1 _27108_ (.A(net2224),
    .B(net5224),
    .Y(_19808_));
 sg13g2_a21oi_1 _27109_ (.A1(net5224),
    .A2(_19807_),
    .Y(_00336_),
    .B1(_19808_));
 sg13g2_and2_1 _27110_ (.A(\shift_reg[94] ),
    .B(net5475),
    .X(_19809_));
 sg13g2_a21oi_1 _27111_ (.A1(net1266),
    .A2(net5524),
    .Y(_19810_),
    .B1(_19809_));
 sg13g2_nor2_1 _27112_ (.A(net1374),
    .B(net5224),
    .Y(_19811_));
 sg13g2_a21oi_1 _27113_ (.A1(net5224),
    .A2(_19810_),
    .Y(_00337_),
    .B1(_19811_));
 sg13g2_and2_1 _27114_ (.A(net1775),
    .B(net5471),
    .X(_19812_));
 sg13g2_a21oi_1 _27115_ (.A1(net1415),
    .A2(net5520),
    .Y(_19813_),
    .B1(_19812_));
 sg13g2_nor2_1 _27116_ (.A(net2223),
    .B(net5221),
    .Y(_19814_));
 sg13g2_a21oi_1 _27117_ (.A1(net5221),
    .A2(_19813_),
    .Y(_00338_),
    .B1(_19814_));
 sg13g2_and2_1 _27118_ (.A(\shift_reg[96] ),
    .B(net5472),
    .X(_19815_));
 sg13g2_a21oi_1 _27119_ (.A1(net1121),
    .A2(net5520),
    .Y(_19816_),
    .B1(_19815_));
 sg13g2_nor2_1 _27120_ (.A(net1950),
    .B(net5222),
    .Y(_19817_));
 sg13g2_a21oi_1 _27121_ (.A1(net5222),
    .A2(_19816_),
    .Y(_00339_),
    .B1(_19817_));
 sg13g2_and2_1 _27122_ (.A(\shift_reg[97] ),
    .B(net5472),
    .X(_19818_));
 sg13g2_a21oi_1 _27123_ (.A1(net1185),
    .A2(net5521),
    .Y(_19819_),
    .B1(_19818_));
 sg13g2_nor2_1 _27124_ (.A(net2094),
    .B(net5225),
    .Y(_19820_));
 sg13g2_a21oi_1 _27125_ (.A1(net5224),
    .A2(_19819_),
    .Y(_00340_),
    .B1(_19820_));
 sg13g2_and2_1 _27126_ (.A(net1994),
    .B(net5471),
    .X(_19821_));
 sg13g2_a21oi_1 _27127_ (.A1(net1367),
    .A2(net5520),
    .Y(_19822_),
    .B1(_19821_));
 sg13g2_nor2_1 _27128_ (.A(net2020),
    .B(net5224),
    .Y(_19823_));
 sg13g2_a21oi_1 _27129_ (.A1(net5225),
    .A2(_19822_),
    .Y(_00341_),
    .B1(_19823_));
 sg13g2_and2_1 _27130_ (.A(net1709),
    .B(net5472),
    .X(_19824_));
 sg13g2_a21oi_1 _27131_ (.A1(net1095),
    .A2(net5520),
    .Y(_19825_),
    .B1(_19824_));
 sg13g2_nor2_1 _27132_ (.A(net2333),
    .B(net5219),
    .Y(_19826_));
 sg13g2_a21oi_1 _27133_ (.A1(net5222),
    .A2(_19825_),
    .Y(_00342_),
    .B1(_19826_));
 sg13g2_and2_1 _27134_ (.A(\shift_reg[100] ),
    .B(net5471),
    .X(_19827_));
 sg13g2_a21oi_1 _27135_ (.A1(net1110),
    .A2(net5520),
    .Y(_19828_),
    .B1(_19827_));
 sg13g2_nor2_1 _27136_ (.A(net1988),
    .B(net5226),
    .Y(_19829_));
 sg13g2_a21oi_1 _27137_ (.A1(net5226),
    .A2(_19828_),
    .Y(_00343_),
    .B1(_19829_));
 sg13g2_and2_1 _27138_ (.A(\shift_reg[101] ),
    .B(net5474),
    .X(_19830_));
 sg13g2_a21oi_1 _27139_ (.A1(net1280),
    .A2(net5523),
    .Y(_19831_),
    .B1(_19830_));
 sg13g2_nor2_1 _27140_ (.A(net1936),
    .B(net5224),
    .Y(_19832_));
 sg13g2_a21oi_1 _27141_ (.A1(net5224),
    .A2(_19831_),
    .Y(_00344_),
    .B1(_19832_));
 sg13g2_and2_1 _27142_ (.A(net1374),
    .B(net5474),
    .X(_19833_));
 sg13g2_a21oi_1 _27143_ (.A1(net1184),
    .A2(net5524),
    .Y(_19834_),
    .B1(_19833_));
 sg13g2_nor2_1 _27144_ (.A(net2275),
    .B(net5225),
    .Y(_19835_));
 sg13g2_a21oi_1 _27145_ (.A1(net5225),
    .A2(_19834_),
    .Y(_00345_),
    .B1(_19835_));
 sg13g2_and2_1 _27146_ (.A(\shift_reg[103] ),
    .B(net5471),
    .X(_19836_));
 sg13g2_a21oi_1 _27147_ (.A1(net1433),
    .A2(net5523),
    .Y(_19837_),
    .B1(_19836_));
 sg13g2_nor2_1 _27148_ (.A(net2023),
    .B(net5226),
    .Y(_19838_));
 sg13g2_a21oi_1 _27149_ (.A1(net5226),
    .A2(_19837_),
    .Y(_00346_),
    .B1(_19838_));
 sg13g2_and2_1 _27150_ (.A(net1950),
    .B(net5473),
    .X(_01855_));
 sg13g2_a21oi_1 _27151_ (.A1(net1272),
    .A2(net5522),
    .Y(_01856_),
    .B1(_01855_));
 sg13g2_nor2_1 _27152_ (.A(net2100),
    .B(net5220),
    .Y(_01857_));
 sg13g2_a21oi_1 _27153_ (.A1(net5220),
    .A2(_01856_),
    .Y(_00347_),
    .B1(_01857_));
 sg13g2_and2_1 _27154_ (.A(\shift_reg[105] ),
    .B(net5474),
    .X(_01858_));
 sg13g2_a21oi_1 _27155_ (.A1(net1315),
    .A2(net5523),
    .Y(_01859_),
    .B1(_01858_));
 sg13g2_nor2_1 _27156_ (.A(net2010),
    .B(net5227),
    .Y(_01860_));
 sg13g2_a21oi_1 _27157_ (.A1(net5227),
    .A2(_01859_),
    .Y(_00348_),
    .B1(_01860_));
 sg13g2_and2_1 _27158_ (.A(\shift_reg[106] ),
    .B(net5474),
    .X(_01861_));
 sg13g2_a21oi_1 _27159_ (.A1(net1160),
    .A2(net5523),
    .Y(_01862_),
    .B1(_01861_));
 sg13g2_nor2_1 _27160_ (.A(net1733),
    .B(net5227),
    .Y(_01863_));
 sg13g2_a21oi_1 _27161_ (.A1(net5227),
    .A2(_01862_),
    .Y(_00349_),
    .B1(_01863_));
 sg13g2_and2_1 _27162_ (.A(\shift_reg[107] ),
    .B(net5473),
    .X(_01864_));
 sg13g2_a21oi_1 _27163_ (.A1(net1112),
    .A2(net5522),
    .Y(_01865_),
    .B1(_01864_));
 sg13g2_nor2_1 _27164_ (.A(net2004),
    .B(net5219),
    .Y(_01866_));
 sg13g2_a21oi_1 _27165_ (.A1(net5219),
    .A2(_01865_),
    .Y(_00350_),
    .B1(_01866_));
 sg13g2_and2_1 _27166_ (.A(\shift_reg[108] ),
    .B(net5474),
    .X(_01867_));
 sg13g2_a21oi_1 _27167_ (.A1(net1139),
    .A2(net5523),
    .Y(_01868_),
    .B1(_01867_));
 sg13g2_nor2_1 _27168_ (.A(net1584),
    .B(net5227),
    .Y(_01869_));
 sg13g2_a21oi_1 _27169_ (.A1(net5227),
    .A2(_01868_),
    .Y(_00351_),
    .B1(_01869_));
 sg13g2_and2_1 _27170_ (.A(net1936),
    .B(net5474),
    .X(_01870_));
 sg13g2_a21oi_1 _27171_ (.A1(net1300),
    .A2(net5523),
    .Y(_01871_),
    .B1(_01870_));
 sg13g2_nor2_1 _27172_ (.A(net2267),
    .B(net5218),
    .Y(_01872_));
 sg13g2_a21oi_1 _27173_ (.A1(net5216),
    .A2(_01871_),
    .Y(_00352_),
    .B1(_01872_));
 sg13g2_and2_1 _27174_ (.A(\shift_reg[110] ),
    .B(net5474),
    .X(_01873_));
 sg13g2_a21oi_1 _27175_ (.A1(net1268),
    .A2(net5523),
    .Y(_01874_),
    .B1(_01873_));
 sg13g2_nor2_1 _27176_ (.A(net1784),
    .B(net5227),
    .Y(_01875_));
 sg13g2_a21oi_1 _27177_ (.A1(net5227),
    .A2(_01874_),
    .Y(_00353_),
    .B1(_01875_));
 sg13g2_and2_1 _27178_ (.A(\shift_reg[111] ),
    .B(net5474),
    .X(_01876_));
 sg13g2_a21oi_1 _27179_ (.A1(net1213),
    .A2(net5523),
    .Y(_01877_),
    .B1(_01876_));
 sg13g2_nor2_1 _27180_ (.A(net1890),
    .B(net5216),
    .Y(_01878_));
 sg13g2_a21oi_1 _27181_ (.A1(net5216),
    .A2(_01877_),
    .Y(_00354_),
    .B1(_01878_));
 sg13g2_and2_1 _27182_ (.A(\shift_reg[112] ),
    .B(net5470),
    .X(_01879_));
 sg13g2_a21oi_1 _27183_ (.A1(net1304),
    .A2(net5518),
    .Y(_01880_),
    .B1(_01879_));
 sg13g2_nor2_1 _27184_ (.A(net1800),
    .B(net5216),
    .Y(_01881_));
 sg13g2_a21oi_1 _27185_ (.A1(net5216),
    .A2(_01880_),
    .Y(_00355_),
    .B1(_01881_));
 sg13g2_and2_1 _27186_ (.A(net2010),
    .B(net5470),
    .X(_01882_));
 sg13g2_a21oi_1 _27187_ (.A1(net1294),
    .A2(net5518),
    .Y(_01883_),
    .B1(_01882_));
 sg13g2_nor2_1 _27188_ (.A(net2165),
    .B(net5216),
    .Y(_01884_));
 sg13g2_a21oi_1 _27189_ (.A1(net5216),
    .A2(_01883_),
    .Y(_00356_),
    .B1(_01884_));
 sg13g2_and2_1 _27190_ (.A(net1733),
    .B(net5470),
    .X(_01885_));
 sg13g2_a21oi_1 _27191_ (.A1(net1316),
    .A2(net5519),
    .Y(_01886_),
    .B1(_01885_));
 sg13g2_nor2_1 _27192_ (.A(net2113),
    .B(net5217),
    .Y(_01887_));
 sg13g2_a21oi_1 _27193_ (.A1(net5217),
    .A2(_01886_),
    .Y(_00357_),
    .B1(_01887_));
 sg13g2_and2_1 _27194_ (.A(\shift_reg[115] ),
    .B(net5470),
    .X(_01888_));
 sg13g2_a21oi_1 _27195_ (.A1(\inv_result[107] ),
    .A2(net5519),
    .Y(_01889_),
    .B1(_01888_));
 sg13g2_nor2_1 _27196_ (.A(net1477),
    .B(net5213),
    .Y(_01890_));
 sg13g2_a21oi_1 _27197_ (.A1(net5213),
    .A2(_01889_),
    .Y(_00358_),
    .B1(_01890_));
 sg13g2_and2_1 _27198_ (.A(\shift_reg[116] ),
    .B(net5470),
    .X(_01891_));
 sg13g2_a21oi_1 _27199_ (.A1(net1373),
    .A2(net5519),
    .Y(_01892_),
    .B1(_01891_));
 sg13g2_nor2_1 _27200_ (.A(net1471),
    .B(net5217),
    .Y(_01893_));
 sg13g2_a21oi_1 _27201_ (.A1(net5217),
    .A2(_01892_),
    .Y(_00359_),
    .B1(_01893_));
 sg13g2_and2_1 _27202_ (.A(\shift_reg[117] ),
    .B(net5470),
    .X(_01894_));
 sg13g2_a21oi_1 _27203_ (.A1(\inv_result[109] ),
    .A2(net5519),
    .Y(_01895_),
    .B1(_01894_));
 sg13g2_nor2_1 _27204_ (.A(net1413),
    .B(net5217),
    .Y(_01896_));
 sg13g2_a21oi_1 _27205_ (.A1(net5217),
    .A2(_01895_),
    .Y(_00360_),
    .B1(_01896_));
 sg13g2_and2_1 _27206_ (.A(net1784),
    .B(net5470),
    .X(_01897_));
 sg13g2_a21oi_1 _27207_ (.A1(net1201),
    .A2(net5519),
    .Y(_01898_),
    .B1(_01897_));
 sg13g2_nor2_1 _27208_ (.A(net1964),
    .B(net5217),
    .Y(_01899_));
 sg13g2_a21oi_1 _27209_ (.A1(net5217),
    .A2(_01898_),
    .Y(_00361_),
    .B1(_01899_));
 sg13g2_and2_1 _27210_ (.A(\shift_reg[119] ),
    .B(net5469),
    .X(_01900_));
 sg13g2_a21oi_1 _27211_ (.A1(net1138),
    .A2(net5519),
    .Y(_01901_),
    .B1(_01900_));
 sg13g2_nor2_1 _27212_ (.A(net1389),
    .B(net5212),
    .Y(_01902_));
 sg13g2_a21oi_1 _27213_ (.A1(net5212),
    .A2(_01901_),
    .Y(_00362_),
    .B1(_01902_));
 sg13g2_and2_1 _27214_ (.A(net1800),
    .B(net5467),
    .X(_01903_));
 sg13g2_a21oi_1 _27215_ (.A1(net1191),
    .A2(net5517),
    .Y(_01904_),
    .B1(_01903_));
 sg13g2_nor2_1 _27216_ (.A(net2362),
    .B(net5213),
    .Y(_01905_));
 sg13g2_a21oi_1 _27217_ (.A1(net5213),
    .A2(_01904_),
    .Y(_00363_),
    .B1(_01905_));
 sg13g2_and2_1 _27218_ (.A(net2165),
    .B(net5467),
    .X(_01906_));
 sg13g2_a21oi_1 _27219_ (.A1(net1169),
    .A2(net5517),
    .Y(_01907_),
    .B1(_01906_));
 sg13g2_nor2_1 _27220_ (.A(net2200),
    .B(net5213),
    .Y(_01908_));
 sg13g2_a21oi_1 _27221_ (.A1(net5213),
    .A2(_01907_),
    .Y(_00364_),
    .B1(_01908_));
 sg13g2_and2_1 _27222_ (.A(\shift_reg[122] ),
    .B(net5467),
    .X(_01909_));
 sg13g2_a21oi_1 _27223_ (.A1(net1277),
    .A2(net5517),
    .Y(_01910_),
    .B1(_01909_));
 sg13g2_nor2_1 _27224_ (.A(net1790),
    .B(net5211),
    .Y(_01911_));
 sg13g2_a21oi_1 _27225_ (.A1(net5211),
    .A2(_01910_),
    .Y(_00365_),
    .B1(_01911_));
 sg13g2_and2_1 _27226_ (.A(net1477),
    .B(net5468),
    .X(_01912_));
 sg13g2_a21oi_1 _27227_ (.A1(net1252),
    .A2(net5517),
    .Y(_01913_),
    .B1(_01912_));
 sg13g2_nor2_1 _27228_ (.A(net2222),
    .B(net5212),
    .Y(_01914_));
 sg13g2_a21oi_1 _27229_ (.A1(net5212),
    .A2(_01913_),
    .Y(_00366_),
    .B1(_01914_));
 sg13g2_and2_1 _27230_ (.A(net1471),
    .B(net5467),
    .X(_01915_));
 sg13g2_a21oi_1 _27231_ (.A1(net1410),
    .A2(net5517),
    .Y(_01916_),
    .B1(_01915_));
 sg13g2_nor2_1 _27232_ (.A(net1959),
    .B(net5211),
    .Y(_01917_));
 sg13g2_a21oi_1 _27233_ (.A1(net5211),
    .A2(_01916_),
    .Y(_00367_),
    .B1(_01917_));
 sg13g2_and2_1 _27234_ (.A(net1413),
    .B(net5467),
    .X(_01918_));
 sg13g2_a21oi_1 _27235_ (.A1(net1350),
    .A2(net5517),
    .Y(_01919_),
    .B1(_01918_));
 sg13g2_nor2_1 _27236_ (.A(net2155),
    .B(net5211),
    .Y(_01920_));
 sg13g2_a21oi_1 _27237_ (.A1(net5211),
    .A2(_01919_),
    .Y(_00368_),
    .B1(_01920_));
 sg13g2_and2_1 _27238_ (.A(\shift_reg[126] ),
    .B(net5467),
    .X(_01921_));
 sg13g2_a21oi_1 _27239_ (.A1(net1333),
    .A2(net5514),
    .Y(_01922_),
    .B1(_01921_));
 sg13g2_nor2_1 _27240_ (.A(net1398),
    .B(net5209),
    .Y(_01923_));
 sg13g2_a21oi_1 _27241_ (.A1(net5209),
    .A2(_01922_),
    .Y(_00369_),
    .B1(_01923_));
 sg13g2_and2_1 _27242_ (.A(net1389),
    .B(net5467),
    .X(_01924_));
 sg13g2_a21oi_1 _27243_ (.A1(net1418),
    .A2(net5516),
    .Y(_01925_),
    .B1(_01924_));
 sg13g2_nor2_1 _27244_ (.A(net1701),
    .B(net5211),
    .Y(_01926_));
 sg13g2_a21oi_1 _27245_ (.A1(net5211),
    .A2(_01925_),
    .Y(_00370_),
    .B1(_01926_));
 sg13g2_and2_1 _27246_ (.A(\shift_reg[128] ),
    .B(net5465),
    .X(_01927_));
 sg13g2_a21oi_1 _27247_ (.A1(net1187),
    .A2(net5514),
    .Y(_01928_),
    .B1(_01927_));
 sg13g2_nor2_1 _27248_ (.A(net1938),
    .B(net5209),
    .Y(_01929_));
 sg13g2_a21oi_1 _27249_ (.A1(net5210),
    .A2(_01928_),
    .Y(_00371_),
    .B1(_01929_));
 sg13g2_and2_1 _27250_ (.A(\shift_reg[129] ),
    .B(net5465),
    .X(_01930_));
 sg13g2_a21oi_1 _27251_ (.A1(\inv_result[121] ),
    .A2(net5513),
    .Y(_01931_),
    .B1(_01930_));
 sg13g2_nor2_1 _27252_ (.A(net2044),
    .B(net5207),
    .Y(_01932_));
 sg13g2_a21oi_1 _27253_ (.A1(net5208),
    .A2(_01931_),
    .Y(_00372_),
    .B1(_01932_));
 sg13g2_and2_1 _27254_ (.A(net1790),
    .B(net5467),
    .X(_01933_));
 sg13g2_a21oi_1 _27255_ (.A1(net1497),
    .A2(net5514),
    .Y(_01934_),
    .B1(_01933_));
 sg13g2_nor2_1 _27256_ (.A(net2432),
    .B(net5209),
    .Y(_01935_));
 sg13g2_a21oi_1 _27257_ (.A1(net5210),
    .A2(_01934_),
    .Y(_00373_),
    .B1(_01935_));
 sg13g2_and2_1 _27258_ (.A(net2222),
    .B(net5465),
    .X(_01936_));
 sg13g2_a21oi_1 _27259_ (.A1(net1624),
    .A2(net5514),
    .Y(_01937_),
    .B1(_01936_));
 sg13g2_nor2_1 _27260_ (.A(net2367),
    .B(net5207),
    .Y(_01938_));
 sg13g2_a21oi_1 _27261_ (.A1(net5207),
    .A2(_01937_),
    .Y(_00374_),
    .B1(_01938_));
 sg13g2_and2_1 _27262_ (.A(net1959),
    .B(net5465),
    .X(_01939_));
 sg13g2_a21oi_1 _27263_ (.A1(net1198),
    .A2(net5514),
    .Y(_01940_),
    .B1(_01939_));
 sg13g2_nor2_1 _27264_ (.A(net2184),
    .B(net5208),
    .Y(_01941_));
 sg13g2_a21oi_1 _27265_ (.A1(net5208),
    .A2(_01940_),
    .Y(_00375_),
    .B1(_01941_));
 sg13g2_and2_1 _27266_ (.A(\shift_reg[133] ),
    .B(net5464),
    .X(_01942_));
 sg13g2_a21oi_1 _27267_ (.A1(net1317),
    .A2(net5513),
    .Y(_01943_),
    .B1(_01942_));
 sg13g2_nor2_1 _27268_ (.A(net2128),
    .B(net5207),
    .Y(_01944_));
 sg13g2_a21oi_1 _27269_ (.A1(net5207),
    .A2(_01943_),
    .Y(_00376_),
    .B1(_01944_));
 sg13g2_and2_1 _27270_ (.A(net1398),
    .B(net5465),
    .X(_01945_));
 sg13g2_a21oi_1 _27271_ (.A1(net2141),
    .A2(net5514),
    .Y(_01946_),
    .B1(_01945_));
 sg13g2_nor2_1 _27272_ (.A(net2291),
    .B(net5209),
    .Y(_01947_));
 sg13g2_a21oi_1 _27273_ (.A1(net5209),
    .A2(_01946_),
    .Y(_00377_),
    .B1(_01947_));
 sg13g2_and2_1 _27274_ (.A(net1701),
    .B(net5464),
    .X(_01948_));
 sg13g2_a21oi_1 _27275_ (.A1(net1831),
    .A2(net5513),
    .Y(_01949_),
    .B1(_01948_));
 sg13g2_nor2_1 _27276_ (.A(net2386),
    .B(net5207),
    .Y(_01950_));
 sg13g2_a21oi_1 _27277_ (.A1(net5208),
    .A2(_01949_),
    .Y(_00378_),
    .B1(_01950_));
 sg13g2_and2_1 _27278_ (.A(\shift_reg[136] ),
    .B(net5464),
    .X(_01951_));
 sg13g2_a21oi_1 _27279_ (.A1(\inv_result[128] ),
    .A2(net5513),
    .Y(_01952_),
    .B1(_01951_));
 sg13g2_nor2_1 _27280_ (.A(net1361),
    .B(net5207),
    .Y(_01953_));
 sg13g2_a21oi_1 _27281_ (.A1(net5207),
    .A2(_01952_),
    .Y(_00379_),
    .B1(_01953_));
 sg13g2_and2_1 _27282_ (.A(\shift_reg[137] ),
    .B(net5464),
    .X(_01954_));
 sg13g2_a21oi_1 _27283_ (.A1(net1382),
    .A2(net5513),
    .Y(_01955_),
    .B1(_01954_));
 sg13g2_nor2_1 _27284_ (.A(net1670),
    .B(net5203),
    .Y(_01956_));
 sg13g2_a21oi_1 _27285_ (.A1(net5203),
    .A2(_01955_),
    .Y(_00380_),
    .B1(_01956_));
 sg13g2_and2_1 _27286_ (.A(\shift_reg[138] ),
    .B(net5461),
    .X(_01957_));
 sg13g2_a21oi_1 _27287_ (.A1(\inv_result[130] ),
    .A2(net5510),
    .Y(_01958_),
    .B1(_01957_));
 sg13g2_nor2_1 _27288_ (.A(net1566),
    .B(net5203),
    .Y(_01959_));
 sg13g2_a21oi_1 _27289_ (.A1(net5203),
    .A2(_01958_),
    .Y(_00381_),
    .B1(_01959_));
 sg13g2_and2_1 _27290_ (.A(\shift_reg[139] ),
    .B(net5464),
    .X(_01960_));
 sg13g2_a21oi_1 _27291_ (.A1(\inv_result[131] ),
    .A2(net5513),
    .Y(_01961_),
    .B1(_01960_));
 sg13g2_nor2_1 _27292_ (.A(net1946),
    .B(net5203),
    .Y(_01962_));
 sg13g2_a21oi_1 _27293_ (.A1(net5203),
    .A2(_01961_),
    .Y(_00382_),
    .B1(_01962_));
 sg13g2_and2_1 _27294_ (.A(\shift_reg[140] ),
    .B(net5464),
    .X(_01963_));
 sg13g2_a21oi_1 _27295_ (.A1(net1772),
    .A2(net5513),
    .Y(_01964_),
    .B1(_01963_));
 sg13g2_nor2_1 _27296_ (.A(net2142),
    .B(net5203),
    .Y(_01965_));
 sg13g2_a21oi_1 _27297_ (.A1(net5203),
    .A2(_01964_),
    .Y(_00383_),
    .B1(_01965_));
 sg13g2_and2_1 _27298_ (.A(\shift_reg[141] ),
    .B(net5464),
    .X(_01966_));
 sg13g2_a21oi_1 _27299_ (.A1(net1258),
    .A2(net5513),
    .Y(_01967_),
    .B1(_01966_));
 sg13g2_nor2_1 _27300_ (.A(net1871),
    .B(net5204),
    .Y(_01968_));
 sg13g2_a21oi_1 _27301_ (.A1(net5204),
    .A2(_01967_),
    .Y(_00384_),
    .B1(_01968_));
 sg13g2_and2_1 _27302_ (.A(\shift_reg[142] ),
    .B(net5461),
    .X(_01969_));
 sg13g2_a21oi_1 _27303_ (.A1(net1628),
    .A2(net5510),
    .Y(_01970_),
    .B1(_01969_));
 sg13g2_nor2_1 _27304_ (.A(net2232),
    .B(net5202),
    .Y(_01971_));
 sg13g2_a21oi_1 _27305_ (.A1(net5202),
    .A2(_01970_),
    .Y(_00385_),
    .B1(_01971_));
 sg13g2_and2_1 _27306_ (.A(net2386),
    .B(net5461),
    .X(_01972_));
 sg13g2_a21oi_1 _27307_ (.A1(net1645),
    .A2(net5510),
    .Y(_01973_),
    .B1(_01972_));
 sg13g2_nor2_1 _27308_ (.A(net2568),
    .B(net5202),
    .Y(_01974_));
 sg13g2_a21oi_1 _27309_ (.A1(net5202),
    .A2(_01973_),
    .Y(_00386_),
    .B1(_01974_));
 sg13g2_and2_1 _27310_ (.A(net1361),
    .B(net5464),
    .X(_01975_));
 sg13g2_a21oi_1 _27311_ (.A1(net1730),
    .A2(net5511),
    .Y(_01976_),
    .B1(_01975_));
 sg13g2_nor2_1 _27312_ (.A(net2380),
    .B(net5204),
    .Y(_01977_));
 sg13g2_a21oi_1 _27313_ (.A1(net5204),
    .A2(_01976_),
    .Y(_00387_),
    .B1(_01977_));
 sg13g2_and2_1 _27314_ (.A(net1670),
    .B(net5461),
    .X(_01978_));
 sg13g2_a21oi_1 _27315_ (.A1(\inv_result[137] ),
    .A2(net5511),
    .Y(_01979_),
    .B1(_01978_));
 sg13g2_nor2_1 _27316_ (.A(net1898),
    .B(net5202),
    .Y(_01980_));
 sg13g2_a21oi_1 _27317_ (.A1(net5202),
    .A2(_01979_),
    .Y(_00388_),
    .B1(_01980_));
 sg13g2_and2_1 _27318_ (.A(net1566),
    .B(net5461),
    .X(_01981_));
 sg13g2_a21oi_1 _27319_ (.A1(net2043),
    .A2(net5510),
    .Y(_01982_),
    .B1(_01981_));
 sg13g2_nor2_1 _27320_ (.A(net2518),
    .B(net5202),
    .Y(_01983_));
 sg13g2_a21oi_1 _27321_ (.A1(net5202),
    .A2(_01982_),
    .Y(_00389_),
    .B1(_01983_));
 sg13g2_and2_1 _27322_ (.A(\shift_reg[147] ),
    .B(net5462),
    .X(_01984_));
 sg13g2_a21oi_1 _27323_ (.A1(\inv_result[139] ),
    .A2(net5511),
    .Y(_01985_),
    .B1(_01984_));
 sg13g2_nor2_1 _27324_ (.A(net1766),
    .B(net5200),
    .Y(_01986_));
 sg13g2_a21oi_1 _27325_ (.A1(net5200),
    .A2(_01985_),
    .Y(_00390_),
    .B1(_01986_));
 sg13g2_and2_1 _27326_ (.A(net2142),
    .B(net5461),
    .X(_01987_));
 sg13g2_a21oi_1 _27327_ (.A1(net1189),
    .A2(net5511),
    .Y(_01988_),
    .B1(_01987_));
 sg13g2_nor2_1 _27328_ (.A(net2226),
    .B(net5200),
    .Y(_01989_));
 sg13g2_a21oi_1 _27329_ (.A1(net5200),
    .A2(_01988_),
    .Y(_00391_),
    .B1(_01989_));
 sg13g2_and2_1 _27330_ (.A(\shift_reg[149] ),
    .B(net5461),
    .X(_01990_));
 sg13g2_a21oi_1 _27331_ (.A1(\inv_result[141] ),
    .A2(net5509),
    .Y(_01991_),
    .B1(_01990_));
 sg13g2_nor2_1 _27332_ (.A(net1445),
    .B(net5199),
    .Y(_01992_));
 sg13g2_a21oi_1 _27333_ (.A1(net5199),
    .A2(_01991_),
    .Y(_00392_),
    .B1(_01992_));
 sg13g2_and2_1 _27334_ (.A(\shift_reg[150] ),
    .B(net5463),
    .X(_01993_));
 sg13g2_a21oi_1 _27335_ (.A1(net1338),
    .A2(net5509),
    .Y(_01994_),
    .B1(_01993_));
 sg13g2_nor2_1 _27336_ (.A(net2053),
    .B(net5199),
    .Y(_01995_));
 sg13g2_a21oi_1 _27337_ (.A1(net5199),
    .A2(_01994_),
    .Y(_00393_),
    .B1(_01995_));
 sg13g2_and2_1 _27338_ (.A(\shift_reg[151] ),
    .B(net5460),
    .X(_01996_));
 sg13g2_a21oi_1 _27339_ (.A1(net1305),
    .A2(net5509),
    .Y(_01997_),
    .B1(_01996_));
 sg13g2_nor2_1 _27340_ (.A(net1400),
    .B(net5199),
    .Y(_01998_));
 sg13g2_a21oi_1 _27341_ (.A1(net5199),
    .A2(_01997_),
    .Y(_00394_),
    .B1(_01998_));
 sg13g2_and2_1 _27342_ (.A(\shift_reg[152] ),
    .B(net5461),
    .X(_01999_));
 sg13g2_a21oi_1 _27343_ (.A1(net1190),
    .A2(net5509),
    .Y(_02000_),
    .B1(_01999_));
 sg13g2_nor2_1 _27344_ (.A(net2194),
    .B(net5199),
    .Y(_02001_));
 sg13g2_a21oi_1 _27345_ (.A1(net5199),
    .A2(_02000_),
    .Y(_00395_),
    .B1(_02001_));
 sg13g2_and2_1 _27346_ (.A(net1898),
    .B(net5463),
    .X(_02002_));
 sg13g2_a21oi_1 _27347_ (.A1(net1236),
    .A2(net5509),
    .Y(_02003_),
    .B1(_02002_));
 sg13g2_nor2_1 _27348_ (.A(net2188),
    .B(net5200),
    .Y(_02004_));
 sg13g2_a21oi_1 _27349_ (.A1(net5200),
    .A2(_02003_),
    .Y(_00396_),
    .B1(_02004_));
 sg13g2_and2_1 _27350_ (.A(\shift_reg[154] ),
    .B(net5456),
    .X(_02005_));
 sg13g2_a21oi_1 _27351_ (.A1(net1202),
    .A2(net5505),
    .Y(_02006_),
    .B1(_02005_));
 sg13g2_nor2_1 _27352_ (.A(net1408),
    .B(net5195),
    .Y(_02007_));
 sg13g2_a21oi_1 _27353_ (.A1(net5195),
    .A2(_02006_),
    .Y(_00397_),
    .B1(_02007_));
 sg13g2_and2_1 _27354_ (.A(\shift_reg[155] ),
    .B(net5457),
    .X(_02008_));
 sg13g2_a21oi_1 _27355_ (.A1(net1165),
    .A2(net5506),
    .Y(_02009_),
    .B1(_02008_));
 sg13g2_nor2_1 _27356_ (.A(net1307),
    .B(net5195),
    .Y(_02010_));
 sg13g2_a21oi_1 _27357_ (.A1(net5195),
    .A2(_02009_),
    .Y(_00398_),
    .B1(_02010_));
 sg13g2_and2_1 _27358_ (.A(\shift_reg[156] ),
    .B(net5456),
    .X(_02011_));
 sg13g2_a21oi_1 _27359_ (.A1(net1761),
    .A2(net5506),
    .Y(_02012_),
    .B1(_02011_));
 sg13g2_nor2_1 _27360_ (.A(net1867),
    .B(net5194),
    .Y(_02013_));
 sg13g2_a21oi_1 _27361_ (.A1(net5194),
    .A2(_02012_),
    .Y(_00399_),
    .B1(_02013_));
 sg13g2_and2_1 _27362_ (.A(net1445),
    .B(net5457),
    .X(_02014_));
 sg13g2_a21oi_1 _27363_ (.A1(net1319),
    .A2(net5506),
    .Y(_02015_),
    .B1(_02014_));
 sg13g2_nor2_1 _27364_ (.A(net1998),
    .B(net5194),
    .Y(_02016_));
 sg13g2_a21oi_1 _27365_ (.A1(net5194),
    .A2(_02015_),
    .Y(_00400_),
    .B1(_02016_));
 sg13g2_and2_1 _27366_ (.A(\shift_reg[158] ),
    .B(net5456),
    .X(_02017_));
 sg13g2_a21oi_1 _27367_ (.A1(net1220),
    .A2(net5506),
    .Y(_02018_),
    .B1(_02017_));
 sg13g2_nor2_1 _27368_ (.A(net1391),
    .B(net5193),
    .Y(_02019_));
 sg13g2_a21oi_1 _27369_ (.A1(net5193),
    .A2(_02018_),
    .Y(_00401_),
    .B1(_02019_));
 sg13g2_and2_1 _27370_ (.A(net1400),
    .B(net5463),
    .X(_02020_));
 sg13g2_a21oi_1 _27371_ (.A1(net1335),
    .A2(net5505),
    .Y(_02021_),
    .B1(_02020_));
 sg13g2_nor2_1 _27372_ (.A(net2167),
    .B(net5195),
    .Y(_02022_));
 sg13g2_a21oi_1 _27373_ (.A1(net5195),
    .A2(_02021_),
    .Y(_00402_),
    .B1(_02022_));
 sg13g2_and2_1 _27374_ (.A(net2194),
    .B(net5457),
    .X(_02023_));
 sg13g2_a21oi_1 _27375_ (.A1(net1107),
    .A2(net5506),
    .Y(_02024_),
    .B1(_02023_));
 sg13g2_nor2_1 _27376_ (.A(net2272),
    .B(net5193),
    .Y(_02025_));
 sg13g2_a21oi_1 _27377_ (.A1(net5193),
    .A2(_02024_),
    .Y(_00403_),
    .B1(_02025_));
 sg13g2_and2_1 _27378_ (.A(\shift_reg[161] ),
    .B(net5457),
    .X(_02026_));
 sg13g2_a21oi_1 _27379_ (.A1(net1102),
    .A2(net5505),
    .Y(_02027_),
    .B1(_02026_));
 sg13g2_nor2_1 _27380_ (.A(net2081),
    .B(net5193),
    .Y(_02028_));
 sg13g2_a21oi_1 _27381_ (.A1(net5193),
    .A2(_02027_),
    .Y(_00404_),
    .B1(_02028_));
 sg13g2_and2_1 _27382_ (.A(net1408),
    .B(net5456),
    .X(_02029_));
 sg13g2_a21oi_1 _27383_ (.A1(net1221),
    .A2(net5505),
    .Y(_02030_),
    .B1(_02029_));
 sg13g2_nor2_1 _27384_ (.A(net2339),
    .B(net5193),
    .Y(_02031_));
 sg13g2_a21oi_1 _27385_ (.A1(net5193),
    .A2(_02030_),
    .Y(_00405_),
    .B1(_02031_));
 sg13g2_and2_1 _27386_ (.A(net1307),
    .B(net5456),
    .X(_02032_));
 sg13g2_a21oi_1 _27387_ (.A1(\inv_result[155] ),
    .A2(net5505),
    .Y(_02033_),
    .B1(_02032_));
 sg13g2_nor2_1 _27388_ (.A(net2012),
    .B(net5188),
    .Y(_02034_));
 sg13g2_a21oi_1 _27389_ (.A1(net5188),
    .A2(_02033_),
    .Y(_00406_),
    .B1(_02034_));
 sg13g2_and2_1 _27390_ (.A(net1867),
    .B(net5456),
    .X(_02035_));
 sg13g2_a21oi_1 _27391_ (.A1(net1256),
    .A2(net5505),
    .Y(_02036_),
    .B1(_02035_));
 sg13g2_nor2_1 _27392_ (.A(net1902),
    .B(net5188),
    .Y(_02037_));
 sg13g2_a21oi_1 _27393_ (.A1(net5189),
    .A2(_02036_),
    .Y(_00407_),
    .B1(_02037_));
 sg13g2_and2_1 _27394_ (.A(net1998),
    .B(net5456),
    .X(_02038_));
 sg13g2_a21oi_1 _27395_ (.A1(net2132),
    .A2(net5505),
    .Y(_02039_),
    .B1(_02038_));
 sg13g2_nor2_1 _27396_ (.A(net2340),
    .B(net5188),
    .Y(_02040_));
 sg13g2_a21oi_1 _27397_ (.A1(net5188),
    .A2(_02039_),
    .Y(_00408_),
    .B1(_02040_));
 sg13g2_and2_1 _27398_ (.A(net1391),
    .B(net5456),
    .X(_02041_));
 sg13g2_a21oi_1 _27399_ (.A1(net1254),
    .A2(net5505),
    .Y(_02042_),
    .B1(_02041_));
 sg13g2_nor2_1 _27400_ (.A(net2058),
    .B(net5187),
    .Y(_02043_));
 sg13g2_a21oi_1 _27401_ (.A1(net5190),
    .A2(_02042_),
    .Y(_00409_),
    .B1(_02043_));
 sg13g2_and2_1 _27402_ (.A(net2167),
    .B(net5454),
    .X(_02044_));
 sg13g2_a21oi_1 _27403_ (.A1(net1322),
    .A2(net5503),
    .Y(_02045_),
    .B1(_02044_));
 sg13g2_nor2_1 _27404_ (.A(net2357),
    .B(net5189),
    .Y(_02046_));
 sg13g2_a21oi_1 _27405_ (.A1(net5189),
    .A2(_02045_),
    .Y(_00410_),
    .B1(_02046_));
 sg13g2_and2_1 _27406_ (.A(\shift_reg[168] ),
    .B(net5455),
    .X(_02047_));
 sg13g2_a21oi_1 _27407_ (.A1(net1088),
    .A2(net5503),
    .Y(_02048_),
    .B1(_02047_));
 sg13g2_nor2_1 _27408_ (.A(net1762),
    .B(net5188),
    .Y(_02049_));
 sg13g2_a21oi_1 _27409_ (.A1(net5188),
    .A2(_02048_),
    .Y(_00411_),
    .B1(_02049_));
 sg13g2_and2_1 _27410_ (.A(\shift_reg[169] ),
    .B(net5455),
    .X(_02050_));
 sg13g2_a21oi_1 _27411_ (.A1(net1232),
    .A2(net5504),
    .Y(_02051_),
    .B1(_02050_));
 sg13g2_nor2_1 _27412_ (.A(net1751),
    .B(net5187),
    .Y(_02052_));
 sg13g2_a21oi_1 _27413_ (.A1(net5187),
    .A2(_02051_),
    .Y(_00412_),
    .B1(_02052_));
 sg13g2_and2_1 _27414_ (.A(\shift_reg[170] ),
    .B(net5455),
    .X(_02053_));
 sg13g2_a21oi_1 _27415_ (.A1(net1156),
    .A2(net5504),
    .Y(_02054_),
    .B1(_02053_));
 sg13g2_nor2_1 _27416_ (.A(net1370),
    .B(net5187),
    .Y(_02055_));
 sg13g2_a21oi_1 _27417_ (.A1(net5187),
    .A2(_02054_),
    .Y(_00413_),
    .B1(_02055_));
 sg13g2_and2_1 _27418_ (.A(\shift_reg[171] ),
    .B(net5454),
    .X(_02056_));
 sg13g2_a21oi_1 _27419_ (.A1(net1109),
    .A2(net5503),
    .Y(_02057_),
    .B1(_02056_));
 sg13g2_nor2_1 _27420_ (.A(net2008),
    .B(net5190),
    .Y(_02058_));
 sg13g2_a21oi_1 _27421_ (.A1(net5188),
    .A2(_02057_),
    .Y(_00414_),
    .B1(_02058_));
 sg13g2_and2_1 _27422_ (.A(\shift_reg[172] ),
    .B(net5454),
    .X(_02059_));
 sg13g2_a21oi_1 _27423_ (.A1(net1229),
    .A2(net5504),
    .Y(_02060_),
    .B1(_02059_));
 sg13g2_nor2_1 _27424_ (.A(net1614),
    .B(net5187),
    .Y(_02061_));
 sg13g2_a21oi_1 _27425_ (.A1(net5187),
    .A2(_02060_),
    .Y(_00415_),
    .B1(_02061_));
 sg13g2_and2_1 _27426_ (.A(\shift_reg[173] ),
    .B(net5454),
    .X(_02062_));
 sg13g2_a21oi_1 _27427_ (.A1(net1101),
    .A2(net5503),
    .Y(_02063_),
    .B1(_02062_));
 sg13g2_nor2_1 _27428_ (.A(net2323),
    .B(net5187),
    .Y(_02064_));
 sg13g2_a21oi_1 _27429_ (.A1(net5191),
    .A2(_02063_),
    .Y(_00416_),
    .B1(_02064_));
 sg13g2_and2_1 _27430_ (.A(net2058),
    .B(net5454),
    .X(_02065_));
 sg13g2_a21oi_1 _27431_ (.A1(net1255),
    .A2(net5503),
    .Y(_02066_),
    .B1(_02065_));
 sg13g2_nor2_1 _27432_ (.A(net2147),
    .B(net5181),
    .Y(_02067_));
 sg13g2_a21oi_1 _27433_ (.A1(net5181),
    .A2(_02066_),
    .Y(_00417_),
    .B1(_02067_));
 sg13g2_and2_1 _27434_ (.A(\shift_reg[175] ),
    .B(net5454),
    .X(_02068_));
 sg13g2_a21oi_1 _27435_ (.A1(net1233),
    .A2(net5504),
    .Y(_02069_),
    .B1(_02068_));
 sg13g2_nor2_1 _27436_ (.A(net1601),
    .B(net5183),
    .Y(_02070_));
 sg13g2_a21oi_1 _27437_ (.A1(net5184),
    .A2(_02069_),
    .Y(_00418_),
    .B1(_02070_));
 sg13g2_and2_1 _27438_ (.A(\shift_reg[176] ),
    .B(net5454),
    .X(_02071_));
 sg13g2_a21oi_1 _27439_ (.A1(net1135),
    .A2(net5504),
    .Y(_02072_),
    .B1(_02071_));
 sg13g2_nor2_1 _27440_ (.A(net1393),
    .B(net5184),
    .Y(_02073_));
 sg13g2_a21oi_1 _27441_ (.A1(net5184),
    .A2(_02072_),
    .Y(_00419_),
    .B1(_02073_));
 sg13g2_and2_1 _27442_ (.A(net1751),
    .B(net5451),
    .X(_02074_));
 sg13g2_a21oi_1 _27443_ (.A1(net1336),
    .A2(net5500),
    .Y(_02075_),
    .B1(_02074_));
 sg13g2_nor2_1 _27444_ (.A(net1972),
    .B(net5181),
    .Y(_02076_));
 sg13g2_a21oi_1 _27445_ (.A1(net5181),
    .A2(_02075_),
    .Y(_00420_),
    .B1(_02076_));
 sg13g2_and2_1 _27446_ (.A(net1370),
    .B(net5454),
    .X(_02077_));
 sg13g2_a21oi_1 _27447_ (.A1(net1278),
    .A2(net5501),
    .Y(_02078_),
    .B1(_02077_));
 sg13g2_nor2_1 _27448_ (.A(net1796),
    .B(net5184),
    .Y(_02079_));
 sg13g2_a21oi_1 _27449_ (.A1(net5184),
    .A2(_02078_),
    .Y(_00421_),
    .B1(_02079_));
 sg13g2_and2_1 _27450_ (.A(net2008),
    .B(net5455),
    .X(_02080_));
 sg13g2_a21oi_1 _27451_ (.A1(net1276),
    .A2(net5503),
    .Y(_02081_),
    .B1(_02080_));
 sg13g2_nor2_1 _27452_ (.A(net2190),
    .B(net5181),
    .Y(_02082_));
 sg13g2_a21oi_1 _27453_ (.A1(net5181),
    .A2(_02081_),
    .Y(_00422_),
    .B1(_02082_));
 sg13g2_and2_1 _27454_ (.A(net1614),
    .B(net5452),
    .X(_02083_));
 sg13g2_a21oi_1 _27455_ (.A1(net1342),
    .A2(net5501),
    .Y(_02084_),
    .B1(_02083_));
 sg13g2_nor2_1 _27456_ (.A(net2244),
    .B(net5183),
    .Y(_02085_));
 sg13g2_a21oi_1 _27457_ (.A1(net5183),
    .A2(_02084_),
    .Y(_00423_),
    .B1(_02085_));
 sg13g2_and2_1 _27458_ (.A(\shift_reg[181] ),
    .B(net5451),
    .X(_02086_));
 sg13g2_a21oi_1 _27459_ (.A1(net1269),
    .A2(net5501),
    .Y(_02087_),
    .B1(_02086_));
 sg13g2_nor2_1 _27460_ (.A(net1881),
    .B(net5182),
    .Y(_02088_));
 sg13g2_a21oi_1 _27461_ (.A1(net5182),
    .A2(_02087_),
    .Y(_00424_),
    .B1(_02088_));
 sg13g2_and2_1 _27462_ (.A(net2147),
    .B(net5451),
    .X(_02089_));
 sg13g2_a21oi_1 _27463_ (.A1(net1444),
    .A2(net5501),
    .Y(_02090_),
    .B1(_02089_));
 sg13g2_nor2_1 _27464_ (.A(net2309),
    .B(net5182),
    .Y(_02091_));
 sg13g2_a21oi_1 _27465_ (.A1(net5182),
    .A2(_02090_),
    .Y(_00425_),
    .B1(_02091_));
 sg13g2_and2_1 _27466_ (.A(net1601),
    .B(net5451),
    .X(_02092_));
 sg13g2_a21oi_1 _27467_ (.A1(net1496),
    .A2(net5501),
    .Y(_02093_),
    .B1(_02092_));
 sg13g2_nor2_1 _27468_ (.A(net2395),
    .B(net5183),
    .Y(_02094_));
 sg13g2_a21oi_1 _27469_ (.A1(net5183),
    .A2(_02093_),
    .Y(_00426_),
    .B1(_02094_));
 sg13g2_and2_1 _27470_ (.A(net1393),
    .B(net5452),
    .X(_02095_));
 sg13g2_a21oi_1 _27471_ (.A1(net1340),
    .A2(net5501),
    .Y(_02096_),
    .B1(_02095_));
 sg13g2_nor2_1 _27472_ (.A(net1713),
    .B(net5183),
    .Y(_02097_));
 sg13g2_a21oi_1 _27473_ (.A1(net5183),
    .A2(_02096_),
    .Y(_00427_),
    .B1(_02097_));
 sg13g2_and2_1 _27474_ (.A(\shift_reg[185] ),
    .B(net5451),
    .X(_02098_));
 sg13g2_a21oi_1 _27475_ (.A1(net1108),
    .A2(net5500),
    .Y(_02099_),
    .B1(_02098_));
 sg13g2_nor2_1 _27476_ (.A(net1862),
    .B(net5176),
    .Y(_02100_));
 sg13g2_a21oi_1 _27477_ (.A1(net5176),
    .A2(_02099_),
    .Y(_00428_),
    .B1(_02100_));
 sg13g2_and2_1 _27478_ (.A(\shift_reg[186] ),
    .B(net5452),
    .X(_02101_));
 sg13g2_a21oi_1 _27479_ (.A1(net1289),
    .A2(net5501),
    .Y(_02102_),
    .B1(_02101_));
 sg13g2_nor2_1 _27480_ (.A(net1658),
    .B(net5177),
    .Y(_02103_));
 sg13g2_a21oi_1 _27481_ (.A1(net5183),
    .A2(_02102_),
    .Y(_00429_),
    .B1(_02103_));
 sg13g2_and2_1 _27482_ (.A(\shift_reg[187] ),
    .B(net5452),
    .X(_02104_));
 sg13g2_a21oi_1 _27483_ (.A1(net1349),
    .A2(net5500),
    .Y(_02105_),
    .B1(_02104_));
 sg13g2_nor2_1 _27484_ (.A(net2107),
    .B(net5177),
    .Y(_02106_));
 sg13g2_a21oi_1 _27485_ (.A1(net5177),
    .A2(_02105_),
    .Y(_00430_),
    .B1(_02106_));
 sg13g2_and2_1 _27486_ (.A(\shift_reg[188] ),
    .B(net5450),
    .X(_02107_));
 sg13g2_a21oi_1 _27487_ (.A1(net1320),
    .A2(net5497),
    .Y(_02108_),
    .B1(_02107_));
 sg13g2_nor2_1 _27488_ (.A(net2124),
    .B(net5177),
    .Y(_02109_));
 sg13g2_a21oi_1 _27489_ (.A1(net5177),
    .A2(_02108_),
    .Y(_00431_),
    .B1(_02109_));
 sg13g2_and2_1 _27490_ (.A(net1881),
    .B(net5449),
    .X(_02110_));
 sg13g2_a21oi_1 _27491_ (.A1(net1157),
    .A2(net5498),
    .Y(_02111_),
    .B1(_02110_));
 sg13g2_nor2_1 _27492_ (.A(net2017),
    .B(net5176),
    .Y(_02112_));
 sg13g2_a21oi_1 _27493_ (.A1(net5176),
    .A2(_02111_),
    .Y(_00432_),
    .B1(_02112_));
 sg13g2_and2_1 _27494_ (.A(\shift_reg[190] ),
    .B(net5451),
    .X(_02113_));
 sg13g2_a21oi_1 _27495_ (.A1(\inv_result[182] ),
    .A2(net5500),
    .Y(_02114_),
    .B1(_02113_));
 sg13g2_nor2_1 _27496_ (.A(net1453),
    .B(net5176),
    .Y(_02115_));
 sg13g2_a21oi_1 _27497_ (.A1(net5176),
    .A2(_02114_),
    .Y(_00433_),
    .B1(_02115_));
 sg13g2_and2_1 _27498_ (.A(\shift_reg[191] ),
    .B(net5450),
    .X(_02116_));
 sg13g2_a21oi_1 _27499_ (.A1(net1348),
    .A2(net5499),
    .Y(_02117_),
    .B1(_02116_));
 sg13g2_nor2_1 _27500_ (.A(net2358),
    .B(net5178),
    .Y(_02118_));
 sg13g2_a21oi_1 _27501_ (.A1(net5177),
    .A2(_02117_),
    .Y(_00434_),
    .B1(_02118_));
 sg13g2_and2_1 _27502_ (.A(net1713),
    .B(net5450),
    .X(_02119_));
 sg13g2_a21oi_1 _27503_ (.A1(net1137),
    .A2(net5499),
    .Y(_02120_),
    .B1(_02119_));
 sg13g2_nor2_1 _27504_ (.A(net2459),
    .B(net5177),
    .Y(_02121_));
 sg13g2_a21oi_1 _27505_ (.A1(net5177),
    .A2(_02120_),
    .Y(_00435_),
    .B1(_02121_));
 sg13g2_and2_1 _27506_ (.A(\shift_reg[193] ),
    .B(net5449),
    .X(_02122_));
 sg13g2_a21oi_1 _27507_ (.A1(\inv_result[185] ),
    .A2(net5498),
    .Y(_02123_),
    .B1(_02122_));
 sg13g2_nor2_1 _27508_ (.A(net1835),
    .B(net5174),
    .Y(_02124_));
 sg13g2_a21oi_1 _27509_ (.A1(net5174),
    .A2(_02123_),
    .Y(_00436_),
    .B1(_02124_));
 sg13g2_and2_1 _27510_ (.A(net1658),
    .B(net5450),
    .X(_02125_));
 sg13g2_a21oi_1 _27511_ (.A1(net1239),
    .A2(net5499),
    .Y(_02126_),
    .B1(_02125_));
 sg13g2_nor2_1 _27512_ (.A(net1692),
    .B(net5178),
    .Y(_02127_));
 sg13g2_a21oi_1 _27513_ (.A1(net5178),
    .A2(_02126_),
    .Y(_00437_),
    .B1(_02127_));
 sg13g2_and2_1 _27514_ (.A(\shift_reg[195] ),
    .B(net5450),
    .X(_02128_));
 sg13g2_a21oi_1 _27515_ (.A1(\inv_result[187] ),
    .A2(net5498),
    .Y(_02129_),
    .B1(_02128_));
 sg13g2_nor2_1 _27516_ (.A(net1719),
    .B(net5178),
    .Y(_02130_));
 sg13g2_a21oi_1 _27517_ (.A1(net5178),
    .A2(_02129_),
    .Y(_00438_),
    .B1(_02130_));
 sg13g2_and2_1 _27518_ (.A(\shift_reg[196] ),
    .B(net5450),
    .X(_02131_));
 sg13g2_a21oi_1 _27519_ (.A1(net1328),
    .A2(net5498),
    .Y(_02132_),
    .B1(_02131_));
 sg13g2_nor2_1 _27520_ (.A(net1847),
    .B(net5170),
    .Y(_02133_));
 sg13g2_a21oi_1 _27521_ (.A1(net5170),
    .A2(_02132_),
    .Y(_00439_),
    .B1(_02133_));
 sg13g2_and2_1 _27522_ (.A(\shift_reg[197] ),
    .B(net5449),
    .X(_02134_));
 sg13g2_a21oi_1 _27523_ (.A1(net1347),
    .A2(net5498),
    .Y(_02135_),
    .B1(_02134_));
 sg13g2_nor2_1 _27524_ (.A(net1921),
    .B(net5174),
    .Y(_02136_));
 sg13g2_a21oi_1 _27525_ (.A1(net5174),
    .A2(_02135_),
    .Y(_00440_),
    .B1(_02136_));
 sg13g2_and2_1 _27526_ (.A(net1453),
    .B(net5449),
    .X(_02137_));
 sg13g2_a21oi_1 _27527_ (.A1(net1337),
    .A2(net5498),
    .Y(_02138_),
    .B1(_02137_));
 sg13g2_nor2_1 _27528_ (.A(net2452),
    .B(net5174),
    .Y(_02139_));
 sg13g2_a21oi_1 _27529_ (.A1(net5179),
    .A2(_02138_),
    .Y(_00441_),
    .B1(_02139_));
 sg13g2_and2_1 _27530_ (.A(net2358),
    .B(net5450),
    .X(_02140_));
 sg13g2_a21oi_1 _27531_ (.A1(\inv_result[191] ),
    .A2(net5499),
    .Y(_02141_),
    .B1(_02140_));
 sg13g2_nor2_1 _27532_ (.A(net2411),
    .B(net5178),
    .Y(_02142_));
 sg13g2_a21oi_1 _27533_ (.A1(net5178),
    .A2(_02141_),
    .Y(_00442_),
    .B1(_02142_));
 sg13g2_and2_1 _27534_ (.A(\shift_reg[200] ),
    .B(net5446),
    .X(_02143_));
 sg13g2_a21oi_1 _27535_ (.A1(net1363),
    .A2(net5496),
    .Y(_02144_),
    .B1(_02143_));
 sg13g2_nor2_1 _27536_ (.A(net2121),
    .B(net5173),
    .Y(_02145_));
 sg13g2_a21oi_1 _27537_ (.A1(net5173),
    .A2(_02144_),
    .Y(_00443_),
    .B1(_02145_));
 sg13g2_and2_1 _27538_ (.A(\shift_reg[201] ),
    .B(net5445),
    .X(_02146_));
 sg13g2_a21oi_1 _27539_ (.A1(net1094),
    .A2(net5495),
    .Y(_02147_),
    .B1(_02146_));
 sg13g2_nor2_1 _27540_ (.A(net1786),
    .B(net5171),
    .Y(_02148_));
 sg13g2_a21oi_1 _27541_ (.A1(net5171),
    .A2(_02147_),
    .Y(_00444_),
    .B1(_02148_));
 sg13g2_and2_1 _27542_ (.A(\shift_reg[202] ),
    .B(net5446),
    .X(_02149_));
 sg13g2_a21oi_1 _27543_ (.A1(\inv_result[194] ),
    .A2(net5496),
    .Y(_02150_),
    .B1(_02149_));
 sg13g2_nor2_1 _27544_ (.A(net1543),
    .B(net5173),
    .Y(_02151_));
 sg13g2_a21oi_1 _27545_ (.A1(net5173),
    .A2(_02150_),
    .Y(_00445_),
    .B1(_02151_));
 sg13g2_and2_1 _27546_ (.A(\shift_reg[203] ),
    .B(net5446),
    .X(_02152_));
 sg13g2_a21oi_1 _27547_ (.A1(net1286),
    .A2(net5496),
    .Y(_02153_),
    .B1(_02152_));
 sg13g2_nor2_1 _27548_ (.A(net1518),
    .B(net5173),
    .Y(_02154_));
 sg13g2_a21oi_1 _27549_ (.A1(net5186),
    .A2(_02153_),
    .Y(_00446_),
    .B1(_02154_));
 sg13g2_and2_1 _27550_ (.A(\shift_reg[204] ),
    .B(net5445),
    .X(_02155_));
 sg13g2_a21oi_1 _27551_ (.A1(net1226),
    .A2(net5495),
    .Y(_02156_),
    .B1(_02155_));
 sg13g2_nor2_1 _27552_ (.A(net1845),
    .B(net5171),
    .Y(_02157_));
 sg13g2_a21oi_1 _27553_ (.A1(net5171),
    .A2(_02156_),
    .Y(_00447_),
    .B1(_02157_));
 sg13g2_and2_1 _27554_ (.A(net1921),
    .B(net5446),
    .X(_02158_));
 sg13g2_a21oi_1 _27555_ (.A1(net1235),
    .A2(net5495),
    .Y(_02159_),
    .B1(_02158_));
 sg13g2_nor2_1 _27556_ (.A(net1942),
    .B(net5172),
    .Y(_02160_));
 sg13g2_a21oi_1 _27557_ (.A1(net5172),
    .A2(_02159_),
    .Y(_00448_),
    .B1(_02160_));
 sg13g2_and2_1 _27558_ (.A(\shift_reg[206] ),
    .B(net5445),
    .X(_02161_));
 sg13g2_a21oi_1 _27559_ (.A1(net2112),
    .A2(net5495),
    .Y(_02162_),
    .B1(_02161_));
 sg13g2_nor2_1 _27560_ (.A(net2170),
    .B(net5165),
    .Y(_02163_));
 sg13g2_a21oi_1 _27561_ (.A1(net5165),
    .A2(_02162_),
    .Y(_00449_),
    .B1(_02163_));
 sg13g2_and2_1 _27562_ (.A(\shift_reg[207] ),
    .B(net5446),
    .X(_02164_));
 sg13g2_a21oi_1 _27563_ (.A1(net1314),
    .A2(net5496),
    .Y(_02165_),
    .B1(_02164_));
 sg13g2_nor2_1 _27564_ (.A(net1425),
    .B(net5168),
    .Y(_02166_));
 sg13g2_a21oi_1 _27565_ (.A1(net5168),
    .A2(_02165_),
    .Y(_00450_),
    .B1(_02166_));
 sg13g2_and2_1 _27566_ (.A(net2121),
    .B(net5447),
    .X(_02167_));
 sg13g2_a21oi_1 _27567_ (.A1(net2172),
    .A2(net5496),
    .Y(_02168_),
    .B1(_02167_));
 sg13g2_nor2_1 _27568_ (.A(net2336),
    .B(net5168),
    .Y(_02169_));
 sg13g2_a21oi_1 _27569_ (.A1(net5168),
    .A2(_02168_),
    .Y(_00451_),
    .B1(_02169_));
 sg13g2_and2_1 _27570_ (.A(\shift_reg[209] ),
    .B(net5445),
    .X(_02170_));
 sg13g2_a21oi_1 _27571_ (.A1(\inv_result[201] ),
    .A2(net5495),
    .Y(_02171_),
    .B1(_02170_));
 sg13g2_nor2_1 _27572_ (.A(net1668),
    .B(net5165),
    .Y(_02172_));
 sg13g2_a21oi_1 _27573_ (.A1(net5165),
    .A2(_02171_),
    .Y(_00452_),
    .B1(_02172_));
 sg13g2_and2_1 _27574_ (.A(net1543),
    .B(net5446),
    .X(_02173_));
 sg13g2_a21oi_1 _27575_ (.A1(net1180),
    .A2(net5496),
    .Y(_02174_),
    .B1(_02173_));
 sg13g2_nor2_1 _27576_ (.A(net1997),
    .B(net5167),
    .Y(_02175_));
 sg13g2_a21oi_1 _27577_ (.A1(net5167),
    .A2(_02174_),
    .Y(_00453_),
    .B1(_02175_));
 sg13g2_and2_1 _27578_ (.A(net1518),
    .B(net5447),
    .X(_02176_));
 sg13g2_a21oi_1 _27579_ (.A1(\inv_result[203] ),
    .A2(net5502),
    .Y(_02177_),
    .B1(_02176_));
 sg13g2_nor2_1 _27580_ (.A(net2101),
    .B(net5168),
    .Y(_02178_));
 sg13g2_a21oi_1 _27581_ (.A1(net5168),
    .A2(_02177_),
    .Y(_00454_),
    .B1(_02178_));
 sg13g2_and2_1 _27582_ (.A(net1845),
    .B(net5445),
    .X(_02179_));
 sg13g2_a21oi_1 _27583_ (.A1(net1129),
    .A2(net5495),
    .Y(_02180_),
    .B1(_02179_));
 sg13g2_nor2_1 _27584_ (.A(net2203),
    .B(net5168),
    .Y(_02181_));
 sg13g2_a21oi_1 _27585_ (.A1(net5168),
    .A2(_02180_),
    .Y(_00455_),
    .B1(_02181_));
 sg13g2_and2_1 _27586_ (.A(\shift_reg[213] ),
    .B(net5445),
    .X(_02182_));
 sg13g2_a21oi_1 _27587_ (.A1(\inv_result[205] ),
    .A2(net5495),
    .Y(_02183_),
    .B1(_02182_));
 sg13g2_nor2_1 _27588_ (.A(net1451),
    .B(net5167),
    .Y(_02184_));
 sg13g2_a21oi_1 _27589_ (.A1(net5165),
    .A2(_02183_),
    .Y(_00456_),
    .B1(_02184_));
 sg13g2_and2_1 _27590_ (.A(\shift_reg[214] ),
    .B(net5444),
    .X(_02185_));
 sg13g2_a21oi_1 _27591_ (.A1(net1234),
    .A2(net5494),
    .Y(_02186_),
    .B1(_02185_));
 sg13g2_nor2_1 _27592_ (.A(net1434),
    .B(net5167),
    .Y(_02187_));
 sg13g2_a21oi_1 _27593_ (.A1(net5167),
    .A2(_02186_),
    .Y(_00457_),
    .B1(_02187_));
 sg13g2_and2_1 _27594_ (.A(net1425),
    .B(net5444),
    .X(_02188_));
 sg13g2_a21oi_1 _27595_ (.A1(net1136),
    .A2(net5494),
    .Y(_02189_),
    .B1(_02188_));
 sg13g2_nor2_1 _27596_ (.A(net1788),
    .B(net5167),
    .Y(_02190_));
 sg13g2_a21oi_1 _27597_ (.A1(net5167),
    .A2(_02189_),
    .Y(_00458_),
    .B1(_02190_));
 sg13g2_and2_1 _27598_ (.A(\shift_reg[216] ),
    .B(net5440),
    .X(_02191_));
 sg13g2_a21oi_1 _27599_ (.A1(net1200),
    .A2(net5489),
    .Y(_02192_),
    .B1(_02191_));
 sg13g2_nor2_1 _27600_ (.A(net2056),
    .B(net5161),
    .Y(_02193_));
 sg13g2_a21oi_1 _27601_ (.A1(net5161),
    .A2(_02192_),
    .Y(_00459_),
    .B1(_02193_));
 sg13g2_and2_1 _27602_ (.A(net1668),
    .B(net5443),
    .X(_02194_));
 sg13g2_a21oi_1 _27603_ (.A1(net1545),
    .A2(net5490),
    .Y(_02195_),
    .B1(_02194_));
 sg13g2_nor2_1 _27604_ (.A(net1973),
    .B(net5159),
    .Y(_02196_));
 sg13g2_a21oi_1 _27605_ (.A1(net5159),
    .A2(_02195_),
    .Y(_00460_),
    .B1(_02196_));
 sg13g2_and2_1 _27606_ (.A(\shift_reg[218] ),
    .B(net5444),
    .X(_02197_));
 sg13g2_a21oi_1 _27607_ (.A1(net1302),
    .A2(net5489),
    .Y(_02198_),
    .B1(_02197_));
 sg13g2_nor2_1 _27608_ (.A(net1431),
    .B(net5161),
    .Y(_02199_));
 sg13g2_a21oi_1 _27609_ (.A1(net5161),
    .A2(_02198_),
    .Y(_00461_),
    .B1(_02199_));
 sg13g2_and2_1 _27610_ (.A(net2101),
    .B(net5447),
    .X(_02200_));
 sg13g2_a21oi_1 _27611_ (.A1(net1103),
    .A2(net5491),
    .Y(_02201_),
    .B1(_02200_));
 sg13g2_nor2_1 _27612_ (.A(net2106),
    .B(net5167),
    .Y(_02202_));
 sg13g2_a21oi_1 _27613_ (.A1(net5161),
    .A2(_02201_),
    .Y(_00462_),
    .B1(_02202_));
 sg13g2_and2_1 _27614_ (.A(\shift_reg[220] ),
    .B(net5444),
    .X(_02203_));
 sg13g2_a21oi_1 _27615_ (.A1(net1275),
    .A2(net5491),
    .Y(_02204_),
    .B1(_02203_));
 sg13g2_nor2_1 _27616_ (.A(net1808),
    .B(net5162),
    .Y(_02205_));
 sg13g2_a21oi_1 _27617_ (.A1(net5161),
    .A2(_02204_),
    .Y(_00463_),
    .B1(_02205_));
 sg13g2_and2_1 _27618_ (.A(\shift_reg[221] ),
    .B(net5447),
    .X(_02206_));
 sg13g2_a21oi_1 _27619_ (.A1(net1104),
    .A2(net5490),
    .Y(_02207_),
    .B1(_02206_));
 sg13g2_nor2_1 _27620_ (.A(net1429),
    .B(net5160),
    .Y(_02208_));
 sg13g2_a21oi_1 _27621_ (.A1(net5159),
    .A2(_02207_),
    .Y(_00464_),
    .B1(_02208_));
 sg13g2_and2_1 _27622_ (.A(net1434),
    .B(net5444),
    .X(_02209_));
 sg13g2_a21oi_1 _27623_ (.A1(net1285),
    .A2(net5490),
    .Y(_02210_),
    .B1(_02209_));
 sg13g2_nor2_1 _27624_ (.A(net2047),
    .B(net5160),
    .Y(_02211_));
 sg13g2_a21oi_1 _27625_ (.A1(net5160),
    .A2(_02210_),
    .Y(_00465_),
    .B1(_02211_));
 sg13g2_and2_1 _27626_ (.A(net1788),
    .B(net5440),
    .X(_02212_));
 sg13g2_a21oi_1 _27627_ (.A1(net1123),
    .A2(net5489),
    .Y(_02213_),
    .B1(_02212_));
 sg13g2_nor2_1 _27628_ (.A(net2041),
    .B(net5160),
    .Y(_02214_));
 sg13g2_a21oi_1 _27629_ (.A1(net5160),
    .A2(_02213_),
    .Y(_00466_),
    .B1(_02214_));
 sg13g2_and2_1 _27630_ (.A(net2056),
    .B(net5441),
    .X(_02215_));
 sg13g2_a21oi_1 _27631_ (.A1(net1248),
    .A2(net5489),
    .Y(_02216_),
    .B1(_02215_));
 sg13g2_nor2_1 _27632_ (.A(net2241),
    .B(net5160),
    .Y(_02217_));
 sg13g2_a21oi_1 _27633_ (.A1(net5160),
    .A2(_02216_),
    .Y(_00467_),
    .B1(_02217_));
 sg13g2_and2_1 _27634_ (.A(\shift_reg[225] ),
    .B(net5441),
    .X(_02218_));
 sg13g2_a21oi_1 _27635_ (.A1(net1127),
    .A2(net5490),
    .Y(_02219_),
    .B1(_02218_));
 sg13g2_nor2_1 _27636_ (.A(net1948),
    .B(net5159),
    .Y(_02220_));
 sg13g2_a21oi_1 _27637_ (.A1(net5159),
    .A2(_02219_),
    .Y(_00468_),
    .B1(_02220_));
 sg13g2_and2_1 _27638_ (.A(net1431),
    .B(net5440),
    .X(_02221_));
 sg13g2_a21oi_1 _27639_ (.A1(net1284),
    .A2(net5489),
    .Y(_02222_),
    .B1(_02221_));
 sg13g2_nor2_1 _27640_ (.A(net2403),
    .B(net5160),
    .Y(_02223_));
 sg13g2_a21oi_1 _27641_ (.A1(net5161),
    .A2(_02222_),
    .Y(_00469_),
    .B1(_02223_));
 sg13g2_and2_1 _27642_ (.A(net2106),
    .B(net5440),
    .X(_02224_));
 sg13g2_a21oi_1 _27643_ (.A1(\inv_result[219] ),
    .A2(net5489),
    .Y(_02225_),
    .B1(_02224_));
 sg13g2_nor2_1 _27644_ (.A(net2643),
    .B(net5156),
    .Y(_02226_));
 sg13g2_a21oi_1 _27645_ (.A1(net5156),
    .A2(_02225_),
    .Y(_00470_),
    .B1(_02226_));
 sg13g2_and2_1 _27646_ (.A(net1808),
    .B(net5440),
    .X(_02227_));
 sg13g2_a21oi_1 _27647_ (.A1(net1283),
    .A2(net5489),
    .Y(_02228_),
    .B1(_02227_));
 sg13g2_nor2_1 _27648_ (.A(net2000),
    .B(net5156),
    .Y(_02229_));
 sg13g2_a21oi_1 _27649_ (.A1(net5156),
    .A2(_02228_),
    .Y(_00471_),
    .B1(_02229_));
 sg13g2_and2_1 _27650_ (.A(net1429),
    .B(net5440),
    .X(_02230_));
 sg13g2_a21oi_1 _27651_ (.A1(net1209),
    .A2(net5490),
    .Y(_02231_),
    .B1(_02230_));
 sg13g2_nor2_1 _27652_ (.A(net1487),
    .B(net5157),
    .Y(_02232_));
 sg13g2_a21oi_1 _27653_ (.A1(net5157),
    .A2(_02231_),
    .Y(_00472_),
    .B1(_02232_));
 sg13g2_and2_1 _27654_ (.A(\shift_reg[230] ),
    .B(net5440),
    .X(_02233_));
 sg13g2_a21oi_1 _27655_ (.A1(net1351),
    .A2(net5487),
    .Y(_02234_),
    .B1(_02233_));
 sg13g2_nor2_1 _27656_ (.A(net1980),
    .B(net5155),
    .Y(_02235_));
 sg13g2_a21oi_1 _27657_ (.A1(net5155),
    .A2(_02234_),
    .Y(_00473_),
    .B1(_02235_));
 sg13g2_and2_1 _27658_ (.A(\shift_reg[231] ),
    .B(net5440),
    .X(_02236_));
 sg13g2_a21oi_1 _27659_ (.A1(net1357),
    .A2(net5489),
    .Y(_02237_),
    .B1(_02236_));
 sg13g2_nor2_1 _27660_ (.A(net1427),
    .B(net5156),
    .Y(_02238_));
 sg13g2_a21oi_1 _27661_ (.A1(net5156),
    .A2(_02237_),
    .Y(_00474_),
    .B1(_02238_));
 sg13g2_and2_1 _27662_ (.A(\shift_reg[232] ),
    .B(net5439),
    .X(_02239_));
 sg13g2_a21oi_1 _27663_ (.A1(net1100),
    .A2(net5488),
    .Y(_02240_),
    .B1(_02239_));
 sg13g2_nor2_1 _27664_ (.A(net1828),
    .B(net5156),
    .Y(_02241_));
 sg13g2_a21oi_1 _27665_ (.A1(net5156),
    .A2(_02240_),
    .Y(_00475_),
    .B1(_02241_));
 sg13g2_and2_1 _27666_ (.A(net1948),
    .B(net5438),
    .X(_02242_));
 sg13g2_a21oi_1 _27667_ (.A1(net1134),
    .A2(net5487),
    .Y(_02243_),
    .B1(_02242_));
 sg13g2_nor2_1 _27668_ (.A(net2193),
    .B(net5155),
    .Y(_02244_));
 sg13g2_a21oi_1 _27669_ (.A1(net5155),
    .A2(_02243_),
    .Y(_00476_),
    .B1(_02244_));
 sg13g2_and2_1 _27670_ (.A(\shift_reg[234] ),
    .B(net5437),
    .X(_02245_));
 sg13g2_a21oi_1 _27671_ (.A1(net1122),
    .A2(net5486),
    .Y(_02246_),
    .B1(_02245_));
 sg13g2_nor2_1 _27672_ (.A(net1502),
    .B(net5152),
    .Y(_02247_));
 sg13g2_a21oi_1 _27673_ (.A1(net5152),
    .A2(_02246_),
    .Y(_00477_),
    .B1(_02247_));
 sg13g2_and2_1 _27674_ (.A(\shift_reg[235] ),
    .B(net5439),
    .X(_02248_));
 sg13g2_a21oi_1 _27675_ (.A1(net1106),
    .A2(net5488),
    .Y(_02249_),
    .B1(_02248_));
 sg13g2_nor2_1 _27676_ (.A(net1345),
    .B(net5157),
    .Y(_02250_));
 sg13g2_a21oi_1 _27677_ (.A1(net5157),
    .A2(_02249_),
    .Y(_00478_),
    .B1(_02250_));
 sg13g2_and2_1 _27678_ (.A(\shift_reg[236] ),
    .B(net5439),
    .X(_02251_));
 sg13g2_a21oi_1 _27679_ (.A1(net1293),
    .A2(net5486),
    .Y(_02252_),
    .B1(_02251_));
 sg13g2_nor2_1 _27680_ (.A(net1404),
    .B(net5152),
    .Y(_02253_));
 sg13g2_a21oi_1 _27681_ (.A1(net5152),
    .A2(_02252_),
    .Y(_00479_),
    .B1(_02253_));
 sg13g2_and2_1 _27682_ (.A(net1487),
    .B(net5439),
    .X(_02254_));
 sg13g2_a21oi_1 _27683_ (.A1(net1099),
    .A2(net5488),
    .Y(_02255_),
    .B1(_02254_));
 sg13g2_nor2_1 _27684_ (.A(net2567),
    .B(net5157),
    .Y(_02256_));
 sg13g2_a21oi_1 _27685_ (.A1(net5157),
    .A2(_02255_),
    .Y(_00480_),
    .B1(_02256_));
 sg13g2_and2_1 _27686_ (.A(net1980),
    .B(net5438),
    .X(_02257_));
 sg13g2_a21oi_1 _27687_ (.A1(net1321),
    .A2(net5486),
    .Y(_02258_),
    .B1(_02257_));
 sg13g2_nor2_1 _27688_ (.A(net2149),
    .B(net5149),
    .Y(_02259_));
 sg13g2_a21oi_1 _27689_ (.A1(net5149),
    .A2(_02258_),
    .Y(_00481_),
    .B1(_02259_));
 sg13g2_and2_1 _27690_ (.A(net1427),
    .B(net5439),
    .X(_02260_));
 sg13g2_a21oi_1 _27691_ (.A1(net1334),
    .A2(net5488),
    .Y(_02261_),
    .B1(_02260_));
 sg13g2_nor2_1 _27692_ (.A(net1611),
    .B(net5150),
    .Y(_02262_));
 sg13g2_a21oi_1 _27693_ (.A1(net5150),
    .A2(_02261_),
    .Y(_00482_),
    .B1(_02262_));
 sg13g2_and2_1 _27694_ (.A(net1828),
    .B(net5437),
    .X(_02263_));
 sg13g2_a21oi_1 _27695_ (.A1(net1318),
    .A2(net5483),
    .Y(_02264_),
    .B1(_02263_));
 sg13g2_nor2_1 _27696_ (.A(net2542),
    .B(net5147),
    .Y(_02265_));
 sg13g2_a21oi_1 _27697_ (.A1(net5147),
    .A2(_02264_),
    .Y(_00483_),
    .B1(_02265_));
 sg13g2_and2_1 _27698_ (.A(\shift_reg[241] ),
    .B(net5437),
    .X(_02266_));
 sg13g2_a21oi_1 _27699_ (.A1(net1251),
    .A2(net5480),
    .Y(_02267_),
    .B1(_02266_));
 sg13g2_nor2_1 _27700_ (.A(net1976),
    .B(net5136),
    .Y(_02268_));
 sg13g2_a21oi_1 _27701_ (.A1(net5136),
    .A2(_02267_),
    .Y(_00484_),
    .B1(_02268_));
 sg13g2_and2_1 _27702_ (.A(net1502),
    .B(net5437),
    .X(_02269_));
 sg13g2_a21oi_1 _27703_ (.A1(net1208),
    .A2(net5483),
    .Y(_02270_),
    .B1(_02269_));
 sg13g2_nor2_1 _27704_ (.A(net2174),
    .B(net5148),
    .Y(_02271_));
 sg13g2_a21oi_1 _27705_ (.A1(net5148),
    .A2(_02270_),
    .Y(_00485_),
    .B1(_02271_));
 sg13g2_and2_1 _27706_ (.A(net1345),
    .B(net5439),
    .X(_02272_));
 sg13g2_a21oi_1 _27707_ (.A1(net2521),
    .A2(net5483),
    .Y(_02273_),
    .B1(_02272_));
 sg13g2_nor2_1 _27708_ (.A(net2795),
    .B(net5148),
    .Y(_02274_));
 sg13g2_a21oi_1 _27709_ (.A1(net5148),
    .A2(_02273_),
    .Y(_00486_),
    .B1(_02274_));
 sg13g2_and2_1 _27710_ (.A(net1404),
    .B(net5437),
    .X(_02275_));
 sg13g2_a21oi_1 _27711_ (.A1(net2592),
    .A2(net5486),
    .Y(_02276_),
    .B1(_02275_));
 sg13g2_nor2_1 _27712_ (.A(net2868),
    .B(net5158),
    .Y(_02277_));
 sg13g2_a21oi_1 _27713_ (.A1(net5152),
    .A2(_02276_),
    .Y(_00487_),
    .B1(_02277_));
 sg13g2_and2_1 _27714_ (.A(\shift_reg[245] ),
    .B(net5435),
    .X(_02278_));
 sg13g2_a21oi_1 _27715_ (.A1(\inv_result[237] ),
    .A2(net5479),
    .Y(_02279_),
    .B1(_02278_));
 sg13g2_nor2_1 _27716_ (.A(net2303),
    .B(net5144),
    .Y(_02280_));
 sg13g2_a21oi_1 _27717_ (.A1(net5144),
    .A2(_02279_),
    .Y(_00488_),
    .B1(_02280_));
 sg13g2_and2_1 _27718_ (.A(\shift_reg[246] ),
    .B(net5435),
    .X(_02281_));
 sg13g2_a21oi_1 _27719_ (.A1(net1098),
    .A2(net5479),
    .Y(_02282_),
    .B1(_02281_));
 sg13g2_nor2_1 _27720_ (.A(net1402),
    .B(net5136),
    .Y(_02283_));
 sg13g2_a21oi_1 _27721_ (.A1(net5137),
    .A2(_02282_),
    .Y(_00489_),
    .B1(_02283_));
 sg13g2_and2_1 _27722_ (.A(net1611),
    .B(net5435),
    .X(_02284_));
 sg13g2_a21oi_1 _27723_ (.A1(net1281),
    .A2(net5479),
    .Y(_02285_),
    .B1(_02284_));
 sg13g2_nor2_1 _27724_ (.A(net2660),
    .B(net5136),
    .Y(_02286_));
 sg13g2_a21oi_1 _27725_ (.A1(net5137),
    .A2(_02285_),
    .Y(_00490_),
    .B1(_02286_));
 sg13g2_and2_1 _27726_ (.A(\shift_reg[248] ),
    .B(net5433),
    .X(_02287_));
 sg13g2_a21oi_1 _27727_ (.A1(\inv_result[240] ),
    .A2(net5477),
    .Y(_02288_),
    .B1(_02287_));
 sg13g2_nor2_1 _27728_ (.A(net1141),
    .B(net5134),
    .Y(_02289_));
 sg13g2_a21oi_1 _27729_ (.A1(net5134),
    .A2(_02288_),
    .Y(_00491_),
    .B1(_02289_));
 sg13g2_and2_1 _27730_ (.A(\shift_reg[249] ),
    .B(net5433),
    .X(_02290_));
 sg13g2_a21oi_1 _27731_ (.A1(\inv_result[241] ),
    .A2(net5478),
    .Y(_02291_),
    .B1(_02290_));
 sg13g2_nor2_1 _27732_ (.A(net1242),
    .B(net5134),
    .Y(_02292_));
 sg13g2_a21oi_1 _27733_ (.A1(net5134),
    .A2(_02291_),
    .Y(_00492_),
    .B1(_02292_));
 sg13g2_and2_1 _27734_ (.A(\shift_reg[250] ),
    .B(net5435),
    .X(_02293_));
 sg13g2_a21oi_1 _27735_ (.A1(\inv_result[242] ),
    .A2(net5479),
    .Y(_02294_),
    .B1(_02293_));
 sg13g2_nor2_1 _27736_ (.A(net1230),
    .B(net5135),
    .Y(_02295_));
 sg13g2_a21oi_1 _27737_ (.A1(net5135),
    .A2(_02294_),
    .Y(_00493_),
    .B1(_02295_));
 sg13g2_and2_1 _27738_ (.A(\shift_reg[251] ),
    .B(net5432),
    .X(_02296_));
 sg13g2_a21oi_1 _27739_ (.A1(\inv_result[243] ),
    .A2(net5477),
    .Y(_02297_),
    .B1(_02296_));
 sg13g2_nor2_1 _27740_ (.A(net1192),
    .B(net5135),
    .Y(_02298_));
 sg13g2_a21oi_1 _27741_ (.A1(net5135),
    .A2(_02297_),
    .Y(_00494_),
    .B1(_02298_));
 sg13g2_and2_1 _27742_ (.A(\shift_reg[252] ),
    .B(net5433),
    .X(_02299_));
 sg13g2_a21oi_1 _27743_ (.A1(net1174),
    .A2(net5479),
    .Y(_02300_),
    .B1(_02299_));
 sg13g2_nor2_1 _27744_ (.A(net1194),
    .B(net5136),
    .Y(_02301_));
 sg13g2_a21oi_1 _27745_ (.A1(net5136),
    .A2(_02300_),
    .Y(_00495_),
    .B1(_02301_));
 sg13g2_and2_1 _27746_ (.A(\shift_reg[253] ),
    .B(net5433),
    .X(_02302_));
 sg13g2_a21oi_1 _27747_ (.A1(net1120),
    .A2(net5479),
    .Y(_02303_),
    .B1(_02302_));
 sg13g2_nor2_1 _27748_ (.A(net1204),
    .B(net5136),
    .Y(_02304_));
 sg13g2_a21oi_1 _27749_ (.A1(net5136),
    .A2(_02303_),
    .Y(_00496_),
    .B1(_02304_));
 sg13g2_and2_1 _27750_ (.A(\shift_reg[254] ),
    .B(net5433),
    .X(_02305_));
 sg13g2_a21oi_1 _27751_ (.A1(net1082),
    .A2(net5477),
    .Y(_02306_),
    .B1(_02305_));
 sg13g2_nor2_1 _27752_ (.A(net1323),
    .B(net5134),
    .Y(_02307_));
 sg13g2_a21oi_1 _27753_ (.A1(net5134),
    .A2(_02306_),
    .Y(_00497_),
    .B1(_02307_));
 sg13g2_and2_1 _27754_ (.A(\shift_reg[255] ),
    .B(net5432),
    .X(_02308_));
 sg13g2_a21oi_1 _27755_ (.A1(\inv_result[247] ),
    .A2(net5477),
    .Y(_02309_),
    .B1(_02308_));
 sg13g2_nor2_1 _27756_ (.A(net1150),
    .B(net5134),
    .Y(_02310_));
 sg13g2_a21oi_1 _27757_ (.A1(net5134),
    .A2(_02309_),
    .Y(_00498_),
    .B1(_02310_));
 sg13g2_and2_1 _27758_ (.A(\shift_reg[256] ),
    .B(net5432),
    .X(_02311_));
 sg13g2_a21oi_1 _27759_ (.A1(\inv_result[248] ),
    .A2(net5478),
    .Y(_02312_),
    .B1(_02311_));
 sg13g2_nor2_1 _27760_ (.A(net1113),
    .B(net5140),
    .Y(_02313_));
 sg13g2_a21oi_1 _27761_ (.A1(net5138),
    .A2(_02312_),
    .Y(_00499_),
    .B1(_02313_));
 sg13g2_and2_1 _27762_ (.A(\shift_reg[257] ),
    .B(net5432),
    .X(_02314_));
 sg13g2_a21oi_1 _27763_ (.A1(net1211),
    .A2(net5477),
    .Y(_02315_),
    .B1(_02314_));
 sg13g2_nor2_1 _27764_ (.A(net1240),
    .B(net5139),
    .Y(_02316_));
 sg13g2_a21oi_1 _27765_ (.A1(net5139),
    .A2(_02315_),
    .Y(_00500_),
    .B1(_02316_));
 sg13g2_and2_1 _27766_ (.A(\shift_reg[258] ),
    .B(net5432),
    .X(_02317_));
 sg13g2_a21oi_1 _27767_ (.A1(net1089),
    .A2(net5478),
    .Y(_02318_),
    .B1(_02317_));
 sg13g2_nor2_1 _27768_ (.A(net1130),
    .B(net5141),
    .Y(_02319_));
 sg13g2_a21oi_1 _27769_ (.A1(net5140),
    .A2(_02318_),
    .Y(_00501_),
    .B1(_02319_));
 sg13g2_and2_1 _27770_ (.A(\shift_reg[259] ),
    .B(net5432),
    .X(_02320_));
 sg13g2_a21oi_1 _27771_ (.A1(net1119),
    .A2(net5477),
    .Y(_02321_),
    .B1(_02320_));
 sg13g2_nor2_1 _27772_ (.A(net1163),
    .B(net5139),
    .Y(_02322_));
 sg13g2_a21oi_1 _27773_ (.A1(net5138),
    .A2(_02321_),
    .Y(_00502_),
    .B1(_02322_));
 sg13g2_and2_1 _27774_ (.A(net1194),
    .B(net5433),
    .X(_02323_));
 sg13g2_a21oi_2 _27775_ (.B1(_02323_),
    .Y(_02324_),
    .A2(net5479),
    .A1(net1170));
 sg13g2_nor2_1 _27776_ (.A(net1210),
    .B(net5141),
    .Y(_02325_));
 sg13g2_a21oi_1 _27777_ (.A1(net5141),
    .A2(_02324_),
    .Y(_00503_),
    .B1(_02325_));
 sg13g2_and2_1 _27778_ (.A(net1204),
    .B(net5433),
    .X(_02326_));
 sg13g2_a21oi_2 _27779_ (.B1(_02326_),
    .Y(_02327_),
    .A2(net5479),
    .A1(\inv_result[253] ));
 sg13g2_nor2_1 _27780_ (.A(net1217),
    .B(net5140),
    .Y(_02328_));
 sg13g2_a21oi_1 _27781_ (.A1(net5140),
    .A2(_02327_),
    .Y(_00504_),
    .B1(_02328_));
 sg13g2_and2_1 _27782_ (.A(\shift_reg[262] ),
    .B(net5432),
    .X(_02329_));
 sg13g2_a21oi_1 _27783_ (.A1(\inv_result[254] ),
    .A2(net5477),
    .Y(_02330_),
    .B1(_02329_));
 sg13g2_nor2_1 _27784_ (.A(net1115),
    .B(net5138),
    .Y(_02331_));
 sg13g2_a21oi_1 _27785_ (.A1(net5138),
    .A2(_02330_),
    .Y(_00505_),
    .B1(_02331_));
 sg13g2_and2_1 _27786_ (.A(\shift_reg[263] ),
    .B(net5432),
    .X(_02332_));
 sg13g2_a21oi_1 _27787_ (.A1(\inv_result[255] ),
    .A2(net5477),
    .Y(_02333_),
    .B1(_02332_));
 sg13g2_nor2_1 _27788_ (.A(net1117),
    .B(net5138),
    .Y(_02334_));
 sg13g2_a21oi_1 _27789_ (.A1(net5138),
    .A2(_02333_),
    .Y(_00506_),
    .B1(_02334_));
 sg13g2_nor3_1 _27790_ (.A(_14811_),
    .B(_14814_),
    .C(_14816_),
    .Y(_02335_));
 sg13g2_nor2_1 _27791_ (.A(net2393),
    .B(_02335_),
    .Y(_02336_));
 sg13g2_nor2_1 _27792_ (.A(net5482),
    .B(net2394),
    .Y(_00507_));
 sg13g2_nand2_1 _27793_ (.Y(_02337_),
    .A(net2316),
    .B(net4143));
 sg13g2_o21ai_1 _27794_ (.B1(_02337_),
    .Y(_00508_),
    .A1(_18908_),
    .A2(net5532));
 sg13g2_nor2_1 _27795_ (.A(net5829),
    .B(net4389),
    .Y(_02338_));
 sg13g2_xnor2_1 _27796_ (.Y(_02339_),
    .A(net3389),
    .B(_02338_));
 sg13g2_nand2_1 _27797_ (.Y(_02340_),
    .A(net5632),
    .B(_02339_));
 sg13g2_o21ai_1 _27798_ (.B1(_02340_),
    .Y(_00509_),
    .A1(_14249_),
    .A2(_19028_));
 sg13g2_nand3_1 _27799_ (.B(net5627),
    .C(_19025_),
    .A(net5881),
    .Y(_02341_));
 sg13g2_nand3_1 _27800_ (.B(net3439),
    .C(net5881),
    .A(net5829),
    .Y(_02342_));
 sg13g2_nand3_1 _27801_ (.B(net5881),
    .C(_19007_),
    .A(net3439),
    .Y(_02343_));
 sg13g2_o21ai_1 _27802_ (.B1(_02342_),
    .Y(_02344_),
    .A1(net4450),
    .A2(_02343_));
 sg13g2_a21o_1 _27803_ (.A2(net3389),
    .A1(\u_inv.counter[0] ),
    .B1(net5881),
    .X(_02345_));
 sg13g2_nor4_1 _27804_ (.A(_14249_),
    .B(net5881),
    .C(net4450),
    .D(_19008_),
    .Y(_02346_));
 sg13g2_o21ai_1 _27805_ (.B1(net5632),
    .Y(_02347_),
    .A1(_02345_),
    .A2(_02346_));
 sg13g2_o21ai_1 _27806_ (.B1(_02341_),
    .Y(_00510_),
    .A1(_02344_),
    .A2(_02347_));
 sg13g2_and2_1 _27807_ (.A(net3371),
    .B(_02344_),
    .X(_02348_));
 sg13g2_nor2_1 _27808_ (.A(net5627),
    .B(_02348_),
    .Y(_02349_));
 sg13g2_o21ai_1 _27809_ (.B1(_02349_),
    .Y(_02350_),
    .A1(net3371),
    .A2(_02344_));
 sg13g2_o21ai_1 _27810_ (.B1(_02350_),
    .Y(_00511_),
    .A1(_14250_),
    .A2(_19028_));
 sg13g2_a21oi_1 _27811_ (.A1(net5632),
    .A2(_02348_),
    .Y(_02351_),
    .B1(net2844));
 sg13g2_nand3_1 _27812_ (.B(net5632),
    .C(_02348_),
    .A(net2844),
    .Y(_02352_));
 sg13g2_inv_1 _27813_ (.Y(_02353_),
    .A(_02352_));
 sg13g2_nand4_1 _27814_ (.B(\u_inv.counter[2] ),
    .C(\u_inv.counter[3] ),
    .A(\u_inv.counter[1] ),
    .Y(_02354_),
    .D(\u_inv.counter[4] ));
 sg13g2_nor3_1 _27815_ (.A(_20877_[0]),
    .B(net2845),
    .C(_02353_),
    .Y(_00512_));
 sg13g2_a21oi_1 _27816_ (.A1(_19025_),
    .A2(_02352_),
    .Y(_02355_),
    .B1(_14253_));
 sg13g2_nand3_1 _27817_ (.B(net3072),
    .C(\u_inv.counter[4] ),
    .A(net3440),
    .Y(_02356_));
 sg13g2_a21o_1 _27818_ (.A2(_02343_),
    .A1(_02342_),
    .B1(_02356_),
    .X(_02357_));
 sg13g2_a21oi_1 _27819_ (.A1(_14253_),
    .A2(_02352_),
    .Y(_00513_),
    .B1(_02355_));
 sg13g2_nor2_2 _27820_ (.A(_14822_),
    .B(_02354_),
    .Y(_02358_));
 sg13g2_nand2_1 _27821_ (.Y(_02359_),
    .A(net5829),
    .B(_02358_));
 sg13g2_o21ai_1 _27822_ (.B1(_14252_),
    .Y(_02360_),
    .A1(_02342_),
    .A2(_02356_));
 sg13g2_xnor2_1 _27823_ (.Y(_02361_),
    .A(_14252_),
    .B(_02357_));
 sg13g2_nand3_1 _27824_ (.B(_02359_),
    .C(_02360_),
    .A(net4450),
    .Y(_02362_));
 sg13g2_o21ai_1 _27825_ (.B1(_02362_),
    .Y(_02363_),
    .A1(net4450),
    .A2(_02361_));
 sg13g2_nand2_1 _27826_ (.Y(_02364_),
    .A(net5632),
    .B(_02363_));
 sg13g2_o21ai_1 _27827_ (.B1(_02364_),
    .Y(_00514_),
    .A1(_14252_),
    .A2(_19028_));
 sg13g2_nor2_1 _27828_ (.A(_14251_),
    .B(_19028_),
    .Y(_02365_));
 sg13g2_a21oi_1 _27829_ (.A1(net5829),
    .A2(_02358_),
    .Y(_02366_),
    .B1(net3431));
 sg13g2_nand3_1 _27830_ (.B(net3431),
    .C(_02358_),
    .A(net5829),
    .Y(_02367_));
 sg13g2_nand2b_1 _27831_ (.Y(_02368_),
    .B(_02367_),
    .A_N(_02366_));
 sg13g2_xnor2_1 _27832_ (.Y(_02369_),
    .A(\u_inv.counter[7] ),
    .B(_02358_));
 sg13g2_mux2_1 _27833_ (.A0(_02368_),
    .A1(_02369_),
    .S(_19007_),
    .X(_02370_));
 sg13g2_nand2b_1 _27834_ (.Y(_02371_),
    .B(_02370_),
    .A_N(net4450));
 sg13g2_a21oi_1 _27835_ (.A1(net4450),
    .A2(_02368_),
    .Y(_02372_),
    .B1(net5627));
 sg13g2_a21o_1 _27836_ (.A2(_02372_),
    .A1(_02371_),
    .B1(_02365_),
    .X(_00515_));
 sg13g2_nor2_1 _27837_ (.A(_14254_),
    .B(_20877_[0]),
    .Y(_02373_));
 sg13g2_nor3_1 _27838_ (.A(_14251_),
    .B(_14252_),
    .C(_02357_),
    .Y(_02374_));
 sg13g2_o21ai_1 _27839_ (.B1(net5632),
    .Y(_02375_),
    .A1(net4450),
    .A2(_02374_));
 sg13g2_a21oi_1 _27840_ (.A1(net4450),
    .A2(_02367_),
    .Y(_02376_),
    .B1(_02375_));
 sg13g2_mux2_1 _27841_ (.A0(_02373_),
    .A1(_14254_),
    .S(_02376_),
    .X(_00516_));
 sg13g2_nand2_1 _27842_ (.Y(_02377_),
    .A(\u_inv.counter[8] ),
    .B(net5632));
 sg13g2_nor4_1 _27843_ (.A(_14251_),
    .B(_14822_),
    .C(_02354_),
    .D(_02377_),
    .Y(_02378_));
 sg13g2_o21ai_1 _27844_ (.B1(net2633),
    .Y(_02379_),
    .A1(_02367_),
    .A2(_02377_));
 sg13g2_nor3_1 _27845_ (.A(net2633),
    .B(_02367_),
    .C(_02377_),
    .Y(_02380_));
 sg13g2_a21oi_1 _27846_ (.A1(net4389),
    .A2(_02378_),
    .Y(_02381_),
    .B1(_02380_));
 sg13g2_o21ai_1 _27847_ (.B1(_02381_),
    .Y(_00517_),
    .A1(_20877_[0]),
    .A2(net2634));
 sg13g2_a21oi_2 _27848_ (.B1(_19016_),
    .Y(_02382_),
    .A2(_14811_),
    .A1(inv_done));
 sg13g2_nand2_2 _27849_ (.Y(_02383_),
    .A(_19014_),
    .B(_19015_));
 sg13g2_nor2_1 _27850_ (.A(\u_inv.d_reg[231] ),
    .B(\u_inv.d_reg[230] ),
    .Y(_02384_));
 sg13g2_nand2_1 _27851_ (.Y(_02385_),
    .A(_14664_),
    .B(_14665_));
 sg13g2_nand3_1 _27852_ (.B(_14664_),
    .C(_14665_),
    .A(_14663_),
    .Y(_02386_));
 sg13g2_nor4_1 _27853_ (.A(\u_inv.d_reg[159] ),
    .B(\u_inv.d_reg[158] ),
    .C(\u_inv.d_reg[147] ),
    .D(_02386_),
    .Y(_02387_));
 sg13g2_nor2_1 _27854_ (.A(\u_inv.d_reg[149] ),
    .B(\u_inv.d_reg[148] ),
    .Y(_02388_));
 sg13g2_nor3_1 _27855_ (.A(\u_inv.d_reg[150] ),
    .B(\u_inv.d_reg[149] ),
    .C(\u_inv.d_reg[148] ),
    .Y(_02389_));
 sg13g2_and2_1 _27856_ (.A(_14658_),
    .B(_02389_),
    .X(_02390_));
 sg13g2_nor2_1 _27857_ (.A(\u_inv.d_reg[153] ),
    .B(\u_inv.d_reg[152] ),
    .Y(_02391_));
 sg13g2_nand2_1 _27858_ (.Y(_02392_),
    .A(_02390_),
    .B(_02391_));
 sg13g2_nor2_1 _27859_ (.A(\u_inv.d_reg[156] ),
    .B(\u_inv.d_reg[155] ),
    .Y(_02393_));
 sg13g2_nand4_1 _27860_ (.B(_14655_),
    .C(_02391_),
    .A(_14652_),
    .Y(_02394_),
    .D(_02393_));
 sg13g2_inv_1 _27861_ (.Y(_02395_),
    .A(_02394_));
 sg13g2_nand3_1 _27862_ (.B(_02390_),
    .C(_02395_),
    .A(_02387_),
    .Y(_02396_));
 sg13g2_nand2_1 _27863_ (.Y(_02397_),
    .A(_14552_),
    .B(_14808_));
 sg13g2_nor2_1 _27864_ (.A(\u_inv.d_reg[2] ),
    .B(_02397_),
    .Y(_02398_));
 sg13g2_or4_1 _27865_ (.A(\u_inv.d_reg[0] ),
    .B(\u_inv.d_reg[3] ),
    .C(\u_inv.d_reg[2] ),
    .D(\u_inv.d_reg[1] ),
    .X(_02399_));
 sg13g2_inv_1 _27866_ (.Y(_02400_),
    .A(_02399_));
 sg13g2_nand2b_1 _27867_ (.Y(_02401_),
    .B(_14805_),
    .A_N(_02399_));
 sg13g2_or4_1 _27868_ (.A(\u_inv.d_reg[6] ),
    .B(\u_inv.d_reg[5] ),
    .C(\u_inv.d_reg[4] ),
    .D(_02399_),
    .X(_02402_));
 sg13g2_nor3_1 _27869_ (.A(\u_inv.d_reg[8] ),
    .B(\u_inv.d_reg[7] ),
    .C(_02402_),
    .Y(_02403_));
 sg13g2_or4_1 _27870_ (.A(\u_inv.d_reg[9] ),
    .B(\u_inv.d_reg[8] ),
    .C(\u_inv.d_reg[7] ),
    .D(_02402_),
    .X(_02404_));
 sg13g2_nand2b_2 _27871_ (.Y(_02405_),
    .B(_14799_),
    .A_N(_02404_));
 sg13g2_or4_1 _27872_ (.A(\u_inv.d_reg[12] ),
    .B(net5874),
    .C(\u_inv.d_reg[10] ),
    .D(_02404_),
    .X(_02406_));
 sg13g2_nor3_1 _27873_ (.A(\u_inv.d_reg[14] ),
    .B(\u_inv.d_reg[13] ),
    .C(_02406_),
    .Y(_02407_));
 sg13g2_or4_1 _27874_ (.A(\u_inv.d_reg[15] ),
    .B(\u_inv.d_reg[14] ),
    .C(\u_inv.d_reg[13] ),
    .D(_02406_),
    .X(_02408_));
 sg13g2_nor3_1 _27875_ (.A(\u_inv.d_reg[17] ),
    .B(net5873),
    .C(_02408_),
    .Y(_02409_));
 sg13g2_or4_1 _27876_ (.A(\u_inv.d_reg[18] ),
    .B(\u_inv.d_reg[17] ),
    .C(\u_inv.d_reg[16] ),
    .D(_02408_),
    .X(_02410_));
 sg13g2_nor3_1 _27877_ (.A(\u_inv.d_reg[20] ),
    .B(\u_inv.d_reg[19] ),
    .C(_02410_),
    .Y(_02411_));
 sg13g2_or4_1 _27878_ (.A(\u_inv.d_reg[21] ),
    .B(\u_inv.d_reg[20] ),
    .C(\u_inv.d_reg[19] ),
    .D(_02410_),
    .X(_02412_));
 sg13g2_nor3_1 _27879_ (.A(\u_inv.d_reg[23] ),
    .B(\u_inv.d_reg[22] ),
    .C(_02412_),
    .Y(_02413_));
 sg13g2_or4_1 _27880_ (.A(\u_inv.d_reg[24] ),
    .B(\u_inv.d_reg[23] ),
    .C(\u_inv.d_reg[22] ),
    .D(_02412_),
    .X(_02414_));
 sg13g2_nor3_1 _27881_ (.A(\u_inv.d_reg[26] ),
    .B(\u_inv.d_reg[25] ),
    .C(_02414_),
    .Y(_02415_));
 sg13g2_nor4_2 _27882_ (.A(\u_inv.d_reg[27] ),
    .B(\u_inv.d_reg[26] ),
    .C(\u_inv.d_reg[25] ),
    .Y(_02416_),
    .D(_02414_));
 sg13g2_nor2_1 _27883_ (.A(\u_inv.d_reg[29] ),
    .B(\u_inv.d_reg[28] ),
    .Y(_02417_));
 sg13g2_nand2_1 _27884_ (.Y(_02418_),
    .A(_02416_),
    .B(_02417_));
 sg13g2_nand4_1 _27885_ (.B(_14779_),
    .C(_02416_),
    .A(_14778_),
    .Y(_02419_),
    .D(_02417_));
 sg13g2_nor2_1 _27886_ (.A(\u_inv.d_reg[33] ),
    .B(\u_inv.d_reg[32] ),
    .Y(_02420_));
 sg13g2_nand2b_2 _27887_ (.Y(_02421_),
    .B(_02420_),
    .A_N(_02419_));
 sg13g2_nand2_1 _27888_ (.Y(_02422_),
    .A(_14772_),
    .B(_14773_));
 sg13g2_nor2_1 _27889_ (.A(\u_inv.d_reg[38] ),
    .B(_02422_),
    .Y(_02423_));
 sg13g2_inv_1 _27890_ (.Y(_02424_),
    .A(_02423_));
 sg13g2_nor3_1 _27891_ (.A(\u_inv.d_reg[39] ),
    .B(\u_inv.d_reg[35] ),
    .C(\u_inv.d_reg[34] ),
    .Y(_02425_));
 sg13g2_nand3_1 _27892_ (.B(_02423_),
    .C(_02425_),
    .A(_02420_),
    .Y(_02426_));
 sg13g2_or4_1 _27893_ (.A(\u_inv.d_reg[41] ),
    .B(\u_inv.d_reg[40] ),
    .C(_02419_),
    .D(_02426_),
    .X(_02427_));
 sg13g2_nor4_1 _27894_ (.A(\u_inv.d_reg[43] ),
    .B(\u_inv.d_reg[42] ),
    .C(\u_inv.d_reg[41] ),
    .D(\u_inv.d_reg[40] ),
    .Y(_02428_));
 sg13g2_inv_1 _27895_ (.Y(_02429_),
    .A(_02428_));
 sg13g2_or3_1 _27896_ (.A(_02419_),
    .B(_02426_),
    .C(_02429_),
    .X(_02430_));
 sg13g2_nor3_1 _27897_ (.A(\u_inv.d_reg[45] ),
    .B(\u_inv.d_reg[44] ),
    .C(_02430_),
    .Y(_02431_));
 sg13g2_nand4_1 _27898_ (.B(_14763_),
    .C(_14764_),
    .A(_14762_),
    .Y(_02432_),
    .D(_14765_));
 sg13g2_or4_1 _27899_ (.A(_02419_),
    .B(_02426_),
    .C(_02429_),
    .D(_02432_),
    .X(_02433_));
 sg13g2_nand3b_1 _27900_ (.B(_14761_),
    .C(_14760_),
    .Y(_02434_),
    .A_N(_02433_));
 sg13g2_nand4_1 _27901_ (.B(_14759_),
    .C(_14760_),
    .A(_14758_),
    .Y(_02435_),
    .D(_14761_));
 sg13g2_or2_1 _27902_ (.X(_02436_),
    .B(_02435_),
    .A(_02433_));
 sg13g2_nand2_1 _27903_ (.Y(_02437_),
    .A(_14756_),
    .B(_14757_));
 sg13g2_or2_1 _27904_ (.X(_02438_),
    .B(_02437_),
    .A(_02436_));
 sg13g2_nand2_1 _27905_ (.Y(_02439_),
    .A(_14754_),
    .B(_14755_));
 sg13g2_or4_1 _27906_ (.A(_02433_),
    .B(_02435_),
    .C(_02437_),
    .D(_02439_),
    .X(_02440_));
 sg13g2_nor3_1 _27907_ (.A(\u_inv.d_reg[57] ),
    .B(\u_inv.d_reg[56] ),
    .C(_02440_),
    .Y(_02441_));
 sg13g2_nand4_1 _27908_ (.B(_14751_),
    .C(_14752_),
    .A(_14750_),
    .Y(_02442_),
    .D(_14753_));
 sg13g2_or2_1 _27909_ (.X(_02443_),
    .B(_02442_),
    .A(_02440_));
 sg13g2_nand2_1 _27910_ (.Y(_02444_),
    .A(_14748_),
    .B(_14749_));
 sg13g2_or2_1 _27911_ (.X(_02445_),
    .B(_02444_),
    .A(_02443_));
 sg13g2_nand2_1 _27912_ (.Y(_02446_),
    .A(_14746_),
    .B(_14747_));
 sg13g2_or4_1 _27913_ (.A(_02440_),
    .B(_02442_),
    .C(_02444_),
    .D(_02446_),
    .X(_02447_));
 sg13g2_nand2_1 _27914_ (.Y(_02448_),
    .A(_14744_),
    .B(_14745_));
 sg13g2_nand4_1 _27915_ (.B(_14743_),
    .C(_14744_),
    .A(_14742_),
    .Y(_02449_),
    .D(_14745_));
 sg13g2_or2_1 _27916_ (.X(_02450_),
    .B(_02449_),
    .A(_02447_));
 sg13g2_nand2_1 _27917_ (.Y(_02451_),
    .A(_14740_),
    .B(_14741_));
 sg13g2_or2_1 _27918_ (.X(_02452_),
    .B(_02451_),
    .A(_02450_));
 sg13g2_nand2_1 _27919_ (.Y(_02453_),
    .A(_14738_),
    .B(_14739_));
 sg13g2_or4_1 _27920_ (.A(_02447_),
    .B(_02449_),
    .C(_02451_),
    .D(_02453_),
    .X(_02454_));
 sg13g2_nand2_1 _27921_ (.Y(_02455_),
    .A(_14736_),
    .B(_14737_));
 sg13g2_nand4_1 _27922_ (.B(_14735_),
    .C(_14736_),
    .A(_14734_),
    .Y(_02456_),
    .D(_14737_));
 sg13g2_nand4_1 _27923_ (.B(_14731_),
    .C(_14732_),
    .A(_14730_),
    .Y(_02457_),
    .D(_14733_));
 sg13g2_nor3_2 _27924_ (.A(_02454_),
    .B(_02456_),
    .C(_02457_),
    .Y(_02458_));
 sg13g2_nor2_1 _27925_ (.A(\u_inv.d_reg[81] ),
    .B(\u_inv.d_reg[80] ),
    .Y(_02459_));
 sg13g2_nor3_1 _27926_ (.A(\u_inv.d_reg[82] ),
    .B(\u_inv.d_reg[81] ),
    .C(\u_inv.d_reg[80] ),
    .Y(_02460_));
 sg13g2_and2_1 _27927_ (.A(_14726_),
    .B(_02460_),
    .X(_02461_));
 sg13g2_nand2_1 _27928_ (.Y(_02462_),
    .A(_14725_),
    .B(_02461_));
 sg13g2_nor2_1 _27929_ (.A(\u_inv.d_reg[85] ),
    .B(_02462_),
    .Y(_02463_));
 sg13g2_nand3_1 _27930_ (.B(_14723_),
    .C(_02463_),
    .A(_14722_),
    .Y(_02464_));
 sg13g2_nor4_2 _27931_ (.A(_02454_),
    .B(_02456_),
    .C(_02457_),
    .Y(_02465_),
    .D(_02464_));
 sg13g2_nand2_1 _27932_ (.Y(_02466_),
    .A(_14720_),
    .B(_14721_));
 sg13g2_nor3_2 _27933_ (.A(\u_inv.d_reg[91] ),
    .B(net5871),
    .C(_02466_),
    .Y(_02467_));
 sg13g2_nor4_1 _27934_ (.A(\u_inv.d_reg[95] ),
    .B(\u_inv.d_reg[94] ),
    .C(\u_inv.d_reg[93] ),
    .D(\u_inv.d_reg[92] ),
    .Y(_02468_));
 sg13g2_nand3_1 _27935_ (.B(_02467_),
    .C(_02468_),
    .A(_02465_),
    .Y(_02469_));
 sg13g2_nor4_1 _27936_ (.A(\u_inv.d_reg[99] ),
    .B(net5870),
    .C(\u_inv.d_reg[97] ),
    .D(\u_inv.d_reg[96] ),
    .Y(_02470_));
 sg13g2_nand4_1 _27937_ (.B(_02467_),
    .C(_02468_),
    .A(_02465_),
    .Y(_02471_),
    .D(_02470_));
 sg13g2_nand2_1 _27938_ (.Y(_02472_),
    .A(_14708_),
    .B(_14709_));
 sg13g2_nor2_1 _27939_ (.A(_02471_),
    .B(_02472_),
    .Y(_02473_));
 sg13g2_nand2_1 _27940_ (.Y(_02474_),
    .A(_14706_),
    .B(_14707_));
 sg13g2_nand3_1 _27941_ (.B(_14707_),
    .C(_02473_),
    .A(_14706_),
    .Y(_02475_));
 sg13g2_nand2_1 _27942_ (.Y(_02476_),
    .A(_14704_),
    .B(_14705_));
 sg13g2_nor4_1 _27943_ (.A(_02471_),
    .B(_02472_),
    .C(_02474_),
    .D(_02476_),
    .Y(_02477_));
 sg13g2_nor4_1 _27944_ (.A(\u_inv.d_reg[107] ),
    .B(\u_inv.d_reg[106] ),
    .C(_02475_),
    .D(_02476_),
    .Y(_02478_));
 sg13g2_nor4_1 _27945_ (.A(\u_inv.d_reg[111] ),
    .B(\u_inv.d_reg[110] ),
    .C(\u_inv.d_reg[109] ),
    .D(\u_inv.d_reg[108] ),
    .Y(_02479_));
 sg13g2_nand4_1 _27946_ (.B(_14703_),
    .C(_02477_),
    .A(_14702_),
    .Y(_02480_),
    .D(_02479_));
 sg13g2_nand4_1 _27947_ (.B(_14695_),
    .C(_14696_),
    .A(_14694_),
    .Y(_02481_),
    .D(_14697_));
 sg13g2_or2_1 _27948_ (.X(_02482_),
    .B(_02481_),
    .A(_02480_));
 sg13g2_nand2_1 _27949_ (.Y(_02483_),
    .A(_14692_),
    .B(_14693_));
 sg13g2_or2_1 _27950_ (.X(_02484_),
    .B(_02483_),
    .A(_02482_));
 sg13g2_nand2_1 _27951_ (.Y(_02485_),
    .A(_14690_),
    .B(_14691_));
 sg13g2_nor4_2 _27952_ (.A(_02485_),
    .B(_02481_),
    .C(_02483_),
    .Y(_02486_),
    .D(_02480_));
 sg13g2_nor2_1 _27953_ (.A(\u_inv.d_reg[121] ),
    .B(\u_inv.d_reg[120] ),
    .Y(_02487_));
 sg13g2_nor3_1 _27954_ (.A(\u_inv.d_reg[122] ),
    .B(\u_inv.d_reg[121] ),
    .C(\u_inv.d_reg[120] ),
    .Y(_02488_));
 sg13g2_nand2_1 _27955_ (.Y(_02489_),
    .A(_14686_),
    .B(_02488_));
 sg13g2_nand3_1 _27956_ (.B(_14686_),
    .C(_02488_),
    .A(_14685_),
    .Y(_02490_));
 sg13g2_nor4_2 _27957_ (.A(\u_inv.d_reg[127] ),
    .B(\u_inv.d_reg[126] ),
    .C(\u_inv.d_reg[125] ),
    .Y(_02491_),
    .D(_02490_));
 sg13g2_nand2_2 _27958_ (.Y(_02492_),
    .A(net1073),
    .B(_02491_));
 sg13g2_nand2_1 _27959_ (.Y(_02493_),
    .A(_14680_),
    .B(_14681_));
 sg13g2_nand3_1 _27960_ (.B(_14680_),
    .C(_14681_),
    .A(_14679_),
    .Y(_02494_));
 sg13g2_nor3_1 _27961_ (.A(\u_inv.d_reg[142] ),
    .B(\u_inv.d_reg[141] ),
    .C(net5869),
    .Y(_02495_));
 sg13g2_nand2_1 _27962_ (.Y(_02496_),
    .A(_14672_),
    .B(_14673_));
 sg13g2_nand3_1 _27963_ (.B(_14672_),
    .C(_14673_),
    .A(_14671_),
    .Y(_02497_));
 sg13g2_nand2_1 _27964_ (.Y(_02498_),
    .A(_14676_),
    .B(_14677_));
 sg13g2_nor3_1 _27965_ (.A(\u_inv.d_reg[135] ),
    .B(\u_inv.d_reg[134] ),
    .C(_02498_),
    .Y(_02499_));
 sg13g2_nor2_1 _27966_ (.A(\u_inv.d_reg[139] ),
    .B(_02497_),
    .Y(_02500_));
 sg13g2_nor2_2 _27967_ (.A(\u_inv.d_reg[131] ),
    .B(_02494_),
    .Y(_02501_));
 sg13g2_and2_1 _27968_ (.A(_14666_),
    .B(_02495_),
    .X(_02502_));
 sg13g2_nand4_1 _27969_ (.B(_02500_),
    .C(_02501_),
    .A(_02499_),
    .Y(_02503_),
    .D(_02502_));
 sg13g2_or2_1 _27970_ (.X(_02504_),
    .B(_02503_),
    .A(_02492_));
 sg13g2_or3_1 _27971_ (.A(_02396_),
    .B(_02492_),
    .C(_02503_),
    .X(_02505_));
 sg13g2_nor4_1 _27972_ (.A(\u_inv.d_reg[171] ),
    .B(\u_inv.d_reg[170] ),
    .C(\u_inv.d_reg[169] ),
    .D(\u_inv.d_reg[168] ),
    .Y(_02506_));
 sg13g2_nor3_1 _27973_ (.A(\u_inv.d_reg[167] ),
    .B(\u_inv.d_reg[166] ),
    .C(\u_inv.d_reg[163] ),
    .Y(_02507_));
 sg13g2_nor3_1 _27974_ (.A(\u_inv.d_reg[162] ),
    .B(\u_inv.d_reg[161] ),
    .C(net5868),
    .Y(_02508_));
 sg13g2_nand4_1 _27975_ (.B(_14645_),
    .C(_02507_),
    .A(_14644_),
    .Y(_02509_),
    .D(_02508_));
 sg13g2_nand4_1 _27976_ (.B(_14636_),
    .C(_14637_),
    .A(_14635_),
    .Y(_02510_),
    .D(_02506_));
 sg13g2_or4_1 _27977_ (.A(\u_inv.d_reg[175] ),
    .B(_02505_),
    .C(_02509_),
    .D(_02510_),
    .X(_02511_));
 sg13g2_nand3_1 _27978_ (.B(_14629_),
    .C(_14630_),
    .A(_14628_),
    .Y(_02512_));
 sg13g2_nor2_1 _27979_ (.A(\u_inv.d_reg[182] ),
    .B(_02512_),
    .Y(_02513_));
 sg13g2_inv_1 _27980_ (.Y(_02514_),
    .A(_02513_));
 sg13g2_nand2_2 _27981_ (.Y(_02515_),
    .A(_14632_),
    .B(_14633_));
 sg13g2_nor2_1 _27982_ (.A(\u_inv.d_reg[178] ),
    .B(_02515_),
    .Y(_02516_));
 sg13g2_nor4_1 _27983_ (.A(\u_inv.d_reg[183] ),
    .B(\u_inv.d_reg[178] ),
    .C(_02514_),
    .D(_02515_),
    .Y(_02517_));
 sg13g2_nor2b_1 _27984_ (.A(_02511_),
    .B_N(_02517_),
    .Y(_02518_));
 sg13g2_nand2b_1 _27985_ (.Y(_02519_),
    .B(_02517_),
    .A_N(_02511_));
 sg13g2_nor2_1 _27986_ (.A(\u_inv.d_reg[185] ),
    .B(net5866),
    .Y(_02520_));
 sg13g2_nor4_2 _27987_ (.A(\u_inv.d_reg[186] ),
    .B(\u_inv.d_reg[185] ),
    .C(\u_inv.d_reg[184] ),
    .Y(_02521_),
    .D(_02519_));
 sg13g2_nor3_1 _27988_ (.A(\u_inv.d_reg[189] ),
    .B(\u_inv.d_reg[188] ),
    .C(\u_inv.d_reg[187] ),
    .Y(_02522_));
 sg13g2_nand4_1 _27989_ (.B(_14619_),
    .C(_02521_),
    .A(_14618_),
    .Y(_02523_),
    .D(_02522_));
 sg13g2_nor3_1 _27990_ (.A(\u_inv.d_reg[194] ),
    .B(\u_inv.d_reg[193] ),
    .C(\u_inv.d_reg[192] ),
    .Y(_02524_));
 sg13g2_inv_1 _27991_ (.Y(_02525_),
    .A(_02524_));
 sg13g2_nand4_1 _27992_ (.B(_14613_),
    .C(_14614_),
    .A(_14612_),
    .Y(_02526_),
    .D(_02524_));
 sg13g2_or4_1 _27993_ (.A(\u_inv.d_reg[199] ),
    .B(\u_inv.d_reg[198] ),
    .C(_02523_),
    .D(_02526_),
    .X(_02527_));
 sg13g2_nand2_1 _27994_ (.Y(_02528_),
    .A(_14608_),
    .B(_14609_));
 sg13g2_nand3_1 _27995_ (.B(_14608_),
    .C(_14609_),
    .A(_14607_),
    .Y(_02529_));
 sg13g2_nand2b_1 _27996_ (.Y(_02530_),
    .B(_14606_),
    .A_N(_02529_));
 sg13g2_nand2b_1 _27997_ (.Y(_02531_),
    .B(_14605_),
    .A_N(_02530_));
 sg13g2_nand2b_1 _27998_ (.Y(_02532_),
    .B(_14604_),
    .A_N(_02531_));
 sg13g2_nor4_2 _27999_ (.A(\u_inv.d_reg[207] ),
    .B(\u_inv.d_reg[206] ),
    .C(_02527_),
    .Y(_02533_),
    .D(_02532_));
 sg13g2_nand4_1 _28000_ (.B(_14599_),
    .C(_14600_),
    .A(_14598_),
    .Y(_02534_),
    .D(_14601_));
 sg13g2_nor3_1 _28001_ (.A(\u_inv.d_reg[213] ),
    .B(\u_inv.d_reg[212] ),
    .C(_02534_),
    .Y(_02535_));
 sg13g2_nand2_1 _28002_ (.Y(_02536_),
    .A(_02533_),
    .B(_02535_));
 sg13g2_nand4_1 _28003_ (.B(_14595_),
    .C(_02533_),
    .A(_14594_),
    .Y(_02537_),
    .D(_02535_));
 sg13g2_nand3_1 _28004_ (.B(_14589_),
    .C(_14590_),
    .A(_14588_),
    .Y(_02538_));
 sg13g2_nand2b_1 _28005_ (.Y(_02539_),
    .B(_14587_),
    .A_N(_02538_));
 sg13g2_nand2_1 _28006_ (.Y(_02540_),
    .A(_14592_),
    .B(_14593_));
 sg13g2_nand3_1 _28007_ (.B(_14592_),
    .C(_14593_),
    .A(_14591_),
    .Y(_02541_));
 sg13g2_or4_1 _28008_ (.A(\u_inv.d_reg[223] ),
    .B(_02537_),
    .C(_02539_),
    .D(_02541_),
    .X(_02542_));
 sg13g2_nand4_1 _28009_ (.B(_14581_),
    .C(_14582_),
    .A(_14580_),
    .Y(_02543_),
    .D(_14583_));
 sg13g2_nor4_2 _28010_ (.A(\u_inv.d_reg[225] ),
    .B(\u_inv.d_reg[224] ),
    .C(_02542_),
    .Y(_02544_),
    .D(_02543_));
 sg13g2_nand2_1 _28011_ (.Y(_02545_),
    .A(_02384_),
    .B(_02544_));
 sg13g2_nor4_1 _28012_ (.A(\u_inv.d_reg[235] ),
    .B(\u_inv.d_reg[234] ),
    .C(\u_inv.d_reg[233] ),
    .D(\u_inv.d_reg[232] ),
    .Y(_02546_));
 sg13g2_nand3_1 _28013_ (.B(_02544_),
    .C(_02546_),
    .A(_02384_),
    .Y(_02547_));
 sg13g2_nor4_1 _28014_ (.A(\u_inv.d_reg[239] ),
    .B(\u_inv.d_reg[238] ),
    .C(\u_inv.d_reg[237] ),
    .D(\u_inv.d_reg[236] ),
    .Y(_02548_));
 sg13g2_nand2b_2 _28015_ (.Y(_02549_),
    .B(_02548_),
    .A_N(_02547_));
 sg13g2_nor4_1 _28016_ (.A(\u_inv.d_reg[243] ),
    .B(\u_inv.d_reg[242] ),
    .C(\u_inv.d_reg[241] ),
    .D(net5865),
    .Y(_02550_));
 sg13g2_nand2b_1 _28017_ (.Y(_02551_),
    .B(_02550_),
    .A_N(_02549_));
 sg13g2_nand3b_1 _28018_ (.B(_14565_),
    .C(_14564_),
    .Y(_02552_),
    .A_N(_02551_));
 sg13g2_nand3b_1 _28019_ (.B(_14563_),
    .C(_14562_),
    .Y(_02553_),
    .A_N(_02552_));
 sg13g2_and2_1 _28020_ (.A(net5830),
    .B(_02553_),
    .X(_02554_));
 sg13g2_nand4_1 _28021_ (.B(_14559_),
    .C(_14560_),
    .A(_14558_),
    .Y(_02555_),
    .D(_14561_));
 sg13g2_nand2b_1 _28022_ (.Y(_02556_),
    .B(_14557_),
    .A_N(_02555_));
 sg13g2_or4_1 _28023_ (.A(\u_inv.d_reg[255] ),
    .B(\u_inv.d_reg[254] ),
    .C(\u_inv.d_reg[253] ),
    .D(_02556_),
    .X(_02557_));
 sg13g2_o21ai_1 _28024_ (.B1(net5831),
    .Y(_02558_),
    .A1(_02553_),
    .A2(_02557_));
 sg13g2_xnor2_1 _28025_ (.Y(_02559_),
    .A(\u_inv.d_reg[256] ),
    .B(_02558_));
 sg13g2_xnor2_1 _28026_ (.Y(_02560_),
    .A(_02558_),
    .B(_14553_));
 sg13g2_o21ai_1 _28027_ (.B1(net5830),
    .Y(_02561_),
    .A1(_02553_),
    .A2(_02556_));
 sg13g2_o21ai_1 _28028_ (.B1(net5830),
    .Y(_02562_),
    .A1(\u_inv.d_reg[254] ),
    .A2(\u_inv.d_reg[253] ));
 sg13g2_nand2_1 _28029_ (.Y(_02563_),
    .A(_02561_),
    .B(_02562_));
 sg13g2_xnor2_1 _28030_ (.Y(_02564_),
    .A(\u_inv.d_reg[255] ),
    .B(_02563_));
 sg13g2_nor3_1 _28031_ (.A(\u_inv.d_reg[249] ),
    .B(\u_inv.d_reg[248] ),
    .C(_02553_),
    .Y(_02565_));
 sg13g2_nor2_1 _28032_ (.A(net5635),
    .B(_02565_),
    .Y(_02566_));
 sg13g2_xnor2_1 _28033_ (.Y(_02567_),
    .A(\u_inv.d_reg[250] ),
    .B(_02566_));
 sg13g2_inv_1 _28034_ (.Y(_02568_),
    .A(_02567_));
 sg13g2_and2_1 _28035_ (.A(net5830),
    .B(_02551_),
    .X(_02569_));
 sg13g2_nor2_1 _28036_ (.A(net5865),
    .B(_02549_),
    .Y(_02570_));
 sg13g2_nor4_1 _28037_ (.A(\u_inv.d_reg[242] ),
    .B(\u_inv.d_reg[241] ),
    .C(net5865),
    .D(_02549_),
    .Y(_02571_));
 sg13g2_o21ai_1 _28038_ (.B1(_02569_),
    .Y(_02572_),
    .A1(_14566_),
    .A2(_02571_));
 sg13g2_o21ai_1 _28039_ (.B1(_02572_),
    .Y(_02573_),
    .A1(net5831),
    .A2(_14566_));
 sg13g2_nor3_1 _28040_ (.A(\u_inv.d_reg[237] ),
    .B(\u_inv.d_reg[236] ),
    .C(_02547_),
    .Y(_02574_));
 sg13g2_nor2_1 _28041_ (.A(net5635),
    .B(_02574_),
    .Y(_02575_));
 sg13g2_xnor2_1 _28042_ (.Y(_02576_),
    .A(_14571_),
    .B(_02575_));
 sg13g2_nand2_1 _28043_ (.Y(_02577_),
    .A(net5833),
    .B(_02547_));
 sg13g2_inv_1 _28044_ (.Y(_02578_),
    .A(_02577_));
 sg13g2_nand4_1 _28045_ (.B(_14577_),
    .C(_02384_),
    .A(_14576_),
    .Y(_02579_),
    .D(_02544_));
 sg13g2_o21ai_1 _28046_ (.B1(\u_inv.d_reg[235] ),
    .Y(_02580_),
    .A1(\u_inv.d_reg[234] ),
    .A2(_02579_));
 sg13g2_a22oi_1 _28047_ (.Y(_02581_),
    .B1(_02578_),
    .B2(_02580_),
    .A2(\u_inv.d_reg[235] ),
    .A1(net5635));
 sg13g2_nor2_1 _28048_ (.A(net5635),
    .B(_02570_),
    .Y(_02582_));
 sg13g2_xnor2_1 _28049_ (.Y(_02583_),
    .A(\u_inv.d_reg[241] ),
    .B(_02582_));
 sg13g2_nor2_1 _28050_ (.A(_02581_),
    .B(_02583_),
    .Y(_02584_));
 sg13g2_nand2_1 _28051_ (.Y(_02585_),
    .A(net5830),
    .B(_02552_));
 sg13g2_o21ai_1 _28052_ (.B1(net5830),
    .Y(_02586_),
    .A1(\u_inv.d_reg[246] ),
    .A2(_02552_));
 sg13g2_xnor2_1 _28053_ (.Y(_02587_),
    .A(\u_inv.d_reg[247] ),
    .B(_02586_));
 sg13g2_xnor2_1 _28054_ (.Y(_02588_),
    .A(\u_inv.d_reg[248] ),
    .B(_02554_));
 sg13g2_nor2b_1 _28055_ (.A(_02588_),
    .B_N(_02587_),
    .Y(_02589_));
 sg13g2_nand4_1 _28056_ (.B(_02576_),
    .C(_02584_),
    .A(_02573_),
    .Y(_02590_),
    .D(_02589_));
 sg13g2_xnor2_1 _28057_ (.Y(_02591_),
    .A(\u_inv.d_reg[246] ),
    .B(_02585_));
 sg13g2_nand2_1 _28058_ (.Y(_02592_),
    .A(net5831),
    .B(_02549_));
 sg13g2_a21oi_1 _28059_ (.A1(_14571_),
    .A2(_02574_),
    .Y(_02593_),
    .B1(_14570_));
 sg13g2_nand2_1 _28060_ (.Y(_02594_),
    .A(net5635),
    .B(\u_inv.d_reg[239] ));
 sg13g2_o21ai_1 _28061_ (.B1(_02594_),
    .Y(_02595_),
    .A1(_02592_),
    .A2(_02593_));
 sg13g2_a21oi_1 _28062_ (.A1(_14568_),
    .A2(_02570_),
    .Y(_02596_),
    .B1(net5635));
 sg13g2_xnor2_1 _28063_ (.Y(_02597_),
    .A(_14567_),
    .B(_02596_));
 sg13g2_nand3_1 _28064_ (.B(_02595_),
    .C(_02597_),
    .A(_02591_),
    .Y(_02598_));
 sg13g2_nor3_1 _28065_ (.A(\u_inv.d_reg[225] ),
    .B(\u_inv.d_reg[224] ),
    .C(_02542_),
    .Y(_02599_));
 sg13g2_and2_1 _28066_ (.A(net5835),
    .B(_02542_),
    .X(_02600_));
 sg13g2_nor2_1 _28067_ (.A(net5636),
    .B(_02599_),
    .Y(_02601_));
 sg13g2_a21oi_1 _28068_ (.A1(net5832),
    .A2(\u_inv.d_reg[226] ),
    .Y(_02602_),
    .B1(_02601_));
 sg13g2_xnor2_1 _28069_ (.Y(_02603_),
    .A(\u_inv.d_reg[227] ),
    .B(_02602_));
 sg13g2_xnor2_1 _28070_ (.Y(_02604_),
    .A(_14582_),
    .B(_02602_));
 sg13g2_nor2_2 _28071_ (.A(net5638),
    .B(_02533_),
    .Y(_02605_));
 sg13g2_a21oi_1 _28072_ (.A1(net5836),
    .A2(_02534_),
    .Y(_02606_),
    .B1(_02605_));
 sg13g2_xnor2_1 _28073_ (.Y(_02607_),
    .A(\u_inv.d_reg[212] ),
    .B(_02606_));
 sg13g2_o21ai_1 _28074_ (.B1(_02606_),
    .Y(_02608_),
    .A1(net5637),
    .A2(_14597_));
 sg13g2_xnor2_1 _28075_ (.Y(_02609_),
    .A(_14596_),
    .B(_02608_));
 sg13g2_nand2_2 _28076_ (.Y(_02610_),
    .A(_02607_),
    .B(_02609_));
 sg13g2_nor2_1 _28077_ (.A(net5636),
    .B(_02544_),
    .Y(_02611_));
 sg13g2_xnor2_1 _28078_ (.Y(_02612_),
    .A(\u_inv.d_reg[230] ),
    .B(_02611_));
 sg13g2_or2_1 _28079_ (.X(_02613_),
    .B(_02541_),
    .A(_02537_));
 sg13g2_o21ai_1 _28080_ (.B1(net5835),
    .Y(_02614_),
    .A1(_02538_),
    .A2(_02613_));
 sg13g2_o21ai_1 _28081_ (.B1(net5835),
    .Y(_02615_),
    .A1(_02539_),
    .A2(_02613_));
 sg13g2_xnor2_1 _28082_ (.Y(_02616_),
    .A(_14586_),
    .B(_02615_));
 sg13g2_xnor2_1 _28083_ (.Y(_02617_),
    .A(\u_inv.d_reg[222] ),
    .B(_02614_));
 sg13g2_inv_2 _28084_ (.Y(_02618_),
    .A(_02617_));
 sg13g2_nor4_2 _28085_ (.A(_02610_),
    .B(_02612_),
    .C(_02616_),
    .Y(_02619_),
    .D(_02618_));
 sg13g2_o21ai_1 _28086_ (.B1(net5832),
    .Y(_02620_),
    .A1(\u_inv.d_reg[227] ),
    .A2(\u_inv.d_reg[226] ));
 sg13g2_nor2b_1 _28087_ (.A(_02601_),
    .B_N(_02620_),
    .Y(_02621_));
 sg13g2_xnor2_1 _28088_ (.Y(_02622_),
    .A(\u_inv.d_reg[228] ),
    .B(_02621_));
 sg13g2_xnor2_1 _28089_ (.Y(_02623_),
    .A(_14573_),
    .B(_02577_));
 sg13g2_inv_1 _28090_ (.Y(_02624_),
    .A(_02623_));
 sg13g2_nand4_1 _28091_ (.B(_02619_),
    .C(_02622_),
    .A(_02603_),
    .Y(_02625_),
    .D(_02624_));
 sg13g2_xnor2_1 _28092_ (.Y(_02626_),
    .A(\u_inv.d_reg[226] ),
    .B(_02601_));
 sg13g2_a21oi_1 _28093_ (.A1(_14579_),
    .A2(_02544_),
    .Y(_02627_),
    .B1(net5636));
 sg13g2_xnor2_1 _28094_ (.Y(_02628_),
    .A(\u_inv.d_reg[231] ),
    .B(_02627_));
 sg13g2_nand2_1 _28095_ (.Y(_02629_),
    .A(net5831),
    .B(_02545_));
 sg13g2_xnor2_1 _28096_ (.Y(_02630_),
    .A(\u_inv.d_reg[232] ),
    .B(_02629_));
 sg13g2_nor2b_1 _28097_ (.A(_02628_),
    .B_N(_02630_),
    .Y(_02631_));
 sg13g2_nand2b_1 _28098_ (.Y(_02632_),
    .B(_02631_),
    .A_N(_02626_));
 sg13g2_nand2_1 _28099_ (.Y(_02633_),
    .A(net5837),
    .B(_02537_));
 sg13g2_xnor2_1 _28100_ (.Y(_02634_),
    .A(_14593_),
    .B(_02633_));
 sg13g2_inv_1 _28101_ (.Y(_02635_),
    .A(_02634_));
 sg13g2_and2_1 _28102_ (.A(net5845),
    .B(_02523_),
    .X(_02636_));
 sg13g2_o21ai_1 _28103_ (.B1(net5841),
    .Y(_02637_),
    .A1(_02523_),
    .A2(_02525_));
 sg13g2_o21ai_1 _28104_ (.B1(net5841),
    .Y(_02638_),
    .A1(_02523_),
    .A2(_02526_));
 sg13g2_inv_1 _28105_ (.Y(_02639_),
    .A(_02638_));
 sg13g2_a21oi_1 _28106_ (.A1(net5842),
    .A2(\u_inv.d_reg[198] ),
    .Y(_02640_),
    .B1(_02639_));
 sg13g2_xnor2_1 _28107_ (.Y(_02641_),
    .A(\u_inv.d_reg[199] ),
    .B(_02640_));
 sg13g2_nand3_1 _28108_ (.B(_14601_),
    .C(_02533_),
    .A(_14600_),
    .Y(_02642_));
 sg13g2_nand2_1 _28109_ (.Y(_02643_),
    .A(net5836),
    .B(_02642_));
 sg13g2_xnor2_1 _28110_ (.Y(_02644_),
    .A(\u_inv.d_reg[210] ),
    .B(_02643_));
 sg13g2_nand2_1 _28111_ (.Y(_02645_),
    .A(net5837),
    .B(_02536_));
 sg13g2_o21ai_1 _28112_ (.B1(net5836),
    .Y(_02646_),
    .A1(\u_inv.d_reg[214] ),
    .A2(_02536_));
 sg13g2_xnor2_1 _28113_ (.Y(_02647_),
    .A(_14594_),
    .B(_02646_));
 sg13g2_inv_1 _28114_ (.Y(_02648_),
    .A(_02647_));
 sg13g2_nand4_1 _28115_ (.B(_02641_),
    .C(_02644_),
    .A(_02635_),
    .Y(_02649_),
    .D(_02648_));
 sg13g2_nor2_1 _28116_ (.A(net5638),
    .B(_02521_),
    .Y(_02650_));
 sg13g2_a21oi_1 _28117_ (.A1(net5846),
    .A2(\u_inv.d_reg[187] ),
    .Y(_02651_),
    .B1(_02650_));
 sg13g2_o21ai_1 _28118_ (.B1(_02651_),
    .Y(_02652_),
    .A1(net5638),
    .A2(_14621_));
 sg13g2_xnor2_1 _28119_ (.Y(_02653_),
    .A(_14620_),
    .B(_02652_));
 sg13g2_xnor2_1 _28120_ (.Y(_02654_),
    .A(\u_inv.d_reg[188] ),
    .B(_02651_));
 sg13g2_nand2_1 _28121_ (.Y(_02655_),
    .A(_02653_),
    .B(_02654_));
 sg13g2_and2_1 _28122_ (.A(net5841),
    .B(_02527_),
    .X(_02656_));
 sg13g2_o21ai_1 _28123_ (.B1(net5841),
    .Y(_02657_),
    .A1(_02527_),
    .A2(_02528_));
 sg13g2_xnor2_1 _28124_ (.Y(_02658_),
    .A(_14607_),
    .B(_02657_));
 sg13g2_xnor2_1 _28125_ (.Y(_02659_),
    .A(\u_inv.d_reg[208] ),
    .B(_02605_));
 sg13g2_o21ai_1 _28126_ (.B1(net5845),
    .Y(_02660_),
    .A1(\u_inv.d_reg[192] ),
    .A2(_02523_));
 sg13g2_inv_1 _28127_ (.Y(_02661_),
    .A(_02660_));
 sg13g2_a21oi_1 _28128_ (.A1(net5845),
    .A2(\u_inv.d_reg[193] ),
    .Y(_02662_),
    .B1(_02661_));
 sg13g2_xnor2_1 _28129_ (.Y(_02663_),
    .A(\u_inv.d_reg[194] ),
    .B(_02662_));
 sg13g2_inv_1 _28130_ (.Y(_02664_),
    .A(_02663_));
 sg13g2_nor4_1 _28131_ (.A(_02655_),
    .B(_02658_),
    .C(_02659_),
    .D(_02664_),
    .Y(_02665_));
 sg13g2_o21ai_1 _28132_ (.B1(net5841),
    .Y(_02666_),
    .A1(_02527_),
    .A2(_02529_));
 sg13g2_xnor2_1 _28133_ (.Y(_02667_),
    .A(_14606_),
    .B(_02666_));
 sg13g2_o21ai_1 _28134_ (.B1(net5841),
    .Y(_02668_),
    .A1(\u_inv.d_reg[200] ),
    .A2(_02527_));
 sg13g2_xnor2_1 _28135_ (.Y(_02669_),
    .A(_14608_),
    .B(_02668_));
 sg13g2_nor2_1 _28136_ (.A(_02667_),
    .B(_02669_),
    .Y(_02670_));
 sg13g2_nand3_1 _28137_ (.B(_02491_),
    .C(_02501_),
    .A(net1073),
    .Y(_02671_));
 sg13g2_nand4_1 _28138_ (.B(_02491_),
    .C(_02499_),
    .A(net1073),
    .Y(_02672_),
    .D(_02501_));
 sg13g2_nor3_1 _28139_ (.A(\u_inv.d_reg[139] ),
    .B(_02497_),
    .C(_02672_),
    .Y(_02673_));
 sg13g2_nor2_2 _28140_ (.A(net5642),
    .B(_02673_),
    .Y(_02674_));
 sg13g2_a21o_1 _28141_ (.A2(_02673_),
    .A1(_02495_),
    .B1(net5642),
    .X(_02675_));
 sg13g2_xnor2_1 _28142_ (.Y(_02676_),
    .A(\u_inv.d_reg[143] ),
    .B(_02675_));
 sg13g2_o21ai_1 _28143_ (.B1(net5853),
    .Y(_02677_),
    .A1(\u_inv.d_reg[141] ),
    .A2(net5869));
 sg13g2_nor2b_1 _28144_ (.A(_02674_),
    .B_N(_02677_),
    .Y(_02678_));
 sg13g2_xnor2_1 _28145_ (.Y(_02679_),
    .A(_14667_),
    .B(_02678_));
 sg13g2_nand2b_2 _28146_ (.Y(_02680_),
    .B(_02676_),
    .A_N(_02679_));
 sg13g2_nor3_1 _28147_ (.A(\u_inv.d_reg[161] ),
    .B(net5868),
    .C(_02505_),
    .Y(_02681_));
 sg13g2_or2_1 _28148_ (.X(_02682_),
    .B(_02509_),
    .A(_02505_));
 sg13g2_nor3_1 _28149_ (.A(\u_inv.d_reg[169] ),
    .B(\u_inv.d_reg[168] ),
    .C(_02682_),
    .Y(_02683_));
 sg13g2_nor2_1 _28150_ (.A(net5640),
    .B(_02683_),
    .Y(_02684_));
 sg13g2_xnor2_1 _28151_ (.Y(_02685_),
    .A(\u_inv.d_reg[170] ),
    .B(_02684_));
 sg13g2_xnor2_1 _28152_ (.Y(_02686_),
    .A(\u_inv.d_reg[192] ),
    .B(_02636_));
 sg13g2_xnor2_1 _28153_ (.Y(_02687_),
    .A(_14617_),
    .B(_02636_));
 sg13g2_nand2_1 _28154_ (.Y(_02688_),
    .A(net5853),
    .B(_02672_));
 sg13g2_o21ai_1 _28155_ (.B1(net5853),
    .Y(_02689_),
    .A1(\u_inv.d_reg[136] ),
    .A2(_02672_));
 sg13g2_xnor2_1 _28156_ (.Y(_02690_),
    .A(\u_inv.d_reg[137] ),
    .B(_02689_));
 sg13g2_xnor2_1 _28157_ (.Y(_02691_),
    .A(_14672_),
    .B(_02689_));
 sg13g2_nor2_1 _28158_ (.A(net5639),
    .B(_02518_),
    .Y(_02692_));
 sg13g2_xnor2_1 _28159_ (.Y(_02693_),
    .A(net5866),
    .B(_02692_));
 sg13g2_and2_1 _28160_ (.A(net5851),
    .B(_02671_),
    .X(_02694_));
 sg13g2_o21ai_1 _28161_ (.B1(net5852),
    .Y(_02695_),
    .A1(\u_inv.d_reg[132] ),
    .A2(_02671_));
 sg13g2_xnor2_1 _28162_ (.Y(_02696_),
    .A(\u_inv.d_reg[133] ),
    .B(_02695_));
 sg13g2_xnor2_1 _28163_ (.Y(_02697_),
    .A(\u_inv.d_reg[132] ),
    .B(_02694_));
 sg13g2_nand2b_2 _28164_ (.Y(_02698_),
    .B(_02696_),
    .A_N(_02697_));
 sg13g2_nand2_1 _28165_ (.Y(_02699_),
    .A(net5849),
    .B(_02505_));
 sg13g2_nor2_1 _28166_ (.A(net5640),
    .B(_02681_),
    .Y(_02700_));
 sg13g2_xnor2_1 _28167_ (.Y(_02701_),
    .A(\u_inv.d_reg[162] ),
    .B(_02700_));
 sg13g2_nor4_1 _28168_ (.A(_02691_),
    .B(_02693_),
    .C(_02698_),
    .D(_02701_),
    .Y(_02702_));
 sg13g2_o21ai_1 _28169_ (.B1(net5853),
    .Y(_02703_),
    .A1(_02386_),
    .A2(_02504_));
 sg13g2_xnor2_1 _28170_ (.Y(_02704_),
    .A(_14662_),
    .B(_02703_));
 sg13g2_nand2_1 _28171_ (.Y(_02705_),
    .A(net5853),
    .B(_02504_));
 sg13g2_o21ai_1 _28172_ (.B1(net5853),
    .Y(_02706_),
    .A1(_02385_),
    .A2(_02504_));
 sg13g2_xnor2_1 _28173_ (.Y(_02707_),
    .A(_14663_),
    .B(_02706_));
 sg13g2_or2_1 _28174_ (.X(_02708_),
    .B(_02707_),
    .A(_02704_));
 sg13g2_nor3_1 _28175_ (.A(\u_inv.d_reg[147] ),
    .B(_02386_),
    .C(_02504_),
    .Y(_02709_));
 sg13g2_or3_1 _28176_ (.A(\u_inv.d_reg[147] ),
    .B(_02386_),
    .C(_02504_),
    .X(_02710_));
 sg13g2_nand2_1 _28177_ (.Y(_02711_),
    .A(net5855),
    .B(_02710_));
 sg13g2_xnor2_1 _28178_ (.Y(_02712_),
    .A(_14661_),
    .B(_02711_));
 sg13g2_inv_1 _28179_ (.Y(_02713_),
    .A(_02712_));
 sg13g2_nand2_1 _28180_ (.Y(_02714_),
    .A(net5848),
    .B(_02511_));
 sg13g2_o21ai_1 _28181_ (.B1(_02714_),
    .Y(_02715_),
    .A1(net5640),
    .A2(_02516_));
 sg13g2_xnor2_1 _28182_ (.Y(_02716_),
    .A(\u_inv.d_reg[179] ),
    .B(_02715_));
 sg13g2_o21ai_1 _28183_ (.B1(net5848),
    .Y(_02717_),
    .A1(_02511_),
    .A2(_02515_));
 sg13g2_xnor2_1 _28184_ (.Y(_02718_),
    .A(_14631_),
    .B(_02717_));
 sg13g2_nor4_1 _28185_ (.A(_02708_),
    .B(_02712_),
    .C(_02716_),
    .D(_02718_),
    .Y(_02719_));
 sg13g2_o21ai_1 _28186_ (.B1(net5849),
    .Y(_02720_),
    .A1(_02392_),
    .A2(_02710_));
 sg13g2_o21ai_1 _28187_ (.B1(_02720_),
    .Y(_02721_),
    .A1(net5641),
    .A2(_14655_));
 sg13g2_xnor2_1 _28188_ (.Y(_02722_),
    .A(\u_inv.d_reg[155] ),
    .B(_02721_));
 sg13g2_inv_1 _28189_ (.Y(_02723_),
    .A(_02722_));
 sg13g2_a21o_1 _28190_ (.A2(_02522_),
    .A1(_02521_),
    .B1(net5638),
    .X(_02724_));
 sg13g2_inv_1 _28191_ (.Y(_02725_),
    .A(_02724_));
 sg13g2_xnor2_1 _28192_ (.Y(_02726_),
    .A(\u_inv.d_reg[190] ),
    .B(_02724_));
 sg13g2_nand4_1 _28193_ (.B(_02719_),
    .C(_02723_),
    .A(_02702_),
    .Y(_02727_),
    .D(_02726_));
 sg13g2_nor4_2 _28194_ (.A(_02680_),
    .B(_02685_),
    .C(_02686_),
    .Y(_02728_),
    .D(_02727_));
 sg13g2_o21ai_1 _28195_ (.B1(net5843),
    .Y(_02729_),
    .A1(_02527_),
    .A2(_02532_));
 sg13g2_inv_1 _28196_ (.Y(_02730_),
    .A(_02729_));
 sg13g2_xnor2_1 _28197_ (.Y(_02731_),
    .A(_14603_),
    .B(_02729_));
 sg13g2_xnor2_1 _28198_ (.Y(_02732_),
    .A(_14614_),
    .B(_02637_));
 sg13g2_a21o_2 _28199_ (.A2(_02681_),
    .A1(_14647_),
    .B1(net5641),
    .X(_02733_));
 sg13g2_nand2_1 _28200_ (.Y(_02734_),
    .A(net5849),
    .B(\u_inv.d_reg[163] ));
 sg13g2_nand2_1 _28201_ (.Y(_02735_),
    .A(_02733_),
    .B(_02734_));
 sg13g2_xnor2_1 _28202_ (.Y(_02736_),
    .A(net5867),
    .B(_02735_));
 sg13g2_a21oi_1 _28203_ (.A1(net5849),
    .A2(net5867),
    .Y(_02737_),
    .B1(_02735_));
 sg13g2_xnor2_1 _28204_ (.Y(_02738_),
    .A(\u_inv.d_reg[165] ),
    .B(_02737_));
 sg13g2_nand2b_2 _28205_ (.Y(_02739_),
    .B(_02738_),
    .A_N(_02736_));
 sg13g2_o21ai_1 _28206_ (.B1(net5841),
    .Y(_02740_),
    .A1(_02527_),
    .A2(_02530_));
 sg13g2_xnor2_1 _28207_ (.Y(_02741_),
    .A(\u_inv.d_reg[204] ),
    .B(_02740_));
 sg13g2_nand2b_1 _28208_ (.Y(_02742_),
    .B(_02741_),
    .A_N(_02739_));
 sg13g2_o21ai_1 _28209_ (.B1(net5849),
    .Y(_02743_),
    .A1(\u_inv.d_reg[165] ),
    .A2(net5867));
 sg13g2_nand3_1 _28210_ (.B(_02734_),
    .C(_02743_),
    .A(_02733_),
    .Y(_02744_));
 sg13g2_a21o_1 _28211_ (.A2(\u_inv.d_reg[166] ),
    .A1(net5849),
    .B1(_02744_),
    .X(_02745_));
 sg13g2_xnor2_1 _28212_ (.Y(_02746_),
    .A(_14642_),
    .B(_02745_));
 sg13g2_nand2_1 _28213_ (.Y(_02747_),
    .A(net5848),
    .B(_02682_));
 sg13g2_o21ai_1 _28214_ (.B1(_02747_),
    .Y(_02748_),
    .A1(net5640),
    .A2(_02506_));
 sg13g2_o21ai_1 _28215_ (.B1(net5848),
    .Y(_02749_),
    .A1(_02510_),
    .A2(_02682_));
 sg13g2_xnor2_1 _28216_ (.Y(_02750_),
    .A(\u_inv.d_reg[175] ),
    .B(_02749_));
 sg13g2_o21ai_1 _28217_ (.B1(net5848),
    .Y(_02751_),
    .A1(\u_inv.d_reg[173] ),
    .A2(\u_inv.d_reg[172] ));
 sg13g2_nand2b_1 _28218_ (.Y(_02752_),
    .B(_02751_),
    .A_N(_02748_));
 sg13g2_xnor2_1 _28219_ (.Y(_02753_),
    .A(_14635_),
    .B(_02752_));
 sg13g2_a21oi_1 _28220_ (.A1(net5848),
    .A2(\u_inv.d_reg[172] ),
    .Y(_02754_),
    .B1(_02748_));
 sg13g2_xnor2_1 _28221_ (.Y(_02755_),
    .A(\u_inv.d_reg[173] ),
    .B(_02754_));
 sg13g2_nand4_1 _28222_ (.B(_02750_),
    .C(_02753_),
    .A(_02746_),
    .Y(_02756_),
    .D(_02755_));
 sg13g2_nor4_1 _28223_ (.A(_02731_),
    .B(_02732_),
    .C(_02742_),
    .D(_02756_),
    .Y(_02757_));
 sg13g2_nand4_1 _28224_ (.B(_02670_),
    .C(_02728_),
    .A(_02665_),
    .Y(_02758_),
    .D(_02757_));
 sg13g2_o21ai_1 _28225_ (.B1(net5835),
    .Y(_02759_),
    .A1(\u_inv.d_reg[219] ),
    .A2(_02613_));
 sg13g2_inv_1 _28226_ (.Y(_02760_),
    .A(_02759_));
 sg13g2_xnor2_1 _28227_ (.Y(_02761_),
    .A(_14589_),
    .B(_02759_));
 sg13g2_o21ai_1 _28228_ (.B1(net5835),
    .Y(_02762_),
    .A1(\u_inv.d_reg[224] ),
    .A2(_02542_));
 sg13g2_xnor2_1 _28229_ (.Y(_02763_),
    .A(\u_inv.d_reg[225] ),
    .B(_02762_));
 sg13g2_inv_1 _28230_ (.Y(_02764_),
    .A(_02763_));
 sg13g2_nor4_1 _28231_ (.A(_02649_),
    .B(_02758_),
    .C(_02761_),
    .D(_02764_),
    .Y(_02765_));
 sg13g2_o21ai_1 _28232_ (.B1(net5837),
    .Y(_02766_),
    .A1(_02537_),
    .A2(_02540_));
 sg13g2_xnor2_1 _28233_ (.Y(_02767_),
    .A(_14591_),
    .B(_02766_));
 sg13g2_o21ai_1 _28234_ (.B1(\u_inv.d_reg[211] ),
    .Y(_02768_),
    .A1(\u_inv.d_reg[210] ),
    .A2(_02642_));
 sg13g2_nand2b_1 _28235_ (.Y(_02769_),
    .B(_02768_),
    .A_N(_02606_));
 sg13g2_o21ai_1 _28236_ (.B1(_02769_),
    .Y(_02770_),
    .A1(net5836),
    .A2(_14598_));
 sg13g2_inv_1 _28237_ (.Y(_02771_),
    .A(_02770_));
 sg13g2_nand2_1 _28238_ (.Y(_02772_),
    .A(\u_inv.d_reg[219] ),
    .B(_02613_));
 sg13g2_a22oi_1 _28239_ (.Y(_02773_),
    .B1(_02760_),
    .B2(_02772_),
    .A2(\u_inv.d_reg[219] ),
    .A1(net5637));
 sg13g2_o21ai_1 _28240_ (.B1(net5837),
    .Y(_02774_),
    .A1(\u_inv.d_reg[216] ),
    .A2(_02537_));
 sg13g2_xnor2_1 _28241_ (.Y(_02775_),
    .A(_14592_),
    .B(_02774_));
 sg13g2_inv_1 _28242_ (.Y(_02776_),
    .A(_02775_));
 sg13g2_nor4_1 _28243_ (.A(_02767_),
    .B(_02771_),
    .C(_02773_),
    .D(_02775_),
    .Y(_02777_));
 sg13g2_nand2_1 _28244_ (.Y(_02778_),
    .A(net5841),
    .B(\u_inv.d_reg[195] ));
 sg13g2_and2_1 _28245_ (.A(_02637_),
    .B(_02778_),
    .X(_02779_));
 sg13g2_inv_1 _28246_ (.Y(_02780_),
    .A(_02779_));
 sg13g2_xnor2_1 _28247_ (.Y(_02781_),
    .A(\u_inv.d_reg[196] ),
    .B(_02779_));
 sg13g2_a21oi_1 _28248_ (.A1(net5842),
    .A2(\u_inv.d_reg[196] ),
    .Y(_02782_),
    .B1(_02780_));
 sg13g2_xnor2_1 _28249_ (.Y(_02783_),
    .A(\u_inv.d_reg[197] ),
    .B(_02782_));
 sg13g2_nor2_1 _28250_ (.A(net5641),
    .B(_02393_),
    .Y(_02784_));
 sg13g2_nor2_1 _28251_ (.A(_02721_),
    .B(_02784_),
    .Y(_02785_));
 sg13g2_xnor2_1 _28252_ (.Y(_02786_),
    .A(_14652_),
    .B(_02785_));
 sg13g2_a21o_2 _28253_ (.A2(_02709_),
    .A1(_02390_),
    .B1(net5641),
    .X(_02787_));
 sg13g2_o21ai_1 _28254_ (.B1(_02787_),
    .Y(_02788_),
    .A1(net5641),
    .A2(_02395_));
 sg13g2_xnor2_1 _28255_ (.Y(_02789_),
    .A(_14651_),
    .B(_02788_));
 sg13g2_xnor2_1 _28256_ (.Y(_02790_),
    .A(\u_inv.d_reg[158] ),
    .B(_02788_));
 sg13g2_a21oi_1 _28257_ (.A1(net5849),
    .A2(\u_inv.d_reg[155] ),
    .Y(_02791_),
    .B1(_02721_));
 sg13g2_xnor2_1 _28258_ (.Y(_02792_),
    .A(_14653_),
    .B(_02791_));
 sg13g2_nor3_2 _28259_ (.A(_02786_),
    .B(_02790_),
    .C(_02792_),
    .Y(_02793_));
 sg13g2_a21oi_1 _28260_ (.A1(net5840),
    .A2(\u_inv.d_reg[206] ),
    .Y(_02794_),
    .B1(_02730_));
 sg13g2_xnor2_1 _28261_ (.Y(_02795_),
    .A(\u_inv.d_reg[207] ),
    .B(_02794_));
 sg13g2_nand4_1 _28262_ (.B(_02783_),
    .C(_02793_),
    .A(_02781_),
    .Y(_02796_),
    .D(_02795_));
 sg13g2_xnor2_1 _28263_ (.Y(_02797_),
    .A(_14643_),
    .B(_02744_));
 sg13g2_xnor2_1 _28264_ (.Y(_02798_),
    .A(_14669_),
    .B(_02674_));
 sg13g2_xnor2_1 _28265_ (.Y(_02799_),
    .A(net5869),
    .B(_02674_));
 sg13g2_a21oi_1 _28266_ (.A1(net5848),
    .A2(\u_inv.d_reg[179] ),
    .Y(_02800_),
    .B1(_02715_));
 sg13g2_xnor2_1 _28267_ (.Y(_02801_),
    .A(\u_inv.d_reg[180] ),
    .B(_02800_));
 sg13g2_xnor2_1 _28268_ (.Y(_02802_),
    .A(\u_inv.d_reg[176] ),
    .B(_02714_));
 sg13g2_o21ai_1 _28269_ (.B1(net5850),
    .Y(_02803_),
    .A1(\u_inv.d_reg[176] ),
    .A2(_02511_));
 sg13g2_xnor2_1 _28270_ (.Y(_02804_),
    .A(\u_inv.d_reg[177] ),
    .B(_02803_));
 sg13g2_and4_1 _28271_ (.A(_02798_),
    .B(_02801_),
    .C(_02802_),
    .D(_02804_),
    .X(_02805_));
 sg13g2_xnor2_1 _28272_ (.Y(_02806_),
    .A(\u_inv.d_reg[172] ),
    .B(_02748_));
 sg13g2_a21oi_1 _28273_ (.A1(_14639_),
    .A2(_02683_),
    .Y(_02807_),
    .B1(net5640));
 sg13g2_xnor2_1 _28274_ (.Y(_02808_),
    .A(\u_inv.d_reg[171] ),
    .B(_02807_));
 sg13g2_nor2_1 _28275_ (.A(_02806_),
    .B(_02808_),
    .Y(_02809_));
 sg13g2_nand3_1 _28276_ (.B(_02805_),
    .C(_02809_),
    .A(_02797_),
    .Y(_02810_));
 sg13g2_o21ai_1 _28277_ (.B1(net5846),
    .Y(_02811_),
    .A1(net5866),
    .A2(_02519_));
 sg13g2_xnor2_1 _28278_ (.Y(_02812_),
    .A(_14624_),
    .B(_02811_));
 sg13g2_a21oi_1 _28279_ (.A1(net5850),
    .A2(_02512_),
    .Y(_02813_),
    .B1(_02715_));
 sg13g2_xnor2_1 _28280_ (.Y(_02814_),
    .A(\u_inv.d_reg[182] ),
    .B(_02813_));
 sg13g2_xnor2_1 _28281_ (.Y(_02815_),
    .A(_14627_),
    .B(_02813_));
 sg13g2_xnor2_1 _28282_ (.Y(_02816_),
    .A(_14655_),
    .B(_02720_));
 sg13g2_a21oi_1 _28283_ (.A1(net5850),
    .A2(_02514_),
    .Y(_02817_),
    .B1(_02715_));
 sg13g2_xnor2_1 _28284_ (.Y(_02818_),
    .A(_14626_),
    .B(_02817_));
 sg13g2_nor4_1 _28285_ (.A(_02812_),
    .B(_02815_),
    .C(_02816_),
    .D(_02818_),
    .Y(_02819_));
 sg13g2_o21ai_1 _28286_ (.B1(net5851),
    .Y(_02820_),
    .A1(_02498_),
    .A2(_02671_));
 sg13g2_xnor2_1 _28287_ (.Y(_02821_),
    .A(\u_inv.d_reg[134] ),
    .B(_02820_));
 sg13g2_xnor2_1 _28288_ (.Y(_02822_),
    .A(\u_inv.d_reg[136] ),
    .B(_02688_));
 sg13g2_o21ai_1 _28289_ (.B1(net5849),
    .Y(_02823_),
    .A1(net5868),
    .A2(_02505_));
 sg13g2_xnor2_1 _28290_ (.Y(_02824_),
    .A(\u_inv.d_reg[161] ),
    .B(_02823_));
 sg13g2_nand3_1 _28291_ (.B(_02822_),
    .C(_02824_),
    .A(_02821_),
    .Y(_02825_));
 sg13g2_a21oi_2 _28292_ (.B1(net5647),
    .Y(_02826_),
    .A2(_02491_),
    .A1(net1073));
 sg13g2_a21oi_1 _28293_ (.A1(net5857),
    .A2(_02493_),
    .Y(_02827_),
    .B1(_02826_));
 sg13g2_xnor2_1 _28294_ (.Y(_02828_),
    .A(_14679_),
    .B(_02827_));
 sg13g2_a21oi_1 _28295_ (.A1(net5857),
    .A2(_02494_),
    .Y(_02829_),
    .B1(_02826_));
 sg13g2_xnor2_1 _28296_ (.Y(_02830_),
    .A(_14678_),
    .B(_02829_));
 sg13g2_nor2_1 _28297_ (.A(_02828_),
    .B(_02830_),
    .Y(_02831_));
 sg13g2_o21ai_1 _28298_ (.B1(net5853),
    .Y(_02832_),
    .A1(\u_inv.d_reg[144] ),
    .A2(_02504_));
 sg13g2_xnor2_1 _28299_ (.Y(_02833_),
    .A(\u_inv.d_reg[145] ),
    .B(_02832_));
 sg13g2_nand2_1 _28300_ (.Y(_02834_),
    .A(_02831_),
    .B(_02833_));
 sg13g2_xnor2_1 _28301_ (.Y(_02835_),
    .A(\u_inv.d_reg[160] ),
    .B(_02699_));
 sg13g2_nor2_2 _28302_ (.A(net5647),
    .B(net1073),
    .Y(_02836_));
 sg13g2_a21oi_1 _28303_ (.A1(net5856),
    .A2(_02490_),
    .Y(_02837_),
    .B1(_02836_));
 sg13g2_xnor2_1 _28304_ (.Y(_02838_),
    .A(\u_inv.d_reg[125] ),
    .B(_02837_));
 sg13g2_o21ai_1 _28305_ (.B1(net5856),
    .Y(_02839_),
    .A1(\u_inv.d_reg[125] ),
    .A2(_02490_));
 sg13g2_nor2b_1 _28306_ (.A(_02836_),
    .B_N(_02839_),
    .Y(_02840_));
 sg13g2_xnor2_1 _28307_ (.Y(_02841_),
    .A(\u_inv.d_reg[126] ),
    .B(_02840_));
 sg13g2_xnor2_1 _28308_ (.Y(_02842_),
    .A(_14681_),
    .B(_02826_));
 sg13g2_nand4_1 _28309_ (.B(_02838_),
    .C(_02841_),
    .A(_02835_),
    .Y(_02843_),
    .D(_02842_));
 sg13g2_o21ai_1 _28310_ (.B1(_02840_),
    .Y(_02844_),
    .A1(net5647),
    .A2(_14683_));
 sg13g2_xnor2_1 _28311_ (.Y(_02845_),
    .A(_14682_),
    .B(_02844_));
 sg13g2_a21oi_1 _28312_ (.A1(net5857),
    .A2(\u_inv.d_reg[128] ),
    .Y(_02846_),
    .B1(_02826_));
 sg13g2_xnor2_1 _28313_ (.Y(_02847_),
    .A(\u_inv.d_reg[129] ),
    .B(_02846_));
 sg13g2_inv_2 _28314_ (.Y(_02848_),
    .A(_02847_));
 sg13g2_xnor2_1 _28315_ (.Y(_02849_),
    .A(_14665_),
    .B(_02705_));
 sg13g2_nor2_1 _28316_ (.A(_02848_),
    .B(_02849_),
    .Y(_02850_));
 sg13g2_a21oi_1 _28317_ (.A1(net1073),
    .A2(_02487_),
    .Y(_02851_),
    .B1(net5647));
 sg13g2_xnor2_1 _28318_ (.Y(_02852_),
    .A(\u_inv.d_reg[122] ),
    .B(_02851_));
 sg13g2_nand2_1 _28319_ (.Y(_02853_),
    .A(net5859),
    .B(_02484_));
 sg13g2_xnor2_1 _28320_ (.Y(_02854_),
    .A(_14691_),
    .B(_02853_));
 sg13g2_inv_1 _28321_ (.Y(_02855_),
    .A(_02854_));
 sg13g2_nand2_1 _28322_ (.Y(_02856_),
    .A(net5859),
    .B(_02480_));
 sg13g2_o21ai_1 _28323_ (.B1(net5859),
    .Y(_02857_),
    .A1(\u_inv.d_reg[112] ),
    .A2(_02480_));
 sg13g2_o21ai_1 _28324_ (.B1(net5859),
    .Y(_02858_),
    .A1(\u_inv.d_reg[114] ),
    .A2(\u_inv.d_reg[113] ));
 sg13g2_nand2_1 _28325_ (.Y(_02859_),
    .A(_02857_),
    .B(_02858_));
 sg13g2_xnor2_1 _28326_ (.Y(_02860_),
    .A(_14694_),
    .B(_02859_));
 sg13g2_o21ai_1 _28327_ (.B1(_02857_),
    .Y(_02861_),
    .A1(net5647),
    .A2(_14696_));
 sg13g2_xnor2_1 _28328_ (.Y(_02862_),
    .A(_14695_),
    .B(_02861_));
 sg13g2_nand2b_2 _28329_ (.Y(_02863_),
    .B(net5862),
    .A_N(_02478_));
 sg13g2_xnor2_1 _28330_ (.Y(_02864_),
    .A(_14701_),
    .B(_02863_));
 sg13g2_nand2_1 _28331_ (.Y(_02865_),
    .A(net5861),
    .B(_02469_));
 sg13g2_o21ai_1 _28332_ (.B1(_02865_),
    .Y(_02866_),
    .A1(net5645),
    .A2(_14713_));
 sg13g2_o21ai_1 _28333_ (.B1(net5860),
    .Y(_02867_),
    .A1(net5870),
    .A2(\u_inv.d_reg[97] ));
 sg13g2_nor2b_1 _28334_ (.A(_02866_),
    .B_N(_02867_),
    .Y(_02868_));
 sg13g2_xnor2_1 _28335_ (.Y(_02869_),
    .A(\u_inv.d_reg[99] ),
    .B(_02868_));
 sg13g2_nor2_1 _28336_ (.A(net5645),
    .B(_02473_),
    .Y(_02870_));
 sg13g2_xnor2_1 _28337_ (.Y(_02871_),
    .A(\u_inv.d_reg[102] ),
    .B(_02870_));
 sg13g2_inv_1 _28338_ (.Y(_02872_),
    .A(_02871_));
 sg13g2_a21oi_1 _28339_ (.A1(net5860),
    .A2(\u_inv.d_reg[97] ),
    .Y(_02873_),
    .B1(_02866_));
 sg13g2_xnor2_1 _28340_ (.Y(_02874_),
    .A(net5870),
    .B(_02873_));
 sg13g2_nand3_1 _28341_ (.B(_02872_),
    .C(_02874_),
    .A(_02869_),
    .Y(_02875_));
 sg13g2_a21o_1 _28342_ (.A2(_02467_),
    .A1(_02465_),
    .B1(net5643),
    .X(_02876_));
 sg13g2_xnor2_1 _28343_ (.Y(_02877_),
    .A(\u_inv.d_reg[92] ),
    .B(_02876_));
 sg13g2_o21ai_1 _28344_ (.B1(_02876_),
    .Y(_02878_),
    .A1(net5644),
    .A2(_14717_));
 sg13g2_xnor2_1 _28345_ (.Y(_02879_),
    .A(_14716_),
    .B(_02878_));
 sg13g2_a21oi_1 _28346_ (.A1(net5861),
    .A2(\u_inv.d_reg[93] ),
    .Y(_02880_),
    .B1(_02878_));
 sg13g2_xnor2_1 _28347_ (.Y(_02881_),
    .A(_14715_),
    .B(_02880_));
 sg13g2_xnor2_1 _28348_ (.Y(_02882_),
    .A(\u_inv.d_reg[94] ),
    .B(_02880_));
 sg13g2_nand3_1 _28349_ (.B(_02879_),
    .C(_02882_),
    .A(_02877_),
    .Y(_02883_));
 sg13g2_o21ai_1 _28350_ (.B1(net5861),
    .Y(_02884_),
    .A1(\u_inv.d_reg[94] ),
    .A2(\u_inv.d_reg[93] ));
 sg13g2_nor2b_1 _28351_ (.A(_02878_),
    .B_N(_02884_),
    .Y(_02885_));
 sg13g2_xnor2_1 _28352_ (.Y(_02886_),
    .A(_14714_),
    .B(_02885_));
 sg13g2_xnor2_1 _28353_ (.Y(_02887_),
    .A(\u_inv.d_reg[97] ),
    .B(_02866_));
 sg13g2_inv_1 _28354_ (.Y(_02888_),
    .A(_02887_));
 sg13g2_or2_1 _28355_ (.X(_02889_),
    .B(_02887_),
    .A(_02886_));
 sg13g2_nor2_1 _28356_ (.A(net5644),
    .B(_02465_),
    .Y(_02890_));
 sg13g2_a21oi_1 _28357_ (.A1(net5861),
    .A2(_02466_),
    .Y(_02891_),
    .B1(_02890_));
 sg13g2_o21ai_1 _28358_ (.B1(_02891_),
    .Y(_02892_),
    .A1(net5645),
    .A2(_14719_));
 sg13g2_xnor2_1 _28359_ (.Y(_02893_),
    .A(_14718_),
    .B(_02892_));
 sg13g2_a21oi_1 _28360_ (.A1(_14721_),
    .A2(_02465_),
    .Y(_02894_),
    .B1(net5644));
 sg13g2_xnor2_1 _28361_ (.Y(_02895_),
    .A(_14720_),
    .B(_02894_));
 sg13g2_xnor2_1 _28362_ (.Y(_02896_),
    .A(\u_inv.d_reg[88] ),
    .B(_02890_));
 sg13g2_nor2b_1 _28363_ (.A(_02896_),
    .B_N(_02895_),
    .Y(_02897_));
 sg13g2_xnor2_1 _28364_ (.Y(_02898_),
    .A(_14713_),
    .B(_02865_));
 sg13g2_inv_1 _28365_ (.Y(_02899_),
    .A(_02898_));
 sg13g2_a21o_1 _28366_ (.A2(_02463_),
    .A1(_02458_),
    .B1(net5643),
    .X(_02900_));
 sg13g2_o21ai_1 _28367_ (.B1(_02900_),
    .Y(_02901_),
    .A1(net5643),
    .A2(_14723_));
 sg13g2_xnor2_1 _28368_ (.Y(_02902_),
    .A(\u_inv.d_reg[87] ),
    .B(_02901_));
 sg13g2_nor2_1 _28369_ (.A(net5643),
    .B(_02458_),
    .Y(_02903_));
 sg13g2_a21oi_1 _28370_ (.A1(_02458_),
    .A2(_02460_),
    .Y(_02904_),
    .B1(net5643));
 sg13g2_xnor2_1 _28371_ (.Y(_02905_),
    .A(\u_inv.d_reg[83] ),
    .B(_02904_));
 sg13g2_a21oi_1 _28372_ (.A1(_02458_),
    .A2(_02459_),
    .Y(_02906_),
    .B1(net5643));
 sg13g2_xnor2_1 _28373_ (.Y(_02907_),
    .A(\u_inv.d_reg[82] ),
    .B(_02906_));
 sg13g2_nor3_1 _28374_ (.A(_02902_),
    .B(_02905_),
    .C(_02907_),
    .Y(_02908_));
 sg13g2_xnor2_1 _28375_ (.Y(_02909_),
    .A(net5871),
    .B(_02891_));
 sg13g2_a21oi_1 _28376_ (.A1(net5861),
    .A2(_02462_),
    .Y(_02910_),
    .B1(_02903_));
 sg13g2_xnor2_1 _28377_ (.Y(_02911_),
    .A(\u_inv.d_reg[85] ),
    .B(_02910_));
 sg13g2_a21oi_1 _28378_ (.A1(_02458_),
    .A2(_02461_),
    .Y(_02912_),
    .B1(net5643));
 sg13g2_xnor2_1 _28379_ (.Y(_02913_),
    .A(_14725_),
    .B(_02912_));
 sg13g2_nand2_1 _28380_ (.Y(_02914_),
    .A(_02911_),
    .B(_02913_));
 sg13g2_nand4_1 _28381_ (.B(_02909_),
    .C(_02911_),
    .A(_02908_),
    .Y(_02915_),
    .D(_02913_));
 sg13g2_o21ai_1 _28382_ (.B1(net5860),
    .Y(_02916_),
    .A1(_02454_),
    .A2(_02456_));
 sg13g2_o21ai_1 _28383_ (.B1(_02916_),
    .Y(_02917_),
    .A1(net5646),
    .A2(_14733_));
 sg13g2_a21oi_1 _28384_ (.A1(net5860),
    .A2(net5872),
    .Y(_02918_),
    .B1(_02917_));
 sg13g2_xnor2_1 _28385_ (.Y(_02919_),
    .A(\u_inv.d_reg[78] ),
    .B(_02918_));
 sg13g2_nand2_1 _28386_ (.Y(_02920_),
    .A(net5860),
    .B(_02454_));
 sg13g2_o21ai_1 _28387_ (.B1(net5860),
    .Y(_02921_),
    .A1(_02454_),
    .A2(_02455_));
 sg13g2_xnor2_1 _28388_ (.Y(_02922_),
    .A(_14735_),
    .B(_02921_));
 sg13g2_xnor2_1 _28389_ (.Y(_02923_),
    .A(\u_inv.d_reg[74] ),
    .B(_02921_));
 sg13g2_xnor2_1 _28390_ (.Y(_02924_),
    .A(_14733_),
    .B(_02916_));
 sg13g2_and2_1 _28391_ (.A(net5856),
    .B(_02447_),
    .X(_02925_));
 sg13g2_o21ai_1 _28392_ (.B1(net5858),
    .Y(_02926_),
    .A1(_02447_),
    .A2(_02448_));
 sg13g2_xnor2_1 _28393_ (.Y(_02927_),
    .A(_14743_),
    .B(_02926_));
 sg13g2_o21ai_1 _28394_ (.B1(net5856),
    .Y(_02928_),
    .A1(\u_inv.d_reg[64] ),
    .A2(_02447_));
 sg13g2_xnor2_1 _28395_ (.Y(_02929_),
    .A(_14744_),
    .B(_02928_));
 sg13g2_nand2_1 _28396_ (.Y(_02930_),
    .A(net5856),
    .B(_02445_));
 sg13g2_xnor2_1 _28397_ (.Y(_02931_),
    .A(_14747_),
    .B(_02930_));
 sg13g2_nor2_1 _28398_ (.A(net5642),
    .B(_02441_),
    .Y(_02932_));
 sg13g2_a21oi_1 _28399_ (.A1(_14751_),
    .A2(_02441_),
    .Y(_02933_),
    .B1(net5642));
 sg13g2_xnor2_1 _28400_ (.Y(_02934_),
    .A(\u_inv.d_reg[59] ),
    .B(_02933_));
 sg13g2_nand2_1 _28401_ (.Y(_02935_),
    .A(net5851),
    .B(_02440_));
 sg13g2_o21ai_1 _28402_ (.B1(net5851),
    .Y(_02936_),
    .A1(\u_inv.d_reg[56] ),
    .A2(_02440_));
 sg13g2_xnor2_1 _28403_ (.Y(_02937_),
    .A(_14752_),
    .B(_02936_));
 sg13g2_xnor2_1 _28404_ (.Y(_02938_),
    .A(_14753_),
    .B(_02935_));
 sg13g2_nor2_1 _28405_ (.A(_02937_),
    .B(_02938_),
    .Y(_02939_));
 sg13g2_xnor2_1 _28406_ (.Y(_02940_),
    .A(_14751_),
    .B(_02932_));
 sg13g2_inv_1 _28407_ (.Y(_02941_),
    .A(_02940_));
 sg13g2_o21ai_1 _28408_ (.B1(net5851),
    .Y(_02942_),
    .A1(\u_inv.d_reg[54] ),
    .A2(_02438_));
 sg13g2_xnor2_1 _28409_ (.Y(_02943_),
    .A(_14754_),
    .B(_02942_));
 sg13g2_inv_2 _28410_ (.Y(_02944_),
    .A(_02943_));
 sg13g2_nand2_1 _28411_ (.Y(_02945_),
    .A(net5851),
    .B(_02438_));
 sg13g2_xnor2_1 _28412_ (.Y(_02946_),
    .A(_14755_),
    .B(_02945_));
 sg13g2_o21ai_1 _28413_ (.B1(net5851),
    .Y(_02947_),
    .A1(\u_inv.d_reg[52] ),
    .A2(_02436_));
 sg13g2_xnor2_1 _28414_ (.Y(_02948_),
    .A(_14756_),
    .B(_02947_));
 sg13g2_nand2_1 _28415_ (.Y(_02949_),
    .A(net5851),
    .B(_02436_));
 sg13g2_xnor2_1 _28416_ (.Y(_02950_),
    .A(\u_inv.d_reg[52] ),
    .B(_02949_));
 sg13g2_xnor2_1 _28417_ (.Y(_02951_),
    .A(_14757_),
    .B(_02949_));
 sg13g2_o21ai_1 _28418_ (.B1(net5852),
    .Y(_02952_),
    .A1(\u_inv.d_reg[50] ),
    .A2(_02434_));
 sg13g2_xnor2_1 _28419_ (.Y(_02953_),
    .A(\u_inv.d_reg[51] ),
    .B(_02952_));
 sg13g2_nand2_1 _28420_ (.Y(_02954_),
    .A(net5852),
    .B(_02434_));
 sg13g2_xnor2_1 _28421_ (.Y(_02955_),
    .A(_14759_),
    .B(_02954_));
 sg13g2_nand2_1 _28422_ (.Y(_02956_),
    .A(net5852),
    .B(_02433_));
 sg13g2_o21ai_1 _28423_ (.B1(net5852),
    .Y(_02957_),
    .A1(\u_inv.d_reg[48] ),
    .A2(_02433_));
 sg13g2_xnor2_1 _28424_ (.Y(_02958_),
    .A(\u_inv.d_reg[49] ),
    .B(_02957_));
 sg13g2_xnor2_1 _28425_ (.Y(_02959_),
    .A(_14760_),
    .B(_02957_));
 sg13g2_nor2_1 _28426_ (.A(_02955_),
    .B(_02959_),
    .Y(_02960_));
 sg13g2_xnor2_1 _28427_ (.Y(_02961_),
    .A(\u_inv.d_reg[48] ),
    .B(_02956_));
 sg13g2_nand2_1 _28428_ (.Y(_02962_),
    .A(net5846),
    .B(_02430_));
 sg13g2_o21ai_1 _28429_ (.B1(net5846),
    .Y(_02963_),
    .A1(\u_inv.d_reg[44] ),
    .A2(_02430_));
 sg13g2_xnor2_1 _28430_ (.Y(_02964_),
    .A(_14764_),
    .B(_02963_));
 sg13g2_nor2_1 _28431_ (.A(net5640),
    .B(_02431_),
    .Y(_02965_));
 sg13g2_xnor2_1 _28432_ (.Y(_02966_),
    .A(\u_inv.d_reg[46] ),
    .B(_02965_));
 sg13g2_nand3b_1 _28433_ (.B(_14775_),
    .C(_14774_),
    .Y(_02967_),
    .A_N(_02421_));
 sg13g2_nand2_1 _28434_ (.Y(_02968_),
    .A(net5844),
    .B(_02967_));
 sg13g2_o21ai_1 _28435_ (.B1(net5844),
    .Y(_02969_),
    .A1(_02424_),
    .A2(_02967_));
 sg13g2_xnor2_1 _28436_ (.Y(_02970_),
    .A(_14770_),
    .B(_02969_));
 sg13g2_nand2_1 _28437_ (.Y(_02971_),
    .A(net5844),
    .B(_02419_));
 sg13g2_xnor2_1 _28438_ (.Y(_02972_),
    .A(_14777_),
    .B(_02971_));
 sg13g2_inv_1 _28439_ (.Y(_02973_),
    .A(_02972_));
 sg13g2_a21oi_1 _28440_ (.A1(_14781_),
    .A2(_02416_),
    .Y(_02974_),
    .B1(net5638));
 sg13g2_xnor2_1 _28441_ (.Y(_02975_),
    .A(_14780_),
    .B(_02974_));
 sg13g2_nor2_1 _28442_ (.A(net5638),
    .B(_02416_),
    .Y(_02976_));
 sg13g2_xnor2_1 _28443_ (.Y(_02977_),
    .A(_14781_),
    .B(_02976_));
 sg13g2_nor2_1 _28444_ (.A(net5637),
    .B(_02407_),
    .Y(_02978_));
 sg13g2_xnor2_1 _28445_ (.Y(_02979_),
    .A(_14794_),
    .B(_02978_));
 sg13g2_o21ai_1 _28446_ (.B1(net5834),
    .Y(_02980_),
    .A1(\u_inv.d_reg[13] ),
    .A2(_02406_));
 sg13g2_xnor2_1 _28447_ (.Y(_02981_),
    .A(_14795_),
    .B(_02980_));
 sg13g2_nor2_1 _28448_ (.A(net5637),
    .B(_02403_),
    .Y(_02982_));
 sg13g2_xnor2_1 _28449_ (.Y(_02983_),
    .A(_14800_),
    .B(_02982_));
 sg13g2_o21ai_1 _28450_ (.B1(net5834),
    .Y(_02984_),
    .A1(\u_inv.d_reg[7] ),
    .A2(_02402_));
 sg13g2_xnor2_1 _28451_ (.Y(_02985_),
    .A(\u_inv.d_reg[8] ),
    .B(_02984_));
 sg13g2_nor2_1 _28452_ (.A(net5636),
    .B(_02398_),
    .Y(_02986_));
 sg13g2_xnor2_1 _28453_ (.Y(_02987_),
    .A(\u_inv.d_reg[3] ),
    .B(_02986_));
 sg13g2_nand2_1 _28454_ (.Y(_02988_),
    .A(net5832),
    .B(\u_inv.d_reg[0] ));
 sg13g2_xnor2_1 _28455_ (.Y(_02989_),
    .A(_14808_),
    .B(_02988_));
 sg13g2_nor2_1 _28456_ (.A(_14552_),
    .B(_02989_),
    .Y(_02990_));
 sg13g2_nand2_1 _28457_ (.Y(_02991_),
    .A(net5832),
    .B(_02397_));
 sg13g2_xnor2_1 _28458_ (.Y(_02992_),
    .A(\u_inv.d_reg[2] ),
    .B(_02991_));
 sg13g2_nand2_1 _28459_ (.Y(_02993_),
    .A(_02990_),
    .B(_02992_));
 sg13g2_or2_1 _28460_ (.X(_02994_),
    .B(_02993_),
    .A(_02987_));
 sg13g2_nand2_1 _28461_ (.Y(_02995_),
    .A(net5832),
    .B(_02399_));
 sg13g2_xnor2_1 _28462_ (.Y(_02996_),
    .A(_14805_),
    .B(_02995_));
 sg13g2_inv_1 _28463_ (.Y(_02997_),
    .A(_02996_));
 sg13g2_o21ai_1 _28464_ (.B1(net5832),
    .Y(_02998_),
    .A1(\u_inv.d_reg[4] ),
    .A2(_02399_));
 sg13g2_xnor2_1 _28465_ (.Y(_02999_),
    .A(_14804_),
    .B(_02998_));
 sg13g2_a21oi_1 _28466_ (.A1(_02994_),
    .A2(_02996_),
    .Y(_03000_),
    .B1(_02999_));
 sg13g2_o21ai_1 _28467_ (.B1(net5833),
    .Y(_03001_),
    .A1(\u_inv.d_reg[5] ),
    .A2(_02401_));
 sg13g2_xnor2_1 _28468_ (.Y(_03002_),
    .A(\u_inv.d_reg[6] ),
    .B(_03001_));
 sg13g2_nor2_1 _28469_ (.A(_03000_),
    .B(_03002_),
    .Y(_03003_));
 sg13g2_nand2_1 _28470_ (.Y(_03004_),
    .A(net5834),
    .B(_02402_));
 sg13g2_xnor2_1 _28471_ (.Y(_03005_),
    .A(\u_inv.d_reg[7] ),
    .B(_03004_));
 sg13g2_xnor2_1 _28472_ (.Y(_03006_),
    .A(_14802_),
    .B(_03004_));
 sg13g2_nand2_1 _28473_ (.Y(_03007_),
    .A(_03003_),
    .B(_03006_));
 sg13g2_nor3_1 _28474_ (.A(_02983_),
    .B(_02985_),
    .C(_03007_),
    .Y(_03008_));
 sg13g2_nand2_1 _28475_ (.Y(_03009_),
    .A(net5834),
    .B(_02406_));
 sg13g2_xnor2_1 _28476_ (.Y(_03010_),
    .A(_14796_),
    .B(_03009_));
 sg13g2_o21ai_1 _28477_ (.B1(net5834),
    .Y(_03011_),
    .A1(net5874),
    .A2(_02405_));
 sg13g2_xnor2_1 _28478_ (.Y(_03012_),
    .A(_14797_),
    .B(_03011_));
 sg13g2_nand3_1 _28479_ (.B(net5874),
    .C(_02405_),
    .A(net5834),
    .Y(_03013_));
 sg13g2_a21o_1 _28480_ (.A2(_02405_),
    .A1(net5834),
    .B1(net5874),
    .X(_03014_));
 sg13g2_nand2_1 _28481_ (.Y(_03015_),
    .A(_03013_),
    .B(_03014_));
 sg13g2_nand2_1 _28482_ (.Y(_03016_),
    .A(net5834),
    .B(_02404_));
 sg13g2_xnor2_1 _28483_ (.Y(_03017_),
    .A(\u_inv.d_reg[10] ),
    .B(_03016_));
 sg13g2_nand3_1 _28484_ (.B(_03014_),
    .C(_03017_),
    .A(_03013_),
    .Y(_03018_));
 sg13g2_nor3_1 _28485_ (.A(_03010_),
    .B(_03012_),
    .C(_03018_),
    .Y(_03019_));
 sg13g2_nand2_1 _28486_ (.Y(_03020_),
    .A(_02979_),
    .B(_03019_));
 sg13g2_or3_1 _28487_ (.A(_02981_),
    .B(_03008_),
    .C(_03020_),
    .X(_03021_));
 sg13g2_inv_2 _28488_ (.Y(_03022_),
    .A(_03021_));
 sg13g2_nand2b_1 _28489_ (.Y(_03023_),
    .B(net5840),
    .A_N(_02415_));
 sg13g2_xnor2_1 _28490_ (.Y(_03024_),
    .A(\u_inv.d_reg[27] ),
    .B(_03023_));
 sg13g2_xnor2_1 _28491_ (.Y(_03025_),
    .A(_14782_),
    .B(_03023_));
 sg13g2_nand2_1 _28492_ (.Y(_03026_),
    .A(net5840),
    .B(_02414_));
 sg13g2_xnor2_1 _28493_ (.Y(_03027_),
    .A(_14784_),
    .B(_03026_));
 sg13g2_o21ai_1 _28494_ (.B1(net5840),
    .Y(_03028_),
    .A1(\u_inv.d_reg[22] ),
    .A2(_02412_));
 sg13g2_xnor2_1 _28495_ (.Y(_03029_),
    .A(\u_inv.d_reg[23] ),
    .B(_03028_));
 sg13g2_nand2b_1 _28496_ (.Y(_03030_),
    .B(net5840),
    .A_N(_02411_));
 sg13g2_xnor2_1 _28497_ (.Y(_03031_),
    .A(\u_inv.d_reg[21] ),
    .B(_03030_));
 sg13g2_xnor2_1 _28498_ (.Y(_03032_),
    .A(_14788_),
    .B(_03030_));
 sg13g2_nand2_1 _28499_ (.Y(_03033_),
    .A(net5836),
    .B(_02410_));
 sg13g2_xnor2_1 _28500_ (.Y(_03034_),
    .A(_14790_),
    .B(_03033_));
 sg13g2_o21ai_1 _28501_ (.B1(net5836),
    .Y(_03035_),
    .A1(net5873),
    .A2(_02408_));
 sg13g2_xnor2_1 _28502_ (.Y(_03036_),
    .A(\u_inv.d_reg[17] ),
    .B(_03035_));
 sg13g2_xnor2_1 _28503_ (.Y(_03037_),
    .A(_14792_),
    .B(_03035_));
 sg13g2_nand2_1 _28504_ (.Y(_03038_),
    .A(net5836),
    .B(_02408_));
 sg13g2_xnor2_1 _28505_ (.Y(_03039_),
    .A(net5873),
    .B(_03038_));
 sg13g2_xnor2_1 _28506_ (.Y(_03040_),
    .A(_14793_),
    .B(_03038_));
 sg13g2_nor2_1 _28507_ (.A(_03037_),
    .B(_03040_),
    .Y(_03041_));
 sg13g2_nor2_1 _28508_ (.A(net5637),
    .B(_02409_),
    .Y(_03042_));
 sg13g2_xnor2_1 _28509_ (.Y(_03043_),
    .A(\u_inv.d_reg[18] ),
    .B(_03042_));
 sg13g2_or4_1 _28510_ (.A(_03034_),
    .B(_03037_),
    .C(_03040_),
    .D(_03043_),
    .X(_03044_));
 sg13g2_o21ai_1 _28511_ (.B1(net5836),
    .Y(_03045_),
    .A1(\u_inv.d_reg[19] ),
    .A2(_02410_));
 sg13g2_xnor2_1 _28512_ (.Y(_03046_),
    .A(_14789_),
    .B(_03045_));
 sg13g2_nor3_1 _28513_ (.A(_03032_),
    .B(_03044_),
    .C(_03046_),
    .Y(_03047_));
 sg13g2_nand2_1 _28514_ (.Y(_03048_),
    .A(net5840),
    .B(_02412_));
 sg13g2_xnor2_1 _28515_ (.Y(_03049_),
    .A(\u_inv.d_reg[22] ),
    .B(_03048_));
 sg13g2_xnor2_1 _28516_ (.Y(_03050_),
    .A(_14787_),
    .B(_03048_));
 sg13g2_nand3_1 _28517_ (.B(_03047_),
    .C(_03049_),
    .A(_03029_),
    .Y(_03051_));
 sg13g2_inv_1 _28518_ (.Y(_03052_),
    .A(_03051_));
 sg13g2_nor2_1 _28519_ (.A(net5638),
    .B(_02413_),
    .Y(_03053_));
 sg13g2_xnor2_1 _28520_ (.Y(_03054_),
    .A(\u_inv.d_reg[24] ),
    .B(_03053_));
 sg13g2_or2_1 _28521_ (.X(_03055_),
    .B(_03054_),
    .A(_03027_));
 sg13g2_nor2_1 _28522_ (.A(_03051_),
    .B(_03055_),
    .Y(_03056_));
 sg13g2_o21ai_1 _28523_ (.B1(net5840),
    .Y(_03057_),
    .A1(\u_inv.d_reg[25] ),
    .A2(_02414_));
 sg13g2_xnor2_1 _28524_ (.Y(_03058_),
    .A(_14783_),
    .B(_03057_));
 sg13g2_nor4_1 _28525_ (.A(_03025_),
    .B(_03051_),
    .C(_03055_),
    .D(_03058_),
    .Y(_03059_));
 sg13g2_nand4_1 _28526_ (.B(_02977_),
    .C(_03022_),
    .A(_02975_),
    .Y(_03060_),
    .D(_03059_));
 sg13g2_o21ai_1 _28527_ (.B1(net5842),
    .Y(_03061_),
    .A1(\u_inv.d_reg[30] ),
    .A2(_02418_));
 sg13g2_xnor2_1 _28528_ (.Y(_03062_),
    .A(_14778_),
    .B(_03061_));
 sg13g2_nand2_1 _28529_ (.Y(_03063_),
    .A(net5842),
    .B(_02418_));
 sg13g2_xnor2_1 _28530_ (.Y(_03064_),
    .A(_14779_),
    .B(_03063_));
 sg13g2_nor3_1 _28531_ (.A(_03060_),
    .B(_03062_),
    .C(_03064_),
    .Y(_03065_));
 sg13g2_nand2b_1 _28532_ (.Y(_03066_),
    .B(_02972_),
    .A_N(_03065_));
 sg13g2_o21ai_1 _28533_ (.B1(net5844),
    .Y(_03067_),
    .A1(\u_inv.d_reg[32] ),
    .A2(_02419_));
 sg13g2_xnor2_1 _28534_ (.Y(_03068_),
    .A(\u_inv.d_reg[33] ),
    .B(_03067_));
 sg13g2_nand3_1 _28535_ (.B(\u_inv.d_reg[34] ),
    .C(_02421_),
    .A(net5844),
    .Y(_03069_));
 sg13g2_a21o_1 _28536_ (.A2(_02421_),
    .A1(net5845),
    .B1(\u_inv.d_reg[34] ),
    .X(_03070_));
 sg13g2_nand2_2 _28537_ (.Y(_03071_),
    .A(_03069_),
    .B(_03070_));
 sg13g2_inv_1 _28538_ (.Y(_03072_),
    .A(_03071_));
 sg13g2_o21ai_1 _28539_ (.B1(net5844),
    .Y(_03073_),
    .A1(\u_inv.d_reg[34] ),
    .A2(_02421_));
 sg13g2_xnor2_1 _28540_ (.Y(_03074_),
    .A(_14774_),
    .B(_03073_));
 sg13g2_o21ai_1 _28541_ (.B1(net5846),
    .Y(_03075_),
    .A1(_02419_),
    .A2(_02426_));
 sg13g2_xnor2_1 _28542_ (.Y(_03076_),
    .A(_14769_),
    .B(_03075_));
 sg13g2_nor2_1 _28543_ (.A(_03074_),
    .B(_03076_),
    .Y(_03077_));
 sg13g2_nand4_1 _28544_ (.B(_03068_),
    .C(_03072_),
    .A(_03066_),
    .Y(_03078_),
    .D(_03077_));
 sg13g2_o21ai_1 _28545_ (.B1(net5844),
    .Y(_03079_),
    .A1(_02422_),
    .A2(_02967_));
 sg13g2_xnor2_1 _28546_ (.Y(_03080_),
    .A(_14771_),
    .B(_03079_));
 sg13g2_o21ai_1 _28547_ (.B1(net5846),
    .Y(_03081_),
    .A1(\u_inv.d_reg[42] ),
    .A2(_02427_));
 sg13g2_xnor2_1 _28548_ (.Y(_03082_),
    .A(_14766_),
    .B(_03081_));
 sg13g2_inv_1 _28549_ (.Y(_03083_),
    .A(_03082_));
 sg13g2_nor4_2 _28550_ (.A(_02970_),
    .B(_03078_),
    .C(_03080_),
    .Y(_03084_),
    .D(_03082_));
 sg13g2_nand2b_1 _28551_ (.Y(_03085_),
    .B(_03084_),
    .A_N(_02966_));
 sg13g2_a21oi_1 _28552_ (.A1(_14763_),
    .A2(_02431_),
    .Y(_03086_),
    .B1(net5640));
 sg13g2_xnor2_1 _28553_ (.Y(_03087_),
    .A(\u_inv.d_reg[47] ),
    .B(_03086_));
 sg13g2_inv_1 _28554_ (.Y(_03088_),
    .A(_03087_));
 sg13g2_xnor2_1 _28555_ (.Y(_03089_),
    .A(_14765_),
    .B(_02962_));
 sg13g2_o21ai_1 _28556_ (.B1(net5844),
    .Y(_03090_),
    .A1(\u_inv.d_reg[36] ),
    .A2(_02967_));
 sg13g2_xnor2_1 _28557_ (.Y(_03091_),
    .A(_14772_),
    .B(_03090_));
 sg13g2_o21ai_1 _28558_ (.B1(_03075_),
    .Y(_03092_),
    .A1(net5638),
    .A2(_14769_));
 sg13g2_xnor2_1 _28559_ (.Y(_03093_),
    .A(_14768_),
    .B(_03092_));
 sg13g2_xnor2_1 _28560_ (.Y(_03094_),
    .A(_14773_),
    .B(_02968_));
 sg13g2_nand2_1 _28561_ (.Y(_03095_),
    .A(net5846),
    .B(_02427_));
 sg13g2_xnor2_1 _28562_ (.Y(_03096_),
    .A(\u_inv.d_reg[42] ),
    .B(_03095_));
 sg13g2_xnor2_1 _28563_ (.Y(_03097_),
    .A(_14767_),
    .B(_03095_));
 sg13g2_nand2_1 _28564_ (.Y(_03098_),
    .A(_03093_),
    .B(_03096_));
 sg13g2_or4_1 _28565_ (.A(_03089_),
    .B(_03091_),
    .C(_03094_),
    .D(_03098_),
    .X(_03099_));
 sg13g2_nor4_2 _28566_ (.A(_02964_),
    .B(_03085_),
    .C(_03087_),
    .Y(_03100_),
    .D(_03099_));
 sg13g2_nand4_1 _28567_ (.B(_02960_),
    .C(_02961_),
    .A(_02953_),
    .Y(_03101_),
    .D(_03100_));
 sg13g2_nor4_1 _28568_ (.A(_02946_),
    .B(_02948_),
    .C(_02951_),
    .D(_03101_),
    .Y(_03102_));
 sg13g2_nand4_1 _28569_ (.B(_02940_),
    .C(_02944_),
    .A(_02939_),
    .Y(_03103_),
    .D(_03102_));
 sg13g2_or4_1 _28570_ (.A(_02929_),
    .B(_02931_),
    .C(_02934_),
    .D(_03103_),
    .X(_03104_));
 sg13g2_nand2_1 _28571_ (.Y(_03105_),
    .A(net5858),
    .B(_02452_));
 sg13g2_xnor2_1 _28572_ (.Y(_03106_),
    .A(_14739_),
    .B(_03105_));
 sg13g2_inv_2 _28573_ (.Y(_03107_),
    .A(_03106_));
 sg13g2_xnor2_1 _28574_ (.Y(_03108_),
    .A(\u_inv.d_reg[64] ),
    .B(_02925_));
 sg13g2_nand2_1 _28575_ (.Y(_03109_),
    .A(net5856),
    .B(_02443_));
 sg13g2_o21ai_1 _28576_ (.B1(net5856),
    .Y(_03110_),
    .A1(\u_inv.d_reg[60] ),
    .A2(_02443_));
 sg13g2_xnor2_1 _28577_ (.Y(_03111_),
    .A(_14748_),
    .B(_03110_));
 sg13g2_xnor2_1 _28578_ (.Y(_03112_),
    .A(_14749_),
    .B(_03109_));
 sg13g2_or2_1 _28579_ (.X(_03113_),
    .B(_03112_),
    .A(_03111_));
 sg13g2_o21ai_1 _28580_ (.B1(net5856),
    .Y(_03114_),
    .A1(\u_inv.d_reg[62] ),
    .A2(_02445_));
 sg13g2_xnor2_1 _28581_ (.Y(_03115_),
    .A(\u_inv.d_reg[63] ),
    .B(_03114_));
 sg13g2_nor2_1 _28582_ (.A(_03108_),
    .B(_03113_),
    .Y(_03116_));
 sg13g2_nand3_1 _28583_ (.B(_03115_),
    .C(_03116_),
    .A(_03107_),
    .Y(_03117_));
 sg13g2_nor4_2 _28584_ (.A(_02924_),
    .B(_02927_),
    .C(_03104_),
    .Y(_03118_),
    .D(_03117_));
 sg13g2_o21ai_1 _28585_ (.B1(net5860),
    .Y(_03119_),
    .A1(\u_inv.d_reg[78] ),
    .A2(\u_inv.d_reg[77] ));
 sg13g2_nor2b_1 _28586_ (.A(_02917_),
    .B_N(_03119_),
    .Y(_03120_));
 sg13g2_xnor2_1 _28587_ (.Y(_03121_),
    .A(\u_inv.d_reg[79] ),
    .B(_03120_));
 sg13g2_xnor2_1 _28588_ (.Y(_03122_),
    .A(_14723_),
    .B(_02900_));
 sg13g2_nor2b_1 _28589_ (.A(_03122_),
    .B_N(_03121_),
    .Y(_03123_));
 sg13g2_nand4_1 _28590_ (.B(_02923_),
    .C(_03118_),
    .A(_02919_),
    .Y(_03124_),
    .D(_03123_));
 sg13g2_a21oi_1 _28591_ (.A1(_14729_),
    .A2(_02458_),
    .Y(_03125_),
    .B1(net5643));
 sg13g2_xnor2_1 _28592_ (.Y(_03126_),
    .A(\u_inv.d_reg[81] ),
    .B(_03125_));
 sg13g2_xnor2_1 _28593_ (.Y(_03127_),
    .A(\u_inv.d_reg[80] ),
    .B(_02903_));
 sg13g2_or2_1 _28594_ (.X(_03128_),
    .B(_03127_),
    .A(_03126_));
 sg13g2_o21ai_1 _28595_ (.B1(_02921_),
    .Y(_03129_),
    .A1(net5646),
    .A2(_14735_));
 sg13g2_xnor2_1 _28596_ (.Y(_03130_),
    .A(_14734_),
    .B(_03129_));
 sg13g2_a21o_1 _28597_ (.A2(_02926_),
    .A1(_14743_),
    .B1(net5647),
    .X(_03131_));
 sg13g2_xnor2_1 _28598_ (.Y(_03132_),
    .A(_14742_),
    .B(_03131_));
 sg13g2_o21ai_1 _28599_ (.B1(net5858),
    .Y(_03133_),
    .A1(\u_inv.d_reg[70] ),
    .A2(_02452_));
 sg13g2_xnor2_1 _28600_ (.Y(_03134_),
    .A(\u_inv.d_reg[71] ),
    .B(_03133_));
 sg13g2_nand2_1 _28601_ (.Y(_03135_),
    .A(net5858),
    .B(_02450_));
 sg13g2_o21ai_1 _28602_ (.B1(net5858),
    .Y(_03136_),
    .A1(\u_inv.d_reg[68] ),
    .A2(_02450_));
 sg13g2_xnor2_1 _28603_ (.Y(_03137_),
    .A(_14740_),
    .B(_03136_));
 sg13g2_inv_1 _28604_ (.Y(_03138_),
    .A(_03137_));
 sg13g2_xnor2_1 _28605_ (.Y(_03139_),
    .A(_14741_),
    .B(_03135_));
 sg13g2_nor2_1 _28606_ (.A(_03137_),
    .B(_03139_),
    .Y(_03140_));
 sg13g2_nor2b_1 _28607_ (.A(_03132_),
    .B_N(_03134_),
    .Y(_03141_));
 sg13g2_xnor2_1 _28608_ (.Y(_03142_),
    .A(net5872),
    .B(_02917_));
 sg13g2_o21ai_1 _28609_ (.B1(net5860),
    .Y(_03143_),
    .A1(\u_inv.d_reg[72] ),
    .A2(_02454_));
 sg13g2_xnor2_1 _28610_ (.Y(_03144_),
    .A(\u_inv.d_reg[73] ),
    .B(_03143_));
 sg13g2_inv_1 _28611_ (.Y(_03145_),
    .A(_03144_));
 sg13g2_xnor2_1 _28612_ (.Y(_03146_),
    .A(\u_inv.d_reg[72] ),
    .B(_02920_));
 sg13g2_nand2_1 _28613_ (.Y(_03147_),
    .A(_03144_),
    .B(_03146_));
 sg13g2_nor2_1 _28614_ (.A(_03142_),
    .B(_03147_),
    .Y(_03148_));
 sg13g2_nand4_1 _28615_ (.B(_03140_),
    .C(_03141_),
    .A(_03130_),
    .Y(_03149_),
    .D(_03148_));
 sg13g2_nor4_1 _28616_ (.A(_02915_),
    .B(_03124_),
    .C(_03128_),
    .D(_03149_),
    .Y(_03150_));
 sg13g2_nand4_1 _28617_ (.B(_02897_),
    .C(_02899_),
    .A(_02893_),
    .Y(_03151_),
    .D(_03150_));
 sg13g2_nor4_1 _28618_ (.A(_02875_),
    .B(_02883_),
    .C(_02889_),
    .D(_03151_),
    .Y(_03152_));
 sg13g2_nand2_1 _28619_ (.Y(_03153_),
    .A(net5862),
    .B(_02475_));
 sg13g2_o21ai_1 _28620_ (.B1(net5862),
    .Y(_03154_),
    .A1(\u_inv.d_reg[104] ),
    .A2(_02475_));
 sg13g2_xnor2_1 _28621_ (.Y(_03155_),
    .A(\u_inv.d_reg[105] ),
    .B(_03154_));
 sg13g2_inv_1 _28622_ (.Y(_03156_),
    .A(_03155_));
 sg13g2_nand2b_1 _28623_ (.Y(_03157_),
    .B(net5862),
    .A_N(_02477_));
 sg13g2_xnor2_1 _28624_ (.Y(_03158_),
    .A(\u_inv.d_reg[106] ),
    .B(_03157_));
 sg13g2_xnor2_1 _28625_ (.Y(_03159_),
    .A(_14703_),
    .B(_03157_));
 sg13g2_a21oi_1 _28626_ (.A1(_14703_),
    .A2(_02477_),
    .Y(_03160_),
    .B1(net5646));
 sg13g2_xnor2_1 _28627_ (.Y(_03161_),
    .A(\u_inv.d_reg[107] ),
    .B(_03160_));
 sg13g2_xnor2_1 _28628_ (.Y(_03162_),
    .A(_14705_),
    .B(_03153_));
 sg13g2_a21oi_1 _28629_ (.A1(_14707_),
    .A2(_02473_),
    .Y(_03163_),
    .B1(net5645));
 sg13g2_xnor2_1 _28630_ (.Y(_03164_),
    .A(\u_inv.d_reg[103] ),
    .B(_03163_));
 sg13g2_nand2_1 _28631_ (.Y(_03165_),
    .A(net5863),
    .B(_02471_));
 sg13g2_o21ai_1 _28632_ (.B1(net5862),
    .Y(_03166_),
    .A1(\u_inv.d_reg[100] ),
    .A2(_02471_));
 sg13g2_xnor2_1 _28633_ (.Y(_03167_),
    .A(\u_inv.d_reg[101] ),
    .B(_03166_));
 sg13g2_xnor2_1 _28634_ (.Y(_03168_),
    .A(\u_inv.d_reg[100] ),
    .B(_03165_));
 sg13g2_nand2_1 _28635_ (.Y(_03169_),
    .A(_03167_),
    .B(_03168_));
 sg13g2_nor4_1 _28636_ (.A(_03161_),
    .B(_03162_),
    .C(_03164_),
    .D(_03169_),
    .Y(_03170_));
 sg13g2_nand4_1 _28637_ (.B(_03155_),
    .C(_03158_),
    .A(_03152_),
    .Y(_03171_),
    .D(_03170_));
 sg13g2_nand2_1 _28638_ (.Y(_03172_),
    .A(net5862),
    .B(\u_inv.d_reg[108] ));
 sg13g2_nand2_1 _28639_ (.Y(_03173_),
    .A(_02863_),
    .B(_03172_));
 sg13g2_xnor2_1 _28640_ (.Y(_03174_),
    .A(\u_inv.d_reg[109] ),
    .B(_03173_));
 sg13g2_xnor2_1 _28641_ (.Y(_03175_),
    .A(_14697_),
    .B(_02856_));
 sg13g2_nor4_1 _28642_ (.A(_02864_),
    .B(_03171_),
    .C(_03174_),
    .D(_03175_),
    .Y(_03176_));
 sg13g2_nand4_1 _28643_ (.B(_02860_),
    .C(_02862_),
    .A(_02855_),
    .Y(_03177_),
    .D(_03176_));
 sg13g2_a21oi_1 _28644_ (.A1(net5857),
    .A2(_02489_),
    .Y(_03178_),
    .B1(_02836_));
 sg13g2_xnor2_1 _28645_ (.Y(_03179_),
    .A(_14685_),
    .B(_03178_));
 sg13g2_xnor2_1 _28646_ (.Y(_03180_),
    .A(\u_inv.d_reg[124] ),
    .B(_03178_));
 sg13g2_a21oi_1 _28647_ (.A1(net1073),
    .A2(_02488_),
    .Y(_03181_),
    .B1(net5647));
 sg13g2_xnor2_1 _28648_ (.Y(_03182_),
    .A(\u_inv.d_reg[123] ),
    .B(_03181_));
 sg13g2_nor4_1 _28649_ (.A(_02852_),
    .B(_03177_),
    .C(_03179_),
    .D(_03182_),
    .Y(_03183_));
 sg13g2_a21oi_1 _28650_ (.A1(_14689_),
    .A2(net1073),
    .Y(_03184_),
    .B1(net5647));
 sg13g2_xnor2_1 _28651_ (.Y(_03185_),
    .A(\u_inv.d_reg[121] ),
    .B(_03184_));
 sg13g2_xnor2_1 _28652_ (.Y(_03186_),
    .A(\u_inv.d_reg[120] ),
    .B(_02836_));
 sg13g2_or2_1 _28653_ (.X(_03187_),
    .B(_03186_),
    .A(_03185_));
 sg13g2_nand2_1 _28654_ (.Y(_03188_),
    .A(net5859),
    .B(_02482_));
 sg13g2_o21ai_1 _28655_ (.B1(net5859),
    .Y(_03189_),
    .A1(\u_inv.d_reg[116] ),
    .A2(_02482_));
 sg13g2_xnor2_1 _28656_ (.Y(_03190_),
    .A(\u_inv.d_reg[117] ),
    .B(_03189_));
 sg13g2_xnor2_1 _28657_ (.Y(_03191_),
    .A(\u_inv.d_reg[116] ),
    .B(_03188_));
 sg13g2_nand2_1 _28658_ (.Y(_03192_),
    .A(_03190_),
    .B(_03191_));
 sg13g2_o21ai_1 _28659_ (.B1(net5859),
    .Y(_03193_),
    .A1(\u_inv.d_reg[118] ),
    .A2(_02484_));
 sg13g2_xnor2_1 _28660_ (.Y(_03194_),
    .A(\u_inv.d_reg[119] ),
    .B(_03193_));
 sg13g2_a21oi_1 _28661_ (.A1(net5862),
    .A2(\u_inv.d_reg[109] ),
    .Y(_03195_),
    .B1(_03173_));
 sg13g2_xnor2_1 _28662_ (.Y(_03196_),
    .A(\u_inv.d_reg[110] ),
    .B(_03195_));
 sg13g2_o21ai_1 _28663_ (.B1(net5862),
    .Y(_03197_),
    .A1(\u_inv.d_reg[110] ),
    .A2(\u_inv.d_reg[109] ));
 sg13g2_nand3_1 _28664_ (.B(_03172_),
    .C(_03197_),
    .A(_02863_),
    .Y(_03198_));
 sg13g2_xnor2_1 _28665_ (.Y(_03199_),
    .A(\u_inv.d_reg[111] ),
    .B(_03198_));
 sg13g2_xnor2_1 _28666_ (.Y(_03200_),
    .A(_14696_),
    .B(_02857_));
 sg13g2_inv_1 _28667_ (.Y(_03201_),
    .A(_03200_));
 sg13g2_nor2_1 _28668_ (.A(_03199_),
    .B(_03200_),
    .Y(_03202_));
 sg13g2_nand3_1 _28669_ (.B(_03196_),
    .C(_03202_),
    .A(_03194_),
    .Y(_03203_));
 sg13g2_nor3_1 _28670_ (.A(_03187_),
    .B(_03192_),
    .C(_03203_),
    .Y(_03204_));
 sg13g2_nand4_1 _28671_ (.B(_02850_),
    .C(_03183_),
    .A(_02845_),
    .Y(_03205_),
    .D(_03204_));
 sg13g2_nor4_2 _28672_ (.A(_02825_),
    .B(_02834_),
    .C(_02843_),
    .Y(_03206_),
    .D(_03205_));
 sg13g2_a21o_1 _28673_ (.A2(_02820_),
    .A1(_14675_),
    .B1(net5642),
    .X(_03207_));
 sg13g2_xnor2_1 _28674_ (.Y(_03208_),
    .A(_14674_),
    .B(_03207_));
 sg13g2_a21oi_1 _28675_ (.A1(_02518_),
    .A2(_02520_),
    .Y(_03209_),
    .B1(net5639));
 sg13g2_xnor2_1 _28676_ (.Y(_03210_),
    .A(\u_inv.d_reg[186] ),
    .B(_03209_));
 sg13g2_inv_1 _28677_ (.Y(_03211_),
    .A(_03210_));
 sg13g2_nor2_1 _28678_ (.A(_03208_),
    .B(_03210_),
    .Y(_03212_));
 sg13g2_a21oi_1 _28679_ (.A1(_02389_),
    .A2(_02709_),
    .Y(_03213_),
    .B1(net5641));
 sg13g2_xnor2_1 _28680_ (.Y(_03214_),
    .A(_14658_),
    .B(_03213_));
 sg13g2_o21ai_1 _28681_ (.B1(net5855),
    .Y(_03215_),
    .A1(\u_inv.d_reg[148] ),
    .A2(_02710_));
 sg13g2_xnor2_1 _28682_ (.Y(_03216_),
    .A(\u_inv.d_reg[149] ),
    .B(_03215_));
 sg13g2_xnor2_1 _28683_ (.Y(_03217_),
    .A(\u_inv.d_reg[152] ),
    .B(_02787_));
 sg13g2_xnor2_1 _28684_ (.Y(_03218_),
    .A(_14622_),
    .B(_02650_));
 sg13g2_nand4_1 _28685_ (.B(_03216_),
    .C(_03217_),
    .A(_03214_),
    .Y(_03219_),
    .D(_03218_));
 sg13g2_a21oi_1 _28686_ (.A1(_02388_),
    .A2(_02709_),
    .Y(_03220_),
    .B1(net5642));
 sg13g2_xnor2_1 _28687_ (.Y(_03221_),
    .A(\u_inv.d_reg[150] ),
    .B(_03220_));
 sg13g2_o21ai_1 _28688_ (.B1(_02787_),
    .Y(_03222_),
    .A1(net5641),
    .A2(_14657_));
 sg13g2_xnor2_1 _28689_ (.Y(_03223_),
    .A(_14656_),
    .B(_03222_));
 sg13g2_nand2b_1 _28690_ (.Y(_03224_),
    .B(_03223_),
    .A_N(_03221_));
 sg13g2_o21ai_1 _28691_ (.B1(net5854),
    .Y(_03225_),
    .A1(_02497_),
    .A2(_02672_));
 sg13g2_xnor2_1 _28692_ (.Y(_03226_),
    .A(\u_inv.d_reg[139] ),
    .B(_03225_));
 sg13g2_o21ai_1 _28693_ (.B1(net5854),
    .Y(_03227_),
    .A1(_02496_),
    .A2(_02672_));
 sg13g2_xnor2_1 _28694_ (.Y(_03228_),
    .A(\u_inv.d_reg[138] ),
    .B(_03227_));
 sg13g2_nand2_2 _28695_ (.Y(_03229_),
    .A(_03226_),
    .B(_03228_));
 sg13g2_xnor2_1 _28696_ (.Y(_03230_),
    .A(_14646_),
    .B(_02733_));
 sg13g2_nor4_2 _28697_ (.A(_03219_),
    .B(_03224_),
    .C(_03229_),
    .Y(_03231_),
    .D(_03230_));
 sg13g2_nand4_1 _28698_ (.B(_03206_),
    .C(_03212_),
    .A(_02819_),
    .Y(_03232_),
    .D(_03231_));
 sg13g2_a21oi_1 _28699_ (.A1(net5847),
    .A2(\u_inv.d_reg[190] ),
    .Y(_03233_),
    .B1(_02725_));
 sg13g2_xnor2_1 _28700_ (.Y(_03234_),
    .A(_14618_),
    .B(_03233_));
 sg13g2_o21ai_1 _28701_ (.B1(net5850),
    .Y(_03235_),
    .A1(\u_inv.d_reg[158] ),
    .A2(_02788_));
 sg13g2_xnor2_1 _28702_ (.Y(_03236_),
    .A(\u_inv.d_reg[159] ),
    .B(_03235_));
 sg13g2_a21oi_1 _28703_ (.A1(_14629_),
    .A2(_02800_),
    .Y(_03237_),
    .B1(net5640));
 sg13g2_xnor2_1 _28704_ (.Y(_03238_),
    .A(_14628_),
    .B(_03237_));
 sg13g2_and2_1 _28705_ (.A(_03236_),
    .B(_03238_),
    .X(_03239_));
 sg13g2_o21ai_1 _28706_ (.B1(net5853),
    .Y(_03240_),
    .A1(net5869),
    .A2(_02674_));
 sg13g2_xnor2_1 _28707_ (.Y(_03241_),
    .A(_14668_),
    .B(_03240_));
 sg13g2_xnor2_1 _28708_ (.Y(_03242_),
    .A(\u_inv.d_reg[141] ),
    .B(_03240_));
 sg13g2_o21ai_1 _28709_ (.B1(net5848),
    .Y(_03243_),
    .A1(\u_inv.d_reg[168] ),
    .A2(_02682_));
 sg13g2_xnor2_1 _28710_ (.Y(_03244_),
    .A(\u_inv.d_reg[169] ),
    .B(_03243_));
 sg13g2_xnor2_1 _28711_ (.Y(_03245_),
    .A(\u_inv.d_reg[168] ),
    .B(_02747_));
 sg13g2_nand3_1 _28712_ (.B(_03244_),
    .C(_03245_),
    .A(_03242_),
    .Y(_03246_));
 sg13g2_xnor2_1 _28713_ (.Y(_03247_),
    .A(\u_inv.d_reg[200] ),
    .B(_02656_));
 sg13g2_xnor2_1 _28714_ (.Y(_03248_),
    .A(_14616_),
    .B(_02660_));
 sg13g2_nor3_1 _28715_ (.A(_03246_),
    .B(_03247_),
    .C(_03248_),
    .Y(_03249_));
 sg13g2_nand3b_1 _28716_ (.B(_03239_),
    .C(_03249_),
    .Y(_03250_),
    .A_N(_03234_));
 sg13g2_nor4_2 _28717_ (.A(_02796_),
    .B(_02810_),
    .C(_03232_),
    .Y(_03251_),
    .D(_03250_));
 sg13g2_xnor2_1 _28718_ (.Y(_03252_),
    .A(\u_inv.d_reg[224] ),
    .B(_02600_));
 sg13g2_a21oi_1 _28719_ (.A1(net5843),
    .A2(\u_inv.d_reg[208] ),
    .Y(_03253_),
    .B1(_02605_));
 sg13g2_xnor2_1 _28720_ (.Y(_03254_),
    .A(_14600_),
    .B(_03253_));
 sg13g2_xnor2_1 _28721_ (.Y(_03255_),
    .A(_14595_),
    .B(_02645_));
 sg13g2_o21ai_1 _28722_ (.B1(net5843),
    .Y(_03256_),
    .A1(_02527_),
    .A2(_02531_));
 sg13g2_xnor2_1 _28723_ (.Y(_03257_),
    .A(net3438),
    .B(_03256_));
 sg13g2_xnor2_1 _28724_ (.Y(_03258_),
    .A(\u_inv.d_reg[198] ),
    .B(_02638_));
 sg13g2_nand2_2 _28725_ (.Y(_03259_),
    .A(_03257_),
    .B(_03258_));
 sg13g2_nor4_1 _28726_ (.A(_03252_),
    .B(_03254_),
    .C(_03255_),
    .D(_03259_),
    .Y(_03260_));
 sg13g2_nand4_1 _28727_ (.B(_02777_),
    .C(_03251_),
    .A(_02765_),
    .Y(_03261_),
    .D(_03260_));
 sg13g2_xnor2_1 _28728_ (.Y(_03262_),
    .A(_14565_),
    .B(_02569_));
 sg13g2_a21oi_1 _28729_ (.A1(net5835),
    .A2(\u_inv.d_reg[220] ),
    .Y(_03263_),
    .B1(_02760_));
 sg13g2_xnor2_1 _28730_ (.Y(_03264_),
    .A(\u_inv.d_reg[221] ),
    .B(_03263_));
 sg13g2_nand2_1 _28731_ (.Y(_03265_),
    .A(net5832),
    .B(\u_inv.d_reg[228] ));
 sg13g2_and2_1 _28732_ (.A(_02621_),
    .B(_03265_),
    .X(_03266_));
 sg13g2_xnor2_1 _28733_ (.Y(_03267_),
    .A(\u_inv.d_reg[229] ),
    .B(_03266_));
 sg13g2_o21ai_1 _28734_ (.B1(net5831),
    .Y(_03268_),
    .A1(\u_inv.d_reg[232] ),
    .A2(_02545_));
 sg13g2_xnor2_1 _28735_ (.Y(_03269_),
    .A(\u_inv.d_reg[233] ),
    .B(_03268_));
 sg13g2_nand4_1 _28736_ (.B(_03264_),
    .C(_03267_),
    .A(_03262_),
    .Y(_03270_),
    .D(_03269_));
 sg13g2_nor4_1 _28737_ (.A(_02625_),
    .B(_02632_),
    .C(_03261_),
    .D(_03270_),
    .Y(_03271_));
 sg13g2_o21ai_1 _28738_ (.B1(net5830),
    .Y(_03272_),
    .A1(\u_inv.d_reg[244] ),
    .A2(_02551_));
 sg13g2_xnor2_1 _28739_ (.Y(_03273_),
    .A(\u_inv.d_reg[245] ),
    .B(_03272_));
 sg13g2_xnor2_1 _28740_ (.Y(_03274_),
    .A(net3442),
    .B(_02592_));
 sg13g2_o21ai_1 _28741_ (.B1(net5833),
    .Y(_03275_),
    .A1(\u_inv.d_reg[236] ),
    .A2(_02547_));
 sg13g2_xnor2_1 _28742_ (.Y(_03276_),
    .A(_14572_),
    .B(_03275_));
 sg13g2_nand2_1 _28743_ (.Y(_03277_),
    .A(net5831),
    .B(_02579_));
 sg13g2_xnor2_1 _28744_ (.Y(_03278_),
    .A(_14575_),
    .B(_03277_));
 sg13g2_nor2_1 _28745_ (.A(_03276_),
    .B(_03278_),
    .Y(_03279_));
 sg13g2_nand4_1 _28746_ (.B(_03273_),
    .C(_03274_),
    .A(_03271_),
    .Y(_03280_),
    .D(_03279_));
 sg13g2_or3_1 _28747_ (.A(_02590_),
    .B(_02598_),
    .C(_03280_),
    .X(_03281_));
 sg13g2_o21ai_1 _28748_ (.B1(_02561_),
    .Y(_03282_),
    .A1(net5635),
    .A2(_14556_));
 sg13g2_xnor2_1 _28749_ (.Y(_03283_),
    .A(_14555_),
    .B(_03282_));
 sg13g2_o21ai_1 _28750_ (.B1(net5831),
    .Y(_03284_),
    .A1(_02553_),
    .A2(_02555_));
 sg13g2_a21oi_1 _28751_ (.A1(_14559_),
    .A2(_02565_),
    .Y(_03285_),
    .B1(_14558_));
 sg13g2_nand2_1 _28752_ (.Y(_03286_),
    .A(net5635),
    .B(\u_inv.d_reg[251] ));
 sg13g2_o21ai_1 _28753_ (.B1(_03286_),
    .Y(_03287_),
    .A1(_03284_),
    .A2(_03285_));
 sg13g2_xnor2_1 _28754_ (.Y(_03288_),
    .A(\u_inv.d_reg[253] ),
    .B(_02561_));
 sg13g2_inv_1 _28755_ (.Y(_03289_),
    .A(_03288_));
 sg13g2_xnor2_1 _28756_ (.Y(_03290_),
    .A(_14557_),
    .B(_03284_));
 sg13g2_nor2_1 _28757_ (.A(_03289_),
    .B(_03290_),
    .Y(_03291_));
 sg13g2_o21ai_1 _28758_ (.B1(net5830),
    .Y(_03292_),
    .A1(\u_inv.d_reg[248] ),
    .A2(_02553_));
 sg13g2_xnor2_1 _28759_ (.Y(_03293_),
    .A(\u_inv.d_reg[249] ),
    .B(_03292_));
 sg13g2_and2_1 _28760_ (.A(net4483),
    .B(_03293_),
    .X(_03294_));
 sg13g2_nand4_1 _28761_ (.B(_03287_),
    .C(_03291_),
    .A(_03283_),
    .Y(_03295_),
    .D(_03294_));
 sg13g2_nor4_2 _28762_ (.A(_02564_),
    .B(_02567_),
    .C(_03295_),
    .Y(_03296_),
    .D(_03281_));
 sg13g2_inv_2 _28763_ (.Y(_03297_),
    .A(net4472));
 sg13g2_and2_1 _28764_ (.A(_02741_),
    .B(_03257_),
    .X(_03298_));
 sg13g2_nand2_1 _28765_ (.Y(_03299_),
    .A(_03262_),
    .B(_03273_));
 sg13g2_nand2_1 _28766_ (.Y(_03300_),
    .A(_02622_),
    .B(_03267_));
 sg13g2_nor2_2 _28767_ (.A(net4502),
    .B(net4473),
    .Y(_03301_));
 sg13g2_nand2_2 _28768_ (.Y(_03302_),
    .A(net4485),
    .B(net4470));
 sg13g2_xnor2_1 _28769_ (.Y(_03303_),
    .A(_14552_),
    .B(net4454));
 sg13g2_nand2_1 _28770_ (.Y(_03304_),
    .A(net1249),
    .B(net5107));
 sg13g2_o21ai_1 _28771_ (.B1(_03304_),
    .Y(_00518_),
    .A1(net5108),
    .A2(_03303_));
 sg13g2_a21oi_1 _28772_ (.A1(_14552_),
    .A2(_14808_),
    .Y(_03305_),
    .B1(_02990_));
 sg13g2_o21ai_1 _28773_ (.B1(net5232),
    .Y(_03306_),
    .A1(net4485),
    .A2(_03305_));
 sg13g2_a21oi_1 _28774_ (.A1(net4472),
    .A2(_03305_),
    .Y(_03307_),
    .B1(_03306_));
 sg13g2_o21ai_1 _28775_ (.B1(_03307_),
    .Y(_03308_),
    .A1(_02989_),
    .A2(net4374));
 sg13g2_o21ai_1 _28776_ (.B1(_03308_),
    .Y(_03309_),
    .A1(net2750),
    .A2(net5239));
 sg13g2_inv_1 _28777_ (.Y(_00519_),
    .A(_03309_));
 sg13g2_a21oi_1 _28778_ (.A1(_02990_),
    .A2(net4472),
    .Y(_03310_),
    .B1(_02992_));
 sg13g2_nor2_1 _28779_ (.A(_02993_),
    .B(net4470),
    .Y(_03311_));
 sg13g2_o21ai_1 _28780_ (.B1(net4486),
    .Y(_03312_),
    .A1(_03310_),
    .A2(_03311_));
 sg13g2_a21oi_1 _28781_ (.A1(_02397_),
    .A2(_02992_),
    .Y(_03313_),
    .B1(_02398_));
 sg13g2_a21oi_1 _28782_ (.A1(net4501),
    .A2(_03313_),
    .Y(_03314_),
    .B1(net5108));
 sg13g2_a22oi_1 _28783_ (.Y(_03315_),
    .B1(_03312_),
    .B2(_03314_),
    .A2(net5108),
    .A1(net2602));
 sg13g2_inv_1 _28784_ (.Y(_00520_),
    .A(_03315_));
 sg13g2_xnor2_1 _28785_ (.Y(_03316_),
    .A(_02987_),
    .B(_03311_));
 sg13g2_nand2_1 _28786_ (.Y(_03317_),
    .A(net4486),
    .B(_03316_));
 sg13g2_o21ai_1 _28787_ (.B1(_02399_),
    .Y(_03318_),
    .A1(_02398_),
    .A2(_02987_));
 sg13g2_a21oi_1 _28788_ (.A1(net4501),
    .A2(_03318_),
    .Y(_03319_),
    .B1(net5108));
 sg13g2_a22oi_1 _28789_ (.Y(_00521_),
    .B1(_03317_),
    .B2(_03319_),
    .A2(net5117),
    .A1(_14514_));
 sg13g2_nand2_1 _28790_ (.Y(_03320_),
    .A(_02994_),
    .B(net4472));
 sg13g2_a21oi_1 _28791_ (.A1(_02996_),
    .A2(_03320_),
    .Y(_03321_),
    .B1(net4505));
 sg13g2_o21ai_1 _28792_ (.B1(_03321_),
    .Y(_03322_),
    .A1(_02996_),
    .A2(_03320_));
 sg13g2_a21oi_1 _28793_ (.A1(_02399_),
    .A2(_02997_),
    .Y(_03323_),
    .B1(net4486));
 sg13g2_a21oi_1 _28794_ (.A1(_02401_),
    .A2(_03323_),
    .Y(_03324_),
    .B1(net5108));
 sg13g2_nand2_1 _28795_ (.Y(_03325_),
    .A(_03322_),
    .B(_03324_));
 sg13g2_o21ai_1 _28796_ (.B1(_03325_),
    .Y(_03326_),
    .A1(net2505),
    .A2(net5232));
 sg13g2_inv_1 _28797_ (.Y(_00522_),
    .A(_03326_));
 sg13g2_nor2_1 _28798_ (.A(net1325),
    .B(net5232),
    .Y(_03327_));
 sg13g2_a21oi_1 _28799_ (.A1(_02994_),
    .A2(_02996_),
    .Y(_03328_),
    .B1(net4501));
 sg13g2_o21ai_1 _28800_ (.B1(net4375),
    .Y(_03329_),
    .A1(_03323_),
    .A2(_03328_));
 sg13g2_xnor2_1 _28801_ (.Y(_03330_),
    .A(_02999_),
    .B(_03329_));
 sg13g2_a21oi_1 _28802_ (.A1(net5239),
    .A2(_03330_),
    .Y(_00523_),
    .B1(_03327_));
 sg13g2_nor2_1 _28803_ (.A(net1206),
    .B(net5241),
    .Y(_03331_));
 sg13g2_o21ai_1 _28804_ (.B1(_02999_),
    .Y(_03332_),
    .A1(_02400_),
    .A2(_02996_));
 sg13g2_a221oi_1 _28805_ (.B2(_02999_),
    .C1(net4455),
    .B1(_03323_),
    .A1(net4486),
    .Y(_03333_),
    .A2(_03000_));
 sg13g2_xnor2_1 _28806_ (.Y(_03334_),
    .A(_03002_),
    .B(_03333_));
 sg13g2_a21oi_1 _28807_ (.A1(net5232),
    .A2(_03334_),
    .Y(_00524_),
    .B1(_03331_));
 sg13g2_nand2_1 _28808_ (.Y(_03335_),
    .A(_03002_),
    .B(_03332_));
 sg13g2_nor2_1 _28809_ (.A(net4486),
    .B(_03335_),
    .Y(_03336_));
 sg13g2_a21oi_1 _28810_ (.A1(_03003_),
    .A2(net4473),
    .Y(_03337_),
    .B1(_03336_));
 sg13g2_xnor2_1 _28811_ (.Y(_03338_),
    .A(_03006_),
    .B(_03337_));
 sg13g2_nand2_1 _28812_ (.Y(_03339_),
    .A(net1111),
    .B(net5108));
 sg13g2_o21ai_1 _28813_ (.B1(_03339_),
    .Y(_00525_),
    .A1(net5108),
    .A2(_03338_));
 sg13g2_nor2_1 _28814_ (.A(net1257),
    .B(net5240),
    .Y(_03340_));
 sg13g2_nor2_1 _28815_ (.A(_03006_),
    .B(_03335_),
    .Y(_03341_));
 sg13g2_nand2_1 _28816_ (.Y(_03342_),
    .A(net4501),
    .B(_03341_));
 sg13g2_nand2b_1 _28817_ (.Y(_03343_),
    .B(net4473),
    .A_N(_03007_));
 sg13g2_nand2_1 _28818_ (.Y(_03344_),
    .A(_03342_),
    .B(_03343_));
 sg13g2_xnor2_1 _28819_ (.Y(_03345_),
    .A(_02985_),
    .B(_03344_));
 sg13g2_a21oi_1 _28820_ (.A1(net5240),
    .A2(_03345_),
    .Y(_00526_),
    .B1(_03340_));
 sg13g2_nor2_1 _28821_ (.A(net1264),
    .B(net5241),
    .Y(_03346_));
 sg13g2_and4_1 _28822_ (.A(_02985_),
    .B(_03002_),
    .C(_03005_),
    .D(_03332_),
    .X(_03347_));
 sg13g2_nand2_1 _28823_ (.Y(_03348_),
    .A(_02985_),
    .B(_03341_));
 sg13g2_a22oi_1 _28824_ (.Y(_03349_),
    .B1(_03343_),
    .B2(_03348_),
    .A2(_02985_),
    .A1(net4486));
 sg13g2_xnor2_1 _28825_ (.Y(_03350_),
    .A(_02983_),
    .B(_03349_));
 sg13g2_a21oi_1 _28826_ (.A1(net5241),
    .A2(_03350_),
    .Y(_00527_),
    .B1(_03346_));
 sg13g2_a21o_1 _28827_ (.A2(_03347_),
    .A1(_02983_),
    .B1(net4487),
    .X(_03351_));
 sg13g2_nand2b_2 _28828_ (.Y(_03352_),
    .B(net4473),
    .A_N(_03008_));
 sg13g2_inv_1 _28829_ (.Y(_03353_),
    .A(_03352_));
 sg13g2_nand2_1 _28830_ (.Y(_03354_),
    .A(_03351_),
    .B(_03352_));
 sg13g2_xnor2_1 _28831_ (.Y(_03355_),
    .A(_03017_),
    .B(_03354_));
 sg13g2_nand2_1 _28832_ (.Y(_03356_),
    .A(net1085),
    .B(net5109));
 sg13g2_o21ai_1 _28833_ (.B1(_03356_),
    .Y(_00528_),
    .A1(net5109),
    .A2(_03355_));
 sg13g2_nor2_1 _28834_ (.A(net1380),
    .B(net5240),
    .Y(_03357_));
 sg13g2_mux2_1 _28835_ (.A0(_03351_),
    .A1(_03352_),
    .S(_03017_),
    .X(_03358_));
 sg13g2_xnor2_1 _28836_ (.Y(_03359_),
    .A(_03015_),
    .B(_03358_));
 sg13g2_a21oi_1 _28837_ (.A1(net5240),
    .A2(_03359_),
    .Y(_00529_),
    .B1(_03357_));
 sg13g2_a221oi_1 _28838_ (.B2(_02983_),
    .C1(_03017_),
    .B1(_03347_),
    .A1(_03013_),
    .Y(_03360_),
    .A2(_03014_));
 sg13g2_nand2_1 _28839_ (.Y(_03361_),
    .A(net4504),
    .B(_03360_));
 sg13g2_or2_1 _28840_ (.X(_03362_),
    .B(_03352_),
    .A(_03018_));
 sg13g2_nand2_1 _28841_ (.Y(_03363_),
    .A(_03361_),
    .B(_03362_));
 sg13g2_xor2_1 _28842_ (.B(_03363_),
    .A(_03012_),
    .X(_03364_));
 sg13g2_nand2_1 _28843_ (.Y(_03365_),
    .A(net1080),
    .B(net5109));
 sg13g2_o21ai_1 _28844_ (.B1(_03365_),
    .Y(_00530_),
    .A1(net5109),
    .A2(_03364_));
 sg13g2_nor2_1 _28845_ (.A(net1353),
    .B(net5240),
    .Y(_03366_));
 sg13g2_nand2_1 _28846_ (.Y(_03367_),
    .A(_03012_),
    .B(_03360_));
 sg13g2_a22oi_1 _28847_ (.Y(_03368_),
    .B1(_03362_),
    .B2(_03367_),
    .A2(_03012_),
    .A1(net4487));
 sg13g2_xor2_1 _28848_ (.B(_03368_),
    .A(_03010_),
    .X(_03369_));
 sg13g2_a21oi_1 _28849_ (.A1(net5240),
    .A2(_03369_),
    .Y(_00531_),
    .B1(_03366_));
 sg13g2_nor2_1 _28850_ (.A(net1372),
    .B(net5240),
    .Y(_03370_));
 sg13g2_nor2b_1 _28851_ (.A(_03367_),
    .B_N(_03010_),
    .Y(_03371_));
 sg13g2_nand2_1 _28852_ (.Y(_03372_),
    .A(_03019_),
    .B(_03353_));
 sg13g2_a22oi_1 _28853_ (.Y(_03373_),
    .B1(_03371_),
    .B2(net4504),
    .A2(_03353_),
    .A1(_03019_));
 sg13g2_xnor2_1 _28854_ (.Y(_03374_),
    .A(_02981_),
    .B(_03373_));
 sg13g2_a21oi_1 _28855_ (.A1(net5240),
    .A2(_03374_),
    .Y(_00532_),
    .B1(_03370_));
 sg13g2_nor2_1 _28856_ (.A(net1177),
    .B(net5241),
    .Y(_03375_));
 sg13g2_nand4_1 _28857_ (.B(_03010_),
    .C(_03012_),
    .A(_02981_),
    .Y(_03376_),
    .D(_03360_));
 sg13g2_a22oi_1 _28858_ (.Y(_03377_),
    .B1(_03372_),
    .B2(_03376_),
    .A2(_02981_),
    .A1(net4487));
 sg13g2_xnor2_1 _28859_ (.Y(_03378_),
    .A(_02979_),
    .B(_03377_));
 sg13g2_a21oi_1 _28860_ (.A1(net5241),
    .A2(_03378_),
    .Y(_00533_),
    .B1(_03375_));
 sg13g2_nor2_1 _28861_ (.A(_02979_),
    .B(_03376_),
    .Y(_03379_));
 sg13g2_and2_1 _28862_ (.A(_03022_),
    .B(net4473),
    .X(_03380_));
 sg13g2_inv_1 _28863_ (.Y(_03381_),
    .A(net4452));
 sg13g2_a21oi_1 _28864_ (.A1(net4503),
    .A2(_03379_),
    .Y(_03382_),
    .B1(net4452));
 sg13g2_xnor2_1 _28865_ (.Y(_03383_),
    .A(_03040_),
    .B(_03382_));
 sg13g2_nand2_1 _28866_ (.Y(_03384_),
    .A(net1087),
    .B(net5109));
 sg13g2_o21ai_1 _28867_ (.B1(_03384_),
    .Y(_00534_),
    .A1(net5109),
    .A2(_03383_));
 sg13g2_nor2_1 _28868_ (.A(net2175),
    .B(net5242),
    .Y(_03385_));
 sg13g2_nand2_1 _28869_ (.Y(_03386_),
    .A(_03040_),
    .B(_03379_));
 sg13g2_a22oi_1 _28870_ (.Y(_03387_),
    .B1(_03381_),
    .B2(_03386_),
    .A2(_03040_),
    .A1(net4488));
 sg13g2_xnor2_1 _28871_ (.Y(_03388_),
    .A(_03036_),
    .B(_03387_));
 sg13g2_a21oi_1 _28872_ (.A1(net5242),
    .A2(_03388_),
    .Y(_00535_),
    .B1(_03385_));
 sg13g2_nor4_1 _28873_ (.A(_02979_),
    .B(_03036_),
    .C(_03039_),
    .D(_03376_),
    .Y(_03389_));
 sg13g2_a22oi_1 _28874_ (.Y(_03390_),
    .B1(_03389_),
    .B2(net4503),
    .A2(net4452),
    .A1(_03041_));
 sg13g2_xnor2_1 _28875_ (.Y(_03391_),
    .A(_03043_),
    .B(_03390_));
 sg13g2_nand2_1 _28876_ (.Y(_03392_),
    .A(net1076),
    .B(net5111));
 sg13g2_o21ai_1 _28877_ (.B1(_03392_),
    .Y(_00536_),
    .A1(net5111),
    .A2(_03391_));
 sg13g2_nor2_1 _28878_ (.A(net1768),
    .B(net5250),
    .Y(_03393_));
 sg13g2_and2_1 _28879_ (.A(_03043_),
    .B(_03389_),
    .X(_03394_));
 sg13g2_a21oi_1 _28880_ (.A1(_03041_),
    .A2(net4452),
    .Y(_03395_),
    .B1(_03394_));
 sg13g2_a21oi_1 _28881_ (.A1(net4488),
    .A2(_03043_),
    .Y(_03396_),
    .B1(_03395_));
 sg13g2_xor2_1 _28882_ (.B(_03396_),
    .A(_03034_),
    .X(_03397_));
 sg13g2_a21oi_1 _28883_ (.A1(net5250),
    .A2(_03397_),
    .Y(_00537_),
    .B1(_03393_));
 sg13g2_nor2_1 _28884_ (.A(net2181),
    .B(net5242),
    .Y(_03398_));
 sg13g2_nand3_1 _28885_ (.B(_03034_),
    .C(_03394_),
    .A(net4503),
    .Y(_03399_));
 sg13g2_nand2b_1 _28886_ (.Y(_03400_),
    .B(net4452),
    .A_N(_03044_));
 sg13g2_nand2_1 _28887_ (.Y(_03401_),
    .A(_03399_),
    .B(_03400_));
 sg13g2_xor2_1 _28888_ (.B(_03401_),
    .A(_03046_),
    .X(_03402_));
 sg13g2_a21oi_1 _28889_ (.A1(net5242),
    .A2(_03402_),
    .Y(_00538_),
    .B1(_03398_));
 sg13g2_nor2_1 _28890_ (.A(net1155),
    .B(net5251),
    .Y(_03403_));
 sg13g2_and3_1 _28891_ (.X(_03404_),
    .A(_03034_),
    .B(_03046_),
    .C(_03394_));
 sg13g2_nand4_1 _28892_ (.B(_03043_),
    .C(_03046_),
    .A(_03034_),
    .Y(_03405_),
    .D(_03389_));
 sg13g2_a22oi_1 _28893_ (.Y(_03406_),
    .B1(_03400_),
    .B2(_03405_),
    .A2(_03046_),
    .A1(net4488));
 sg13g2_xnor2_1 _28894_ (.Y(_03407_),
    .A(_03031_),
    .B(_03406_));
 sg13g2_a21oi_1 _28895_ (.A1(net5251),
    .A2(_03407_),
    .Y(_00539_),
    .B1(_03403_));
 sg13g2_nor2_1 _28896_ (.A(net1386),
    .B(net5250),
    .Y(_03408_));
 sg13g2_nand2_1 _28897_ (.Y(_03409_),
    .A(_03032_),
    .B(_03404_));
 sg13g2_nor2_1 _28898_ (.A(net4489),
    .B(_03409_),
    .Y(_03410_));
 sg13g2_a21oi_1 _28899_ (.A1(_03047_),
    .A2(net4452),
    .Y(_03411_),
    .B1(_03410_));
 sg13g2_xnor2_1 _28900_ (.Y(_03412_),
    .A(_03050_),
    .B(_03411_));
 sg13g2_a21oi_1 _28901_ (.A1(net5250),
    .A2(_03412_),
    .Y(_00540_),
    .B1(_03408_));
 sg13g2_nor2_1 _28902_ (.A(net1228),
    .B(net5251),
    .Y(_03413_));
 sg13g2_nor2_1 _28903_ (.A(_03049_),
    .B(_03409_),
    .Y(_03414_));
 sg13g2_a21oi_1 _28904_ (.A1(_03047_),
    .A2(net4453),
    .Y(_03415_),
    .B1(_03414_));
 sg13g2_a21oi_1 _28905_ (.A1(net4489),
    .A2(_03050_),
    .Y(_03416_),
    .B1(_03415_));
 sg13g2_xnor2_1 _28906_ (.Y(_03417_),
    .A(_03029_),
    .B(_03416_));
 sg13g2_a21oi_1 _28907_ (.A1(net5251),
    .A2(_03417_),
    .Y(_00541_),
    .B1(_03413_));
 sg13g2_nor2_1 _28908_ (.A(net1262),
    .B(net5251),
    .Y(_03418_));
 sg13g2_nor4_1 _28909_ (.A(_03029_),
    .B(_03031_),
    .C(_03049_),
    .D(_03405_),
    .Y(_03419_));
 sg13g2_a22oi_1 _28910_ (.Y(_03420_),
    .B1(_03419_),
    .B2(net4507),
    .A2(net4452),
    .A1(_03052_));
 sg13g2_xnor2_1 _28911_ (.Y(_03421_),
    .A(_03054_),
    .B(_03420_));
 sg13g2_a21oi_1 _28912_ (.A1(net5251),
    .A2(_03421_),
    .Y(_00542_),
    .B1(_03418_));
 sg13g2_nor2_1 _28913_ (.A(net1259),
    .B(net5251),
    .Y(_03422_));
 sg13g2_and2_1 _28914_ (.A(_03054_),
    .B(_03419_),
    .X(_03423_));
 sg13g2_a21oi_1 _28915_ (.A1(_03052_),
    .A2(net4452),
    .Y(_03424_),
    .B1(_03423_));
 sg13g2_a21oi_1 _28916_ (.A1(net4489),
    .A2(_03054_),
    .Y(_03425_),
    .B1(_03424_));
 sg13g2_xor2_1 _28917_ (.B(_03425_),
    .A(_03027_),
    .X(_03426_));
 sg13g2_a21oi_1 _28918_ (.A1(net5252),
    .A2(_03426_),
    .Y(_00543_),
    .B1(_03422_));
 sg13g2_nor2_1 _28919_ (.A(net1175),
    .B(net5251),
    .Y(_03427_));
 sg13g2_and2_1 _28920_ (.A(_03027_),
    .B(_03423_),
    .X(_03428_));
 sg13g2_nand2_1 _28921_ (.Y(_03429_),
    .A(_03056_),
    .B(net4453));
 sg13g2_a22oi_1 _28922_ (.Y(_03430_),
    .B1(_03428_),
    .B2(net4507),
    .A2(net4453),
    .A1(_03056_));
 sg13g2_xnor2_1 _28923_ (.Y(_03431_),
    .A(_03058_),
    .B(_03430_));
 sg13g2_a21oi_1 _28924_ (.A1(net5252),
    .A2(_03431_),
    .Y(_00544_),
    .B1(_03427_));
 sg13g2_nor2_1 _28925_ (.A(net2027),
    .B(net5250),
    .Y(_03432_));
 sg13g2_and2_1 _28926_ (.A(_03058_),
    .B(_03428_),
    .X(_03433_));
 sg13g2_nand4_1 _28927_ (.B(_03054_),
    .C(_03058_),
    .A(_03027_),
    .Y(_03434_),
    .D(_03419_));
 sg13g2_a22oi_1 _28928_ (.Y(_03435_),
    .B1(_03429_),
    .B2(_03434_),
    .A2(_03058_),
    .A1(net4489));
 sg13g2_xnor2_1 _28929_ (.Y(_03436_),
    .A(_03024_),
    .B(_03435_));
 sg13g2_a21oi_1 _28930_ (.A1(net5252),
    .A2(_03436_),
    .Y(_00545_),
    .B1(_03432_));
 sg13g2_nor2_1 _28931_ (.A(net1388),
    .B(net5250),
    .Y(_03437_));
 sg13g2_nand2_1 _28932_ (.Y(_03438_),
    .A(_03025_),
    .B(_03433_));
 sg13g2_nand2_1 _28933_ (.Y(_03439_),
    .A(_03059_),
    .B(net4453));
 sg13g2_o21ai_1 _28934_ (.B1(_03439_),
    .Y(_03440_),
    .A1(net4489),
    .A2(_03438_));
 sg13g2_xnor2_1 _28935_ (.Y(_03441_),
    .A(_02977_),
    .B(_03440_));
 sg13g2_a21oi_1 _28936_ (.A1(net5252),
    .A2(_03441_),
    .Y(_00546_),
    .B1(_03437_));
 sg13g2_nor2_1 _28937_ (.A(net1339),
    .B(net5250),
    .Y(_03442_));
 sg13g2_o21ai_1 _28938_ (.B1(_03439_),
    .Y(_03443_),
    .A1(_02977_),
    .A2(_03438_));
 sg13g2_o21ai_1 _28939_ (.B1(_03443_),
    .Y(_03444_),
    .A1(net4507),
    .A2(_02977_));
 sg13g2_xor2_1 _28940_ (.B(_03444_),
    .A(_02975_),
    .X(_03445_));
 sg13g2_a21oi_1 _28941_ (.A1(net5250),
    .A2(_03445_),
    .Y(_00547_),
    .B1(_03442_));
 sg13g2_nor4_2 _28942_ (.A(_02975_),
    .B(_02977_),
    .C(_03024_),
    .Y(_03446_),
    .D(_03434_));
 sg13g2_nand2_1 _28943_ (.Y(_03447_),
    .A(net4506),
    .B(_03446_));
 sg13g2_nand2b_1 _28944_ (.Y(_03448_),
    .B(net4476),
    .A_N(_03060_));
 sg13g2_nand2_1 _28945_ (.Y(_03449_),
    .A(_03447_),
    .B(_03448_));
 sg13g2_xor2_1 _28946_ (.B(_03449_),
    .A(_03064_),
    .X(_03450_));
 sg13g2_nand2_1 _28947_ (.Y(_03451_),
    .A(net1078),
    .B(net5116));
 sg13g2_o21ai_1 _28948_ (.B1(_03451_),
    .Y(_00548_),
    .A1(net5116),
    .A2(_03450_));
 sg13g2_nor2_1 _28949_ (.A(net1356),
    .B(net5253),
    .Y(_03452_));
 sg13g2_nand2_1 _28950_ (.Y(_03453_),
    .A(_03064_),
    .B(_03446_));
 sg13g2_a22oi_1 _28951_ (.Y(_03454_),
    .B1(_03448_),
    .B2(_03453_),
    .A2(_03064_),
    .A1(net4491));
 sg13g2_xor2_1 _28952_ (.B(_03454_),
    .A(_03062_),
    .X(_03455_));
 sg13g2_a21oi_1 _28953_ (.A1(net5253),
    .A2(_03455_),
    .Y(_00549_),
    .B1(_03452_));
 sg13g2_nand3_1 _28954_ (.B(_03064_),
    .C(_03446_),
    .A(_03062_),
    .Y(_03456_));
 sg13g2_nand2_1 _28955_ (.Y(_03457_),
    .A(net4508),
    .B(_03456_));
 sg13g2_o21ai_1 _28956_ (.B1(_03457_),
    .Y(_03458_),
    .A1(_03065_),
    .A2(net4470));
 sg13g2_xnor2_1 _28957_ (.Y(_03459_),
    .A(_02973_),
    .B(_03458_));
 sg13g2_nand2_1 _28958_ (.Y(_03460_),
    .A(net1079),
    .B(net5113));
 sg13g2_o21ai_1 _28959_ (.B1(_03460_),
    .Y(_00550_),
    .A1(net5113),
    .A2(_03459_));
 sg13g2_nor2_1 _28960_ (.A(net1265),
    .B(net5258),
    .Y(_03461_));
 sg13g2_and2_1 _28961_ (.A(_02973_),
    .B(_03456_),
    .X(_03462_));
 sg13g2_nor2_1 _28962_ (.A(net4490),
    .B(_03462_),
    .Y(_03463_));
 sg13g2_nor2_1 _28963_ (.A(net4474),
    .B(_03463_),
    .Y(_03464_));
 sg13g2_nor2_1 _28964_ (.A(_03068_),
    .B(_03464_),
    .Y(_03465_));
 sg13g2_xor2_1 _28965_ (.B(_03464_),
    .A(_03068_),
    .X(_03466_));
 sg13g2_a21oi_1 _28966_ (.A1(net5257),
    .A2(_03466_),
    .Y(_00551_),
    .B1(_03461_));
 sg13g2_nor2_1 _28967_ (.A(net4474),
    .B(_03465_),
    .Y(_03467_));
 sg13g2_xnor2_1 _28968_ (.Y(_03468_),
    .A(_03071_),
    .B(_03467_));
 sg13g2_nand2_1 _28969_ (.Y(_03469_),
    .A(net1077),
    .B(net5113));
 sg13g2_o21ai_1 _28970_ (.B1(_03469_),
    .Y(_00552_),
    .A1(net5113),
    .A2(_03468_));
 sg13g2_nor2_1 _28971_ (.A(net1144),
    .B(net5258),
    .Y(_03470_));
 sg13g2_a221oi_1 _28972_ (.B2(_02973_),
    .C1(_03068_),
    .B1(_03456_),
    .A1(_03069_),
    .Y(_03471_),
    .A2(_03070_));
 sg13g2_or3_1 _28973_ (.A(_03068_),
    .B(_03072_),
    .C(_03462_),
    .X(_03472_));
 sg13g2_a22oi_1 _28974_ (.Y(_03473_),
    .B1(net4470),
    .B2(_03472_),
    .A2(_03071_),
    .A1(net4490));
 sg13g2_xor2_1 _28975_ (.B(_03473_),
    .A(_03074_),
    .X(_03474_));
 sg13g2_a21oi_1 _28976_ (.A1(net5257),
    .A2(_03474_),
    .Y(_00553_),
    .B1(_03470_));
 sg13g2_nor2_1 _28977_ (.A(net1171),
    .B(net5257),
    .Y(_03475_));
 sg13g2_and2_1 _28978_ (.A(_03074_),
    .B(_03471_),
    .X(_03476_));
 sg13g2_a21oi_1 _28979_ (.A1(net4508),
    .A2(_03476_),
    .Y(_03477_),
    .B1(net4474));
 sg13g2_xnor2_1 _28980_ (.Y(_03478_),
    .A(_03094_),
    .B(_03477_));
 sg13g2_a21oi_1 _28981_ (.A1(net5257),
    .A2(_03478_),
    .Y(_00554_),
    .B1(_03475_));
 sg13g2_nor2_1 _28982_ (.A(net1352),
    .B(net5258),
    .Y(_03479_));
 sg13g2_and2_1 _28983_ (.A(_03094_),
    .B(_03476_),
    .X(_03480_));
 sg13g2_nand2_1 _28984_ (.Y(_03481_),
    .A(net4490),
    .B(_03094_));
 sg13g2_o21ai_1 _28985_ (.B1(_03481_),
    .Y(_03482_),
    .A1(net4474),
    .A2(_03480_));
 sg13g2_xnor2_1 _28986_ (.Y(_03483_),
    .A(_03091_),
    .B(_03482_));
 sg13g2_a21oi_1 _28987_ (.A1(net5258),
    .A2(_03483_),
    .Y(_00555_),
    .B1(_03479_));
 sg13g2_nor2_1 _28988_ (.A(net1176),
    .B(net5257),
    .Y(_03484_));
 sg13g2_and4_1 _28989_ (.A(_03074_),
    .B(_03091_),
    .C(_03094_),
    .D(_03471_),
    .X(_03485_));
 sg13g2_a21oi_1 _28990_ (.A1(net4508),
    .A2(_03485_),
    .Y(_03486_),
    .B1(net4474));
 sg13g2_xnor2_1 _28991_ (.Y(_03487_),
    .A(_03080_),
    .B(_03486_));
 sg13g2_a21oi_1 _28992_ (.A1(net5257),
    .A2(_03487_),
    .Y(_00556_),
    .B1(_03484_));
 sg13g2_nor2_1 _28993_ (.A(net1188),
    .B(net5257),
    .Y(_03488_));
 sg13g2_nand2_1 _28994_ (.Y(_03489_),
    .A(_03080_),
    .B(_03485_));
 sg13g2_a22oi_1 _28995_ (.Y(_03490_),
    .B1(net4470),
    .B2(_03489_),
    .A2(_03080_),
    .A1(net4490));
 sg13g2_xor2_1 _28996_ (.B(_03490_),
    .A(_02970_),
    .X(_03491_));
 sg13g2_a21oi_1 _28997_ (.A1(net5257),
    .A2(_03491_),
    .Y(_00557_),
    .B1(_03488_));
 sg13g2_nor2_1 _28998_ (.A(net1197),
    .B(net5258),
    .Y(_03492_));
 sg13g2_nor2b_1 _28999_ (.A(_03489_),
    .B_N(_02970_),
    .Y(_03493_));
 sg13g2_a21oi_1 _29000_ (.A1(net4508),
    .A2(_03493_),
    .Y(_03494_),
    .B1(net4474));
 sg13g2_xnor2_1 _29001_ (.Y(_03495_),
    .A(_03076_),
    .B(_03494_));
 sg13g2_a21oi_1 _29002_ (.A1(net5258),
    .A2(_03495_),
    .Y(_00558_),
    .B1(_03492_));
 sg13g2_nor2_1 _29003_ (.A(net1246),
    .B(net5259),
    .Y(_03496_));
 sg13g2_nand4_1 _29004_ (.B(_03076_),
    .C(_03080_),
    .A(_02970_),
    .Y(_03497_),
    .D(_03485_));
 sg13g2_a22oi_1 _29005_ (.Y(_03498_),
    .B1(net4470),
    .B2(_03497_),
    .A2(_03076_),
    .A1(net4491));
 sg13g2_xnor2_1 _29006_ (.Y(_03499_),
    .A(_03093_),
    .B(_03498_));
 sg13g2_a21oi_1 _29007_ (.A1(net5259),
    .A2(_03499_),
    .Y(_00559_),
    .B1(_03496_));
 sg13g2_nor2_1 _29008_ (.A(net1358),
    .B(net5265),
    .Y(_03500_));
 sg13g2_nor2_1 _29009_ (.A(_03093_),
    .B(_03497_),
    .Y(_03501_));
 sg13g2_a21oi_1 _29010_ (.A1(net4512),
    .A2(_03501_),
    .Y(_03502_),
    .B1(net4475));
 sg13g2_xnor2_1 _29011_ (.Y(_03503_),
    .A(_03097_),
    .B(_03502_));
 sg13g2_a21oi_1 _29012_ (.A1(net5259),
    .A2(_03503_),
    .Y(_00560_),
    .B1(_03500_));
 sg13g2_nor2_1 _29013_ (.A(net1306),
    .B(net5259),
    .Y(_03504_));
 sg13g2_nor3_1 _29014_ (.A(_03093_),
    .B(_03096_),
    .C(_03497_),
    .Y(_03505_));
 sg13g2_nand2_1 _29015_ (.Y(_03506_),
    .A(net4490),
    .B(_03097_));
 sg13g2_o21ai_1 _29016_ (.B1(_03506_),
    .Y(_03507_),
    .A1(net4475),
    .A2(_03505_));
 sg13g2_xnor2_1 _29017_ (.Y(_03508_),
    .A(_03082_),
    .B(_03507_));
 sg13g2_a21oi_1 _29018_ (.A1(net5259),
    .A2(_03508_),
    .Y(_00561_),
    .B1(_03504_));
 sg13g2_nor2_1 _29019_ (.A(net1290),
    .B(net5267),
    .Y(_03509_));
 sg13g2_nor4_2 _29020_ (.A(_03083_),
    .B(_03093_),
    .C(_03096_),
    .Y(_03510_),
    .D(_03497_));
 sg13g2_a21oi_1 _29021_ (.A1(net4515),
    .A2(_03510_),
    .Y(_03511_),
    .B1(net4479));
 sg13g2_xnor2_1 _29022_ (.Y(_03512_),
    .A(_03089_),
    .B(_03511_));
 sg13g2_a21oi_1 _29023_ (.A1(net5267),
    .A2(_03512_),
    .Y(_00562_),
    .B1(_03509_));
 sg13g2_nor2_1 _29024_ (.A(net1178),
    .B(net5267),
    .Y(_03513_));
 sg13g2_nand2_1 _29025_ (.Y(_03514_),
    .A(_03089_),
    .B(_03510_));
 sg13g2_a22oi_1 _29026_ (.Y(_03515_),
    .B1(net4471),
    .B2(_03514_),
    .A2(_03089_),
    .A1(net4493));
 sg13g2_xor2_1 _29027_ (.B(_03515_),
    .A(_02964_),
    .X(_03516_));
 sg13g2_a21oi_1 _29028_ (.A1(net5267),
    .A2(_03516_),
    .Y(_00563_),
    .B1(_03513_));
 sg13g2_nor2_1 _29029_ (.A(net1186),
    .B(net5273),
    .Y(_03517_));
 sg13g2_nor2b_1 _29030_ (.A(_03514_),
    .B_N(_02964_),
    .Y(_03518_));
 sg13g2_a21oi_1 _29031_ (.A1(net4515),
    .A2(_03518_),
    .Y(_03519_),
    .B1(net4479));
 sg13g2_xnor2_1 _29032_ (.Y(_03520_),
    .A(_02966_),
    .B(_03519_));
 sg13g2_a21oi_1 _29033_ (.A1(net5267),
    .A2(_03520_),
    .Y(_00564_),
    .B1(_03517_));
 sg13g2_nor2_1 _29034_ (.A(net1216),
    .B(net5267),
    .Y(_03521_));
 sg13g2_nand4_1 _29035_ (.B(_02966_),
    .C(_03089_),
    .A(_02964_),
    .Y(_03522_),
    .D(_03510_));
 sg13g2_and2_1 _29036_ (.A(net4493),
    .B(_02966_),
    .X(_03523_));
 sg13g2_a21o_1 _29037_ (.A2(_03522_),
    .A1(net4471),
    .B1(_03523_),
    .X(_03524_));
 sg13g2_xnor2_1 _29038_ (.Y(_03525_),
    .A(_03087_),
    .B(_03524_));
 sg13g2_a21oi_1 _29039_ (.A1(net5267),
    .A2(_03525_),
    .Y(_00565_),
    .B1(_03521_));
 sg13g2_nor2_1 _29040_ (.A(net1279),
    .B(net5274),
    .Y(_03526_));
 sg13g2_nor2_1 _29041_ (.A(_03088_),
    .B(_03522_),
    .Y(_03527_));
 sg13g2_a21oi_1 _29042_ (.A1(net4517),
    .A2(_03527_),
    .Y(_03528_),
    .B1(net4477));
 sg13g2_xor2_1 _29043_ (.B(_03528_),
    .A(_02961_),
    .X(_03529_));
 sg13g2_a21oi_1 _29044_ (.A1(net5274),
    .A2(_03529_),
    .Y(_00566_),
    .B1(_03526_));
 sg13g2_nand2_1 _29045_ (.Y(_03530_),
    .A(net1166),
    .B(net5120));
 sg13g2_nor3_1 _29046_ (.A(_02961_),
    .B(_03088_),
    .C(_03522_),
    .Y(_03531_));
 sg13g2_nor2_1 _29047_ (.A(_02959_),
    .B(_03531_),
    .Y(_03532_));
 sg13g2_nor4_1 _29048_ (.A(_02958_),
    .B(_02961_),
    .C(_03088_),
    .D(_03522_),
    .Y(_03533_));
 sg13g2_nand2b_1 _29049_ (.Y(_03534_),
    .B(net4517),
    .A_N(_03533_));
 sg13g2_a21oi_1 _29050_ (.A1(net4494),
    .A2(_02959_),
    .Y(_03535_),
    .B1(net5120));
 sg13g2_o21ai_1 _29051_ (.B1(_03535_),
    .Y(_03536_),
    .A1(_03532_),
    .A2(_03534_));
 sg13g2_o21ai_1 _29052_ (.B1(_03530_),
    .Y(_00567_),
    .A1(net4477),
    .A2(_03536_));
 sg13g2_nor2_1 _29053_ (.A(net1299),
    .B(net5274),
    .Y(_03537_));
 sg13g2_nand2_1 _29054_ (.Y(_03538_),
    .A(net4379),
    .B(_03534_));
 sg13g2_xnor2_1 _29055_ (.Y(_03539_),
    .A(_02955_),
    .B(_03538_));
 sg13g2_a21oi_1 _29056_ (.A1(net5275),
    .A2(_03539_),
    .Y(_00568_),
    .B1(_03537_));
 sg13g2_nor2_1 _29057_ (.A(net1147),
    .B(net5274),
    .Y(_03540_));
 sg13g2_and2_1 _29058_ (.A(_02955_),
    .B(_03533_),
    .X(_03541_));
 sg13g2_a21oi_1 _29059_ (.A1(net4517),
    .A2(_03541_),
    .Y(_03542_),
    .B1(net4477));
 sg13g2_nor2_1 _29060_ (.A(_02953_),
    .B(_03542_),
    .Y(_03543_));
 sg13g2_xor2_1 _29061_ (.B(_03542_),
    .A(_02953_),
    .X(_03544_));
 sg13g2_a21oi_1 _29062_ (.A1(net5274),
    .A2(_03544_),
    .Y(_00569_),
    .B1(_03540_));
 sg13g2_o21ai_1 _29063_ (.B1(_02950_),
    .Y(_03545_),
    .A1(net4477),
    .A2(_03543_));
 sg13g2_nor3_1 _29064_ (.A(_02950_),
    .B(net4477),
    .C(_03543_),
    .Y(_03546_));
 sg13g2_nor2_1 _29065_ (.A(net5120),
    .B(_03546_),
    .Y(_03547_));
 sg13g2_a22oi_1 _29066_ (.Y(_03548_),
    .B1(_03545_),
    .B2(_03547_),
    .A2(net5120),
    .A1(net2550));
 sg13g2_inv_1 _29067_ (.Y(_00570_),
    .A(_03548_));
 sg13g2_nor2_1 _29068_ (.A(net2287),
    .B(net5274),
    .Y(_03549_));
 sg13g2_nor2_1 _29069_ (.A(_02950_),
    .B(_02953_),
    .Y(_03550_));
 sg13g2_nand2_1 _29070_ (.Y(_03551_),
    .A(_03541_),
    .B(_03550_));
 sg13g2_a22oi_1 _29071_ (.Y(_03552_),
    .B1(net4471),
    .B2(_03551_),
    .A2(_02951_),
    .A1(net4494));
 sg13g2_xor2_1 _29072_ (.B(_03552_),
    .A(_02948_),
    .X(_03553_));
 sg13g2_a21oi_1 _29073_ (.A1(net5274),
    .A2(_03553_),
    .Y(_00571_),
    .B1(_03549_));
 sg13g2_nor2_1 _29074_ (.A(net1167),
    .B(net5275),
    .Y(_03554_));
 sg13g2_and4_1 _29075_ (.A(_02948_),
    .B(_02955_),
    .C(_03533_),
    .D(_03550_),
    .X(_03555_));
 sg13g2_a21oi_1 _29076_ (.A1(net4517),
    .A2(_03555_),
    .Y(_03556_),
    .B1(net4477));
 sg13g2_xnor2_1 _29077_ (.Y(_03557_),
    .A(_02946_),
    .B(_03556_));
 sg13g2_a21oi_1 _29078_ (.A1(net5275),
    .A2(_03557_),
    .Y(_00572_),
    .B1(_03554_));
 sg13g2_nor2_1 _29079_ (.A(net1179),
    .B(net5274),
    .Y(_03558_));
 sg13g2_nor2_1 _29080_ (.A(_02946_),
    .B(net4478),
    .Y(_03559_));
 sg13g2_nor2_1 _29081_ (.A(_03556_),
    .B(_03559_),
    .Y(_03560_));
 sg13g2_xnor2_1 _29082_ (.Y(_03561_),
    .A(_02944_),
    .B(_03560_));
 sg13g2_a21oi_1 _29083_ (.A1(net5275),
    .A2(_03561_),
    .Y(_00573_),
    .B1(_03558_));
 sg13g2_and2_1 _29084_ (.A(_02943_),
    .B(_02946_),
    .X(_03562_));
 sg13g2_and2_1 _29085_ (.A(_03555_),
    .B(_03562_),
    .X(_03563_));
 sg13g2_a21oi_1 _29086_ (.A1(net4516),
    .A2(_03563_),
    .Y(_03564_),
    .B1(net4478));
 sg13g2_xnor2_1 _29087_ (.Y(_03565_),
    .A(_02938_),
    .B(_03564_));
 sg13g2_nand2_1 _29088_ (.Y(_03566_),
    .A(net1090),
    .B(net5120));
 sg13g2_o21ai_1 _29089_ (.B1(_03566_),
    .Y(_00574_),
    .A1(net5120),
    .A2(_03565_));
 sg13g2_nand2_1 _29090_ (.Y(_03567_),
    .A(net1091),
    .B(net5120));
 sg13g2_and2_1 _29091_ (.A(_02937_),
    .B(_02938_),
    .X(_03568_));
 sg13g2_a21o_1 _29092_ (.A2(_03568_),
    .A1(_03563_),
    .B1(net4494),
    .X(_03569_));
 sg13g2_a21oi_1 _29093_ (.A1(_02938_),
    .A2(_03563_),
    .Y(_03570_),
    .B1(_02937_));
 sg13g2_a21oi_1 _29094_ (.A1(net4494),
    .A2(_02937_),
    .Y(_03571_),
    .B1(net5122));
 sg13g2_o21ai_1 _29095_ (.B1(_03571_),
    .Y(_03572_),
    .A1(_03569_),
    .A2(_03570_));
 sg13g2_o21ai_1 _29096_ (.B1(_03567_),
    .Y(_00575_),
    .A1(net4477),
    .A2(_03572_));
 sg13g2_nor2b_1 _29097_ (.A(net4462),
    .B_N(_03569_),
    .Y(_03573_));
 sg13g2_xnor2_1 _29098_ (.Y(_03574_),
    .A(_02940_),
    .B(_03573_));
 sg13g2_nand2_1 _29099_ (.Y(_03575_),
    .A(net1084),
    .B(net5121));
 sg13g2_o21ai_1 _29100_ (.B1(_03575_),
    .Y(_00576_),
    .A1(net5121),
    .A2(_03574_));
 sg13g2_nand2_1 _29101_ (.Y(_03576_),
    .A(net1096),
    .B(net5121));
 sg13g2_and4_1 _29102_ (.A(_02941_),
    .B(_03555_),
    .C(_03562_),
    .D(_03568_),
    .X(_03577_));
 sg13g2_nor2_1 _29103_ (.A(_02934_),
    .B(_03577_),
    .Y(_03578_));
 sg13g2_nand2_1 _29104_ (.Y(_03579_),
    .A(_02934_),
    .B(_03577_));
 sg13g2_nand2_1 _29105_ (.Y(_03580_),
    .A(net4520),
    .B(_03579_));
 sg13g2_a21oi_1 _29106_ (.A1(net4495),
    .A2(_02934_),
    .Y(_03581_),
    .B1(net5122));
 sg13g2_o21ai_1 _29107_ (.B1(_03581_),
    .Y(_03582_),
    .A1(_03578_),
    .A2(_03580_));
 sg13g2_o21ai_1 _29108_ (.B1(_03576_),
    .Y(_00577_),
    .A1(net4481),
    .A2(_03582_));
 sg13g2_nand2_1 _29109_ (.Y(_03583_),
    .A(net4378),
    .B(_03580_));
 sg13g2_xnor2_1 _29110_ (.Y(_03584_),
    .A(_03112_),
    .B(_03583_));
 sg13g2_nand2_1 _29111_ (.Y(_03585_),
    .A(net1086),
    .B(net5121));
 sg13g2_o21ai_1 _29112_ (.B1(_03585_),
    .Y(_00578_),
    .A1(net5122),
    .A2(_03584_));
 sg13g2_nand2_1 _29113_ (.Y(_03586_),
    .A(net1093),
    .B(net5121));
 sg13g2_and2_1 _29114_ (.A(_03111_),
    .B(_03112_),
    .X(_03587_));
 sg13g2_nand3_1 _29115_ (.B(_03577_),
    .C(_03587_),
    .A(_02934_),
    .Y(_03588_));
 sg13g2_and2_1 _29116_ (.A(net4520),
    .B(_03588_),
    .X(_03589_));
 sg13g2_nand2b_1 _29117_ (.Y(_03590_),
    .B(_03579_),
    .A_N(_03111_));
 sg13g2_nand3_1 _29118_ (.B(_03589_),
    .C(_03590_),
    .A(_03113_),
    .Y(_03591_));
 sg13g2_a21oi_1 _29119_ (.A1(net4495),
    .A2(_03111_),
    .Y(_03592_),
    .B1(net5126));
 sg13g2_nand2_1 _29120_ (.Y(_03593_),
    .A(_03591_),
    .B(_03592_));
 sg13g2_o21ai_1 _29121_ (.B1(_03586_),
    .Y(_00579_),
    .A1(net4481),
    .A2(_03593_));
 sg13g2_nor2_1 _29122_ (.A(net4465),
    .B(_03589_),
    .Y(_03594_));
 sg13g2_xor2_1 _29123_ (.B(_03594_),
    .A(_02931_),
    .X(_03595_));
 sg13g2_nor2_1 _29124_ (.A(net1219),
    .B(net5276),
    .Y(_03596_));
 sg13g2_a21oi_1 _29125_ (.A1(net5276),
    .A2(_03595_),
    .Y(_00580_),
    .B1(_03596_));
 sg13g2_nor2_1 _29126_ (.A(net1303),
    .B(net5281),
    .Y(_03597_));
 sg13g2_xnor2_1 _29127_ (.Y(_03598_),
    .A(net4520),
    .B(_02931_));
 sg13g2_nand2_1 _29128_ (.Y(_03599_),
    .A(_03594_),
    .B(_03598_));
 sg13g2_xor2_1 _29129_ (.B(_03599_),
    .A(_03115_),
    .X(_03600_));
 sg13g2_a21oi_1 _29130_ (.A1(net5281),
    .A2(_03600_),
    .Y(_00581_),
    .B1(_03597_));
 sg13g2_nor2_1 _29131_ (.A(net1263),
    .B(net5281),
    .Y(_03601_));
 sg13g2_nor2b_1 _29132_ (.A(_03115_),
    .B_N(_02931_),
    .Y(_03602_));
 sg13g2_and4_1 _29133_ (.A(_02934_),
    .B(_03577_),
    .C(_03587_),
    .D(_03602_),
    .X(_03603_));
 sg13g2_a21oi_1 _29134_ (.A1(net4520),
    .A2(_03603_),
    .Y(_03604_),
    .B1(net4481));
 sg13g2_xnor2_1 _29135_ (.Y(_03605_),
    .A(_03108_),
    .B(_03604_));
 sg13g2_a21oi_1 _29136_ (.A1(net5281),
    .A2(_03605_),
    .Y(_00582_),
    .B1(_03601_));
 sg13g2_nand2_1 _29137_ (.Y(_03606_),
    .A(net1083),
    .B(net5125));
 sg13g2_and2_1 _29138_ (.A(_03108_),
    .B(_03603_),
    .X(_03607_));
 sg13g2_and2_1 _29139_ (.A(_02929_),
    .B(_03108_),
    .X(_03608_));
 sg13g2_and2_1 _29140_ (.A(_03603_),
    .B(_03608_),
    .X(_03609_));
 sg13g2_nor2_1 _29141_ (.A(net4495),
    .B(_03609_),
    .Y(_03610_));
 sg13g2_o21ai_1 _29142_ (.B1(_03610_),
    .Y(_03611_),
    .A1(_02929_),
    .A2(_03607_));
 sg13g2_a21oi_1 _29143_ (.A1(net4495),
    .A2(_02929_),
    .Y(_03612_),
    .B1(net5126));
 sg13g2_nand2_1 _29144_ (.Y(_03613_),
    .A(_03611_),
    .B(_03612_));
 sg13g2_o21ai_1 _29145_ (.B1(_03606_),
    .Y(_00583_),
    .A1(net4481),
    .A2(_03613_));
 sg13g2_nor2_1 _29146_ (.A(net4464),
    .B(_03610_),
    .Y(_03614_));
 sg13g2_xor2_1 _29147_ (.B(_03614_),
    .A(_02927_),
    .X(_03615_));
 sg13g2_nand2_1 _29148_ (.Y(_03616_),
    .A(net1105),
    .B(net5125));
 sg13g2_o21ai_1 _29149_ (.B1(_03616_),
    .Y(_00584_),
    .A1(net5125),
    .A2(_03615_));
 sg13g2_nand2_1 _29150_ (.Y(_03617_),
    .A(net1081),
    .B(net5124));
 sg13g2_a21o_1 _29151_ (.A2(_03614_),
    .A1(_02927_),
    .B1(net4481),
    .X(_03618_));
 sg13g2_xor2_1 _29152_ (.B(_03618_),
    .A(_03132_),
    .X(_03619_));
 sg13g2_o21ai_1 _29153_ (.B1(_03617_),
    .Y(_00585_),
    .A1(net5124),
    .A2(_03619_));
 sg13g2_nor2_1 _29154_ (.A(net1128),
    .B(net5285),
    .Y(_03620_));
 sg13g2_nand3_1 _29155_ (.B(_03132_),
    .C(_03609_),
    .A(_02927_),
    .Y(_03621_));
 sg13g2_a21o_1 _29156_ (.A2(_03621_),
    .A1(net4521),
    .B1(net4464),
    .X(_03622_));
 sg13g2_xnor2_1 _29157_ (.Y(_03623_),
    .A(_03139_),
    .B(_03622_));
 sg13g2_a21oi_1 _29158_ (.A1(net5285),
    .A2(_03623_),
    .Y(_00586_),
    .B1(_03620_));
 sg13g2_nand2_1 _29159_ (.Y(_03624_),
    .A(_03137_),
    .B(_03139_));
 sg13g2_nor2_1 _29160_ (.A(_03621_),
    .B(_03624_),
    .Y(_03625_));
 sg13g2_nor2_1 _29161_ (.A(net4496),
    .B(_03625_),
    .Y(_03626_));
 sg13g2_a21oi_1 _29162_ (.A1(_03138_),
    .A2(_03621_),
    .Y(_03627_),
    .B1(_03140_));
 sg13g2_o21ai_1 _29163_ (.B1(net5288),
    .Y(_03628_),
    .A1(net4521),
    .A2(_03624_));
 sg13g2_a21oi_1 _29164_ (.A1(_03626_),
    .A2(_03627_),
    .Y(_03629_),
    .B1(_03628_));
 sg13g2_nand2_1 _29165_ (.Y(_03630_),
    .A(net4471),
    .B(_03629_));
 sg13g2_a21oi_1 _29166_ (.A1(_03137_),
    .A2(net4464),
    .Y(_03631_),
    .B1(_03630_));
 sg13g2_a21o_1 _29167_ (.A2(net5127),
    .A1(net1309),
    .B1(_03631_),
    .X(_00587_));
 sg13g2_nor2_1 _29168_ (.A(net4464),
    .B(_03626_),
    .Y(_03632_));
 sg13g2_xnor2_1 _29169_ (.Y(_03633_),
    .A(_03107_),
    .B(_03632_));
 sg13g2_nand2_1 _29170_ (.Y(_03634_),
    .A(net1092),
    .B(net5127));
 sg13g2_o21ai_1 _29171_ (.B1(_03634_),
    .Y(_00588_),
    .A1(net5133),
    .A2(_03633_));
 sg13g2_nor2_1 _29172_ (.A(net1168),
    .B(net5284),
    .Y(_03635_));
 sg13g2_xnor2_1 _29173_ (.Y(_03636_),
    .A(net4521),
    .B(_03107_));
 sg13g2_nor3_1 _29174_ (.A(net4464),
    .B(_03626_),
    .C(_03636_),
    .Y(_03637_));
 sg13g2_xnor2_1 _29175_ (.Y(_03638_),
    .A(_03134_),
    .B(_03637_));
 sg13g2_a21oi_1 _29176_ (.A1(net5285),
    .A2(_03638_),
    .Y(_00589_),
    .B1(_03635_));
 sg13g2_nor2_1 _29177_ (.A(net1126),
    .B(net5281),
    .Y(_03639_));
 sg13g2_or2_1 _29178_ (.X(_03640_),
    .B(_03624_),
    .A(_03134_));
 sg13g2_nor3_1 _29179_ (.A(_03107_),
    .B(_03621_),
    .C(_03640_),
    .Y(_03641_));
 sg13g2_a21oi_1 _29180_ (.A1(net4522),
    .A2(_03641_),
    .Y(_03642_),
    .B1(net4480));
 sg13g2_xor2_1 _29181_ (.B(_03642_),
    .A(_03146_),
    .X(_03643_));
 sg13g2_a21oi_1 _29182_ (.A1(net5286),
    .A2(_03643_),
    .Y(_00590_),
    .B1(_03639_));
 sg13g2_nand4_1 _29183_ (.B(_03106_),
    .C(_03132_),
    .A(_02927_),
    .Y(_03644_),
    .D(_03608_));
 sg13g2_nor4_1 _29184_ (.A(_03144_),
    .B(_03146_),
    .C(_03640_),
    .D(_03644_),
    .Y(_03645_));
 sg13g2_and2_1 _29185_ (.A(_03603_),
    .B(_03645_),
    .X(_03646_));
 sg13g2_o21ai_1 _29186_ (.B1(_03147_),
    .Y(_03647_),
    .A1(_03145_),
    .A2(_03641_));
 sg13g2_nor3_1 _29187_ (.A(net4496),
    .B(_03646_),
    .C(_03647_),
    .Y(_03648_));
 sg13g2_o21ai_1 _29188_ (.B1(net5288),
    .Y(_03649_),
    .A1(net4522),
    .A2(_03144_));
 sg13g2_nor3_1 _29189_ (.A(net4480),
    .B(_03648_),
    .C(_03649_),
    .Y(_03650_));
 sg13g2_a21o_1 _29190_ (.A2(net5132),
    .A1(net1526),
    .B1(_03650_),
    .X(_00591_));
 sg13g2_o21ai_1 _29191_ (.B1(net4378),
    .Y(_03651_),
    .A1(net4496),
    .A2(_03646_));
 sg13g2_xnor2_1 _29192_ (.Y(_03652_),
    .A(_02922_),
    .B(_03651_));
 sg13g2_nor2_1 _29193_ (.A(net1996),
    .B(net5288),
    .Y(_03653_));
 sg13g2_a21oi_1 _29194_ (.A1(net5288),
    .A2(_03652_),
    .Y(_00592_),
    .B1(_03653_));
 sg13g2_nor2_1 _29195_ (.A(net1253),
    .B(net5289),
    .Y(_03654_));
 sg13g2_nor2_1 _29196_ (.A(_02923_),
    .B(_03130_),
    .Y(_03655_));
 sg13g2_nand2_1 _29197_ (.Y(_03656_),
    .A(_02922_),
    .B(_03646_));
 sg13g2_nor2_1 _29198_ (.A(_03130_),
    .B(_03656_),
    .Y(_03657_));
 sg13g2_xnor2_1 _29199_ (.Y(_03658_),
    .A(_03130_),
    .B(_03656_));
 sg13g2_a22oi_1 _29200_ (.Y(_03659_),
    .B1(_03658_),
    .B2(net4522),
    .A2(net4468),
    .A1(_03130_));
 sg13g2_a21oi_1 _29201_ (.A1(net5289),
    .A2(_03659_),
    .Y(_00593_),
    .B1(_03654_));
 sg13g2_nor2_1 _29202_ (.A(net1143),
    .B(net5289),
    .Y(_03660_));
 sg13g2_a21oi_1 _29203_ (.A1(net4522),
    .A2(_03657_),
    .Y(_03661_),
    .B1(net4480));
 sg13g2_xnor2_1 _29204_ (.Y(_03662_),
    .A(_02924_),
    .B(_03661_));
 sg13g2_a21oi_1 _29205_ (.A1(net5289),
    .A2(_03662_),
    .Y(_00594_),
    .B1(_03660_));
 sg13g2_nand3_1 _29206_ (.B(_03142_),
    .C(_03657_),
    .A(_02924_),
    .Y(_03663_));
 sg13g2_a21o_1 _29207_ (.A2(_03657_),
    .A1(_02924_),
    .B1(_03142_),
    .X(_03664_));
 sg13g2_nand2_1 _29208_ (.Y(_03665_),
    .A(_03663_),
    .B(_03664_));
 sg13g2_a21oi_1 _29209_ (.A1(net4522),
    .A2(_03665_),
    .Y(_03666_),
    .B1(net5132));
 sg13g2_o21ai_1 _29210_ (.B1(_03666_),
    .Y(_03667_),
    .A1(_03142_),
    .A2(net4378));
 sg13g2_o21ai_1 _29211_ (.B1(_03667_),
    .Y(_03668_),
    .A1(net2770),
    .A2(net5289));
 sg13g2_inv_1 _29212_ (.Y(_00595_),
    .A(_03668_));
 sg13g2_nor2_1 _29213_ (.A(net1207),
    .B(net5289),
    .Y(_03669_));
 sg13g2_a21oi_1 _29214_ (.A1(net4522),
    .A2(_03663_),
    .Y(_03670_),
    .B1(net4468));
 sg13g2_xnor2_1 _29215_ (.Y(_03671_),
    .A(_02919_),
    .B(_03670_));
 sg13g2_a21oi_1 _29216_ (.A1(net5289),
    .A2(_03671_),
    .Y(_00596_),
    .B1(_03669_));
 sg13g2_nor2_1 _29217_ (.A(net1203),
    .B(net5290),
    .Y(_03672_));
 sg13g2_xnor2_1 _29218_ (.Y(_03673_),
    .A(net4496),
    .B(_02919_));
 sg13g2_nand2_1 _29219_ (.Y(_03674_),
    .A(_03670_),
    .B(_03673_));
 sg13g2_xor2_1 _29220_ (.B(_03674_),
    .A(_03121_),
    .X(_03675_));
 sg13g2_a21oi_1 _29221_ (.A1(net5289),
    .A2(_03675_),
    .Y(_00597_),
    .B1(_03672_));
 sg13g2_nand4_1 _29222_ (.B(_03142_),
    .C(_03645_),
    .A(_02924_),
    .Y(_03676_),
    .D(_03655_));
 sg13g2_nor3_2 _29223_ (.A(_02919_),
    .B(_03121_),
    .C(_03676_),
    .Y(_03677_));
 sg13g2_and2_1 _29224_ (.A(_03603_),
    .B(_03677_),
    .X(_03678_));
 sg13g2_a21oi_1 _29225_ (.A1(net4526),
    .A2(_03678_),
    .Y(_03679_),
    .B1(net4480));
 sg13g2_xnor2_1 _29226_ (.Y(_03680_),
    .A(_03127_),
    .B(_03679_));
 sg13g2_nand2_1 _29227_ (.Y(_03681_),
    .A(net1097),
    .B(net5128));
 sg13g2_o21ai_1 _29228_ (.B1(_03681_),
    .Y(_00598_),
    .A1(net5128),
    .A2(_03680_));
 sg13g2_nand2_1 _29229_ (.Y(_03682_),
    .A(_03126_),
    .B(_03127_));
 sg13g2_and3_2 _29230_ (.X(_03683_),
    .A(_03126_),
    .B(_03127_),
    .C(_03678_));
 sg13g2_a21oi_1 _29231_ (.A1(_03127_),
    .A2(_03678_),
    .Y(_03684_),
    .B1(_03126_));
 sg13g2_nor3_1 _29232_ (.A(net4496),
    .B(_03683_),
    .C(_03684_),
    .Y(_03685_));
 sg13g2_and2_1 _29233_ (.A(net4496),
    .B(_03126_),
    .X(_03686_));
 sg13g2_nor4_1 _29234_ (.A(net5131),
    .B(net4480),
    .C(_03685_),
    .D(_03686_),
    .Y(_03687_));
 sg13g2_a21o_1 _29235_ (.A2(net5130),
    .A1(net1832),
    .B1(_03687_),
    .X(_00599_));
 sg13g2_nor2_1 _29236_ (.A(net1282),
    .B(net5287),
    .Y(_03688_));
 sg13g2_o21ai_1 _29237_ (.B1(net4378),
    .Y(_03689_),
    .A1(net4496),
    .A2(_03683_));
 sg13g2_xnor2_1 _29238_ (.Y(_03690_),
    .A(_02907_),
    .B(_03689_));
 sg13g2_a21oi_1 _29239_ (.A1(net5287),
    .A2(_03690_),
    .Y(_00600_),
    .B1(_03688_));
 sg13g2_nand2_1 _29240_ (.Y(_03691_),
    .A(_02905_),
    .B(_02907_));
 sg13g2_nand3_1 _29241_ (.B(_02907_),
    .C(_03683_),
    .A(_02905_),
    .Y(_03692_));
 sg13g2_inv_1 _29242_ (.Y(_03693_),
    .A(_03692_));
 sg13g2_a21oi_1 _29243_ (.A1(_02907_),
    .A2(_03683_),
    .Y(_03694_),
    .B1(_02905_));
 sg13g2_o21ai_1 _29244_ (.B1(net4526),
    .Y(_03695_),
    .A1(_03693_),
    .A2(_03694_));
 sg13g2_o21ai_1 _29245_ (.B1(_03695_),
    .Y(_03696_),
    .A1(_02905_),
    .A2(net4378));
 sg13g2_mux2_1 _29246_ (.A0(net2329),
    .A1(_03696_),
    .S(net5288),
    .X(_00601_));
 sg13g2_nor2_1 _29247_ (.A(net1152),
    .B(net5293),
    .Y(_03697_));
 sg13g2_a21oi_1 _29248_ (.A1(net4527),
    .A2(_03693_),
    .Y(_03698_),
    .B1(net4480));
 sg13g2_xor2_1 _29249_ (.B(_03698_),
    .A(_02913_),
    .X(_03699_));
 sg13g2_a21oi_1 _29250_ (.A1(net5293),
    .A2(_03699_),
    .Y(_00602_),
    .B1(_03697_));
 sg13g2_nand2_1 _29251_ (.Y(_03700_),
    .A(_02911_),
    .B(_03692_));
 sg13g2_or2_1 _29252_ (.X(_03701_),
    .B(_02913_),
    .A(_02911_));
 sg13g2_or2_1 _29253_ (.X(_03702_),
    .B(_03701_),
    .A(_03692_));
 sg13g2_nand3_1 _29254_ (.B(_03700_),
    .C(_03702_),
    .A(_02914_),
    .Y(_03703_));
 sg13g2_a221oi_1 _29255_ (.B2(net4525),
    .C1(net5129),
    .B1(_03703_),
    .A1(_02911_),
    .Y(_03704_),
    .A2(net4466));
 sg13g2_a21oi_1 _29256_ (.A1(_14519_),
    .A2(net5129),
    .Y(_00603_),
    .B1(_03704_));
 sg13g2_a21oi_1 _29257_ (.A1(net4525),
    .A2(_03702_),
    .Y(_03705_),
    .B1(net4466));
 sg13g2_xor2_1 _29258_ (.B(_03705_),
    .A(_03122_),
    .X(_03706_));
 sg13g2_nand2_1 _29259_ (.Y(_03707_),
    .A(net1266),
    .B(net5128));
 sg13g2_o21ai_1 _29260_ (.B1(_03707_),
    .Y(_00604_),
    .A1(net5129),
    .A2(_03706_));
 sg13g2_nor2_1 _29261_ (.A(net1415),
    .B(net5287),
    .Y(_03708_));
 sg13g2_xnor2_1 _29262_ (.Y(_03709_),
    .A(net4525),
    .B(_03122_));
 sg13g2_nand2_1 _29263_ (.Y(_03710_),
    .A(_03705_),
    .B(_03709_));
 sg13g2_xnor2_1 _29264_ (.Y(_03711_),
    .A(_02902_),
    .B(_03710_));
 sg13g2_a21oi_1 _29265_ (.A1(net5287),
    .A2(_03711_),
    .Y(_00605_),
    .B1(_03708_));
 sg13g2_and2_1 _29266_ (.A(_02902_),
    .B(_03122_),
    .X(_03712_));
 sg13g2_nand2b_1 _29267_ (.Y(_03713_),
    .B(_03712_),
    .A_N(_03702_));
 sg13g2_a21oi_1 _29268_ (.A1(net4526),
    .A2(_03713_),
    .Y(_03714_),
    .B1(net4466));
 sg13g2_xor2_1 _29269_ (.B(_03714_),
    .A(_02896_),
    .X(_03715_));
 sg13g2_nand2_1 _29270_ (.Y(_03716_),
    .A(net1121),
    .B(net5128));
 sg13g2_o21ai_1 _29271_ (.B1(_03716_),
    .Y(_00606_),
    .A1(net5129),
    .A2(_03715_));
 sg13g2_nand2_1 _29272_ (.Y(_03717_),
    .A(_02895_),
    .B(_03713_));
 sg13g2_nand3b_1 _29273_ (.B(_02896_),
    .C(_03712_),
    .Y(_03718_),
    .A_N(_02895_));
 sg13g2_nor4_1 _29274_ (.A(_03682_),
    .B(_03691_),
    .C(_03701_),
    .D(_03718_),
    .Y(_03719_));
 sg13g2_nand2_2 _29275_ (.Y(_03720_),
    .A(_03678_),
    .B(_03719_));
 sg13g2_nand3b_1 _29276_ (.B(_03717_),
    .C(_03720_),
    .Y(_03721_),
    .A_N(_02897_));
 sg13g2_a221oi_1 _29277_ (.B2(net4525),
    .C1(net5131),
    .B1(_03721_),
    .A1(_02895_),
    .Y(_03722_),
    .A2(net4466));
 sg13g2_a21oi_1 _29278_ (.A1(_14520_),
    .A2(net5129),
    .Y(_00607_),
    .B1(_03722_));
 sg13g2_a21oi_1 _29279_ (.A1(net4525),
    .A2(_03720_),
    .Y(_03723_),
    .B1(net4466));
 sg13g2_nor2_1 _29280_ (.A(net1367),
    .B(net5287),
    .Y(_03724_));
 sg13g2_xnor2_1 _29281_ (.Y(_03725_),
    .A(_02909_),
    .B(_03723_));
 sg13g2_a21oi_1 _29282_ (.A1(net5287),
    .A2(_03725_),
    .Y(_00608_),
    .B1(_03724_));
 sg13g2_or3_1 _29283_ (.A(_02893_),
    .B(_02909_),
    .C(_03720_),
    .X(_03726_));
 sg13g2_o21ai_1 _29284_ (.B1(_02893_),
    .Y(_03727_),
    .A1(_02909_),
    .A2(_03720_));
 sg13g2_nand2_1 _29285_ (.Y(_03728_),
    .A(_03726_),
    .B(_03727_));
 sg13g2_a221oi_1 _29286_ (.B2(net4525),
    .C1(net5128),
    .B1(_03728_),
    .A1(_02893_),
    .Y(_03729_),
    .A2(net4466));
 sg13g2_a21oi_1 _29287_ (.A1(_14521_),
    .A2(net5128),
    .Y(_00609_),
    .B1(_03729_));
 sg13g2_a21oi_1 _29288_ (.A1(net4525),
    .A2(_03726_),
    .Y(_03730_),
    .B1(net4467));
 sg13g2_xnor2_1 _29289_ (.Y(_03731_),
    .A(_02877_),
    .B(_03730_));
 sg13g2_nand2_1 _29290_ (.Y(_03732_),
    .A(net1110),
    .B(net5129));
 sg13g2_o21ai_1 _29291_ (.B1(_03732_),
    .Y(_00610_),
    .A1(net5128),
    .A2(_03731_));
 sg13g2_nor4_1 _29292_ (.A(_02877_),
    .B(_02879_),
    .C(_02893_),
    .D(_02909_),
    .Y(_03733_));
 sg13g2_nand3_1 _29293_ (.B(_03719_),
    .C(_03733_),
    .A(_03678_),
    .Y(_03734_));
 sg13g2_o21ai_1 _29294_ (.B1(_02879_),
    .Y(_03735_),
    .A1(_02877_),
    .A2(_03726_));
 sg13g2_nand2_1 _29295_ (.Y(_03736_),
    .A(_03734_),
    .B(_03735_));
 sg13g2_a221oi_1 _29296_ (.B2(net4526),
    .C1(net5128),
    .B1(_03736_),
    .A1(_02879_),
    .Y(_03737_),
    .A2(net4466));
 sg13g2_a21oi_1 _29297_ (.A1(_14522_),
    .A2(net5130),
    .Y(_00611_),
    .B1(_03737_));
 sg13g2_nor2_1 _29298_ (.A(net1184),
    .B(net5292),
    .Y(_03738_));
 sg13g2_a21oi_1 _29299_ (.A1(net4525),
    .A2(_03734_),
    .Y(_03739_),
    .B1(net4466));
 sg13g2_xnor2_1 _29300_ (.Y(_03740_),
    .A(_02882_),
    .B(_03739_));
 sg13g2_a21oi_1 _29301_ (.A1(net5293),
    .A2(_03740_),
    .Y(_00612_),
    .B1(_03738_));
 sg13g2_nor2_1 _29302_ (.A(net1433),
    .B(net5287),
    .Y(_03741_));
 sg13g2_xnor2_1 _29303_ (.Y(_03742_),
    .A(net4526),
    .B(_02881_));
 sg13g2_nand2_1 _29304_ (.Y(_03743_),
    .A(_03739_),
    .B(_03742_));
 sg13g2_xnor2_1 _29305_ (.Y(_03744_),
    .A(_02886_),
    .B(_03743_));
 sg13g2_a21oi_1 _29306_ (.A1(net5287),
    .A2(_03744_),
    .Y(_00613_),
    .B1(_03741_));
 sg13g2_nor2_1 _29307_ (.A(net1272),
    .B(net5292),
    .Y(_03745_));
 sg13g2_and4_1 _29308_ (.A(_02881_),
    .B(_02886_),
    .C(_03719_),
    .D(_03733_),
    .X(_03746_));
 sg13g2_and2_1 _29309_ (.A(_03678_),
    .B(_03746_),
    .X(_03747_));
 sg13g2_a21oi_1 _29310_ (.A1(net4524),
    .A2(_03747_),
    .Y(_03748_),
    .B1(net4482));
 sg13g2_xnor2_1 _29311_ (.Y(_03749_),
    .A(_02898_),
    .B(_03748_));
 sg13g2_a21oi_1 _29312_ (.A1(net5292),
    .A2(_03749_),
    .Y(_00614_),
    .B1(_03745_));
 sg13g2_nor2_1 _29313_ (.A(net1315),
    .B(net5293),
    .Y(_03750_));
 sg13g2_nand3_1 _29314_ (.B(_02898_),
    .C(_03747_),
    .A(_02887_),
    .Y(_03751_));
 sg13g2_a21o_1 _29315_ (.A2(_03747_),
    .A1(_02898_),
    .B1(_02887_),
    .X(_03752_));
 sg13g2_nand2_1 _29316_ (.Y(_03753_),
    .A(_03751_),
    .B(_03752_));
 sg13g2_a22oi_1 _29317_ (.Y(_03754_),
    .B1(_03753_),
    .B2(net4524),
    .A2(net4467),
    .A1(_02888_));
 sg13g2_a21oi_1 _29318_ (.A1(net5292),
    .A2(_03754_),
    .Y(_00615_),
    .B1(_03750_));
 sg13g2_a21oi_1 _29319_ (.A1(net4524),
    .A2(_03751_),
    .Y(_03755_),
    .B1(net4467));
 sg13g2_nor2_1 _29320_ (.A(net1160),
    .B(net5293),
    .Y(_03756_));
 sg13g2_xnor2_1 _29321_ (.Y(_03757_),
    .A(_02874_),
    .B(_03755_));
 sg13g2_a21oi_1 _29322_ (.A1(net5293),
    .A2(_03757_),
    .Y(_00616_),
    .B1(_03756_));
 sg13g2_nor2_1 _29323_ (.A(_02869_),
    .B(_02874_),
    .Y(_03758_));
 sg13g2_nor2b_2 _29324_ (.A(_03751_),
    .B_N(_03758_),
    .Y(_03759_));
 sg13g2_o21ai_1 _29325_ (.B1(_02869_),
    .Y(_03760_),
    .A1(_02874_),
    .A2(_03751_));
 sg13g2_nand2b_1 _29326_ (.Y(_03761_),
    .B(_03760_),
    .A_N(_03759_));
 sg13g2_a221oi_1 _29327_ (.B2(net4524),
    .C1(net5130),
    .B1(_03761_),
    .A1(_02869_),
    .Y(_03762_),
    .A2(net4467));
 sg13g2_a21oi_1 _29328_ (.A1(_14523_),
    .A2(net5130),
    .Y(_00617_),
    .B1(_03762_));
 sg13g2_a21oi_1 _29329_ (.A1(net4527),
    .A2(_03759_),
    .Y(_03763_),
    .B1(net4482));
 sg13g2_xor2_1 _29330_ (.B(_03763_),
    .A(_03168_),
    .X(_03764_));
 sg13g2_nand2_1 _29331_ (.Y(_03765_),
    .A(net1139),
    .B(net5130));
 sg13g2_o21ai_1 _29332_ (.B1(_03765_),
    .Y(_00618_),
    .A1(net5130),
    .A2(_03764_));
 sg13g2_nand2b_1 _29333_ (.Y(_03766_),
    .B(_03167_),
    .A_N(_03759_));
 sg13g2_nor2_1 _29334_ (.A(_03167_),
    .B(_03168_),
    .Y(_03767_));
 sg13g2_nand2_1 _29335_ (.Y(_03768_),
    .A(_03758_),
    .B(_03767_));
 sg13g2_inv_1 _29336_ (.Y(_03769_),
    .A(_03768_));
 sg13g2_nand2_1 _29337_ (.Y(_03770_),
    .A(_03759_),
    .B(_03767_));
 sg13g2_nand3_1 _29338_ (.B(_03766_),
    .C(_03770_),
    .A(_03169_),
    .Y(_03771_));
 sg13g2_a221oi_1 _29339_ (.B2(net4524),
    .C1(net5130),
    .B1(_03771_),
    .A1(_03167_),
    .Y(_03772_),
    .A2(net4467));
 sg13g2_a21oi_1 _29340_ (.A1(_14524_),
    .A2(net5130),
    .Y(_00619_),
    .B1(_03772_));
 sg13g2_a21oi_1 _29341_ (.A1(net4524),
    .A2(_03770_),
    .Y(_03773_),
    .B1(net4467));
 sg13g2_xnor2_1 _29342_ (.Y(_03774_),
    .A(_02872_),
    .B(_03773_));
 sg13g2_nor2_1 _29343_ (.A(net1268),
    .B(net5292),
    .Y(_03775_));
 sg13g2_a21oi_1 _29344_ (.A1(net5292),
    .A2(_03774_),
    .Y(_00620_),
    .B1(_03775_));
 sg13g2_nor2_1 _29345_ (.A(net1213),
    .B(net5292),
    .Y(_03776_));
 sg13g2_xnor2_1 _29346_ (.Y(_03777_),
    .A(net4524),
    .B(_02871_));
 sg13g2_nand2_1 _29347_ (.Y(_03778_),
    .A(_03773_),
    .B(_03777_));
 sg13g2_xnor2_1 _29348_ (.Y(_03779_),
    .A(_03164_),
    .B(_03778_));
 sg13g2_a21oi_1 _29349_ (.A1(net5292),
    .A2(_03779_),
    .Y(_00621_),
    .B1(_03776_));
 sg13g2_nand4_1 _29350_ (.B(_02887_),
    .C(_02898_),
    .A(_02871_),
    .Y(_03780_),
    .D(_03164_));
 sg13g2_inv_1 _29351_ (.Y(_03781_),
    .A(_03780_));
 sg13g2_and4_1 _29352_ (.A(_03603_),
    .B(_03677_),
    .C(_03746_),
    .D(_03781_),
    .X(_03782_));
 sg13g2_and2_1 _29353_ (.A(_03769_),
    .B(_03782_),
    .X(_03783_));
 sg13g2_a21oi_1 _29354_ (.A1(net4524),
    .A2(_03783_),
    .Y(_03784_),
    .B1(net4482));
 sg13g2_xnor2_1 _29355_ (.Y(_03785_),
    .A(_03162_),
    .B(_03784_));
 sg13g2_nand2_1 _29356_ (.Y(_03786_),
    .A(net1304),
    .B(net5132));
 sg13g2_o21ai_1 _29357_ (.B1(_03786_),
    .Y(_00622_),
    .A1(net5132),
    .A2(_03785_));
 sg13g2_nand2_1 _29358_ (.Y(_03787_),
    .A(_03162_),
    .B(_03783_));
 sg13g2_and4_1 _29359_ (.A(_03156_),
    .B(_03162_),
    .C(_03769_),
    .D(_03782_),
    .X(_03788_));
 sg13g2_xnor2_1 _29360_ (.Y(_03789_),
    .A(_03155_),
    .B(_03787_));
 sg13g2_a221oi_1 _29361_ (.B2(net4522),
    .C1(net5132),
    .B1(_03789_),
    .A1(_03155_),
    .Y(_03790_),
    .A2(net4468));
 sg13g2_a21oi_1 _29362_ (.A1(_14525_),
    .A2(net5132),
    .Y(_00623_),
    .B1(_03790_));
 sg13g2_nor2_1 _29363_ (.A(net1316),
    .B(net5290),
    .Y(_03791_));
 sg13g2_a21oi_1 _29364_ (.A1(net4522),
    .A2(_03788_),
    .Y(_03792_),
    .B1(net4480));
 sg13g2_xnor2_1 _29365_ (.Y(_03793_),
    .A(_03159_),
    .B(_03792_));
 sg13g2_a21oi_1 _29366_ (.A1(net5290),
    .A2(_03793_),
    .Y(_00624_),
    .B1(_03791_));
 sg13g2_and3_2 _29367_ (.X(_03794_),
    .A(_03159_),
    .B(_03161_),
    .C(_03788_));
 sg13g2_a21oi_1 _29368_ (.A1(_03159_),
    .A2(_03788_),
    .Y(_03795_),
    .B1(_03161_));
 sg13g2_o21ai_1 _29369_ (.B1(net4523),
    .Y(_03796_),
    .A1(_03794_),
    .A2(_03795_));
 sg13g2_o21ai_1 _29370_ (.B1(_03796_),
    .Y(_03797_),
    .A1(_03161_),
    .A2(net4378));
 sg13g2_mux2_1 _29371_ (.A0(net2040),
    .A1(_03797_),
    .S(net5290),
    .X(_00625_));
 sg13g2_nor2_1 _29372_ (.A(net1373),
    .B(net5291),
    .Y(_03798_));
 sg13g2_a21oi_1 _29373_ (.A1(net4523),
    .A2(_03794_),
    .Y(_03799_),
    .B1(net4480));
 sg13g2_xnor2_1 _29374_ (.Y(_03800_),
    .A(_02864_),
    .B(_03799_));
 sg13g2_a21oi_1 _29375_ (.A1(net5291),
    .A2(_03800_),
    .Y(_00626_),
    .B1(_03798_));
 sg13g2_and3_1 _29376_ (.X(_03801_),
    .A(_02864_),
    .B(_03174_),
    .C(_03794_));
 sg13g2_a21oi_1 _29377_ (.A1(_02864_),
    .A2(_03794_),
    .Y(_03802_),
    .B1(_03174_));
 sg13g2_or2_1 _29378_ (.X(_03803_),
    .B(_03802_),
    .A(_03801_));
 sg13g2_a21oi_1 _29379_ (.A1(net4523),
    .A2(_03803_),
    .Y(_03804_),
    .B1(net5132));
 sg13g2_o21ai_1 _29380_ (.B1(_03804_),
    .Y(_03805_),
    .A1(_03174_),
    .A2(_03302_));
 sg13g2_o21ai_1 _29381_ (.B1(_03805_),
    .Y(_03806_),
    .A1(net2397),
    .A2(net5291));
 sg13g2_inv_1 _29382_ (.Y(_00627_),
    .A(_03806_));
 sg13g2_nor2_1 _29383_ (.A(net1201),
    .B(net5291),
    .Y(_03807_));
 sg13g2_o21ai_1 _29384_ (.B1(net4379),
    .Y(_03808_),
    .A1(net4496),
    .A2(_03801_));
 sg13g2_xor2_1 _29385_ (.B(_03808_),
    .A(_03196_),
    .X(_03809_));
 sg13g2_a21oi_1 _29386_ (.A1(net5291),
    .A2(_03809_),
    .Y(_00628_),
    .B1(_03807_));
 sg13g2_nor2_1 _29387_ (.A(net1138),
    .B(net5291),
    .Y(_03810_));
 sg13g2_xnor2_1 _29388_ (.Y(_03811_),
    .A(net4523),
    .B(_03196_));
 sg13g2_nor2_1 _29389_ (.A(_03808_),
    .B(_03811_),
    .Y(_03812_));
 sg13g2_xor2_1 _29390_ (.B(_03812_),
    .A(_03199_),
    .X(_03813_));
 sg13g2_a21oi_1 _29391_ (.A1(net5291),
    .A2(_03813_),
    .Y(_00629_),
    .B1(_03810_));
 sg13g2_nand3_1 _29392_ (.B(_03174_),
    .C(_03199_),
    .A(_02864_),
    .Y(_03814_));
 sg13g2_nor2_1 _29393_ (.A(_03196_),
    .B(_03814_),
    .Y(_03815_));
 sg13g2_and4_1 _29394_ (.A(_03159_),
    .B(_03161_),
    .C(_03788_),
    .D(_03815_),
    .X(_03816_));
 sg13g2_a21o_1 _29395_ (.A2(_03816_),
    .A1(net4521),
    .B1(net4481),
    .X(_03817_));
 sg13g2_xor2_1 _29396_ (.B(_03817_),
    .A(_03175_),
    .X(_03818_));
 sg13g2_nand2_1 _29397_ (.Y(_03819_),
    .A(net1191),
    .B(net5127));
 sg13g2_o21ai_1 _29398_ (.B1(_03819_),
    .Y(_00630_),
    .A1(net5127),
    .A2(_03818_));
 sg13g2_nor2_1 _29399_ (.A(net1169),
    .B(net5284),
    .Y(_03820_));
 sg13g2_nand3_1 _29400_ (.B(_03200_),
    .C(_03816_),
    .A(_03175_),
    .Y(_03821_));
 sg13g2_a21o_1 _29401_ (.A2(_03816_),
    .A1(_03175_),
    .B1(_03200_),
    .X(_03822_));
 sg13g2_nand2_1 _29402_ (.Y(_03823_),
    .A(_03821_),
    .B(_03822_));
 sg13g2_a22oi_1 _29403_ (.Y(_03824_),
    .B1(_03823_),
    .B2(net4521),
    .A2(net4465),
    .A1(_03201_));
 sg13g2_a21oi_1 _29404_ (.A1(net5284),
    .A2(_03824_),
    .Y(_00631_),
    .B1(_03820_));
 sg13g2_nor2_1 _29405_ (.A(net1277),
    .B(net5284),
    .Y(_03825_));
 sg13g2_a21oi_1 _29406_ (.A1(net4521),
    .A2(_03821_),
    .Y(_03826_),
    .B1(net4464));
 sg13g2_xnor2_1 _29407_ (.Y(_03827_),
    .A(_02862_),
    .B(_03826_));
 sg13g2_a21oi_1 _29408_ (.A1(net5284),
    .A2(_03827_),
    .Y(_00632_),
    .B1(_03825_));
 sg13g2_nor2_1 _29409_ (.A(_02862_),
    .B(_03821_),
    .Y(_03828_));
 sg13g2_nand2b_1 _29410_ (.Y(_03829_),
    .B(_03828_),
    .A_N(_02860_));
 sg13g2_xor2_1 _29411_ (.B(_03828_),
    .A(_02860_),
    .X(_03830_));
 sg13g2_a221oi_1 _29412_ (.B2(net4521),
    .C1(net5127),
    .B1(_03830_),
    .A1(_02860_),
    .Y(_03831_),
    .A2(net4464));
 sg13g2_a21oi_1 _29413_ (.A1(_14526_),
    .A2(net5127),
    .Y(_00633_),
    .B1(_03831_));
 sg13g2_nor2_1 _29414_ (.A(net1410),
    .B(net5284),
    .Y(_03832_));
 sg13g2_a21oi_1 _29415_ (.A1(net4521),
    .A2(_03829_),
    .Y(_03833_),
    .B1(net4464));
 sg13g2_xnor2_1 _29416_ (.Y(_03834_),
    .A(_03191_),
    .B(_03833_));
 sg13g2_a21oi_1 _29417_ (.A1(net5284),
    .A2(_03834_),
    .Y(_00634_),
    .B1(_03832_));
 sg13g2_nor4_1 _29418_ (.A(_02860_),
    .B(_02862_),
    .C(_03190_),
    .D(_03191_),
    .Y(_03835_));
 sg13g2_nand4_1 _29419_ (.B(_03200_),
    .C(_03816_),
    .A(_03175_),
    .Y(_03836_),
    .D(_03835_));
 sg13g2_o21ai_1 _29420_ (.B1(_03190_),
    .Y(_03837_),
    .A1(_03191_),
    .A2(_03829_));
 sg13g2_nand2_1 _29421_ (.Y(_03838_),
    .A(_03836_),
    .B(_03837_));
 sg13g2_a221oi_1 _29422_ (.B2(net4528),
    .C1(net5127),
    .B1(_03838_),
    .A1(_03190_),
    .Y(_03839_),
    .A2(net4465));
 sg13g2_a21oi_1 _29423_ (.A1(_14527_),
    .A2(net5127),
    .Y(_00635_),
    .B1(_03839_));
 sg13g2_a21o_1 _29424_ (.A2(_03836_),
    .A1(net4520),
    .B1(net4463),
    .X(_03840_));
 sg13g2_xnor2_1 _29425_ (.Y(_03841_),
    .A(_02854_),
    .B(_03840_));
 sg13g2_nand2_1 _29426_ (.Y(_03842_),
    .A(net1333),
    .B(net5125));
 sg13g2_o21ai_1 _29427_ (.B1(_03842_),
    .Y(_00636_),
    .A1(net5125),
    .A2(_03841_));
 sg13g2_nor2_1 _29428_ (.A(net1418),
    .B(net5285),
    .Y(_03843_));
 sg13g2_xnor2_1 _29429_ (.Y(_03844_),
    .A(net4495),
    .B(_02854_));
 sg13g2_nor2_1 _29430_ (.A(_03840_),
    .B(_03844_),
    .Y(_03845_));
 sg13g2_xnor2_1 _29431_ (.Y(_03846_),
    .A(_03194_),
    .B(_03845_));
 sg13g2_a21oi_1 _29432_ (.A1(net5284),
    .A2(_03846_),
    .Y(_00637_),
    .B1(_03843_));
 sg13g2_nand2b_1 _29433_ (.Y(_03847_),
    .B(_02854_),
    .A_N(_03194_));
 sg13g2_or2_1 _29434_ (.X(_03848_),
    .B(_03847_),
    .A(_03836_));
 sg13g2_a21oi_1 _29435_ (.A1(net4520),
    .A2(_03848_),
    .Y(_03849_),
    .B1(net4465));
 sg13g2_xor2_1 _29436_ (.B(_03849_),
    .A(_03186_),
    .X(_03850_));
 sg13g2_nand2_1 _29437_ (.Y(_03851_),
    .A(net1187),
    .B(net5126));
 sg13g2_o21ai_1 _29438_ (.B1(_03851_),
    .Y(_00638_),
    .A1(net5125),
    .A2(_03850_));
 sg13g2_nand2_1 _29439_ (.Y(_03852_),
    .A(_03185_),
    .B(_03186_));
 sg13g2_or2_1 _29440_ (.X(_03853_),
    .B(_03852_),
    .A(_03848_));
 sg13g2_nand2b_1 _29441_ (.Y(_03854_),
    .B(_03848_),
    .A_N(_03185_));
 sg13g2_nand3_1 _29442_ (.B(_03853_),
    .C(_03854_),
    .A(_03187_),
    .Y(_03855_));
 sg13g2_a21oi_1 _29443_ (.A1(net4520),
    .A2(_03855_),
    .Y(_03856_),
    .B1(net5126));
 sg13g2_o21ai_1 _29444_ (.B1(_03856_),
    .Y(_03857_),
    .A1(_03185_),
    .A2(net4378));
 sg13g2_o21ai_1 _29445_ (.B1(_03857_),
    .Y(_03858_),
    .A1(net3165),
    .A2(net5283));
 sg13g2_inv_1 _29446_ (.Y(_00639_),
    .A(_03858_));
 sg13g2_nor2_1 _29447_ (.A(net1497),
    .B(net5281),
    .Y(_03859_));
 sg13g2_o21ai_1 _29448_ (.B1(net4471),
    .Y(_03860_),
    .A1(net4495),
    .A2(_03853_));
 sg13g2_xor2_1 _29449_ (.B(_03860_),
    .A(_02852_),
    .X(_03861_));
 sg13g2_a21oi_1 _29450_ (.A1(net5281),
    .A2(_03861_),
    .Y(_00640_),
    .B1(_03859_));
 sg13g2_nor2_1 _29451_ (.A(net1624),
    .B(net5283),
    .Y(_03862_));
 sg13g2_o21ai_1 _29452_ (.B1(_03860_),
    .Y(_03863_),
    .A1(net4495),
    .A2(_02852_));
 sg13g2_xnor2_1 _29453_ (.Y(_03864_),
    .A(_03182_),
    .B(_03863_));
 sg13g2_a21oi_1 _29454_ (.A1(net5283),
    .A2(_03864_),
    .Y(_00641_),
    .B1(_03862_));
 sg13g2_nand2_1 _29455_ (.Y(_03865_),
    .A(_02852_),
    .B(_03182_));
 sg13g2_or4_1 _29456_ (.A(_03836_),
    .B(_03847_),
    .C(_03852_),
    .D(_03865_),
    .X(_03866_));
 sg13g2_a21oi_1 _29457_ (.A1(net4519),
    .A2(_03866_),
    .Y(_03867_),
    .B1(net4463));
 sg13g2_xnor2_1 _29458_ (.Y(_03868_),
    .A(_03180_),
    .B(_03867_));
 sg13g2_nand2_1 _29459_ (.Y(_03869_),
    .A(net1198),
    .B(net5124));
 sg13g2_o21ai_1 _29460_ (.B1(_03869_),
    .Y(_00642_),
    .A1(net5124),
    .A2(_03868_));
 sg13g2_nand2b_1 _29461_ (.Y(_03870_),
    .B(_03179_),
    .A_N(_02838_));
 sg13g2_or2_1 _29462_ (.X(_03871_),
    .B(_03870_),
    .A(_03866_));
 sg13g2_o21ai_1 _29463_ (.B1(_02838_),
    .Y(_03872_),
    .A1(_03180_),
    .A2(_03866_));
 sg13g2_nand2_1 _29464_ (.Y(_03873_),
    .A(_03871_),
    .B(_03872_));
 sg13g2_a221oi_1 _29465_ (.B2(net4519),
    .C1(net5124),
    .B1(_03873_),
    .A1(_02838_),
    .Y(_03874_),
    .A2(net4463));
 sg13g2_a21oi_1 _29466_ (.A1(_14528_),
    .A2(net5125),
    .Y(_00643_),
    .B1(_03874_));
 sg13g2_nor2_1 _29467_ (.A(net2141),
    .B(net5282),
    .Y(_03875_));
 sg13g2_a21oi_1 _29468_ (.A1(net4519),
    .A2(_03871_),
    .Y(_03876_),
    .B1(net4463));
 sg13g2_xnor2_1 _29469_ (.Y(_03877_),
    .A(_02841_),
    .B(_03876_));
 sg13g2_a21oi_1 _29470_ (.A1(net5282),
    .A2(_03877_),
    .Y(_00644_),
    .B1(_03875_));
 sg13g2_nor2_1 _29471_ (.A(net1831),
    .B(net5282),
    .Y(_03878_));
 sg13g2_xnor2_1 _29472_ (.Y(_03879_),
    .A(net4495),
    .B(_02841_));
 sg13g2_nand2_1 _29473_ (.Y(_03880_),
    .A(_03876_),
    .B(_03879_));
 sg13g2_xor2_1 _29474_ (.B(_03880_),
    .A(_02845_),
    .X(_03881_));
 sg13g2_a21oi_1 _29475_ (.A1(net5282),
    .A2(_03881_),
    .Y(_00645_),
    .B1(_03878_));
 sg13g2_nor2_1 _29476_ (.A(net2032),
    .B(net5282),
    .Y(_03882_));
 sg13g2_or2_1 _29477_ (.X(_03883_),
    .B(_02845_),
    .A(_02841_));
 sg13g2_or2_1 _29478_ (.X(_03884_),
    .B(_03883_),
    .A(_03871_));
 sg13g2_a21oi_1 _29479_ (.A1(net4519),
    .A2(_03884_),
    .Y(_03885_),
    .B1(net4463));
 sg13g2_xnor2_1 _29480_ (.Y(_03886_),
    .A(_02842_),
    .B(_03885_));
 sg13g2_a21oi_1 _29481_ (.A1(net5282),
    .A2(_03886_),
    .Y(_00646_),
    .B1(_03882_));
 sg13g2_nor2_1 _29482_ (.A(_02842_),
    .B(_03884_),
    .Y(_03887_));
 sg13g2_nand2_1 _29483_ (.Y(_03888_),
    .A(_02848_),
    .B(_03887_));
 sg13g2_xnor2_1 _29484_ (.Y(_03889_),
    .A(_02848_),
    .B(_03887_));
 sg13g2_a221oi_1 _29485_ (.B2(net4519),
    .C1(net5124),
    .B1(_03889_),
    .A1(_02847_),
    .Y(_03890_),
    .A2(net4463));
 sg13g2_a21oi_1 _29486_ (.A1(_14529_),
    .A2(net5124),
    .Y(_00647_),
    .B1(_03890_));
 sg13g2_nor2_1 _29487_ (.A(net2123),
    .B(net5277),
    .Y(_03891_));
 sg13g2_a21oi_1 _29488_ (.A1(net4519),
    .A2(_03888_),
    .Y(_03892_),
    .B1(net4463));
 sg13g2_xor2_1 _29489_ (.B(_03892_),
    .A(_02828_),
    .X(_03893_));
 sg13g2_a21oi_1 _29490_ (.A1(net5277),
    .A2(_03893_),
    .Y(_00648_),
    .B1(_03891_));
 sg13g2_nand2_1 _29491_ (.Y(_03894_),
    .A(_02830_),
    .B(net4463));
 sg13g2_nand2_2 _29492_ (.Y(_03895_),
    .A(_02828_),
    .B(_02830_));
 sg13g2_o21ai_1 _29493_ (.B1(net4519),
    .Y(_03896_),
    .A1(_03888_),
    .A2(_03895_));
 sg13g2_a21oi_1 _29494_ (.A1(_02848_),
    .A2(_03887_),
    .Y(_03897_),
    .B1(_02830_));
 sg13g2_nor3_1 _29495_ (.A(_02831_),
    .B(_03896_),
    .C(_03897_),
    .Y(_03898_));
 sg13g2_o21ai_1 _29496_ (.B1(net5281),
    .Y(_03899_),
    .A1(net4519),
    .A2(_03895_));
 sg13g2_nor3_1 _29497_ (.A(net4481),
    .B(_03898_),
    .C(_03899_),
    .Y(_03900_));
 sg13g2_a22oi_1 _29498_ (.Y(_03901_),
    .B1(_03894_),
    .B2(_03900_),
    .A2(net5124),
    .A1(net2487));
 sg13g2_inv_1 _29499_ (.Y(_00649_),
    .A(_03901_));
 sg13g2_nor2_1 _29500_ (.A(net1772),
    .B(net5282),
    .Y(_03902_));
 sg13g2_nand2_1 _29501_ (.Y(_03903_),
    .A(net4378),
    .B(_03896_));
 sg13g2_xnor2_1 _29502_ (.Y(_03904_),
    .A(_02697_),
    .B(_03903_));
 sg13g2_a21oi_1 _29503_ (.A1(net5282),
    .A2(_03904_),
    .Y(_00650_),
    .B1(_03902_));
 sg13g2_o21ai_1 _29504_ (.B1(_02696_),
    .Y(_03905_),
    .A1(_03888_),
    .A2(_03895_));
 sg13g2_nor4_1 _29505_ (.A(_02696_),
    .B(_02842_),
    .C(_02847_),
    .D(_03895_),
    .Y(_03906_));
 sg13g2_nand2_1 _29506_ (.Y(_03907_),
    .A(_02697_),
    .B(_03906_));
 sg13g2_or2_1 _29507_ (.X(_03908_),
    .B(_03907_),
    .A(_03884_));
 sg13g2_nand3_1 _29508_ (.B(_03905_),
    .C(_03908_),
    .A(_02698_),
    .Y(_03909_));
 sg13g2_a221oi_1 _29509_ (.B2(net4516),
    .C1(net5122),
    .B1(_03909_),
    .A1(_02696_),
    .Y(_03910_),
    .A2(net4462));
 sg13g2_a21oi_1 _29510_ (.A1(_14530_),
    .A2(net5122),
    .Y(_00651_),
    .B1(_03910_));
 sg13g2_nor2_1 _29511_ (.A(net1628),
    .B(net5276),
    .Y(_03911_));
 sg13g2_a21oi_1 _29512_ (.A1(net4516),
    .A2(_03908_),
    .Y(_03912_),
    .B1(net4462));
 sg13g2_xnor2_1 _29513_ (.Y(_03913_),
    .A(_02821_),
    .B(_03912_));
 sg13g2_a21oi_1 _29514_ (.A1(net5277),
    .A2(_03913_),
    .Y(_00652_),
    .B1(_03911_));
 sg13g2_nor2_1 _29515_ (.A(net1645),
    .B(net5276),
    .Y(_03914_));
 sg13g2_xnor2_1 _29516_ (.Y(_03915_),
    .A(net4494),
    .B(_02821_));
 sg13g2_nand2_1 _29517_ (.Y(_03916_),
    .A(_03912_),
    .B(_03915_));
 sg13g2_xnor2_1 _29518_ (.Y(_03917_),
    .A(_03208_),
    .B(_03916_));
 sg13g2_a21oi_1 _29519_ (.A1(net5276),
    .A2(_03917_),
    .Y(_00653_),
    .B1(_03914_));
 sg13g2_nor2b_1 _29520_ (.A(_02821_),
    .B_N(_03208_),
    .Y(_03918_));
 sg13g2_nor2b_1 _29521_ (.A(_03908_),
    .B_N(_03918_),
    .Y(_03919_));
 sg13g2_a21oi_1 _29522_ (.A1(net4516),
    .A2(_03919_),
    .Y(_03920_),
    .B1(net4478));
 sg13g2_xor2_1 _29523_ (.B(_03920_),
    .A(_02822_),
    .X(_03921_));
 sg13g2_nor2_1 _29524_ (.A(net1730),
    .B(net5276),
    .Y(_03922_));
 sg13g2_a21oi_1 _29525_ (.A1(net5276),
    .A2(_03921_),
    .Y(_00654_),
    .B1(_03922_));
 sg13g2_nor2_1 _29526_ (.A(net2052),
    .B(net5278),
    .Y(_03923_));
 sg13g2_nand2b_1 _29527_ (.Y(_03924_),
    .B(_03919_),
    .A_N(_02822_));
 sg13g2_nand2b_1 _29528_ (.Y(_03925_),
    .B(_02691_),
    .A_N(_03924_));
 sg13g2_xnor2_1 _29529_ (.Y(_03926_),
    .A(_02690_),
    .B(_03924_));
 sg13g2_a22oi_1 _29530_ (.Y(_03927_),
    .B1(_03926_),
    .B2(net4516),
    .A2(net4462),
    .A1(_02690_));
 sg13g2_a21oi_1 _29531_ (.A1(net5276),
    .A2(_03927_),
    .Y(_00655_),
    .B1(_03923_));
 sg13g2_nor2_1 _29532_ (.A(net2043),
    .B(net5278),
    .Y(_03928_));
 sg13g2_a21oi_1 _29533_ (.A1(net4516),
    .A2(_03925_),
    .Y(_03929_),
    .B1(net4462));
 sg13g2_xnor2_1 _29534_ (.Y(_03930_),
    .A(_03228_),
    .B(_03929_));
 sg13g2_a21oi_1 _29535_ (.A1(net5278),
    .A2(_03930_),
    .Y(_00656_),
    .B1(_03928_));
 sg13g2_or2_1 _29536_ (.X(_03931_),
    .B(_03228_),
    .A(_03226_));
 sg13g2_nor2_1 _29537_ (.A(_02690_),
    .B(_03931_),
    .Y(_03932_));
 sg13g2_nor2_1 _29538_ (.A(_03925_),
    .B(_03931_),
    .Y(_03933_));
 sg13g2_o21ai_1 _29539_ (.B1(_03226_),
    .Y(_03934_),
    .A1(_03228_),
    .A2(_03925_));
 sg13g2_nand2b_1 _29540_ (.Y(_03935_),
    .B(_03934_),
    .A_N(_03933_));
 sg13g2_a221oi_1 _29541_ (.B2(net4516),
    .C1(net5121),
    .B1(_03935_),
    .A1(_03226_),
    .Y(_03936_),
    .A2(net4462));
 sg13g2_a21oi_1 _29542_ (.A1(_14531_),
    .A2(net5121),
    .Y(_00657_),
    .B1(_03936_));
 sg13g2_nor2_1 _29543_ (.A(net1189),
    .B(net5278),
    .Y(_03937_));
 sg13g2_a21oi_1 _29544_ (.A1(net4518),
    .A2(_03933_),
    .Y(_03938_),
    .B1(net4478));
 sg13g2_xnor2_1 _29545_ (.Y(_03939_),
    .A(_02799_),
    .B(_03938_));
 sg13g2_a21oi_1 _29546_ (.A1(net5278),
    .A2(_03939_),
    .Y(_00658_),
    .B1(_03937_));
 sg13g2_nand3_1 _29547_ (.B(_03241_),
    .C(_03933_),
    .A(_02799_),
    .Y(_03940_));
 sg13g2_a21o_1 _29548_ (.A2(_03933_),
    .A1(_02799_),
    .B1(_03241_),
    .X(_03941_));
 sg13g2_nand2_1 _29549_ (.Y(_03942_),
    .A(_03940_),
    .B(_03941_));
 sg13g2_a21oi_1 _29550_ (.A1(net4516),
    .A2(_03942_),
    .Y(_03943_),
    .B1(net5121));
 sg13g2_o21ai_1 _29551_ (.B1(_03943_),
    .Y(_03944_),
    .A1(_03241_),
    .A2(net4379));
 sg13g2_o21ai_1 _29552_ (.B1(_03944_),
    .Y(_03945_),
    .A1(net2762),
    .A2(net5279));
 sg13g2_inv_1 _29553_ (.Y(_00659_),
    .A(_03945_));
 sg13g2_nor2_1 _29554_ (.A(net1338),
    .B(net5279),
    .Y(_03946_));
 sg13g2_a21oi_1 _29555_ (.A1(net4517),
    .A2(_03940_),
    .Y(_03947_),
    .B1(net4462));
 sg13g2_xor2_1 _29556_ (.B(_03947_),
    .A(_02679_),
    .X(_03948_));
 sg13g2_a21oi_1 _29557_ (.A1(net5279),
    .A2(_03948_),
    .Y(_00660_),
    .B1(_03946_));
 sg13g2_nor2_1 _29558_ (.A(net1305),
    .B(net5279),
    .Y(_03949_));
 sg13g2_xnor2_1 _29559_ (.Y(_03950_),
    .A(net4517),
    .B(_02679_));
 sg13g2_nand2_1 _29560_ (.Y(_03951_),
    .A(_03947_),
    .B(_03950_));
 sg13g2_xor2_1 _29561_ (.B(_03951_),
    .A(_02676_),
    .X(_03952_));
 sg13g2_a21oi_1 _29562_ (.A1(net5279),
    .A2(_03952_),
    .Y(_00661_),
    .B1(_03949_));
 sg13g2_nor2b_1 _29563_ (.A(_02676_),
    .B_N(_02679_),
    .Y(_03953_));
 sg13g2_nor4_1 _29564_ (.A(_02798_),
    .B(_02822_),
    .C(_03242_),
    .D(_03907_),
    .Y(_03954_));
 sg13g2_nand4_1 _29565_ (.B(_03932_),
    .C(_03953_),
    .A(_03918_),
    .Y(_03955_),
    .D(_03954_));
 sg13g2_nor2_2 _29566_ (.A(_03884_),
    .B(_03955_),
    .Y(_03956_));
 sg13g2_or4_1 _29567_ (.A(_03866_),
    .B(_03870_),
    .C(_03883_),
    .D(_03955_),
    .X(_03957_));
 sg13g2_a21oi_1 _29568_ (.A1(net4517),
    .A2(_03956_),
    .Y(_03958_),
    .B1(net4477));
 sg13g2_xnor2_1 _29569_ (.Y(_03959_),
    .A(_02849_),
    .B(_03958_));
 sg13g2_nor2_1 _29570_ (.A(net1190),
    .B(net5279),
    .Y(_03960_));
 sg13g2_a21oi_1 _29571_ (.A1(net5279),
    .A2(_03959_),
    .Y(_00662_),
    .B1(_03960_));
 sg13g2_nand2_1 _29572_ (.Y(_03961_),
    .A(_02849_),
    .B(_03956_));
 sg13g2_nor2b_1 _29573_ (.A(_02833_),
    .B_N(_02849_),
    .Y(_03962_));
 sg13g2_nand2_1 _29574_ (.Y(_03963_),
    .A(_03956_),
    .B(_03962_));
 sg13g2_xnor2_1 _29575_ (.Y(_03964_),
    .A(_02833_),
    .B(_03961_));
 sg13g2_a221oi_1 _29576_ (.B2(net4517),
    .C1(net5120),
    .B1(_03964_),
    .A1(_02833_),
    .Y(_03965_),
    .A2(net4469));
 sg13g2_a21oi_1 _29577_ (.A1(_14532_),
    .A2(net5123),
    .Y(_00663_),
    .B1(_03965_));
 sg13g2_nor2_1 _29578_ (.A(net1202),
    .B(net5271),
    .Y(_03966_));
 sg13g2_a21oi_1 _29579_ (.A1(net4514),
    .A2(_03963_),
    .Y(_03967_),
    .B1(net4460));
 sg13g2_xor2_1 _29580_ (.B(_03967_),
    .A(_02707_),
    .X(_03968_));
 sg13g2_a21oi_1 _29581_ (.A1(net5271),
    .A2(_03968_),
    .Y(_00664_),
    .B1(_03966_));
 sg13g2_nand2_1 _29582_ (.Y(_03969_),
    .A(net1165),
    .B(net5118));
 sg13g2_and2_1 _29583_ (.A(_02704_),
    .B(_02707_),
    .X(_03970_));
 sg13g2_nor2b_1 _29584_ (.A(_03963_),
    .B_N(_03970_),
    .Y(_03971_));
 sg13g2_nor2_1 _29585_ (.A(net4493),
    .B(_03971_),
    .Y(_03972_));
 sg13g2_nand2b_1 _29586_ (.Y(_03973_),
    .B(_03963_),
    .A_N(_02704_));
 sg13g2_nand3_1 _29587_ (.B(_03972_),
    .C(_03973_),
    .A(_02708_),
    .Y(_03974_));
 sg13g2_a21oi_1 _29588_ (.A1(net4493),
    .A2(_02704_),
    .Y(_03975_),
    .B1(net5119));
 sg13g2_nand2_1 _29589_ (.Y(_03976_),
    .A(_03974_),
    .B(_03975_));
 sg13g2_o21ai_1 _29590_ (.B1(_03969_),
    .Y(_00665_),
    .A1(net4479),
    .A2(_03976_));
 sg13g2_nor2_1 _29591_ (.A(net4461),
    .B(_03972_),
    .Y(_03977_));
 sg13g2_xnor2_1 _29592_ (.Y(_03978_),
    .A(_02713_),
    .B(_03977_));
 sg13g2_nor2_1 _29593_ (.A(net1761),
    .B(net5271),
    .Y(_03979_));
 sg13g2_a21oi_1 _29594_ (.A1(net5271),
    .A2(_03978_),
    .Y(_00666_),
    .B1(_03979_));
 sg13g2_nor2_1 _29595_ (.A(net1319),
    .B(net5271),
    .Y(_03980_));
 sg13g2_nand2_1 _29596_ (.Y(_03981_),
    .A(_02712_),
    .B(_03971_));
 sg13g2_xnor2_1 _29597_ (.Y(_03982_),
    .A(_03216_),
    .B(_03981_));
 sg13g2_a22oi_1 _29598_ (.Y(_03983_),
    .B1(_03982_),
    .B2(net4513),
    .A2(net4460),
    .A1(_03216_));
 sg13g2_a21oi_1 _29599_ (.A1(net5272),
    .A2(_03983_),
    .Y(_00667_),
    .B1(_03980_));
 sg13g2_o21ai_1 _29600_ (.B1(net4513),
    .Y(_03984_),
    .A1(_03216_),
    .A2(_03981_));
 sg13g2_nor2b_1 _29601_ (.A(net4460),
    .B_N(_03984_),
    .Y(_03985_));
 sg13g2_xor2_1 _29602_ (.B(_03985_),
    .A(_03221_),
    .X(_03986_));
 sg13g2_nor2_1 _29603_ (.A(net1220),
    .B(net5271),
    .Y(_03987_));
 sg13g2_a21oi_1 _29604_ (.A1(net5271),
    .A2(_03986_),
    .Y(_00668_),
    .B1(_03987_));
 sg13g2_nor2_1 _29605_ (.A(net1335),
    .B(net5272),
    .Y(_03988_));
 sg13g2_xnor2_1 _29606_ (.Y(_03989_),
    .A(net4513),
    .B(_03221_));
 sg13g2_nand2_1 _29607_ (.Y(_03990_),
    .A(_03985_),
    .B(_03989_));
 sg13g2_xor2_1 _29608_ (.B(_03990_),
    .A(_03214_),
    .X(_03991_));
 sg13g2_a21oi_1 _29609_ (.A1(net5271),
    .A2(_03991_),
    .Y(_00669_),
    .B1(_03988_));
 sg13g2_nand3_1 _29610_ (.B(_03962_),
    .C(_03970_),
    .A(_03221_),
    .Y(_03992_));
 sg13g2_nor4_1 _29611_ (.A(_02713_),
    .B(_03214_),
    .C(_03216_),
    .D(_03992_),
    .Y(_03993_));
 sg13g2_nand2_1 _29612_ (.Y(_03994_),
    .A(_03956_),
    .B(_03993_));
 sg13g2_a21oi_1 _29613_ (.A1(net4513),
    .A2(_03994_),
    .Y(_03995_),
    .B1(net4460));
 sg13g2_xnor2_1 _29614_ (.Y(_03996_),
    .A(_03217_),
    .B(_03995_));
 sg13g2_nand2_1 _29615_ (.Y(_03997_),
    .A(net1107),
    .B(net5118));
 sg13g2_o21ai_1 _29616_ (.B1(_03997_),
    .Y(_00670_),
    .A1(net5118),
    .A2(_03996_));
 sg13g2_nor2_1 _29617_ (.A(_03217_),
    .B(_03223_),
    .Y(_03998_));
 sg13g2_nand3_1 _29618_ (.B(_03993_),
    .C(_03998_),
    .A(_03956_),
    .Y(_03999_));
 sg13g2_o21ai_1 _29619_ (.B1(_03223_),
    .Y(_04000_),
    .A1(_03217_),
    .A2(_03994_));
 sg13g2_nand2_1 _29620_ (.Y(_04001_),
    .A(_03999_),
    .B(_04000_));
 sg13g2_a221oi_1 _29621_ (.B2(net4513),
    .C1(net5118),
    .B1(_04001_),
    .A1(_03223_),
    .Y(_04002_),
    .A2(net4460));
 sg13g2_a21oi_1 _29622_ (.A1(_14533_),
    .A2(net5118),
    .Y(_00671_),
    .B1(_04002_));
 sg13g2_nor2_1 _29623_ (.A(net1221),
    .B(net5270),
    .Y(_04003_));
 sg13g2_a21oi_1 _29624_ (.A1(net4514),
    .A2(_03999_),
    .Y(_04004_),
    .B1(net4460));
 sg13g2_xor2_1 _29625_ (.B(_04004_),
    .A(_02816_),
    .X(_04005_));
 sg13g2_a21oi_1 _29626_ (.A1(net5270),
    .A2(_04005_),
    .Y(_00672_),
    .B1(_04003_));
 sg13g2_nor2b_1 _29627_ (.A(_03999_),
    .B_N(_02816_),
    .Y(_04006_));
 sg13g2_and2_1 _29628_ (.A(_02722_),
    .B(_02816_),
    .X(_04007_));
 sg13g2_nor2b_1 _29629_ (.A(_03999_),
    .B_N(_04007_),
    .Y(_04008_));
 sg13g2_xnor2_1 _29630_ (.Y(_04009_),
    .A(_02722_),
    .B(_04006_));
 sg13g2_a21oi_1 _29631_ (.A1(net4513),
    .A2(_04009_),
    .Y(_04010_),
    .B1(net5118));
 sg13g2_o21ai_1 _29632_ (.B1(_04010_),
    .Y(_04011_),
    .A1(_02722_),
    .A2(net4379));
 sg13g2_o21ai_1 _29633_ (.B1(_04011_),
    .Y(_04012_),
    .A1(net2728),
    .A2(net5270));
 sg13g2_inv_1 _29634_ (.Y(_00673_),
    .A(_04012_));
 sg13g2_nor2_1 _29635_ (.A(net1256),
    .B(net5270),
    .Y(_04013_));
 sg13g2_a21oi_1 _29636_ (.A1(net4513),
    .A2(_04008_),
    .Y(_04014_),
    .B1(net4479));
 sg13g2_xnor2_1 _29637_ (.Y(_04015_),
    .A(_02792_),
    .B(_04014_));
 sg13g2_a21oi_1 _29638_ (.A1(net5270),
    .A2(_04015_),
    .Y(_00674_),
    .B1(_04013_));
 sg13g2_and2_1 _29639_ (.A(_02792_),
    .B(_04008_),
    .X(_04016_));
 sg13g2_nand2_1 _29640_ (.Y(_04017_),
    .A(_02786_),
    .B(_04016_));
 sg13g2_nor2_1 _29641_ (.A(net4493),
    .B(_04017_),
    .Y(_04018_));
 sg13g2_nand2b_1 _29642_ (.Y(_04019_),
    .B(net4460),
    .A_N(_02786_));
 sg13g2_nor3_1 _29643_ (.A(net4493),
    .B(_02786_),
    .C(_04016_),
    .Y(_04020_));
 sg13g2_nor3_1 _29644_ (.A(net5118),
    .B(_04018_),
    .C(_04020_),
    .Y(_04021_));
 sg13g2_a22oi_1 _29645_ (.Y(_00675_),
    .B1(_04019_),
    .B2(_04021_),
    .A2(net5118),
    .A1(_14534_));
 sg13g2_nor2_1 _29646_ (.A(net1254),
    .B(net5270),
    .Y(_04022_));
 sg13g2_a21oi_1 _29647_ (.A1(net4514),
    .A2(_04017_),
    .Y(_04023_),
    .B1(net4460));
 sg13g2_xnor2_1 _29648_ (.Y(_04024_),
    .A(_02789_),
    .B(_04023_));
 sg13g2_a21oi_1 _29649_ (.A1(net5272),
    .A2(_04024_),
    .Y(_00676_),
    .B1(_04022_));
 sg13g2_nor2_1 _29650_ (.A(net1322),
    .B(net5270),
    .Y(_04025_));
 sg13g2_o21ai_1 _29651_ (.B1(net4379),
    .Y(_04026_),
    .A1(_02793_),
    .A2(_04018_));
 sg13g2_a21oi_1 _29652_ (.A1(net4513),
    .A2(_02789_),
    .Y(_04027_),
    .B1(_04026_));
 sg13g2_xnor2_1 _29653_ (.Y(_04028_),
    .A(_03236_),
    .B(_04027_));
 sg13g2_a21oi_1 _29654_ (.A1(net5270),
    .A2(_04028_),
    .Y(_00677_),
    .B1(_04025_));
 sg13g2_nand4_1 _29655_ (.B(_03993_),
    .C(_03998_),
    .A(_02790_),
    .Y(_04029_),
    .D(_04007_));
 sg13g2_nand2_1 _29656_ (.Y(_04030_),
    .A(_02786_),
    .B(_02792_));
 sg13g2_or2_1 _29657_ (.X(_04031_),
    .B(_04030_),
    .A(_03236_));
 sg13g2_nor3_2 _29658_ (.A(_03957_),
    .B(_04029_),
    .C(_04031_),
    .Y(_04032_));
 sg13g2_or3_1 _29659_ (.A(_03957_),
    .B(_04029_),
    .C(_04031_),
    .X(_04033_));
 sg13g2_o21ai_1 _29660_ (.B1(net4471),
    .Y(_04034_),
    .A1(net4493),
    .A2(_04033_));
 sg13g2_xnor2_1 _29661_ (.Y(_04035_),
    .A(_02835_),
    .B(_04034_));
 sg13g2_nand2_1 _29662_ (.Y(_04036_),
    .A(net1088),
    .B(net5119));
 sg13g2_o21ai_1 _29663_ (.B1(_04036_),
    .Y(_00678_),
    .A1(net5119),
    .A2(_04035_));
 sg13g2_nor2_1 _29664_ (.A(net1232),
    .B(net5269),
    .Y(_04037_));
 sg13g2_nor2_1 _29665_ (.A(_02835_),
    .B(_04033_),
    .Y(_04038_));
 sg13g2_nor3_1 _29666_ (.A(_02824_),
    .B(_02835_),
    .C(_04033_),
    .Y(_04039_));
 sg13g2_xor2_1 _29667_ (.B(_04038_),
    .A(_02824_),
    .X(_04040_));
 sg13g2_a22oi_1 _29668_ (.Y(_04041_),
    .B1(_04040_),
    .B2(net4515),
    .A2(net4461),
    .A1(_02824_));
 sg13g2_a21oi_1 _29669_ (.A1(net5269),
    .A2(_04041_),
    .Y(_00679_),
    .B1(_04037_));
 sg13g2_a21oi_1 _29670_ (.A1(net4515),
    .A2(_04039_),
    .Y(_04042_),
    .B1(net4479));
 sg13g2_xnor2_1 _29671_ (.Y(_04043_),
    .A(_02701_),
    .B(_04042_));
 sg13g2_nor2_1 _29672_ (.A(net1156),
    .B(net5269),
    .Y(_04044_));
 sg13g2_a21oi_1 _29673_ (.A1(net5269),
    .A2(_04043_),
    .Y(_00680_),
    .B1(_04044_));
 sg13g2_nor2_1 _29674_ (.A(_03230_),
    .B(net4379),
    .Y(_04045_));
 sg13g2_nor2_1 _29675_ (.A(_02824_),
    .B(_02835_),
    .Y(_04046_));
 sg13g2_nand2_1 _29676_ (.Y(_04047_),
    .A(_02701_),
    .B(_04039_));
 sg13g2_nand3_1 _29677_ (.B(_03230_),
    .C(_04046_),
    .A(_02701_),
    .Y(_04048_));
 sg13g2_xnor2_1 _29678_ (.Y(_04049_),
    .A(_03230_),
    .B(_04047_));
 sg13g2_o21ai_1 _29679_ (.B1(net5267),
    .Y(_04050_),
    .A1(net4493),
    .A2(_04049_));
 sg13g2_nor2_1 _29680_ (.A(_04045_),
    .B(_04050_),
    .Y(_04051_));
 sg13g2_a21oi_1 _29681_ (.A1(_14535_),
    .A2(net5119),
    .Y(_00681_),
    .B1(_04051_));
 sg13g2_nor2_1 _29682_ (.A(net1229),
    .B(net5268),
    .Y(_04052_));
 sg13g2_o21ai_1 _29683_ (.B1(net4515),
    .Y(_04053_),
    .A1(_04033_),
    .A2(_04048_));
 sg13g2_nand2_1 _29684_ (.Y(_04054_),
    .A(net4379),
    .B(_04053_));
 sg13g2_xnor2_1 _29685_ (.Y(_04055_),
    .A(_02736_),
    .B(_04054_));
 sg13g2_a21oi_1 _29686_ (.A1(net5268),
    .A2(_04055_),
    .Y(_00682_),
    .B1(_04052_));
 sg13g2_nand2b_1 _29687_ (.Y(_04056_),
    .B(_02736_),
    .A_N(_02738_));
 sg13g2_or3_1 _29688_ (.A(_04033_),
    .B(_04048_),
    .C(_04056_),
    .X(_04057_));
 sg13g2_nand2_1 _29689_ (.Y(_04058_),
    .A(_02739_),
    .B(_04057_));
 sg13g2_a221oi_1 _29690_ (.B2(net4515),
    .C1(net5119),
    .B1(_04058_),
    .A1(_02738_),
    .Y(_04059_),
    .A2(_04054_));
 sg13g2_a21oi_1 _29691_ (.A1(_14536_),
    .A2(net5119),
    .Y(_00683_),
    .B1(_04059_));
 sg13g2_nor2_1 _29692_ (.A(net1255),
    .B(net5268),
    .Y(_04060_));
 sg13g2_a21o_1 _29693_ (.A2(_04057_),
    .A1(net4515),
    .B1(net4461),
    .X(_04061_));
 sg13g2_xor2_1 _29694_ (.B(_04061_),
    .A(_02797_),
    .X(_04062_));
 sg13g2_a21oi_1 _29695_ (.A1(net5268),
    .A2(_04062_),
    .Y(_00684_),
    .B1(_04060_));
 sg13g2_nor2_1 _29696_ (.A(net1233),
    .B(net5268),
    .Y(_04063_));
 sg13g2_xnor2_1 _29697_ (.Y(_04064_),
    .A(net4515),
    .B(_02797_));
 sg13g2_nor2_1 _29698_ (.A(_04061_),
    .B(_04064_),
    .Y(_04065_));
 sg13g2_xnor2_1 _29699_ (.Y(_04066_),
    .A(_02746_),
    .B(_04065_));
 sg13g2_a21oi_1 _29700_ (.A1(net5268),
    .A2(_04066_),
    .Y(_00685_),
    .B1(_04063_));
 sg13g2_nor2_1 _29701_ (.A(net1135),
    .B(net5268),
    .Y(_04067_));
 sg13g2_nor4_1 _29702_ (.A(_02746_),
    .B(_02797_),
    .C(_04048_),
    .D(_04056_),
    .Y(_04068_));
 sg13g2_nand2_1 _29703_ (.Y(_04069_),
    .A(_04032_),
    .B(_04068_));
 sg13g2_a21oi_1 _29704_ (.A1(net4510),
    .A2(_04069_),
    .Y(_04070_),
    .B1(net4457));
 sg13g2_xnor2_1 _29705_ (.Y(_04071_),
    .A(_03245_),
    .B(_04070_));
 sg13g2_a21oi_1 _29706_ (.A1(net5268),
    .A2(_04071_),
    .Y(_00686_),
    .B1(_04067_));
 sg13g2_nor2_1 _29707_ (.A(_03244_),
    .B(_03245_),
    .Y(_04072_));
 sg13g2_nand3_1 _29708_ (.B(_04068_),
    .C(_04072_),
    .A(_04032_),
    .Y(_04073_));
 sg13g2_inv_1 _29709_ (.Y(_04074_),
    .A(_04073_));
 sg13g2_o21ai_1 _29710_ (.B1(_03244_),
    .Y(_04075_),
    .A1(_03245_),
    .A2(_04069_));
 sg13g2_nand2_1 _29711_ (.Y(_04076_),
    .A(_04073_),
    .B(_04075_));
 sg13g2_a221oi_1 _29712_ (.B2(net4509),
    .C1(net5114),
    .B1(_04076_),
    .A1(_03244_),
    .Y(_04077_),
    .A2(net4457));
 sg13g2_a21oi_1 _29713_ (.A1(_14537_),
    .A2(net5114),
    .Y(_00687_),
    .B1(_04077_));
 sg13g2_nor2_1 _29714_ (.A(net1278),
    .B(net5262),
    .Y(_04078_));
 sg13g2_a21oi_1 _29715_ (.A1(net4509),
    .A2(_04073_),
    .Y(_04079_),
    .B1(net4457));
 sg13g2_xor2_1 _29716_ (.B(_04079_),
    .A(_02685_),
    .X(_04080_));
 sg13g2_a21oi_1 _29717_ (.A1(net5263),
    .A2(_04080_),
    .Y(_00688_),
    .B1(_04078_));
 sg13g2_nor2_1 _29718_ (.A(net1276),
    .B(net5262),
    .Y(_04081_));
 sg13g2_a21oi_1 _29719_ (.A1(_02685_),
    .A2(_04074_),
    .Y(_04082_),
    .B1(_02808_));
 sg13g2_and3_1 _29720_ (.X(_04083_),
    .A(_02685_),
    .B(_02808_),
    .C(_04074_));
 sg13g2_a21o_1 _29721_ (.A2(_04083_),
    .A1(net4509),
    .B1(net5114),
    .X(_04084_));
 sg13g2_a21oi_1 _29722_ (.A1(net4509),
    .A2(_04082_),
    .Y(_04085_),
    .B1(_04084_));
 sg13g2_o21ai_1 _29723_ (.B1(_04085_),
    .Y(_04086_),
    .A1(_02808_),
    .A2(net4377));
 sg13g2_nor2b_1 _29724_ (.A(_04081_),
    .B_N(_04086_),
    .Y(_00689_));
 sg13g2_nor2_1 _29725_ (.A(net1342),
    .B(net5263),
    .Y(_04087_));
 sg13g2_a21oi_1 _29726_ (.A1(net4509),
    .A2(_04083_),
    .Y(_04088_),
    .B1(net4475));
 sg13g2_xnor2_1 _29727_ (.Y(_04089_),
    .A(_02806_),
    .B(_04088_));
 sg13g2_a21oi_1 _29728_ (.A1(net5263),
    .A2(_04089_),
    .Y(_00690_),
    .B1(_04087_));
 sg13g2_nand2_1 _29729_ (.Y(_04090_),
    .A(_02806_),
    .B(_04083_));
 sg13g2_xnor2_1 _29730_ (.Y(_04091_),
    .A(_02755_),
    .B(_04090_));
 sg13g2_a221oi_1 _29731_ (.B2(net4509),
    .C1(net5114),
    .B1(_04091_),
    .A1(_02755_),
    .Y(_04092_),
    .A2(net4458));
 sg13g2_a21oi_1 _29732_ (.A1(_14538_),
    .A2(net5115),
    .Y(_00691_),
    .B1(_04092_));
 sg13g2_o21ai_1 _29733_ (.B1(net4509),
    .Y(_04093_),
    .A1(_02755_),
    .A2(_04090_));
 sg13g2_nor2b_1 _29734_ (.A(net4457),
    .B_N(_04093_),
    .Y(_04094_));
 sg13g2_xnor2_1 _29735_ (.Y(_04095_),
    .A(_02753_),
    .B(_04094_));
 sg13g2_nand2_1 _29736_ (.Y(_04096_),
    .A(net1444),
    .B(net5114));
 sg13g2_o21ai_1 _29737_ (.B1(_04096_),
    .Y(_00692_),
    .A1(net5115),
    .A2(_04095_));
 sg13g2_nor2_1 _29738_ (.A(net1496),
    .B(net5262),
    .Y(_04097_));
 sg13g2_xnor2_1 _29739_ (.Y(_04098_),
    .A(net4491),
    .B(_02753_));
 sg13g2_nand2_1 _29740_ (.Y(_04099_),
    .A(_04094_),
    .B(_04098_));
 sg13g2_xor2_1 _29741_ (.B(_04099_),
    .A(_02750_),
    .X(_04100_));
 sg13g2_a21oi_1 _29742_ (.A1(net5262),
    .A2(_04100_),
    .Y(_00693_),
    .B1(_04097_));
 sg13g2_nor2_1 _29743_ (.A(net1340),
    .B(net5262),
    .Y(_04101_));
 sg13g2_nand4_1 _29744_ (.B(_02806_),
    .C(_02808_),
    .A(_02685_),
    .Y(_04102_),
    .D(_04072_));
 sg13g2_nor4_1 _29745_ (.A(_02750_),
    .B(_02753_),
    .C(_02755_),
    .D(_04102_),
    .Y(_04103_));
 sg13g2_and3_2 _29746_ (.X(_04104_),
    .A(_04032_),
    .B(_04068_),
    .C(_04103_));
 sg13g2_inv_1 _29747_ (.Y(_04105_),
    .A(_04104_));
 sg13g2_a21oi_1 _29748_ (.A1(net4511),
    .A2(_04105_),
    .Y(_04106_),
    .B1(net4457));
 sg13g2_xnor2_1 _29749_ (.Y(_04107_),
    .A(_02802_),
    .B(_04106_));
 sg13g2_a21oi_1 _29750_ (.A1(net5263),
    .A2(_04107_),
    .Y(_00694_),
    .B1(_04101_));
 sg13g2_nor2_1 _29751_ (.A(_02802_),
    .B(_02804_),
    .Y(_04108_));
 sg13g2_and2_1 _29752_ (.A(_04104_),
    .B(_04108_),
    .X(_04109_));
 sg13g2_o21ai_1 _29753_ (.B1(_02804_),
    .Y(_04110_),
    .A1(_02802_),
    .A2(_04105_));
 sg13g2_nand2b_1 _29754_ (.Y(_04111_),
    .B(_04110_),
    .A_N(_04109_));
 sg13g2_a221oi_1 _29755_ (.B2(net4510),
    .C1(net5114),
    .B1(_04111_),
    .A1(_02804_),
    .Y(_04112_),
    .A2(net4458));
 sg13g2_a21oi_1 _29756_ (.A1(_14539_),
    .A2(net5113),
    .Y(_00695_),
    .B1(_04112_));
 sg13g2_a21oi_1 _29757_ (.A1(net4510),
    .A2(_04109_),
    .Y(_04113_),
    .B1(net4475));
 sg13g2_xnor2_1 _29758_ (.Y(_04114_),
    .A(_02718_),
    .B(_04113_));
 sg13g2_nor2_1 _29759_ (.A(net1289),
    .B(net5262),
    .Y(_04115_));
 sg13g2_a21oi_1 _29760_ (.A1(net5262),
    .A2(_04114_),
    .Y(_00696_),
    .B1(_04115_));
 sg13g2_nor2_1 _29761_ (.A(net1349),
    .B(net5262),
    .Y(_04116_));
 sg13g2_nand3_1 _29762_ (.B(_02718_),
    .C(_04109_),
    .A(_02716_),
    .Y(_04117_));
 sg13g2_a21o_1 _29763_ (.A2(_04109_),
    .A1(_02718_),
    .B1(_02716_),
    .X(_04118_));
 sg13g2_nand2_1 _29764_ (.Y(_04119_),
    .A(_04117_),
    .B(_04118_));
 sg13g2_a21oi_1 _29765_ (.A1(net4510),
    .A2(_04119_),
    .Y(_04120_),
    .B1(net5114));
 sg13g2_o21ai_1 _29766_ (.B1(_04120_),
    .Y(_04121_),
    .A1(_02716_),
    .A2(net4377));
 sg13g2_nor2b_1 _29767_ (.A(_04116_),
    .B_N(_04121_),
    .Y(_00697_));
 sg13g2_nor2_1 _29768_ (.A(net1320),
    .B(net5260),
    .Y(_04122_));
 sg13g2_a21oi_1 _29769_ (.A1(net4510),
    .A2(_04117_),
    .Y(_04123_),
    .B1(net4457));
 sg13g2_xnor2_1 _29770_ (.Y(_04124_),
    .A(_02801_),
    .B(_04123_));
 sg13g2_a21oi_1 _29771_ (.A1(net5260),
    .A2(_04124_),
    .Y(_00698_),
    .B1(_04122_));
 sg13g2_nor2_1 _29772_ (.A(_02801_),
    .B(_04117_),
    .Y(_04125_));
 sg13g2_nand2b_1 _29773_ (.Y(_04126_),
    .B(_04125_),
    .A_N(_03238_));
 sg13g2_xor2_1 _29774_ (.B(_04125_),
    .A(_03238_),
    .X(_04127_));
 sg13g2_a221oi_1 _29775_ (.B2(net4509),
    .C1(net5114),
    .B1(_04127_),
    .A1(_03238_),
    .Y(_04128_),
    .A2(net4457));
 sg13g2_a21oi_1 _29776_ (.A1(_14540_),
    .A2(net5113),
    .Y(_00699_),
    .B1(_04128_));
 sg13g2_nor2_1 _29777_ (.A(net2422),
    .B(net5259),
    .Y(_04129_));
 sg13g2_a21oi_1 _29778_ (.A1(net4511),
    .A2(_04126_),
    .Y(_04130_),
    .B1(net4457));
 sg13g2_xnor2_1 _29779_ (.Y(_04131_),
    .A(_02814_),
    .B(_04130_));
 sg13g2_a21oi_1 _29780_ (.A1(net5265),
    .A2(_04131_),
    .Y(_00700_),
    .B1(_04129_));
 sg13g2_nor2_1 _29781_ (.A(net1348),
    .B(net5260),
    .Y(_04132_));
 sg13g2_xnor2_1 _29782_ (.Y(_04133_),
    .A(net4491),
    .B(_02814_));
 sg13g2_nand2_1 _29783_ (.Y(_04134_),
    .A(_04130_),
    .B(_04133_));
 sg13g2_xnor2_1 _29784_ (.Y(_04135_),
    .A(_02818_),
    .B(_04134_));
 sg13g2_a21oi_1 _29785_ (.A1(net5264),
    .A2(_04135_),
    .Y(_00701_),
    .B1(_04132_));
 sg13g2_nor2_1 _29786_ (.A(net1137),
    .B(net5260),
    .Y(_04136_));
 sg13g2_nand3_1 _29787_ (.B(_02718_),
    .C(_02818_),
    .A(_02716_),
    .Y(_04137_));
 sg13g2_nand2_1 _29788_ (.Y(_04138_),
    .A(_02815_),
    .B(_04108_));
 sg13g2_nor4_1 _29789_ (.A(_02801_),
    .B(_03238_),
    .C(_04137_),
    .D(_04138_),
    .Y(_04139_));
 sg13g2_and2_1 _29790_ (.A(_04104_),
    .B(_04139_),
    .X(_04140_));
 sg13g2_a21oi_1 _29791_ (.A1(net4508),
    .A2(_04140_),
    .Y(_04141_),
    .B1(net4474));
 sg13g2_xnor2_1 _29792_ (.Y(_04142_),
    .A(_02693_),
    .B(_04141_));
 sg13g2_a21oi_1 _29793_ (.A1(net5260),
    .A2(_04142_),
    .Y(_00702_),
    .B1(_04136_));
 sg13g2_nand2_1 _29794_ (.Y(_04143_),
    .A(_02693_),
    .B(_02812_));
 sg13g2_nand2_1 _29795_ (.Y(_04144_),
    .A(_02693_),
    .B(_04140_));
 sg13g2_nor2b_1 _29796_ (.A(_04144_),
    .B_N(_02812_),
    .Y(_04145_));
 sg13g2_xor2_1 _29797_ (.B(_04144_),
    .A(_02812_),
    .X(_04146_));
 sg13g2_a21oi_1 _29798_ (.A1(net4508),
    .A2(_04146_),
    .Y(_04147_),
    .B1(net5113));
 sg13g2_o21ai_1 _29799_ (.B1(_04147_),
    .Y(_04148_),
    .A1(_02812_),
    .A2(net4377));
 sg13g2_o21ai_1 _29800_ (.B1(_04148_),
    .Y(_04149_),
    .A1(net2672),
    .A2(net5260));
 sg13g2_inv_1 _29801_ (.Y(_00703_),
    .A(_04149_));
 sg13g2_nor2_1 _29802_ (.A(net1239),
    .B(net5260),
    .Y(_04150_));
 sg13g2_a21oi_1 _29803_ (.A1(net4512),
    .A2(_04145_),
    .Y(_04151_),
    .B1(net4475));
 sg13g2_xnor2_1 _29804_ (.Y(_04152_),
    .A(_03210_),
    .B(_04151_));
 sg13g2_a21oi_1 _29805_ (.A1(net5260),
    .A2(_04152_),
    .Y(_00704_),
    .B1(_04150_));
 sg13g2_nand2_1 _29806_ (.Y(_04153_),
    .A(net2640),
    .B(net5113));
 sg13g2_nand2_1 _29807_ (.Y(_04154_),
    .A(_03210_),
    .B(_04145_));
 sg13g2_nor2_1 _29808_ (.A(_03218_),
    .B(_04154_),
    .Y(_04155_));
 sg13g2_nor2_1 _29809_ (.A(net4490),
    .B(_04155_),
    .Y(_04156_));
 sg13g2_nand2_1 _29810_ (.Y(_04157_),
    .A(_03218_),
    .B(_04154_));
 sg13g2_a21oi_1 _29811_ (.A1(_04156_),
    .A2(_04157_),
    .Y(_04158_),
    .B1(net5115));
 sg13g2_o21ai_1 _29812_ (.B1(_04158_),
    .Y(_04159_),
    .A1(net4512),
    .A2(_03218_));
 sg13g2_o21ai_1 _29813_ (.B1(_04153_),
    .Y(_00705_),
    .A1(net4474),
    .A2(_04159_));
 sg13g2_or2_1 _29814_ (.X(_04160_),
    .B(_04156_),
    .A(net4458));
 sg13g2_xor2_1 _29815_ (.B(_04160_),
    .A(_02654_),
    .X(_04161_));
 sg13g2_nor2_1 _29816_ (.A(net1328),
    .B(net5261),
    .Y(_04162_));
 sg13g2_a21oi_1 _29817_ (.A1(net5261),
    .A2(_04161_),
    .Y(_00706_),
    .B1(_04162_));
 sg13g2_nor2_1 _29818_ (.A(_02653_),
    .B(_02654_),
    .Y(_04163_));
 sg13g2_nand2_1 _29819_ (.Y(_04164_),
    .A(_04155_),
    .B(_04163_));
 sg13g2_nand2_1 _29820_ (.Y(_04165_),
    .A(_02655_),
    .B(_04164_));
 sg13g2_a221oi_1 _29821_ (.B2(net4508),
    .C1(net5115),
    .B1(_04165_),
    .A1(_02653_),
    .Y(_04166_),
    .A2(_04160_));
 sg13g2_a21oi_1 _29822_ (.A1(_14541_),
    .A2(net5115),
    .Y(_00707_),
    .B1(_04166_));
 sg13g2_a21oi_1 _29823_ (.A1(net4508),
    .A2(_04164_),
    .Y(_04167_),
    .B1(net4458));
 sg13g2_xnor2_1 _29824_ (.Y(_04168_),
    .A(_02726_),
    .B(_04167_));
 sg13g2_nor2_1 _29825_ (.A(net1337),
    .B(net5261),
    .Y(_04169_));
 sg13g2_a21oi_1 _29826_ (.A1(net5261),
    .A2(_04168_),
    .Y(_00708_),
    .B1(_04169_));
 sg13g2_nor2_1 _29827_ (.A(net3084),
    .B(net5261),
    .Y(_04170_));
 sg13g2_xnor2_1 _29828_ (.Y(_04171_),
    .A(net4490),
    .B(_02726_));
 sg13g2_nand2_1 _29829_ (.Y(_04172_),
    .A(_04167_),
    .B(_04171_));
 sg13g2_xnor2_1 _29830_ (.Y(_04173_),
    .A(_03234_),
    .B(_04172_));
 sg13g2_a21oi_1 _29831_ (.A1(net5258),
    .A2(_04173_),
    .Y(_00709_),
    .B1(_04170_));
 sg13g2_nor4_1 _29832_ (.A(_02726_),
    .B(_03211_),
    .C(_03218_),
    .D(_04143_),
    .Y(_04174_));
 sg13g2_nand4_1 _29833_ (.B(_04140_),
    .C(_04163_),
    .A(_03234_),
    .Y(_04175_),
    .D(_04174_));
 sg13g2_nor2_1 _29834_ (.A(_02687_),
    .B(_04175_),
    .Y(_04176_));
 sg13g2_nand2b_1 _29835_ (.Y(_04177_),
    .B(net4506),
    .A_N(_04176_));
 sg13g2_a21oi_1 _29836_ (.A1(_02687_),
    .A2(_04175_),
    .Y(_04178_),
    .B1(_04177_));
 sg13g2_o21ai_1 _29837_ (.B1(net5258),
    .Y(_04179_),
    .A1(net4506),
    .A2(_02687_));
 sg13g2_nor3_1 _29838_ (.A(net4476),
    .B(_04178_),
    .C(_04179_),
    .Y(_04180_));
 sg13g2_a21o_1 _29839_ (.A2(net5116),
    .A1(net1363),
    .B1(_04180_),
    .X(_00710_));
 sg13g2_nand2_1 _29840_ (.Y(_04181_),
    .A(net4376),
    .B(_04177_));
 sg13g2_xnor2_1 _29841_ (.Y(_04182_),
    .A(_03248_),
    .B(_04181_));
 sg13g2_nand2_1 _29842_ (.Y(_04183_),
    .A(net1094),
    .B(net5116));
 sg13g2_o21ai_1 _29843_ (.B1(_04183_),
    .Y(_00711_),
    .A1(net5116),
    .A2(_04182_));
 sg13g2_nor2_1 _29844_ (.A(net1631),
    .B(net5261),
    .Y(_04184_));
 sg13g2_xnor2_1 _29845_ (.Y(_04185_),
    .A(net4490),
    .B(_03248_));
 sg13g2_nor2_1 _29846_ (.A(_04181_),
    .B(_04185_),
    .Y(_04186_));
 sg13g2_xnor2_1 _29847_ (.Y(_04187_),
    .A(_02663_),
    .B(_04186_));
 sg13g2_a21oi_1 _29848_ (.A1(net5261),
    .A2(_04187_),
    .Y(_00712_),
    .B1(_04184_));
 sg13g2_nor2_1 _29849_ (.A(net1286),
    .B(net5255),
    .Y(_04188_));
 sg13g2_nor2b_1 _29850_ (.A(_02663_),
    .B_N(_03248_),
    .Y(_04189_));
 sg13g2_and2_1 _29851_ (.A(_04176_),
    .B(_04189_),
    .X(_04190_));
 sg13g2_a21oi_1 _29852_ (.A1(net4506),
    .A2(_04190_),
    .Y(_04191_),
    .B1(net4476));
 sg13g2_xnor2_1 _29853_ (.Y(_04192_),
    .A(_02732_),
    .B(_04191_));
 sg13g2_a21oi_1 _29854_ (.A1(net5255),
    .A2(_04192_),
    .Y(_00713_),
    .B1(_04188_));
 sg13g2_and2_1 _29855_ (.A(_02732_),
    .B(_04190_),
    .X(_04193_));
 sg13g2_o21ai_1 _29856_ (.B1(net4376),
    .Y(_04194_),
    .A1(net4489),
    .A2(_04193_));
 sg13g2_nor2_1 _29857_ (.A(net1226),
    .B(net5255),
    .Y(_04195_));
 sg13g2_xor2_1 _29858_ (.B(_04194_),
    .A(_02781_),
    .X(_04196_));
 sg13g2_a21oi_1 _29859_ (.A1(net5255),
    .A2(_04196_),
    .Y(_00714_),
    .B1(_04195_));
 sg13g2_nor2_1 _29860_ (.A(net1235),
    .B(net5255),
    .Y(_04197_));
 sg13g2_nand2b_1 _29861_ (.Y(_04198_),
    .B(_04193_),
    .A_N(_02781_));
 sg13g2_xnor2_1 _29862_ (.Y(_04199_),
    .A(_02783_),
    .B(_04198_));
 sg13g2_a22oi_1 _29863_ (.Y(_04200_),
    .B1(_04199_),
    .B2(net4506),
    .A2(net4459),
    .A1(_02783_));
 sg13g2_a21oi_1 _29864_ (.A1(net5255),
    .A2(_04200_),
    .Y(_00715_),
    .B1(_04197_));
 sg13g2_nor2_1 _29865_ (.A(net2112),
    .B(net5253),
    .Y(_04201_));
 sg13g2_o21ai_1 _29866_ (.B1(net4506),
    .Y(_04202_),
    .A1(_02783_),
    .A2(_04198_));
 sg13g2_nand2_1 _29867_ (.Y(_04203_),
    .A(net4376),
    .B(_04202_));
 sg13g2_xor2_1 _29868_ (.B(_04203_),
    .A(_03258_),
    .X(_04204_));
 sg13g2_a21oi_1 _29869_ (.A1(net5253),
    .A2(_04204_),
    .Y(_00716_),
    .B1(_04201_));
 sg13g2_nor2_1 _29870_ (.A(net1314),
    .B(net5254),
    .Y(_04205_));
 sg13g2_xnor2_1 _29871_ (.Y(_04206_),
    .A(net4507),
    .B(_03258_));
 sg13g2_nor2_1 _29872_ (.A(_04203_),
    .B(_04206_),
    .Y(_04207_));
 sg13g2_xnor2_1 _29873_ (.Y(_04208_),
    .A(_02641_),
    .B(_04207_));
 sg13g2_a21oi_1 _29874_ (.A1(net5254),
    .A2(_04208_),
    .Y(_00717_),
    .B1(_04205_));
 sg13g2_nor2_1 _29875_ (.A(net2172),
    .B(net5253),
    .Y(_04209_));
 sg13g2_nor4_1 _29876_ (.A(_02641_),
    .B(_02781_),
    .C(_02783_),
    .D(_03258_),
    .Y(_04210_));
 sg13g2_and2_1 _29877_ (.A(_04193_),
    .B(_04210_),
    .X(_04211_));
 sg13g2_a21oi_1 _29878_ (.A1(net4506),
    .A2(_04211_),
    .Y(_04212_),
    .B1(net4476));
 sg13g2_xnor2_1 _29879_ (.Y(_04213_),
    .A(_03247_),
    .B(_04212_));
 sg13g2_a21oi_1 _29880_ (.A1(net5253),
    .A2(_04213_),
    .Y(_00718_),
    .B1(_04209_));
 sg13g2_and3_2 _29881_ (.X(_04214_),
    .A(_02669_),
    .B(_03247_),
    .C(_04211_));
 sg13g2_a21oi_1 _29882_ (.A1(_03247_),
    .A2(_04211_),
    .Y(_04215_),
    .B1(_02669_));
 sg13g2_or2_1 _29883_ (.X(_04216_),
    .B(_04215_),
    .A(_04214_));
 sg13g2_a21oi_1 _29884_ (.A1(net4506),
    .A2(_04216_),
    .Y(_04217_),
    .B1(net5116));
 sg13g2_o21ai_1 _29885_ (.B1(_04217_),
    .Y(_04218_),
    .A1(_02669_),
    .A2(net4376));
 sg13g2_o21ai_1 _29886_ (.B1(_04218_),
    .Y(_04219_),
    .A1(net2979),
    .A2(net5254));
 sg13g2_inv_1 _29887_ (.Y(_00719_),
    .A(_04219_));
 sg13g2_nor2_1 _29888_ (.A(net1180),
    .B(net5254),
    .Y(_04220_));
 sg13g2_o21ai_1 _29889_ (.B1(net4376),
    .Y(_04221_),
    .A1(net4491),
    .A2(_04214_));
 sg13g2_xnor2_1 _29890_ (.Y(_04222_),
    .A(_02658_),
    .B(_04221_));
 sg13g2_a21oi_1 _29891_ (.A1(net5254),
    .A2(_04222_),
    .Y(_00720_),
    .B1(_04220_));
 sg13g2_and3_1 _29892_ (.X(_04223_),
    .A(_02658_),
    .B(_02667_),
    .C(_04214_));
 sg13g2_a21oi_1 _29893_ (.A1(_02658_),
    .A2(_04214_),
    .Y(_04224_),
    .B1(_02667_));
 sg13g2_o21ai_1 _29894_ (.B1(net4507),
    .Y(_04225_),
    .A1(_04223_),
    .A2(_04224_));
 sg13g2_and2_1 _29895_ (.A(net5253),
    .B(_04225_),
    .X(_04226_));
 sg13g2_o21ai_1 _29896_ (.B1(_04226_),
    .Y(_04227_),
    .A1(_02667_),
    .A2(net4376));
 sg13g2_o21ai_1 _29897_ (.B1(_04227_),
    .Y(_04228_),
    .A1(net2948),
    .A2(net5254));
 sg13g2_inv_1 _29898_ (.Y(_00721_),
    .A(_04228_));
 sg13g2_nor2_1 _29899_ (.A(net1129),
    .B(net5254),
    .Y(_04229_));
 sg13g2_o21ai_1 _29900_ (.B1(net4376),
    .Y(_04230_),
    .A1(net4491),
    .A2(_04223_));
 sg13g2_xor2_1 _29901_ (.B(_04230_),
    .A(_02741_),
    .X(_04231_));
 sg13g2_a21oi_1 _29902_ (.A1(net5254),
    .A2(_04231_),
    .Y(_00722_),
    .B1(_04229_));
 sg13g2_nor2_1 _29903_ (.A(_02741_),
    .B(_03257_),
    .Y(_04232_));
 sg13g2_and2_1 _29904_ (.A(_04223_),
    .B(_04232_),
    .X(_04233_));
 sg13g2_o21ai_1 _29905_ (.B1(net4507),
    .Y(_04234_),
    .A1(_03298_),
    .A2(_04233_));
 sg13g2_a21oi_1 _29906_ (.A1(_03257_),
    .A2(_04230_),
    .Y(_04235_),
    .B1(net5116));
 sg13g2_a22oi_1 _29907_ (.Y(_00723_),
    .B1(_04234_),
    .B2(_04235_),
    .A2(net5116),
    .A1(_14542_));
 sg13g2_nor2_1 _29908_ (.A(net1234),
    .B(net5256),
    .Y(_04236_));
 sg13g2_o21ai_1 _29909_ (.B1(net4376),
    .Y(_04237_),
    .A1(net4489),
    .A2(_04233_));
 sg13g2_xnor2_1 _29910_ (.Y(_04238_),
    .A(_02731_),
    .B(_04237_));
 sg13g2_a21oi_1 _29911_ (.A1(net5256),
    .A2(_04238_),
    .Y(_00724_),
    .B1(_04236_));
 sg13g2_nor2_1 _29912_ (.A(net1136),
    .B(net5256),
    .Y(_04239_));
 sg13g2_xnor2_1 _29913_ (.Y(_04240_),
    .A(net4489),
    .B(_02731_));
 sg13g2_nor2_1 _29914_ (.A(_04237_),
    .B(_04240_),
    .Y(_04241_));
 sg13g2_xnor2_1 _29915_ (.Y(_04242_),
    .A(_02795_),
    .B(_04241_));
 sg13g2_a21oi_1 _29916_ (.A1(net5256),
    .A2(_04242_),
    .Y(_00725_),
    .B1(_04239_));
 sg13g2_nor2_1 _29917_ (.A(net1200),
    .B(net5247),
    .Y(_04243_));
 sg13g2_nand2b_1 _29918_ (.Y(_04244_),
    .B(_04189_),
    .A_N(_02795_));
 sg13g2_nand4_1 _29919_ (.B(_03247_),
    .C(_04210_),
    .A(_02669_),
    .Y(_04245_),
    .D(_04232_));
 sg13g2_and2_1 _29920_ (.A(_02686_),
    .B(_02732_),
    .X(_04246_));
 sg13g2_nand4_1 _29921_ (.B(_02667_),
    .C(_02731_),
    .A(_02658_),
    .Y(_04247_),
    .D(_04246_));
 sg13g2_nor4_2 _29922_ (.A(_04175_),
    .B(_04244_),
    .C(_04245_),
    .Y(_04248_),
    .D(_04247_));
 sg13g2_a21oi_1 _29923_ (.A1(net4502),
    .A2(_04248_),
    .Y(_04249_),
    .B1(net4473));
 sg13g2_xnor2_1 _29924_ (.Y(_04250_),
    .A(_02659_),
    .B(_04249_));
 sg13g2_a21oi_1 _29925_ (.A1(net5247),
    .A2(_04250_),
    .Y(_00726_),
    .B1(_04243_));
 sg13g2_nand2b_1 _29926_ (.Y(_04251_),
    .B(net4456),
    .A_N(_03254_));
 sg13g2_nand3_1 _29927_ (.B(_03254_),
    .C(_04248_),
    .A(_02659_),
    .Y(_04252_));
 sg13g2_a21o_1 _29928_ (.A2(_04248_),
    .A1(_02659_),
    .B1(_03254_),
    .X(_04253_));
 sg13g2_nand2_1 _29929_ (.Y(_04254_),
    .A(_04252_),
    .B(_04253_));
 sg13g2_a21oi_1 _29930_ (.A1(net4503),
    .A2(_04254_),
    .Y(_04255_),
    .B1(net5111));
 sg13g2_a22oi_1 _29931_ (.Y(_00727_),
    .B1(_04251_),
    .B2(_04255_),
    .A2(net5111),
    .A1(_14543_));
 sg13g2_a21oi_1 _29932_ (.A1(net4503),
    .A2(_04252_),
    .Y(_04256_),
    .B1(net4456));
 sg13g2_xnor2_1 _29933_ (.Y(_04257_),
    .A(_02644_),
    .B(_04256_));
 sg13g2_nor2_1 _29934_ (.A(net1302),
    .B(net5247),
    .Y(_04258_));
 sg13g2_a21oi_1 _29935_ (.A1(net5248),
    .A2(_04257_),
    .Y(_00728_),
    .B1(_04258_));
 sg13g2_nor3_1 _29936_ (.A(_02644_),
    .B(_02770_),
    .C(_04252_),
    .Y(_04259_));
 sg13g2_o21ai_1 _29937_ (.B1(_02770_),
    .Y(_04260_),
    .A1(_02644_),
    .A2(_04252_));
 sg13g2_nand2b_1 _29938_ (.Y(_04261_),
    .B(_04260_),
    .A_N(_04259_));
 sg13g2_a221oi_1 _29939_ (.B2(net4503),
    .C1(net5111),
    .B1(_04261_),
    .A1(_02770_),
    .Y(_04262_),
    .A2(net4456));
 sg13g2_a21oi_1 _29940_ (.A1(_14544_),
    .A2(net5111),
    .Y(_00729_),
    .B1(_04262_));
 sg13g2_nor2_1 _29941_ (.A(net1275),
    .B(net5247),
    .Y(_04263_));
 sg13g2_o21ai_1 _29942_ (.B1(net4375),
    .Y(_04264_),
    .A1(net4487),
    .A2(_04259_));
 sg13g2_xor2_1 _29943_ (.B(_04264_),
    .A(_02607_),
    .X(_04265_));
 sg13g2_a21oi_1 _29944_ (.A1(net5248),
    .A2(_04265_),
    .Y(_00730_),
    .B1(_04263_));
 sg13g2_nor2_1 _29945_ (.A(_02607_),
    .B(_02609_),
    .Y(_04266_));
 sg13g2_nand2_1 _29946_ (.Y(_04267_),
    .A(_04259_),
    .B(_04266_));
 sg13g2_nand2_1 _29947_ (.Y(_04268_),
    .A(_02610_),
    .B(_04267_));
 sg13g2_a221oi_1 _29948_ (.B2(net4502),
    .C1(net5112),
    .B1(_04268_),
    .A1(_02609_),
    .Y(_04269_),
    .A2(_04264_));
 sg13g2_a21oi_1 _29949_ (.A1(_14545_),
    .A2(net5111),
    .Y(_00731_),
    .B1(_04269_));
 sg13g2_a21oi_1 _29950_ (.A1(net4502),
    .A2(_04267_),
    .Y(_04270_),
    .B1(net4456));
 sg13g2_xor2_1 _29951_ (.B(_04270_),
    .A(_03255_),
    .X(_04271_));
 sg13g2_nor2_1 _29952_ (.A(net1285),
    .B(net5247),
    .Y(_04272_));
 sg13g2_a21oi_1 _29953_ (.A1(net5247),
    .A2(_04271_),
    .Y(_00732_),
    .B1(_04272_));
 sg13g2_nor2_1 _29954_ (.A(net1123),
    .B(net5247),
    .Y(_04273_));
 sg13g2_xnor2_1 _29955_ (.Y(_04274_),
    .A(net4502),
    .B(_03255_));
 sg13g2_nand2_1 _29956_ (.Y(_04275_),
    .A(_04270_),
    .B(_04274_));
 sg13g2_xnor2_1 _29957_ (.Y(_04276_),
    .A(_02647_),
    .B(_04275_));
 sg13g2_a21oi_1 _29958_ (.A1(net5247),
    .A2(_04276_),
    .Y(_00733_),
    .B1(_04273_));
 sg13g2_nor2_1 _29959_ (.A(net1248),
    .B(net5246),
    .Y(_04277_));
 sg13g2_nor2b_1 _29960_ (.A(_02644_),
    .B_N(_03255_),
    .Y(_04278_));
 sg13g2_nand4_1 _29961_ (.B(_02659_),
    .C(_03254_),
    .A(_02647_),
    .Y(_04279_),
    .D(_04278_));
 sg13g2_nor4_1 _29962_ (.A(_02607_),
    .B(_02609_),
    .C(_02770_),
    .D(_04279_),
    .Y(_04280_));
 sg13g2_and2_1 _29963_ (.A(_04248_),
    .B(_04280_),
    .X(_04281_));
 sg13g2_o21ai_1 _29964_ (.B1(net4375),
    .Y(_04282_),
    .A1(net4488),
    .A2(_04281_));
 sg13g2_xnor2_1 _29965_ (.Y(_04283_),
    .A(_02634_),
    .B(_04282_));
 sg13g2_a21oi_1 _29966_ (.A1(net5245),
    .A2(_04283_),
    .Y(_00734_),
    .B1(_04277_));
 sg13g2_nor2_1 _29967_ (.A(net1127),
    .B(net5245),
    .Y(_04284_));
 sg13g2_nand3_1 _29968_ (.B(_02775_),
    .C(_04281_),
    .A(_02634_),
    .Y(_04285_));
 sg13g2_a21o_1 _29969_ (.A2(_04281_),
    .A1(_02634_),
    .B1(_02775_),
    .X(_04286_));
 sg13g2_nand2_1 _29970_ (.Y(_04287_),
    .A(_04285_),
    .B(_04286_));
 sg13g2_a22oi_1 _29971_ (.Y(_04288_),
    .B1(_04287_),
    .B2(net4502),
    .A2(net4456),
    .A1(_02776_));
 sg13g2_a21oi_1 _29972_ (.A1(net5245),
    .A2(_04288_),
    .Y(_00735_),
    .B1(_04284_));
 sg13g2_nor2_1 _29973_ (.A(net1284),
    .B(net5245),
    .Y(_04289_));
 sg13g2_a21oi_1 _29974_ (.A1(net4502),
    .A2(_04285_),
    .Y(_04290_),
    .B1(net4459));
 sg13g2_xor2_1 _29975_ (.B(_04290_),
    .A(_02767_),
    .X(_04291_));
 sg13g2_a21oi_1 _29976_ (.A1(net5245),
    .A2(_04291_),
    .Y(_00736_),
    .B1(_04289_));
 sg13g2_nand3_1 _29977_ (.B(_02767_),
    .C(_02775_),
    .A(_02634_),
    .Y(_04292_));
 sg13g2_nor2b_1 _29978_ (.A(_04285_),
    .B_N(_02767_),
    .Y(_04293_));
 sg13g2_and2_1 _29979_ (.A(_02773_),
    .B(_04293_),
    .X(_04294_));
 sg13g2_xnor2_1 _29980_ (.Y(_04295_),
    .A(_02773_),
    .B(_04293_));
 sg13g2_a21oi_1 _29981_ (.A1(net4504),
    .A2(_04295_),
    .Y(_04296_),
    .B1(net5111));
 sg13g2_o21ai_1 _29982_ (.B1(_04296_),
    .Y(_04297_),
    .A1(_02773_),
    .A2(net4375));
 sg13g2_o21ai_1 _29983_ (.B1(_04297_),
    .Y(_04298_),
    .A1(net2775),
    .A2(net5246));
 sg13g2_inv_1 _29984_ (.Y(_00737_),
    .A(_04298_));
 sg13g2_nor2_1 _29985_ (.A(net1283),
    .B(net5246),
    .Y(_04299_));
 sg13g2_o21ai_1 _29986_ (.B1(net4375),
    .Y(_04300_),
    .A1(net4487),
    .A2(_04294_));
 sg13g2_xnor2_1 _29987_ (.Y(_04301_),
    .A(_02761_),
    .B(_04300_));
 sg13g2_a21oi_1 _29988_ (.A1(net5245),
    .A2(_04301_),
    .Y(_00738_),
    .B1(_04299_));
 sg13g2_nor2_1 _29989_ (.A(net1209),
    .B(net5245),
    .Y(_04302_));
 sg13g2_nand2_1 _29990_ (.Y(_04303_),
    .A(_02761_),
    .B(_04294_));
 sg13g2_xnor2_1 _29991_ (.Y(_04304_),
    .A(_03264_),
    .B(_04303_));
 sg13g2_a22oi_1 _29992_ (.Y(_04305_),
    .B1(_04304_),
    .B2(net4504),
    .A2(net4456),
    .A1(_03264_));
 sg13g2_a21oi_1 _29993_ (.A1(net5245),
    .A2(_04305_),
    .Y(_00739_),
    .B1(_04302_));
 sg13g2_nor2_1 _29994_ (.A(net1351),
    .B(net5244),
    .Y(_04306_));
 sg13g2_o21ai_1 _29995_ (.B1(net4504),
    .Y(_04307_),
    .A1(_03264_),
    .A2(_04303_));
 sg13g2_nor2b_1 _29996_ (.A(net4456),
    .B_N(_04307_),
    .Y(_04308_));
 sg13g2_xnor2_1 _29997_ (.Y(_04309_),
    .A(_02617_),
    .B(_04308_));
 sg13g2_a21oi_1 _29998_ (.A1(net5244),
    .A2(_04309_),
    .Y(_00740_),
    .B1(_04306_));
 sg13g2_nor2_1 _29999_ (.A(net1357),
    .B(net5246),
    .Y(_04310_));
 sg13g2_xnor2_1 _30000_ (.Y(_04311_),
    .A(net4504),
    .B(_02618_));
 sg13g2_nand2_1 _30001_ (.Y(_04312_),
    .A(_04308_),
    .B(_04311_));
 sg13g2_xnor2_1 _30002_ (.Y(_04313_),
    .A(_02616_),
    .B(_04312_));
 sg13g2_a21oi_1 _30003_ (.A1(net5244),
    .A2(_04313_),
    .Y(_00741_),
    .B1(_04310_));
 sg13g2_nand4_1 _30004_ (.B(_02618_),
    .C(_02761_),
    .A(_02616_),
    .Y(_04314_),
    .D(_02773_));
 sg13g2_nor3_1 _30005_ (.A(_03264_),
    .B(_04292_),
    .C(_04314_),
    .Y(_04315_));
 sg13g2_nand4_1 _30006_ (.B(_04248_),
    .C(_04280_),
    .A(net4502),
    .Y(_04316_),
    .D(_04315_));
 sg13g2_and2_1 _30007_ (.A(_04281_),
    .B(_04315_),
    .X(_04317_));
 sg13g2_o21ai_1 _30008_ (.B1(net4375),
    .Y(_04318_),
    .A1(net4487),
    .A2(_04317_));
 sg13g2_xnor2_1 _30009_ (.Y(_04319_),
    .A(_03252_),
    .B(_04318_));
 sg13g2_nand2_1 _30010_ (.Y(_04320_),
    .A(net1100),
    .B(net5109));
 sg13g2_o21ai_1 _30011_ (.B1(_04320_),
    .Y(_00742_),
    .A1(net5109),
    .A2(_04319_));
 sg13g2_nor2_1 _30012_ (.A(net1134),
    .B(net5244),
    .Y(_04321_));
 sg13g2_nor2b_2 _30013_ (.A(_02763_),
    .B_N(_03252_),
    .Y(_04322_));
 sg13g2_nor2b_1 _30014_ (.A(_04316_),
    .B_N(_04322_),
    .Y(_04323_));
 sg13g2_and2_1 _30015_ (.A(_04317_),
    .B(_04322_),
    .X(_04324_));
 sg13g2_nor3_1 _30016_ (.A(net4487),
    .B(_02764_),
    .C(_03252_),
    .Y(_04325_));
 sg13g2_a221oi_1 _30017_ (.B2(net4504),
    .C1(_04325_),
    .B1(_04324_),
    .A1(_02763_),
    .Y(_04326_),
    .A2(_04318_));
 sg13g2_a21oi_1 _30018_ (.A1(net5244),
    .A2(_04326_),
    .Y(_00743_),
    .B1(_04321_));
 sg13g2_nor2_1 _30019_ (.A(net1122),
    .B(net5243),
    .Y(_04327_));
 sg13g2_nor2_1 _30020_ (.A(net4473),
    .B(_04323_),
    .Y(_04328_));
 sg13g2_xnor2_1 _30021_ (.Y(_04329_),
    .A(_02626_),
    .B(_04328_));
 sg13g2_a21oi_1 _30022_ (.A1(net5243),
    .A2(_04329_),
    .Y(_00744_),
    .B1(_04327_));
 sg13g2_nand2_1 _30023_ (.Y(_04330_),
    .A(_02626_),
    .B(_04324_));
 sg13g2_nor2_1 _30024_ (.A(_02603_),
    .B(_04330_),
    .Y(_04331_));
 sg13g2_xnor2_1 _30025_ (.Y(_04332_),
    .A(_02603_),
    .B(_04330_));
 sg13g2_a221oi_1 _30026_ (.B2(net4504),
    .C1(net5110),
    .B1(_04332_),
    .A1(_02603_),
    .Y(_04333_),
    .A2(net4456));
 sg13g2_a21oi_1 _30027_ (.A1(_14546_),
    .A2(net5110),
    .Y(_00745_),
    .B1(_04333_));
 sg13g2_nor2_1 _30028_ (.A(net1293),
    .B(net5243),
    .Y(_04334_));
 sg13g2_o21ai_1 _30029_ (.B1(net4375),
    .Y(_04335_),
    .A1(net4487),
    .A2(_04331_));
 sg13g2_xor2_1 _30030_ (.B(_04335_),
    .A(_02622_),
    .X(_04336_));
 sg13g2_a21oi_1 _30031_ (.A1(net5243),
    .A2(_04336_),
    .Y(_00746_),
    .B1(_04334_));
 sg13g2_nor2_1 _30032_ (.A(_02622_),
    .B(_03267_),
    .Y(_04337_));
 sg13g2_nand2_1 _30033_ (.Y(_04338_),
    .A(_04331_),
    .B(_04337_));
 sg13g2_nand2_1 _30034_ (.Y(_04339_),
    .A(_03300_),
    .B(_04338_));
 sg13g2_a221oi_1 _30035_ (.B2(net4501),
    .C1(net5110),
    .B1(_04339_),
    .A1(_03267_),
    .Y(_04340_),
    .A2(_04335_));
 sg13g2_a21oi_1 _30036_ (.A1(_14547_),
    .A2(net5110),
    .Y(_00747_),
    .B1(_04340_));
 sg13g2_nor2_1 _30037_ (.A(net1321),
    .B(net5243),
    .Y(_04341_));
 sg13g2_a21oi_1 _30038_ (.A1(net4501),
    .A2(_04338_),
    .Y(_04342_),
    .B1(net4455));
 sg13g2_xor2_1 _30039_ (.B(_04342_),
    .A(_02612_),
    .X(_04343_));
 sg13g2_a21oi_1 _30040_ (.A1(net5243),
    .A2(_04343_),
    .Y(_00748_),
    .B1(_04341_));
 sg13g2_nor2_1 _30041_ (.A(net1334),
    .B(net5243),
    .Y(_04344_));
 sg13g2_xnor2_1 _30042_ (.Y(_04345_),
    .A(net4501),
    .B(_02612_));
 sg13g2_nand2_1 _30043_ (.Y(_04346_),
    .A(_04342_),
    .B(_04345_));
 sg13g2_xnor2_1 _30044_ (.Y(_04347_),
    .A(_02628_),
    .B(_04346_));
 sg13g2_a21oi_1 _30045_ (.A1(net5243),
    .A2(_04347_),
    .Y(_00749_),
    .B1(_04344_));
 sg13g2_nor2_1 _30046_ (.A(net1318),
    .B(net5232),
    .Y(_04348_));
 sg13g2_and4_1 _30047_ (.A(_02604_),
    .B(_02612_),
    .C(_02626_),
    .D(_02628_),
    .X(_04349_));
 sg13g2_and4_1 _30048_ (.A(_04317_),
    .B(_04322_),
    .C(_04337_),
    .D(_04349_),
    .X(_04350_));
 sg13g2_a21oi_1 _30049_ (.A1(net4500),
    .A2(_04350_),
    .Y(_04351_),
    .B1(net4472));
 sg13g2_xor2_1 _30050_ (.B(_04351_),
    .A(_02630_),
    .X(_04352_));
 sg13g2_a21oi_1 _30051_ (.A1(net5232),
    .A2(_04352_),
    .Y(_00750_),
    .B1(_04348_));
 sg13g2_nor2_1 _30052_ (.A(net1251),
    .B(net5231),
    .Y(_04353_));
 sg13g2_nor2_1 _30053_ (.A(_02630_),
    .B(_03269_),
    .Y(_04354_));
 sg13g2_nor2b_1 _30054_ (.A(_02630_),
    .B_N(_04350_),
    .Y(_04355_));
 sg13g2_nand2_1 _30055_ (.Y(_04356_),
    .A(_04350_),
    .B(_04354_));
 sg13g2_xor2_1 _30056_ (.B(_04355_),
    .A(_03269_),
    .X(_04357_));
 sg13g2_a22oi_1 _30057_ (.Y(_04358_),
    .B1(_04357_),
    .B2(net4500),
    .A2(net4454),
    .A1(_03269_));
 sg13g2_a21oi_1 _30058_ (.A1(net5232),
    .A2(_04358_),
    .Y(_00751_),
    .B1(_04353_));
 sg13g2_a21oi_1 _30059_ (.A1(net4500),
    .A2(_04356_),
    .Y(_04359_),
    .B1(net4454));
 sg13g2_xor2_1 _30060_ (.B(_04359_),
    .A(_03278_),
    .X(_04360_));
 sg13g2_nor2_1 _30061_ (.A(net1208),
    .B(net5233),
    .Y(_04361_));
 sg13g2_a21oi_1 _30062_ (.A1(net5233),
    .A2(_04360_),
    .Y(_00752_),
    .B1(_04361_));
 sg13g2_a21o_1 _30063_ (.A2(_04359_),
    .A1(_03278_),
    .B1(_02581_),
    .X(_04362_));
 sg13g2_and4_1 _30064_ (.A(_02581_),
    .B(_03278_),
    .C(_04350_),
    .D(_04354_),
    .X(_04363_));
 sg13g2_a21oi_1 _30065_ (.A1(net4500),
    .A2(_04363_),
    .Y(_04364_),
    .B1(net5107));
 sg13g2_o21ai_1 _30066_ (.B1(_04364_),
    .Y(_04365_),
    .A1(net4472),
    .A2(_04362_));
 sg13g2_o21ai_1 _30067_ (.B1(_04365_),
    .Y(_04366_),
    .A1(net2521),
    .A2(net5233));
 sg13g2_inv_1 _30068_ (.Y(_00753_),
    .A(_04366_));
 sg13g2_o21ai_1 _30069_ (.B1(net4374),
    .Y(_04367_),
    .A1(net4485),
    .A2(_04363_));
 sg13g2_xnor2_1 _30070_ (.Y(_04368_),
    .A(_02623_),
    .B(_04367_));
 sg13g2_nor2_1 _30071_ (.A(net2592),
    .B(net5238),
    .Y(_04369_));
 sg13g2_a21oi_1 _30072_ (.A1(net5233),
    .A2(_04368_),
    .Y(_00754_),
    .B1(_04369_));
 sg13g2_nand2_1 _30073_ (.Y(_04370_),
    .A(_02623_),
    .B(_03276_));
 sg13g2_nand2_1 _30074_ (.Y(_04371_),
    .A(_02623_),
    .B(_04363_));
 sg13g2_nor2b_1 _30075_ (.A(_04371_),
    .B_N(_03276_),
    .Y(_04372_));
 sg13g2_xor2_1 _30076_ (.B(_04371_),
    .A(_03276_),
    .X(_04373_));
 sg13g2_a21oi_1 _30077_ (.A1(net4499),
    .A2(_04373_),
    .Y(_04374_),
    .B1(net5107));
 sg13g2_o21ai_1 _30078_ (.B1(_04374_),
    .Y(_04375_),
    .A1(_03276_),
    .A2(net4374));
 sg13g2_o21ai_1 _30079_ (.B1(_04375_),
    .Y(_04376_),
    .A1(net2816),
    .A2(net5234));
 sg13g2_inv_1 _30080_ (.Y(_00755_),
    .A(_04376_));
 sg13g2_o21ai_1 _30081_ (.B1(net4374),
    .Y(_04377_),
    .A1(net4484),
    .A2(_04372_));
 sg13g2_xor2_1 _30082_ (.B(_04377_),
    .A(_02576_),
    .X(_04378_));
 sg13g2_nand2_1 _30083_ (.Y(_04379_),
    .A(net1098),
    .B(net5107));
 sg13g2_o21ai_1 _30084_ (.B1(_04379_),
    .Y(_00756_),
    .A1(net5107),
    .A2(_04378_));
 sg13g2_nor2_1 _30085_ (.A(net1281),
    .B(net5233),
    .Y(_04380_));
 sg13g2_xnor2_1 _30086_ (.Y(_04381_),
    .A(net4499),
    .B(_02576_));
 sg13g2_nor2_1 _30087_ (.A(_04377_),
    .B(_04381_),
    .Y(_04382_));
 sg13g2_xnor2_1 _30088_ (.Y(_04383_),
    .A(_02595_),
    .B(_04382_));
 sg13g2_a21oi_1 _30089_ (.A1(net5233),
    .A2(_04383_),
    .Y(_00757_),
    .B1(_04380_));
 sg13g2_nor2_1 _30090_ (.A(net1227),
    .B(net5234),
    .Y(_04384_));
 sg13g2_nor3_1 _30091_ (.A(_02576_),
    .B(_02595_),
    .C(_04370_),
    .Y(_04385_));
 sg13g2_nand2_2 _30092_ (.Y(_04386_),
    .A(_04363_),
    .B(_04385_));
 sg13g2_a21oi_1 _30093_ (.A1(net4498),
    .A2(_04386_),
    .Y(_04387_),
    .B1(net4454));
 sg13g2_nor3_1 _30094_ (.A(net4483),
    .B(_03274_),
    .C(_04386_),
    .Y(_04388_));
 sg13g2_xnor2_1 _30095_ (.Y(_04389_),
    .A(_03274_),
    .B(_04387_));
 sg13g2_a21oi_1 _30096_ (.A1(net5234),
    .A2(_04389_),
    .Y(_00758_),
    .B1(_04384_));
 sg13g2_or2_1 _30097_ (.X(_04390_),
    .B(net5234),
    .A(net3411));
 sg13g2_nor3_1 _30098_ (.A(_02583_),
    .B(net4472),
    .C(_04388_),
    .Y(_04391_));
 sg13g2_nand2b_1 _30099_ (.Y(_04392_),
    .B(_02583_),
    .A_N(_03274_));
 sg13g2_nor2_1 _30100_ (.A(_04386_),
    .B(_04392_),
    .Y(_04393_));
 sg13g2_a21o_1 _30101_ (.A2(_04393_),
    .A1(net4498),
    .B1(net5104),
    .X(_04394_));
 sg13g2_o21ai_1 _30102_ (.B1(_04390_),
    .Y(_04395_),
    .A1(_04391_),
    .A2(_04394_));
 sg13g2_inv_1 _30103_ (.Y(_00759_),
    .A(_04395_));
 sg13g2_nor2_1 _30104_ (.A(net1267),
    .B(net5234),
    .Y(_04396_));
 sg13g2_o21ai_1 _30105_ (.B1(net4374),
    .Y(_04397_),
    .A1(net4483),
    .A2(_04393_));
 sg13g2_xor2_1 _30106_ (.B(_04397_),
    .A(_02597_),
    .X(_04398_));
 sg13g2_a21oi_1 _30107_ (.A1(net5234),
    .A2(_04398_),
    .Y(_00760_),
    .B1(_04396_));
 sg13g2_nor4_1 _30108_ (.A(_02573_),
    .B(_02597_),
    .C(_04386_),
    .D(_04392_),
    .Y(_04399_));
 sg13g2_or4_1 _30109_ (.A(net4483),
    .B(_02597_),
    .C(_04386_),
    .D(_04392_),
    .X(_04400_));
 sg13g2_a22oi_1 _30110_ (.Y(_04401_),
    .B1(_04400_),
    .B2(_02573_),
    .A2(_04399_),
    .A1(net4498));
 sg13g2_nor3_1 _30111_ (.A(net5104),
    .B(net4472),
    .C(_04401_),
    .Y(_04402_));
 sg13g2_a21o_1 _30112_ (.A2(net5104),
    .A1(net1381),
    .B1(_04402_),
    .X(_00761_));
 sg13g2_o21ai_1 _30113_ (.B1(net4374),
    .Y(_04403_),
    .A1(net4483),
    .A2(_04399_));
 sg13g2_xor2_1 _30114_ (.B(_04403_),
    .A(_03262_),
    .X(_04404_));
 sg13g2_nor2_1 _30115_ (.A(net1174),
    .B(net5233),
    .Y(_04405_));
 sg13g2_a21oi_1 _30116_ (.A1(net5233),
    .A2(_04404_),
    .Y(_00762_),
    .B1(_04405_));
 sg13g2_nor2_1 _30117_ (.A(_03262_),
    .B(_03273_),
    .Y(_04406_));
 sg13g2_nand2_1 _30118_ (.Y(_04407_),
    .A(_04399_),
    .B(_04406_));
 sg13g2_nand2_1 _30119_ (.Y(_04408_),
    .A(_03299_),
    .B(_04407_));
 sg13g2_a221oi_1 _30120_ (.B2(net4498),
    .C1(net5105),
    .B1(_04408_),
    .A1(_03273_),
    .Y(_04409_),
    .A2(_04403_));
 sg13g2_a21oi_1 _30121_ (.A1(_14548_),
    .A2(net5105),
    .Y(_00763_),
    .B1(_04409_));
 sg13g2_a21oi_1 _30122_ (.A1(net4498),
    .A2(_04407_),
    .Y(_04410_),
    .B1(net4454));
 sg13g2_xnor2_1 _30123_ (.Y(_04411_),
    .A(_02591_),
    .B(_04410_));
 sg13g2_nand2_1 _30124_ (.Y(_04412_),
    .A(net1082),
    .B(net5104));
 sg13g2_o21ai_1 _30125_ (.B1(_04412_),
    .Y(_00764_),
    .A1(net5104),
    .A2(_04411_));
 sg13g2_nor2_1 _30126_ (.A(net1341),
    .B(net5231),
    .Y(_04413_));
 sg13g2_xnor2_1 _30127_ (.Y(_04414_),
    .A(net4483),
    .B(_02591_));
 sg13g2_nand2_1 _30128_ (.Y(_04415_),
    .A(_04410_),
    .B(_04414_));
 sg13g2_xor2_1 _30129_ (.B(_04415_),
    .A(_02587_),
    .X(_04416_));
 sg13g2_a21oi_1 _30130_ (.A1(net5231),
    .A2(_04416_),
    .Y(_00765_),
    .B1(_04413_));
 sg13g2_nor2_1 _30131_ (.A(net1212),
    .B(net5234),
    .Y(_04417_));
 sg13g2_nor3_1 _30132_ (.A(_02587_),
    .B(_02591_),
    .C(_04407_),
    .Y(_04418_));
 sg13g2_o21ai_1 _30133_ (.B1(net4374),
    .Y(_04419_),
    .A1(net4483),
    .A2(_04418_));
 sg13g2_nand3_1 _30134_ (.B(_02588_),
    .C(_04418_),
    .A(net4498),
    .Y(_04420_));
 sg13g2_xnor2_1 _30135_ (.Y(_04421_),
    .A(_02588_),
    .B(_04419_));
 sg13g2_a21oi_1 _30136_ (.A1(net5234),
    .A2(_04421_),
    .Y(_00766_),
    .B1(_04417_));
 sg13g2_and2_1 _30137_ (.A(_03293_),
    .B(_04420_),
    .X(_04422_));
 sg13g2_nand3b_1 _30138_ (.B(_04418_),
    .C(_02588_),
    .Y(_04423_),
    .A_N(_03293_));
 sg13g2_o21ai_1 _30139_ (.B1(net5231),
    .Y(_04424_),
    .A1(net4484),
    .A2(_04423_));
 sg13g2_a21oi_1 _30140_ (.A1(net4470),
    .A2(_04422_),
    .Y(_04425_),
    .B1(_04424_));
 sg13g2_a21oi_1 _30141_ (.A1(_14549_),
    .A2(net5104),
    .Y(_00767_),
    .B1(_04425_));
 sg13g2_a21oi_1 _30142_ (.A1(net4498),
    .A2(_04423_),
    .Y(_04426_),
    .B1(net4454));
 sg13g2_xnor2_1 _30143_ (.Y(_04427_),
    .A(_02568_),
    .B(_04426_));
 sg13g2_nand2_1 _30144_ (.Y(_04428_),
    .A(net1089),
    .B(net5106));
 sg13g2_o21ai_1 _30145_ (.B1(_04428_),
    .Y(_00768_),
    .A1(net5106),
    .A2(_04427_));
 sg13g2_nand2b_1 _30146_ (.Y(_04429_),
    .B(_02567_),
    .A_N(_04423_));
 sg13g2_nor3_1 _30147_ (.A(_02568_),
    .B(_03287_),
    .C(_04423_),
    .Y(_04430_));
 sg13g2_xnor2_1 _30148_ (.Y(_04431_),
    .A(_03287_),
    .B(_04429_));
 sg13g2_a221oi_1 _30149_ (.B2(net4498),
    .C1(net5104),
    .B1(_04431_),
    .A1(_03287_),
    .Y(_04432_),
    .A2(net4454));
 sg13g2_a21oi_1 _30150_ (.A1(_14550_),
    .A2(net5104),
    .Y(_00769_),
    .B1(_04432_));
 sg13g2_o21ai_1 _30151_ (.B1(net4374),
    .Y(_04433_),
    .A1(net4484),
    .A2(_04430_));
 sg13g2_xnor2_1 _30152_ (.Y(_04434_),
    .A(_03290_),
    .B(_04433_));
 sg13g2_nand2_1 _30153_ (.Y(_04435_),
    .A(net1170),
    .B(net5106));
 sg13g2_o21ai_1 _30154_ (.B1(_04435_),
    .Y(_00770_),
    .A1(net5106),
    .A2(_04434_));
 sg13g2_and3_1 _30155_ (.X(_04436_),
    .A(_03289_),
    .B(_03290_),
    .C(_04430_));
 sg13g2_a21oi_1 _30156_ (.A1(_03290_),
    .A2(_04430_),
    .Y(_04437_),
    .B1(_03289_));
 sg13g2_o21ai_1 _30157_ (.B1(net4499),
    .Y(_04438_),
    .A1(_04436_),
    .A2(_04437_));
 sg13g2_a21oi_1 _30158_ (.A1(_03288_),
    .A2(net4454),
    .Y(_04439_),
    .B1(net5105));
 sg13g2_a22oi_1 _30159_ (.Y(_00771_),
    .B1(_04438_),
    .B2(_04439_),
    .A2(net5105),
    .A1(_14551_));
 sg13g2_nor2_1 _30160_ (.A(net1366),
    .B(net5231),
    .Y(_04440_));
 sg13g2_nor2_1 _30161_ (.A(net4484),
    .B(_04436_),
    .Y(_04441_));
 sg13g2_nor2_1 _30162_ (.A(net4455),
    .B(_04441_),
    .Y(_04442_));
 sg13g2_xnor2_1 _30163_ (.Y(_04443_),
    .A(_03283_),
    .B(_04442_));
 sg13g2_a21oi_1 _30164_ (.A1(net5231),
    .A2(_04443_),
    .Y(_00772_),
    .B1(_04440_));
 sg13g2_nor2_1 _30165_ (.A(net1476),
    .B(net5231),
    .Y(_04444_));
 sg13g2_o21ai_1 _30166_ (.B1(net4470),
    .Y(_04445_),
    .A1(net4483),
    .A2(_03283_));
 sg13g2_nor2b_1 _30167_ (.A(_04441_),
    .B_N(_04445_),
    .Y(_04446_));
 sg13g2_xor2_1 _30168_ (.B(_04446_),
    .A(_02564_),
    .X(_04447_));
 sg13g2_a21oi_1 _30169_ (.A1(net5231),
    .A2(_04447_),
    .Y(_00773_),
    .B1(_04444_));
 sg13g2_xnor2_1 _30170_ (.Y(_04448_),
    .A(\u_inv.d_next[256] ),
    .B(\u_inv.d_reg[256] ));
 sg13g2_xor2_1 _30171_ (.B(\u_inv.d_reg[256] ),
    .A(\u_inv.d_next[256] ),
    .X(_04449_));
 sg13g2_nor2_1 _30172_ (.A(\u_inv.d_next[255] ),
    .B(\u_inv.d_reg[255] ),
    .Y(_04450_));
 sg13g2_nand2_1 _30173_ (.Y(_04451_),
    .A(\u_inv.d_next[255] ),
    .B(\u_inv.d_reg[255] ));
 sg13g2_nor2b_1 _30174_ (.A(_04450_),
    .B_N(_04451_),
    .Y(_04452_));
 sg13g2_nand2b_2 _30175_ (.Y(_04453_),
    .B(_04451_),
    .A_N(_04450_));
 sg13g2_nand2_1 _30176_ (.Y(_04454_),
    .A(\u_inv.d_next[254] ),
    .B(\u_inv.d_reg[254] ));
 sg13g2_xor2_1 _30177_ (.B(\u_inv.d_reg[254] ),
    .A(\u_inv.d_next[254] ),
    .X(_04455_));
 sg13g2_xnor2_1 _30178_ (.Y(_04456_),
    .A(\u_inv.d_next[254] ),
    .B(\u_inv.d_reg[254] ));
 sg13g2_nor2_1 _30179_ (.A(_04452_),
    .B(_04455_),
    .Y(_04457_));
 sg13g2_nor2_1 _30180_ (.A(\u_inv.d_next[253] ),
    .B(\u_inv.d_reg[253] ),
    .Y(_04458_));
 sg13g2_nand2_1 _30181_ (.Y(_04459_),
    .A(\u_inv.d_next[253] ),
    .B(\u_inv.d_reg[253] ));
 sg13g2_nor2b_2 _30182_ (.A(_04458_),
    .B_N(_04459_),
    .Y(_04460_));
 sg13g2_nand2_1 _30183_ (.Y(_04461_),
    .A(\u_inv.d_next[252] ),
    .B(\u_inv.d_reg[252] ));
 sg13g2_xnor2_1 _30184_ (.Y(_04462_),
    .A(\u_inv.d_next[252] ),
    .B(\u_inv.d_reg[252] ));
 sg13g2_inv_1 _30185_ (.Y(_04463_),
    .A(_04462_));
 sg13g2_nor2_1 _30186_ (.A(_04460_),
    .B(_04463_),
    .Y(_04464_));
 sg13g2_inv_1 _30187_ (.Y(_04465_),
    .A(_04464_));
 sg13g2_nand2_1 _30188_ (.Y(_04466_),
    .A(_04457_),
    .B(_04464_));
 sg13g2_nand2_1 _30189_ (.Y(_04467_),
    .A(\u_inv.d_next[250] ),
    .B(\u_inv.d_reg[250] ));
 sg13g2_xor2_1 _30190_ (.B(\u_inv.d_reg[250] ),
    .A(\u_inv.d_next[250] ),
    .X(_04468_));
 sg13g2_nor2_1 _30191_ (.A(\u_inv.d_next[251] ),
    .B(\u_inv.d_reg[251] ),
    .Y(_04469_));
 sg13g2_xor2_1 _30192_ (.B(\u_inv.d_reg[251] ),
    .A(\u_inv.d_next[251] ),
    .X(_04470_));
 sg13g2_nor2_1 _30193_ (.A(_04468_),
    .B(_04470_),
    .Y(_04471_));
 sg13g2_nor2_1 _30194_ (.A(\u_inv.d_next[249] ),
    .B(\u_inv.d_reg[249] ),
    .Y(_04472_));
 sg13g2_nand2_1 _30195_ (.Y(_04473_),
    .A(\u_inv.d_next[249] ),
    .B(\u_inv.d_reg[249] ));
 sg13g2_nor2b_2 _30196_ (.A(_04472_),
    .B_N(_04473_),
    .Y(_04474_));
 sg13g2_nand2b_2 _30197_ (.Y(_04475_),
    .B(_04473_),
    .A_N(_04472_));
 sg13g2_nand2_1 _30198_ (.Y(_04476_),
    .A(\u_inv.d_next[248] ),
    .B(\u_inv.d_reg[248] ));
 sg13g2_xor2_1 _30199_ (.B(\u_inv.d_reg[248] ),
    .A(\u_inv.d_next[248] ),
    .X(_04477_));
 sg13g2_xnor2_1 _30200_ (.Y(_04478_),
    .A(\u_inv.d_next[248] ),
    .B(\u_inv.d_reg[248] ));
 sg13g2_nor2_1 _30201_ (.A(_04474_),
    .B(_04477_),
    .Y(_04479_));
 sg13g2_nand2_1 _30202_ (.Y(_04480_),
    .A(_04471_),
    .B(_04479_));
 sg13g2_inv_1 _30203_ (.Y(_04481_),
    .A(_04480_));
 sg13g2_nor2_1 _30204_ (.A(_04466_),
    .B(_04480_),
    .Y(_04482_));
 sg13g2_nor2_1 _30205_ (.A(\u_inv.d_next[245] ),
    .B(\u_inv.d_reg[245] ),
    .Y(_04483_));
 sg13g2_nand2_1 _30206_ (.Y(_04484_),
    .A(\u_inv.d_next[245] ),
    .B(\u_inv.d_reg[245] ));
 sg13g2_nand2b_2 _30207_ (.Y(_04485_),
    .B(_04484_),
    .A_N(_04483_));
 sg13g2_nand2_1 _30208_ (.Y(_04486_),
    .A(\u_inv.d_next[244] ),
    .B(\u_inv.d_reg[244] ));
 sg13g2_inv_1 _30209_ (.Y(_04487_),
    .A(_04486_));
 sg13g2_or2_1 _30210_ (.X(_04488_),
    .B(\u_inv.d_reg[244] ),
    .A(\u_inv.d_next[244] ));
 sg13g2_nand2_2 _30211_ (.Y(_04489_),
    .A(_04486_),
    .B(_04488_));
 sg13g2_nand2_1 _30212_ (.Y(_04490_),
    .A(_04485_),
    .B(_04489_));
 sg13g2_inv_1 _30213_ (.Y(_04491_),
    .A(_04490_));
 sg13g2_xor2_1 _30214_ (.B(\u_inv.d_reg[246] ),
    .A(\u_inv.d_next[246] ),
    .X(_04492_));
 sg13g2_xor2_1 _30215_ (.B(\u_inv.d_reg[247] ),
    .A(\u_inv.d_next[247] ),
    .X(_04493_));
 sg13g2_xnor2_1 _30216_ (.Y(_04494_),
    .A(\u_inv.d_next[247] ),
    .B(\u_inv.d_reg[247] ));
 sg13g2_nor3_1 _30217_ (.A(_04490_),
    .B(_04492_),
    .C(_04493_),
    .Y(_04495_));
 sg13g2_nor2_1 _30218_ (.A(\u_inv.d_next[243] ),
    .B(\u_inv.d_reg[243] ),
    .Y(_04496_));
 sg13g2_nand2_1 _30219_ (.Y(_04497_),
    .A(\u_inv.d_next[243] ),
    .B(\u_inv.d_reg[243] ));
 sg13g2_nor2b_1 _30220_ (.A(_04496_),
    .B_N(_04497_),
    .Y(_04498_));
 sg13g2_nand2b_2 _30221_ (.Y(_04499_),
    .B(_04497_),
    .A_N(_04496_));
 sg13g2_nand2_1 _30222_ (.Y(_04500_),
    .A(\u_inv.d_next[242] ),
    .B(\u_inv.d_reg[242] ));
 sg13g2_xor2_1 _30223_ (.B(\u_inv.d_reg[242] ),
    .A(\u_inv.d_next[242] ),
    .X(_04501_));
 sg13g2_inv_1 _30224_ (.Y(_04502_),
    .A(_04501_));
 sg13g2_nor2_1 _30225_ (.A(_04498_),
    .B(_04501_),
    .Y(_04503_));
 sg13g2_xnor2_1 _30226_ (.Y(_04504_),
    .A(\u_inv.d_next[241] ),
    .B(\u_inv.d_reg[241] ));
 sg13g2_inv_1 _30227_ (.Y(_04505_),
    .A(_04504_));
 sg13g2_nand2_1 _30228_ (.Y(_04506_),
    .A(\u_inv.d_next[240] ),
    .B(net5865));
 sg13g2_xor2_1 _30229_ (.B(net5865),
    .A(\u_inv.d_next[240] ),
    .X(_04507_));
 sg13g2_nor2_1 _30230_ (.A(_04505_),
    .B(_04507_),
    .Y(_04508_));
 sg13g2_inv_1 _30231_ (.Y(_04509_),
    .A(_04508_));
 sg13g2_and2_1 _30232_ (.A(_04503_),
    .B(_04508_),
    .X(_04510_));
 sg13g2_inv_1 _30233_ (.Y(_04511_),
    .A(_04510_));
 sg13g2_and2_1 _30234_ (.A(_04495_),
    .B(_04510_),
    .X(_04512_));
 sg13g2_inv_1 _30235_ (.Y(_04513_),
    .A(_04512_));
 sg13g2_and2_1 _30236_ (.A(_04482_),
    .B(_04512_),
    .X(_04514_));
 sg13g2_xor2_1 _30237_ (.B(\u_inv.d_reg[239] ),
    .A(\u_inv.d_next[239] ),
    .X(_04515_));
 sg13g2_xnor2_1 _30238_ (.Y(_04516_),
    .A(\u_inv.d_next[239] ),
    .B(\u_inv.d_reg[239] ));
 sg13g2_nand2_1 _30239_ (.Y(_04517_),
    .A(\u_inv.d_next[238] ),
    .B(\u_inv.d_reg[238] ));
 sg13g2_xnor2_1 _30240_ (.Y(_04518_),
    .A(\u_inv.d_next[238] ),
    .B(\u_inv.d_reg[238] ));
 sg13g2_inv_1 _30241_ (.Y(_04519_),
    .A(_04518_));
 sg13g2_nand2_1 _30242_ (.Y(_04520_),
    .A(_04516_),
    .B(_04518_));
 sg13g2_nor2_1 _30243_ (.A(\u_inv.d_next[237] ),
    .B(\u_inv.d_reg[237] ),
    .Y(_04521_));
 sg13g2_nand2_1 _30244_ (.Y(_04522_),
    .A(\u_inv.d_next[237] ),
    .B(\u_inv.d_reg[237] ));
 sg13g2_nand2b_2 _30245_ (.Y(_04523_),
    .B(_04522_),
    .A_N(_04521_));
 sg13g2_nand2_1 _30246_ (.Y(_04524_),
    .A(\u_inv.d_next[236] ),
    .B(\u_inv.d_reg[236] ));
 sg13g2_xor2_1 _30247_ (.B(\u_inv.d_reg[236] ),
    .A(\u_inv.d_next[236] ),
    .X(_04525_));
 sg13g2_xnor2_1 _30248_ (.Y(_04526_),
    .A(\u_inv.d_next[236] ),
    .B(\u_inv.d_reg[236] ));
 sg13g2_nand2_1 _30249_ (.Y(_04527_),
    .A(_04523_),
    .B(_04526_));
 sg13g2_inv_1 _30250_ (.Y(_04528_),
    .A(_04527_));
 sg13g2_nor2_1 _30251_ (.A(_04520_),
    .B(_04527_),
    .Y(_04529_));
 sg13g2_or2_1 _30252_ (.X(_04530_),
    .B(\u_inv.d_reg[235] ),
    .A(\u_inv.d_next[235] ));
 sg13g2_nand2_1 _30253_ (.Y(_04531_),
    .A(\u_inv.d_next[235] ),
    .B(\u_inv.d_reg[235] ));
 sg13g2_and2_1 _30254_ (.A(_04530_),
    .B(_04531_),
    .X(_04532_));
 sg13g2_nand2_1 _30255_ (.Y(_04533_),
    .A(_04530_),
    .B(_04531_));
 sg13g2_nand2_1 _30256_ (.Y(_04534_),
    .A(\u_inv.d_next[234] ),
    .B(\u_inv.d_reg[234] ));
 sg13g2_inv_1 _30257_ (.Y(_04535_),
    .A(_04534_));
 sg13g2_xor2_1 _30258_ (.B(\u_inv.d_reg[234] ),
    .A(\u_inv.d_next[234] ),
    .X(_04536_));
 sg13g2_inv_1 _30259_ (.Y(_04537_),
    .A(_04536_));
 sg13g2_nor2_1 _30260_ (.A(_04532_),
    .B(_04536_),
    .Y(_04538_));
 sg13g2_xor2_1 _30261_ (.B(\u_inv.d_reg[233] ),
    .A(\u_inv.d_next[233] ),
    .X(_04539_));
 sg13g2_xnor2_1 _30262_ (.Y(_04540_),
    .A(\u_inv.d_next[233] ),
    .B(\u_inv.d_reg[233] ));
 sg13g2_xor2_1 _30263_ (.B(\u_inv.d_reg[232] ),
    .A(\u_inv.d_next[232] ),
    .X(_04541_));
 sg13g2_xnor2_1 _30264_ (.Y(_04542_),
    .A(\u_inv.d_next[232] ),
    .B(\u_inv.d_reg[232] ));
 sg13g2_nor2_1 _30265_ (.A(_04539_),
    .B(_04541_),
    .Y(_04543_));
 sg13g2_inv_1 _30266_ (.Y(_04544_),
    .A(_04543_));
 sg13g2_and2_1 _30267_ (.A(_04538_),
    .B(_04543_),
    .X(_04545_));
 sg13g2_inv_1 _30268_ (.Y(_04546_),
    .A(_04545_));
 sg13g2_and2_1 _30269_ (.A(_04529_),
    .B(_04545_),
    .X(_04547_));
 sg13g2_xor2_1 _30270_ (.B(\u_inv.d_reg[229] ),
    .A(\u_inv.d_next[229] ),
    .X(_04548_));
 sg13g2_and2_1 _30271_ (.A(\u_inv.d_next[228] ),
    .B(\u_inv.d_reg[228] ),
    .X(_04549_));
 sg13g2_xor2_1 _30272_ (.B(\u_inv.d_reg[228] ),
    .A(\u_inv.d_next[228] ),
    .X(_04550_));
 sg13g2_nor2_1 _30273_ (.A(_04548_),
    .B(_04550_),
    .Y(_04551_));
 sg13g2_inv_1 _30274_ (.Y(_04552_),
    .A(_04551_));
 sg13g2_nand2_1 _30275_ (.Y(_04553_),
    .A(\u_inv.d_next[230] ),
    .B(\u_inv.d_reg[230] ));
 sg13g2_xnor2_1 _30276_ (.Y(_04554_),
    .A(\u_inv.d_next[230] ),
    .B(\u_inv.d_reg[230] ));
 sg13g2_nor2_1 _30277_ (.A(\u_inv.d_next[231] ),
    .B(\u_inv.d_reg[231] ),
    .Y(_04555_));
 sg13g2_xnor2_1 _30278_ (.Y(_04556_),
    .A(\u_inv.d_next[231] ),
    .B(\u_inv.d_reg[231] ));
 sg13g2_and2_1 _30279_ (.A(_04554_),
    .B(_04556_),
    .X(_04557_));
 sg13g2_nand2_1 _30280_ (.Y(_04558_),
    .A(_04551_),
    .B(_04557_));
 sg13g2_xor2_1 _30281_ (.B(\u_inv.d_reg[227] ),
    .A(\u_inv.d_next[227] ),
    .X(_04559_));
 sg13g2_xnor2_1 _30282_ (.Y(_04560_),
    .A(\u_inv.d_next[227] ),
    .B(\u_inv.d_reg[227] ));
 sg13g2_nand2_1 _30283_ (.Y(_04561_),
    .A(\u_inv.d_next[226] ),
    .B(\u_inv.d_reg[226] ));
 sg13g2_xnor2_1 _30284_ (.Y(_04562_),
    .A(\u_inv.d_next[226] ),
    .B(\u_inv.d_reg[226] ));
 sg13g2_inv_1 _30285_ (.Y(_04563_),
    .A(_04562_));
 sg13g2_nand2_1 _30286_ (.Y(_04564_),
    .A(net5875),
    .B(\u_inv.d_reg[225] ));
 sg13g2_nor2_1 _30287_ (.A(net5875),
    .B(\u_inv.d_reg[225] ),
    .Y(_04565_));
 sg13g2_xor2_1 _30288_ (.B(\u_inv.d_reg[225] ),
    .A(net5875),
    .X(_04566_));
 sg13g2_xnor2_1 _30289_ (.Y(_04567_),
    .A(net5875),
    .B(\u_inv.d_reg[225] ));
 sg13g2_nand2_1 _30290_ (.Y(_04568_),
    .A(\u_inv.d_next[224] ),
    .B(\u_inv.d_reg[224] ));
 sg13g2_xor2_1 _30291_ (.B(\u_inv.d_reg[224] ),
    .A(\u_inv.d_next[224] ),
    .X(_04569_));
 sg13g2_xnor2_1 _30292_ (.Y(_04570_),
    .A(\u_inv.d_next[224] ),
    .B(\u_inv.d_reg[224] ));
 sg13g2_nor2_1 _30293_ (.A(_04566_),
    .B(_04569_),
    .Y(_04571_));
 sg13g2_nand3_1 _30294_ (.B(_04562_),
    .C(_04571_),
    .A(_04560_),
    .Y(_04572_));
 sg13g2_inv_1 _30295_ (.Y(_04573_),
    .A(_04572_));
 sg13g2_nor2_1 _30296_ (.A(_04558_),
    .B(_04572_),
    .Y(_04574_));
 sg13g2_and2_1 _30297_ (.A(_04547_),
    .B(_04574_),
    .X(_04575_));
 sg13g2_nand2_2 _30298_ (.Y(_04576_),
    .A(_04514_),
    .B(_04575_));
 sg13g2_nand2_1 _30299_ (.Y(_04577_),
    .A(\u_inv.d_next[223] ),
    .B(\u_inv.d_reg[223] ));
 sg13g2_xnor2_1 _30300_ (.Y(_04578_),
    .A(\u_inv.d_next[223] ),
    .B(\u_inv.d_reg[223] ));
 sg13g2_nor2_1 _30301_ (.A(_14180_),
    .B(_14587_),
    .Y(_04579_));
 sg13g2_xor2_1 _30302_ (.B(\u_inv.d_reg[222] ),
    .A(\u_inv.d_next[222] ),
    .X(_04580_));
 sg13g2_xnor2_1 _30303_ (.Y(_04581_),
    .A(\u_inv.d_next[222] ),
    .B(\u_inv.d_reg[222] ));
 sg13g2_nand2_1 _30304_ (.Y(_04582_),
    .A(_04578_),
    .B(_04581_));
 sg13g2_xor2_1 _30305_ (.B(\u_inv.d_reg[221] ),
    .A(\u_inv.d_next[221] ),
    .X(_04583_));
 sg13g2_xnor2_1 _30306_ (.Y(_04584_),
    .A(\u_inv.d_next[221] ),
    .B(\u_inv.d_reg[221] ));
 sg13g2_nand2_1 _30307_ (.Y(_04585_),
    .A(\u_inv.d_next[220] ),
    .B(\u_inv.d_reg[220] ));
 sg13g2_xor2_1 _30308_ (.B(\u_inv.d_reg[220] ),
    .A(\u_inv.d_next[220] ),
    .X(_04586_));
 sg13g2_xnor2_1 _30309_ (.Y(_04587_),
    .A(\u_inv.d_next[220] ),
    .B(\u_inv.d_reg[220] ));
 sg13g2_nand2_1 _30310_ (.Y(_04588_),
    .A(_04584_),
    .B(_04587_));
 sg13g2_nor2_1 _30311_ (.A(_04582_),
    .B(_04588_),
    .Y(_04589_));
 sg13g2_nor2_1 _30312_ (.A(\u_inv.d_next[219] ),
    .B(\u_inv.d_reg[219] ),
    .Y(_04590_));
 sg13g2_xor2_1 _30313_ (.B(\u_inv.d_reg[219] ),
    .A(\u_inv.d_next[219] ),
    .X(_04591_));
 sg13g2_xnor2_1 _30314_ (.Y(_04592_),
    .A(\u_inv.d_next[219] ),
    .B(\u_inv.d_reg[219] ));
 sg13g2_nand2_1 _30315_ (.Y(_04593_),
    .A(\u_inv.d_next[218] ),
    .B(\u_inv.d_reg[218] ));
 sg13g2_xor2_1 _30316_ (.B(\u_inv.d_reg[218] ),
    .A(\u_inv.d_next[218] ),
    .X(_04594_));
 sg13g2_xnor2_1 _30317_ (.Y(_04595_),
    .A(\u_inv.d_next[218] ),
    .B(\u_inv.d_reg[218] ));
 sg13g2_nor2_1 _30318_ (.A(_04591_),
    .B(_04594_),
    .Y(_04596_));
 sg13g2_nor2_1 _30319_ (.A(\u_inv.d_next[217] ),
    .B(\u_inv.d_reg[217] ),
    .Y(_04597_));
 sg13g2_nand2_1 _30320_ (.Y(_04598_),
    .A(\u_inv.d_next[217] ),
    .B(\u_inv.d_reg[217] ));
 sg13g2_nor2b_2 _30321_ (.A(_04597_),
    .B_N(_04598_),
    .Y(_04599_));
 sg13g2_nand2_1 _30322_ (.Y(_04600_),
    .A(\u_inv.d_next[216] ),
    .B(\u_inv.d_reg[216] ));
 sg13g2_xor2_1 _30323_ (.B(\u_inv.d_reg[216] ),
    .A(\u_inv.d_next[216] ),
    .X(_04601_));
 sg13g2_xnor2_1 _30324_ (.Y(_04602_),
    .A(\u_inv.d_next[216] ),
    .B(\u_inv.d_reg[216] ));
 sg13g2_nor2_1 _30325_ (.A(_04599_),
    .B(_04601_),
    .Y(_04603_));
 sg13g2_and2_1 _30326_ (.A(_04596_),
    .B(_04603_),
    .X(_04604_));
 sg13g2_nand2_1 _30327_ (.Y(_04605_),
    .A(_04589_),
    .B(_04604_));
 sg13g2_xor2_1 _30328_ (.B(\u_inv.d_reg[213] ),
    .A(\u_inv.d_next[213] ),
    .X(_04606_));
 sg13g2_xnor2_1 _30329_ (.Y(_04607_),
    .A(\u_inv.d_next[213] ),
    .B(\u_inv.d_reg[213] ));
 sg13g2_and2_1 _30330_ (.A(\u_inv.d_next[212] ),
    .B(\u_inv.d_reg[212] ),
    .X(_04608_));
 sg13g2_or2_1 _30331_ (.X(_04609_),
    .B(\u_inv.d_reg[212] ),
    .A(\u_inv.d_next[212] ));
 sg13g2_nand2b_2 _30332_ (.Y(_04610_),
    .B(_04609_),
    .A_N(_04608_));
 sg13g2_and2_1 _30333_ (.A(_04607_),
    .B(_04610_),
    .X(_04611_));
 sg13g2_nand2_1 _30334_ (.Y(_04612_),
    .A(\u_inv.d_next[214] ),
    .B(\u_inv.d_reg[214] ));
 sg13g2_xor2_1 _30335_ (.B(\u_inv.d_reg[214] ),
    .A(\u_inv.d_next[214] ),
    .X(_04613_));
 sg13g2_xnor2_1 _30336_ (.Y(_04614_),
    .A(\u_inv.d_next[214] ),
    .B(\u_inv.d_reg[214] ));
 sg13g2_nor2_1 _30337_ (.A(\u_inv.d_next[215] ),
    .B(\u_inv.d_reg[215] ),
    .Y(_04615_));
 sg13g2_xor2_1 _30338_ (.B(\u_inv.d_reg[215] ),
    .A(\u_inv.d_next[215] ),
    .X(_04616_));
 sg13g2_xnor2_1 _30339_ (.Y(_04617_),
    .A(\u_inv.d_next[215] ),
    .B(\u_inv.d_reg[215] ));
 sg13g2_nor2_1 _30340_ (.A(_04613_),
    .B(_04616_),
    .Y(_04618_));
 sg13g2_nand2_1 _30341_ (.Y(_04619_),
    .A(_04611_),
    .B(_04618_));
 sg13g2_nand2_1 _30342_ (.Y(_04620_),
    .A(\u_inv.d_next[211] ),
    .B(\u_inv.d_reg[211] ));
 sg13g2_nor2_1 _30343_ (.A(\u_inv.d_next[211] ),
    .B(\u_inv.d_reg[211] ),
    .Y(_04621_));
 sg13g2_xnor2_1 _30344_ (.Y(_04622_),
    .A(\u_inv.d_next[211] ),
    .B(\u_inv.d_reg[211] ));
 sg13g2_nand2_1 _30345_ (.Y(_04623_),
    .A(\u_inv.d_next[210] ),
    .B(\u_inv.d_reg[210] ));
 sg13g2_xnor2_1 _30346_ (.Y(_04624_),
    .A(\u_inv.d_next[210] ),
    .B(\u_inv.d_reg[210] ));
 sg13g2_and2_1 _30347_ (.A(_04622_),
    .B(_04624_),
    .X(_04625_));
 sg13g2_xor2_1 _30348_ (.B(\u_inv.d_reg[209] ),
    .A(\u_inv.d_next[209] ),
    .X(_04626_));
 sg13g2_xnor2_1 _30349_ (.Y(_04627_),
    .A(\u_inv.d_next[209] ),
    .B(\u_inv.d_reg[209] ));
 sg13g2_xor2_1 _30350_ (.B(\u_inv.d_reg[208] ),
    .A(\u_inv.d_next[208] ),
    .X(_04628_));
 sg13g2_xnor2_1 _30351_ (.Y(_04629_),
    .A(\u_inv.d_next[208] ),
    .B(\u_inv.d_reg[208] ));
 sg13g2_nand3_1 _30352_ (.B(_04627_),
    .C(_04629_),
    .A(_04625_),
    .Y(_04630_));
 sg13g2_or2_1 _30353_ (.X(_04631_),
    .B(_04630_),
    .A(_04619_));
 sg13g2_nor2_1 _30354_ (.A(_04605_),
    .B(_04631_),
    .Y(_04632_));
 sg13g2_xor2_1 _30355_ (.B(\u_inv.d_reg[207] ),
    .A(\u_inv.d_next[207] ),
    .X(_04633_));
 sg13g2_xnor2_1 _30356_ (.Y(_04634_),
    .A(\u_inv.d_next[207] ),
    .B(\u_inv.d_reg[207] ));
 sg13g2_nand2_1 _30357_ (.Y(_04635_),
    .A(\u_inv.d_next[206] ),
    .B(\u_inv.d_reg[206] ));
 sg13g2_xor2_1 _30358_ (.B(\u_inv.d_reg[206] ),
    .A(\u_inv.d_next[206] ),
    .X(_04636_));
 sg13g2_nor2_1 _30359_ (.A(_04633_),
    .B(_04636_),
    .Y(_04637_));
 sg13g2_nand2_1 _30360_ (.Y(_04638_),
    .A(_14186_),
    .B(_14604_));
 sg13g2_nand2_1 _30361_ (.Y(_04639_),
    .A(\u_inv.d_next[205] ),
    .B(\u_inv.d_reg[205] ));
 sg13g2_nand2_2 _30362_ (.Y(_04640_),
    .A(_04638_),
    .B(_04639_));
 sg13g2_and2_1 _30363_ (.A(\u_inv.d_next[204] ),
    .B(\u_inv.d_reg[204] ),
    .X(_04641_));
 sg13g2_xnor2_1 _30364_ (.Y(_04642_),
    .A(\u_inv.d_next[204] ),
    .B(\u_inv.d_reg[204] ));
 sg13g2_inv_2 _30365_ (.Y(_04643_),
    .A(_04642_));
 sg13g2_and2_1 _30366_ (.A(_04640_),
    .B(_04642_),
    .X(_04644_));
 sg13g2_nand2_1 _30367_ (.Y(_04645_),
    .A(_04637_),
    .B(_04644_));
 sg13g2_xnor2_1 _30368_ (.Y(_04646_),
    .A(\u_inv.d_next[203] ),
    .B(\u_inv.d_reg[203] ));
 sg13g2_nand2_1 _30369_ (.Y(_04647_),
    .A(\u_inv.d_next[202] ),
    .B(\u_inv.d_reg[202] ));
 sg13g2_xnor2_1 _30370_ (.Y(_04648_),
    .A(\u_inv.d_next[202] ),
    .B(\u_inv.d_reg[202] ));
 sg13g2_nand2_1 _30371_ (.Y(_04649_),
    .A(_04646_),
    .B(_04648_));
 sg13g2_nor2_1 _30372_ (.A(\u_inv.d_next[201] ),
    .B(\u_inv.d_reg[201] ),
    .Y(_04650_));
 sg13g2_nand2_1 _30373_ (.Y(_04651_),
    .A(\u_inv.d_next[201] ),
    .B(\u_inv.d_reg[201] ));
 sg13g2_nor2b_2 _30374_ (.A(_04650_),
    .B_N(_04651_),
    .Y(_04652_));
 sg13g2_nand2b_1 _30375_ (.Y(_04653_),
    .B(_04651_),
    .A_N(_04650_));
 sg13g2_nand2_1 _30376_ (.Y(_04654_),
    .A(\u_inv.d_next[200] ),
    .B(\u_inv.d_reg[200] ));
 sg13g2_xor2_1 _30377_ (.B(\u_inv.d_reg[200] ),
    .A(\u_inv.d_next[200] ),
    .X(_04655_));
 sg13g2_or2_1 _30378_ (.X(_04656_),
    .B(_04655_),
    .A(_04652_));
 sg13g2_or2_1 _30379_ (.X(_04657_),
    .B(_04656_),
    .A(_04649_));
 sg13g2_nor2_1 _30380_ (.A(_04645_),
    .B(_04657_),
    .Y(_04658_));
 sg13g2_nor2_1 _30381_ (.A(\u_inv.d_next[197] ),
    .B(\u_inv.d_reg[197] ),
    .Y(_04659_));
 sg13g2_nand2_1 _30382_ (.Y(_04660_),
    .A(\u_inv.d_next[197] ),
    .B(\u_inv.d_reg[197] ));
 sg13g2_nand2b_2 _30383_ (.Y(_04661_),
    .B(_04660_),
    .A_N(_04659_));
 sg13g2_nand2_1 _30384_ (.Y(_04662_),
    .A(\u_inv.d_next[196] ),
    .B(\u_inv.d_reg[196] ));
 sg13g2_xnor2_1 _30385_ (.Y(_04663_),
    .A(\u_inv.d_next[196] ),
    .B(\u_inv.d_reg[196] ));
 sg13g2_nand2_1 _30386_ (.Y(_04664_),
    .A(_04661_),
    .B(_04663_));
 sg13g2_inv_1 _30387_ (.Y(_04665_),
    .A(_04664_));
 sg13g2_xor2_1 _30388_ (.B(\u_inv.d_reg[199] ),
    .A(\u_inv.d_next[199] ),
    .X(_04666_));
 sg13g2_xnor2_1 _30389_ (.Y(_04667_),
    .A(\u_inv.d_next[199] ),
    .B(\u_inv.d_reg[199] ));
 sg13g2_nand2_1 _30390_ (.Y(_04668_),
    .A(\u_inv.d_next[198] ),
    .B(\u_inv.d_reg[198] ));
 sg13g2_xor2_1 _30391_ (.B(\u_inv.d_reg[198] ),
    .A(\u_inv.d_next[198] ),
    .X(_04669_));
 sg13g2_nor3_1 _30392_ (.A(_04664_),
    .B(_04666_),
    .C(_04669_),
    .Y(_04670_));
 sg13g2_xnor2_1 _30393_ (.Y(_04671_),
    .A(\u_inv.d_next[193] ),
    .B(\u_inv.d_reg[193] ));
 sg13g2_nand2_1 _30394_ (.Y(_04672_),
    .A(\u_inv.d_next[192] ),
    .B(\u_inv.d_reg[192] ));
 sg13g2_xnor2_1 _30395_ (.Y(_04673_),
    .A(\u_inv.d_next[192] ),
    .B(\u_inv.d_reg[192] ));
 sg13g2_nand2_1 _30396_ (.Y(_04674_),
    .A(_04671_),
    .B(_04673_));
 sg13g2_xnor2_1 _30397_ (.Y(_04675_),
    .A(\u_inv.d_next[195] ),
    .B(\u_inv.d_reg[195] ));
 sg13g2_nand2_1 _30398_ (.Y(_04676_),
    .A(\u_inv.d_next[194] ),
    .B(\u_inv.d_reg[194] ));
 sg13g2_xnor2_1 _30399_ (.Y(_04677_),
    .A(\u_inv.d_next[194] ),
    .B(\u_inv.d_reg[194] ));
 sg13g2_and2_1 _30400_ (.A(_04675_),
    .B(_04677_),
    .X(_04678_));
 sg13g2_nor2b_1 _30401_ (.A(_04674_),
    .B_N(_04678_),
    .Y(_04679_));
 sg13g2_inv_1 _30402_ (.Y(_04680_),
    .A(_04679_));
 sg13g2_and3_2 _30403_ (.X(_04681_),
    .A(_04658_),
    .B(_04670_),
    .C(_04679_));
 sg13g2_nand2_1 _30404_ (.Y(_04682_),
    .A(_04632_),
    .B(_04681_));
 sg13g2_nor2_1 _30405_ (.A(_04576_),
    .B(_04682_),
    .Y(_04683_));
 sg13g2_inv_1 _30406_ (.Y(_04684_),
    .A(_04683_));
 sg13g2_nor2_1 _30407_ (.A(\u_inv.d_next[191] ),
    .B(\u_inv.d_reg[191] ),
    .Y(_04685_));
 sg13g2_nand2_1 _30408_ (.Y(_04686_),
    .A(\u_inv.d_next[191] ),
    .B(\u_inv.d_reg[191] ));
 sg13g2_nand2b_2 _30409_ (.Y(_04687_),
    .B(_04686_),
    .A_N(_04685_));
 sg13g2_nand2_1 _30410_ (.Y(_04688_),
    .A(\u_inv.d_next[190] ),
    .B(\u_inv.d_reg[190] ));
 sg13g2_xnor2_1 _30411_ (.Y(_04689_),
    .A(\u_inv.d_next[190] ),
    .B(\u_inv.d_reg[190] ));
 sg13g2_nand2_1 _30412_ (.Y(_04690_),
    .A(_04687_),
    .B(_04689_));
 sg13g2_xnor2_1 _30413_ (.Y(_04691_),
    .A(\u_inv.d_next[189] ),
    .B(\u_inv.d_reg[189] ));
 sg13g2_inv_1 _30414_ (.Y(_04692_),
    .A(_04691_));
 sg13g2_nand2_1 _30415_ (.Y(_04693_),
    .A(\u_inv.d_next[188] ),
    .B(\u_inv.d_reg[188] ));
 sg13g2_xnor2_1 _30416_ (.Y(_04694_),
    .A(\u_inv.d_next[188] ),
    .B(\u_inv.d_reg[188] ));
 sg13g2_nand2_1 _30417_ (.Y(_04695_),
    .A(_04691_),
    .B(_04694_));
 sg13g2_nor2_1 _30418_ (.A(_04690_),
    .B(_04695_),
    .Y(_04696_));
 sg13g2_nor2_1 _30419_ (.A(\u_inv.d_next[187] ),
    .B(\u_inv.d_reg[187] ),
    .Y(_04697_));
 sg13g2_xor2_1 _30420_ (.B(\u_inv.d_reg[187] ),
    .A(\u_inv.d_next[187] ),
    .X(_04698_));
 sg13g2_xnor2_1 _30421_ (.Y(_04699_),
    .A(\u_inv.d_next[187] ),
    .B(\u_inv.d_reg[187] ));
 sg13g2_nand2_1 _30422_ (.Y(_04700_),
    .A(\u_inv.d_next[186] ),
    .B(\u_inv.d_reg[186] ));
 sg13g2_xor2_1 _30423_ (.B(\u_inv.d_reg[186] ),
    .A(\u_inv.d_next[186] ),
    .X(_04701_));
 sg13g2_nor2_1 _30424_ (.A(_04698_),
    .B(_04701_),
    .Y(_04702_));
 sg13g2_nor2_1 _30425_ (.A(\u_inv.d_next[185] ),
    .B(\u_inv.d_reg[185] ),
    .Y(_04703_));
 sg13g2_nand2_1 _30426_ (.Y(_04704_),
    .A(\u_inv.d_next[185] ),
    .B(\u_inv.d_reg[185] ));
 sg13g2_nor2b_2 _30427_ (.A(_04703_),
    .B_N(_04704_),
    .Y(_04705_));
 sg13g2_nand2b_1 _30428_ (.Y(_04706_),
    .B(_04704_),
    .A_N(_04703_));
 sg13g2_nand2_1 _30429_ (.Y(_04707_),
    .A(\u_inv.d_next[184] ),
    .B(net5866));
 sg13g2_xor2_1 _30430_ (.B(net5866),
    .A(\u_inv.d_next[184] ),
    .X(_04708_));
 sg13g2_xnor2_1 _30431_ (.Y(_04709_),
    .A(\u_inv.d_next[184] ),
    .B(net5866));
 sg13g2_nor2_1 _30432_ (.A(_04705_),
    .B(_04708_),
    .Y(_04710_));
 sg13g2_and2_1 _30433_ (.A(_04702_),
    .B(_04710_),
    .X(_04711_));
 sg13g2_nand2_2 _30434_ (.Y(_04712_),
    .A(_04696_),
    .B(_04711_));
 sg13g2_xnor2_1 _30435_ (.Y(_04713_),
    .A(\u_inv.d_next[181] ),
    .B(\u_inv.d_reg[181] ));
 sg13g2_and2_1 _30436_ (.A(\u_inv.d_next[180] ),
    .B(\u_inv.d_reg[180] ),
    .X(_04714_));
 sg13g2_xor2_1 _30437_ (.B(\u_inv.d_reg[180] ),
    .A(\u_inv.d_next[180] ),
    .X(_04715_));
 sg13g2_xnor2_1 _30438_ (.Y(_04716_),
    .A(\u_inv.d_next[180] ),
    .B(\u_inv.d_reg[180] ));
 sg13g2_nand2_1 _30439_ (.Y(_04717_),
    .A(_04713_),
    .B(_04716_));
 sg13g2_xor2_1 _30440_ (.B(\u_inv.d_reg[183] ),
    .A(\u_inv.d_next[183] ),
    .X(_04718_));
 sg13g2_xnor2_1 _30441_ (.Y(_04719_),
    .A(\u_inv.d_next[183] ),
    .B(\u_inv.d_reg[183] ));
 sg13g2_nand2_1 _30442_ (.Y(_04720_),
    .A(\u_inv.d_next[182] ),
    .B(\u_inv.d_reg[182] ));
 sg13g2_xor2_1 _30443_ (.B(\u_inv.d_reg[182] ),
    .A(\u_inv.d_next[182] ),
    .X(_04721_));
 sg13g2_nor3_1 _30444_ (.A(_04717_),
    .B(_04718_),
    .C(_04721_),
    .Y(_04722_));
 sg13g2_xnor2_1 _30445_ (.Y(_04723_),
    .A(\u_inv.d_next[179] ),
    .B(\u_inv.d_reg[179] ));
 sg13g2_nand2_1 _30446_ (.Y(_04724_),
    .A(\u_inv.d_next[178] ),
    .B(\u_inv.d_reg[178] ));
 sg13g2_xnor2_1 _30447_ (.Y(_04725_),
    .A(\u_inv.d_next[178] ),
    .B(\u_inv.d_reg[178] ));
 sg13g2_and2_1 _30448_ (.A(_04723_),
    .B(_04725_),
    .X(_04726_));
 sg13g2_xor2_1 _30449_ (.B(\u_inv.d_reg[177] ),
    .A(\u_inv.d_next[177] ),
    .X(_04727_));
 sg13g2_and2_1 _30450_ (.A(\u_inv.d_next[176] ),
    .B(\u_inv.d_reg[176] ),
    .X(_04728_));
 sg13g2_xor2_1 _30451_ (.B(\u_inv.d_reg[176] ),
    .A(\u_inv.d_next[176] ),
    .X(_04729_));
 sg13g2_nor2_1 _30452_ (.A(_04727_),
    .B(_04729_),
    .Y(_04730_));
 sg13g2_or2_1 _30453_ (.X(_04731_),
    .B(_04729_),
    .A(_04727_));
 sg13g2_nand3_1 _30454_ (.B(_04726_),
    .C(_04730_),
    .A(_04722_),
    .Y(_04732_));
 sg13g2_nor2_2 _30455_ (.A(_04712_),
    .B(_04732_),
    .Y(_04733_));
 sg13g2_nor2_1 _30456_ (.A(\u_inv.d_next[175] ),
    .B(\u_inv.d_reg[175] ),
    .Y(_04734_));
 sg13g2_nand2_1 _30457_ (.Y(_04735_),
    .A(\u_inv.d_next[175] ),
    .B(\u_inv.d_reg[175] ));
 sg13g2_nand2b_2 _30458_ (.Y(_04736_),
    .B(_04735_),
    .A_N(_04734_));
 sg13g2_nand2_1 _30459_ (.Y(_04737_),
    .A(\u_inv.d_next[174] ),
    .B(\u_inv.d_reg[174] ));
 sg13g2_xnor2_1 _30460_ (.Y(_04738_),
    .A(\u_inv.d_next[174] ),
    .B(\u_inv.d_reg[174] ));
 sg13g2_and2_1 _30461_ (.A(_04736_),
    .B(_04738_),
    .X(_04739_));
 sg13g2_xor2_1 _30462_ (.B(\u_inv.d_reg[173] ),
    .A(\u_inv.d_next[173] ),
    .X(_04740_));
 sg13g2_xnor2_1 _30463_ (.Y(_04741_),
    .A(\u_inv.d_next[173] ),
    .B(\u_inv.d_reg[173] ));
 sg13g2_nor2_1 _30464_ (.A(_14198_),
    .B(_14637_),
    .Y(_04742_));
 sg13g2_xnor2_1 _30465_ (.Y(_04743_),
    .A(\u_inv.d_next[172] ),
    .B(\u_inv.d_reg[172] ));
 sg13g2_inv_2 _30466_ (.Y(_04744_),
    .A(_04743_));
 sg13g2_nor2_1 _30467_ (.A(_04740_),
    .B(_04744_),
    .Y(_04745_));
 sg13g2_nand2_1 _30468_ (.Y(_04746_),
    .A(_04739_),
    .B(_04745_));
 sg13g2_nor2_1 _30469_ (.A(\u_inv.d_next[171] ),
    .B(\u_inv.d_reg[171] ),
    .Y(_04747_));
 sg13g2_nand2_1 _30470_ (.Y(_04748_),
    .A(\u_inv.d_next[171] ),
    .B(\u_inv.d_reg[171] ));
 sg13g2_nand2b_2 _30471_ (.Y(_04749_),
    .B(_04748_),
    .A_N(_04747_));
 sg13g2_nand2_1 _30472_ (.Y(_04750_),
    .A(\u_inv.d_next[170] ),
    .B(\u_inv.d_reg[170] ));
 sg13g2_xnor2_1 _30473_ (.Y(_04751_),
    .A(\u_inv.d_next[170] ),
    .B(\u_inv.d_reg[170] ));
 sg13g2_nand2_1 _30474_ (.Y(_04752_),
    .A(_04749_),
    .B(_04751_));
 sg13g2_xor2_1 _30475_ (.B(\u_inv.d_reg[169] ),
    .A(\u_inv.d_next[169] ),
    .X(_04753_));
 sg13g2_xor2_1 _30476_ (.B(\u_inv.d_reg[168] ),
    .A(\u_inv.d_next[168] ),
    .X(_04754_));
 sg13g2_or2_1 _30477_ (.X(_04755_),
    .B(_04754_),
    .A(_04753_));
 sg13g2_or2_1 _30478_ (.X(_04756_),
    .B(_04755_),
    .A(_04752_));
 sg13g2_nor2_1 _30479_ (.A(_04746_),
    .B(_04756_),
    .Y(_04757_));
 sg13g2_xor2_1 _30480_ (.B(\u_inv.d_reg[165] ),
    .A(\u_inv.d_next[165] ),
    .X(_04758_));
 sg13g2_xnor2_1 _30481_ (.Y(_04759_),
    .A(\u_inv.d_next[165] ),
    .B(\u_inv.d_reg[165] ));
 sg13g2_and2_1 _30482_ (.A(\u_inv.d_next[164] ),
    .B(net5867),
    .X(_04760_));
 sg13g2_xor2_1 _30483_ (.B(net5867),
    .A(\u_inv.d_next[164] ),
    .X(_04761_));
 sg13g2_xnor2_1 _30484_ (.Y(_04762_),
    .A(\u_inv.d_next[164] ),
    .B(net5867));
 sg13g2_nand2_1 _30485_ (.Y(_04763_),
    .A(_04759_),
    .B(_04762_));
 sg13g2_xor2_1 _30486_ (.B(\u_inv.d_reg[167] ),
    .A(\u_inv.d_next[167] ),
    .X(_04764_));
 sg13g2_xnor2_1 _30487_ (.Y(_04765_),
    .A(\u_inv.d_next[167] ),
    .B(\u_inv.d_reg[167] ));
 sg13g2_nand2_1 _30488_ (.Y(_04766_),
    .A(\u_inv.d_next[166] ),
    .B(\u_inv.d_reg[166] ));
 sg13g2_xor2_1 _30489_ (.B(\u_inv.d_reg[166] ),
    .A(\u_inv.d_next[166] ),
    .X(_04767_));
 sg13g2_xnor2_1 _30490_ (.Y(_04768_),
    .A(\u_inv.d_next[166] ),
    .B(\u_inv.d_reg[166] ));
 sg13g2_nor3_1 _30491_ (.A(_04763_),
    .B(_04764_),
    .C(_04767_),
    .Y(_04769_));
 sg13g2_nor2_1 _30492_ (.A(\u_inv.d_next[163] ),
    .B(\u_inv.d_reg[163] ),
    .Y(_04770_));
 sg13g2_nand2_1 _30493_ (.Y(_04771_),
    .A(\u_inv.d_next[163] ),
    .B(\u_inv.d_reg[163] ));
 sg13g2_xnor2_1 _30494_ (.Y(_04772_),
    .A(\u_inv.d_next[163] ),
    .B(\u_inv.d_reg[163] ));
 sg13g2_nand2_1 _30495_ (.Y(_04773_),
    .A(\u_inv.d_next[162] ),
    .B(\u_inv.d_reg[162] ));
 sg13g2_xor2_1 _30496_ (.B(\u_inv.d_reg[162] ),
    .A(\u_inv.d_next[162] ),
    .X(_04774_));
 sg13g2_xnor2_1 _30497_ (.Y(_04775_),
    .A(\u_inv.d_next[162] ),
    .B(\u_inv.d_reg[162] ));
 sg13g2_nand2_1 _30498_ (.Y(_04776_),
    .A(_04772_),
    .B(_04775_));
 sg13g2_nor2b_1 _30499_ (.A(\u_inv.d_reg[161] ),
    .B_N(\u_inv.d_next[161] ),
    .Y(_04777_));
 sg13g2_nand2b_1 _30500_ (.Y(_04778_),
    .B(\u_inv.d_reg[161] ),
    .A_N(\u_inv.d_next[161] ));
 sg13g2_xnor2_1 _30501_ (.Y(_04779_),
    .A(\u_inv.d_next[161] ),
    .B(\u_inv.d_reg[161] ));
 sg13g2_nand2b_2 _30502_ (.Y(_04780_),
    .B(_04778_),
    .A_N(_04777_));
 sg13g2_nand2_1 _30503_ (.Y(_04781_),
    .A(\u_inv.d_next[160] ),
    .B(net5868));
 sg13g2_xor2_1 _30504_ (.B(net5868),
    .A(\u_inv.d_next[160] ),
    .X(_04782_));
 sg13g2_xnor2_1 _30505_ (.Y(_04783_),
    .A(\u_inv.d_next[160] ),
    .B(net5868));
 sg13g2_nor2_1 _30506_ (.A(_04780_),
    .B(_04782_),
    .Y(_04784_));
 sg13g2_nor3_1 _30507_ (.A(_04776_),
    .B(_04780_),
    .C(_04782_),
    .Y(_04785_));
 sg13g2_and2_1 _30508_ (.A(_04769_),
    .B(_04785_),
    .X(_04786_));
 sg13g2_and2_1 _30509_ (.A(_04757_),
    .B(_04786_),
    .X(_04787_));
 sg13g2_and2_1 _30510_ (.A(_04733_),
    .B(_04787_),
    .X(_04788_));
 sg13g2_nand2_2 _30511_ (.Y(_04789_),
    .A(_04733_),
    .B(_04787_));
 sg13g2_xor2_1 _30512_ (.B(\u_inv.d_reg[159] ),
    .A(\u_inv.d_next[159] ),
    .X(_04790_));
 sg13g2_xnor2_1 _30513_ (.Y(_04791_),
    .A(\u_inv.d_next[159] ),
    .B(\u_inv.d_reg[159] ));
 sg13g2_nand2_1 _30514_ (.Y(_04792_),
    .A(\u_inv.d_next[158] ),
    .B(\u_inv.d_reg[158] ));
 sg13g2_xor2_1 _30515_ (.B(\u_inv.d_reg[158] ),
    .A(\u_inv.d_next[158] ),
    .X(_04793_));
 sg13g2_xnor2_1 _30516_ (.Y(_04794_),
    .A(\u_inv.d_next[158] ),
    .B(\u_inv.d_reg[158] ));
 sg13g2_nand2_1 _30517_ (.Y(_04795_),
    .A(_04791_),
    .B(_04794_));
 sg13g2_xor2_1 _30518_ (.B(\u_inv.d_reg[157] ),
    .A(\u_inv.d_next[157] ),
    .X(_04796_));
 sg13g2_xor2_1 _30519_ (.B(\u_inv.d_reg[156] ),
    .A(\u_inv.d_next[156] ),
    .X(_04797_));
 sg13g2_or2_1 _30520_ (.X(_04798_),
    .B(_04797_),
    .A(_04796_));
 sg13g2_inv_1 _30521_ (.Y(_04799_),
    .A(_04798_));
 sg13g2_nor2_1 _30522_ (.A(_04795_),
    .B(_04798_),
    .Y(_04800_));
 sg13g2_xnor2_1 _30523_ (.Y(_04801_),
    .A(\u_inv.d_next[155] ),
    .B(\u_inv.d_reg[155] ));
 sg13g2_and2_1 _30524_ (.A(\u_inv.d_next[154] ),
    .B(\u_inv.d_reg[154] ),
    .X(_04802_));
 sg13g2_xnor2_1 _30525_ (.Y(_04803_),
    .A(\u_inv.d_next[154] ),
    .B(\u_inv.d_reg[154] ));
 sg13g2_inv_1 _30526_ (.Y(_04804_),
    .A(_04803_));
 sg13g2_nand2_1 _30527_ (.Y(_04805_),
    .A(_04801_),
    .B(_04803_));
 sg13g2_xor2_1 _30528_ (.B(\u_inv.d_reg[153] ),
    .A(\u_inv.d_next[153] ),
    .X(_04806_));
 sg13g2_xor2_1 _30529_ (.B(\u_inv.d_reg[152] ),
    .A(\u_inv.d_next[152] ),
    .X(_04807_));
 sg13g2_or2_1 _30530_ (.X(_04808_),
    .B(_04807_),
    .A(_04806_));
 sg13g2_or4_1 _30531_ (.A(_04795_),
    .B(_04798_),
    .C(_04805_),
    .D(_04808_),
    .X(_04809_));
 sg13g2_nor2_1 _30532_ (.A(\u_inv.d_next[151] ),
    .B(\u_inv.d_reg[151] ),
    .Y(_04810_));
 sg13g2_xor2_1 _30533_ (.B(\u_inv.d_reg[151] ),
    .A(\u_inv.d_next[151] ),
    .X(_04811_));
 sg13g2_xnor2_1 _30534_ (.Y(_04812_),
    .A(\u_inv.d_next[151] ),
    .B(\u_inv.d_reg[151] ));
 sg13g2_nand2_1 _30535_ (.Y(_04813_),
    .A(\u_inv.d_next[150] ),
    .B(\u_inv.d_reg[150] ));
 sg13g2_xor2_1 _30536_ (.B(\u_inv.d_reg[150] ),
    .A(\u_inv.d_next[150] ),
    .X(_04814_));
 sg13g2_xnor2_1 _30537_ (.Y(_04815_),
    .A(\u_inv.d_next[150] ),
    .B(\u_inv.d_reg[150] ));
 sg13g2_nor2_1 _30538_ (.A(_04811_),
    .B(_04814_),
    .Y(_04816_));
 sg13g2_xor2_1 _30539_ (.B(\u_inv.d_reg[149] ),
    .A(\u_inv.d_next[149] ),
    .X(_04817_));
 sg13g2_xnor2_1 _30540_ (.Y(_04818_),
    .A(\u_inv.d_next[149] ),
    .B(\u_inv.d_reg[149] ));
 sg13g2_and2_1 _30541_ (.A(\u_inv.d_next[148] ),
    .B(\u_inv.d_reg[148] ),
    .X(_04819_));
 sg13g2_xor2_1 _30542_ (.B(\u_inv.d_reg[148] ),
    .A(\u_inv.d_next[148] ),
    .X(_04820_));
 sg13g2_nor2_1 _30543_ (.A(_04817_),
    .B(_04820_),
    .Y(_04821_));
 sg13g2_inv_1 _30544_ (.Y(_04822_),
    .A(_04821_));
 sg13g2_nand2_1 _30545_ (.Y(_04823_),
    .A(_04816_),
    .B(_04821_));
 sg13g2_xor2_1 _30546_ (.B(\u_inv.d_reg[147] ),
    .A(\u_inv.d_next[147] ),
    .X(_04824_));
 sg13g2_xnor2_1 _30547_ (.Y(_04825_),
    .A(\u_inv.d_next[147] ),
    .B(\u_inv.d_reg[147] ));
 sg13g2_xor2_1 _30548_ (.B(\u_inv.d_reg[146] ),
    .A(\u_inv.d_next[146] ),
    .X(_04826_));
 sg13g2_nor2_1 _30549_ (.A(_04824_),
    .B(_04826_),
    .Y(_04827_));
 sg13g2_xnor2_1 _30550_ (.Y(_04828_),
    .A(net5876),
    .B(\u_inv.d_reg[145] ));
 sg13g2_xor2_1 _30551_ (.B(\u_inv.d_reg[145] ),
    .A(net5876),
    .X(_04829_));
 sg13g2_nand2_1 _30552_ (.Y(_04830_),
    .A(\u_inv.d_next[144] ),
    .B(\u_inv.d_reg[144] ));
 sg13g2_xor2_1 _30553_ (.B(\u_inv.d_reg[144] ),
    .A(\u_inv.d_next[144] ),
    .X(_04831_));
 sg13g2_nor2_1 _30554_ (.A(_04829_),
    .B(_04831_),
    .Y(_04832_));
 sg13g2_and4_1 _30555_ (.A(_04816_),
    .B(_04821_),
    .C(_04827_),
    .D(_04832_),
    .X(_04833_));
 sg13g2_nor2b_2 _30556_ (.A(_04809_),
    .B_N(_04833_),
    .Y(_04834_));
 sg13g2_nor2b_1 _30557_ (.A(\u_inv.d_reg[136] ),
    .B_N(\u_inv.d_next[136] ),
    .Y(_04835_));
 sg13g2_o21ai_1 _30558_ (.B1(_04835_),
    .Y(_04836_),
    .A1(\u_inv.d_next[137] ),
    .A2(_14672_));
 sg13g2_o21ai_1 _30559_ (.B1(_04836_),
    .Y(_04837_),
    .A1(_14209_),
    .A2(\u_inv.d_reg[137] ));
 sg13g2_inv_1 _30560_ (.Y(_04838_),
    .A(_04837_));
 sg13g2_xnor2_1 _30561_ (.Y(_04839_),
    .A(\u_inv.d_next[141] ),
    .B(\u_inv.d_reg[141] ));
 sg13g2_nand2_1 _30562_ (.Y(_04840_),
    .A(\u_inv.d_next[140] ),
    .B(net5869));
 sg13g2_xnor2_1 _30563_ (.Y(_04841_),
    .A(\u_inv.d_next[140] ),
    .B(net5869));
 sg13g2_and2_1 _30564_ (.A(_04839_),
    .B(_04841_),
    .X(_04842_));
 sg13g2_nor2_1 _30565_ (.A(\u_inv.d_next[143] ),
    .B(\u_inv.d_reg[143] ),
    .Y(_04843_));
 sg13g2_nand2_1 _30566_ (.Y(_04844_),
    .A(\u_inv.d_next[143] ),
    .B(\u_inv.d_reg[143] ));
 sg13g2_nor2b_1 _30567_ (.A(_04843_),
    .B_N(_04844_),
    .Y(_04845_));
 sg13g2_nand2b_2 _30568_ (.Y(_04846_),
    .B(_04844_),
    .A_N(_04843_));
 sg13g2_nand2_1 _30569_ (.Y(_04847_),
    .A(\u_inv.d_next[142] ),
    .B(\u_inv.d_reg[142] ));
 sg13g2_xor2_1 _30570_ (.B(\u_inv.d_reg[142] ),
    .A(\u_inv.d_next[142] ),
    .X(_04848_));
 sg13g2_nand3b_1 _30571_ (.B(_04842_),
    .C(_04846_),
    .Y(_04849_),
    .A_N(_04848_));
 sg13g2_xor2_1 _30572_ (.B(\u_inv.d_reg[139] ),
    .A(\u_inv.d_next[139] ),
    .X(_04850_));
 sg13g2_and2_1 _30573_ (.A(\u_inv.d_next[138] ),
    .B(\u_inv.d_reg[138] ),
    .X(_04851_));
 sg13g2_xor2_1 _30574_ (.B(\u_inv.d_reg[138] ),
    .A(\u_inv.d_next[138] ),
    .X(_04852_));
 sg13g2_or2_1 _30575_ (.X(_04853_),
    .B(_04852_),
    .A(_04850_));
 sg13g2_nor2_1 _30576_ (.A(_14207_),
    .B(\u_inv.d_reg[141] ),
    .Y(_04854_));
 sg13g2_nor2b_1 _30577_ (.A(net5869),
    .B_N(\u_inv.d_next[140] ),
    .Y(_04855_));
 sg13g2_nand2_1 _30578_ (.Y(_04856_),
    .A(\u_inv.d_next[140] ),
    .B(_14669_));
 sg13g2_a21oi_1 _30579_ (.A1(_04839_),
    .A2(_04855_),
    .Y(_04857_),
    .B1(_04854_));
 sg13g2_nand2_1 _30580_ (.Y(_04858_),
    .A(\u_inv.d_next[138] ),
    .B(_14671_));
 sg13g2_nor2_1 _30581_ (.A(_04850_),
    .B(_04858_),
    .Y(_04859_));
 sg13g2_a21oi_1 _30582_ (.A1(\u_inv.d_next[139] ),
    .A2(_14670_),
    .Y(_04860_),
    .B1(_04859_));
 sg13g2_a21o_1 _30583_ (.A2(_14670_),
    .A1(\u_inv.d_next[139] ),
    .B1(_04859_),
    .X(_04861_));
 sg13g2_nor2b_1 _30584_ (.A(\u_inv.d_reg[142] ),
    .B_N(\u_inv.d_next[142] ),
    .Y(_04862_));
 sg13g2_nor2_1 _30585_ (.A(_04848_),
    .B(_04857_),
    .Y(_04863_));
 sg13g2_or2_1 _30586_ (.X(_04864_),
    .B(_04863_),
    .A(_04862_));
 sg13g2_o21ai_1 _30587_ (.B1(_04860_),
    .Y(_04865_),
    .A1(_04838_),
    .A2(_04853_));
 sg13g2_nand2b_1 _30588_ (.Y(_04866_),
    .B(_04865_),
    .A_N(_04849_));
 sg13g2_o21ai_1 _30589_ (.B1(_04866_),
    .Y(_04867_),
    .A1(_14206_),
    .A2(\u_inv.d_reg[143] ));
 sg13g2_a21oi_1 _30590_ (.A1(_04846_),
    .A2(_04864_),
    .Y(_04868_),
    .B1(_04867_));
 sg13g2_xor2_1 _30591_ (.B(\u_inv.d_reg[135] ),
    .A(\u_inv.d_next[135] ),
    .X(_04869_));
 sg13g2_xnor2_1 _30592_ (.Y(_04870_),
    .A(\u_inv.d_next[135] ),
    .B(\u_inv.d_reg[135] ));
 sg13g2_nand2_1 _30593_ (.Y(_04871_),
    .A(\u_inv.d_next[134] ),
    .B(\u_inv.d_reg[134] ));
 sg13g2_xor2_1 _30594_ (.B(\u_inv.d_reg[134] ),
    .A(\u_inv.d_next[134] ),
    .X(_04872_));
 sg13g2_xnor2_1 _30595_ (.Y(_04873_),
    .A(\u_inv.d_next[134] ),
    .B(\u_inv.d_reg[134] ));
 sg13g2_nand2_1 _30596_ (.Y(_04874_),
    .A(_04870_),
    .B(_04873_));
 sg13g2_xnor2_1 _30597_ (.Y(_04875_),
    .A(\u_inv.d_next[133] ),
    .B(\u_inv.d_reg[133] ));
 sg13g2_xor2_1 _30598_ (.B(\u_inv.d_reg[133] ),
    .A(\u_inv.d_next[133] ),
    .X(_04876_));
 sg13g2_nand2_1 _30599_ (.Y(_04877_),
    .A(\u_inv.d_next[132] ),
    .B(\u_inv.d_reg[132] ));
 sg13g2_xor2_1 _30600_ (.B(\u_inv.d_reg[132] ),
    .A(\u_inv.d_next[132] ),
    .X(_04878_));
 sg13g2_inv_1 _30601_ (.Y(_04879_),
    .A(_04878_));
 sg13g2_nor2_1 _30602_ (.A(_04876_),
    .B(_04878_),
    .Y(_04880_));
 sg13g2_nand2b_1 _30603_ (.Y(_04881_),
    .B(_04880_),
    .A_N(_04874_));
 sg13g2_xnor2_1 _30604_ (.Y(_04882_),
    .A(\u_inv.d_next[131] ),
    .B(\u_inv.d_reg[131] ));
 sg13g2_nand2_1 _30605_ (.Y(_04883_),
    .A(\u_inv.d_next[130] ),
    .B(\u_inv.d_reg[130] ));
 sg13g2_xnor2_1 _30606_ (.Y(_04884_),
    .A(\u_inv.d_next[130] ),
    .B(\u_inv.d_reg[130] ));
 sg13g2_and2_1 _30607_ (.A(net5619),
    .B(_04884_),
    .X(_04885_));
 sg13g2_nand2_1 _30608_ (.Y(_04886_),
    .A(net5619),
    .B(_04884_));
 sg13g2_nor2b_1 _30609_ (.A(\u_inv.d_next[129] ),
    .B_N(\u_inv.d_reg[129] ),
    .Y(_04887_));
 sg13g2_nand2b_1 _30610_ (.Y(_04888_),
    .B(\u_inv.d_next[129] ),
    .A_N(\u_inv.d_reg[129] ));
 sg13g2_nand2_1 _30611_ (.Y(_04889_),
    .A(\u_inv.d_next[128] ),
    .B(_14681_));
 sg13g2_nand2_1 _30612_ (.Y(_04890_),
    .A(_04888_),
    .B(_04889_));
 sg13g2_o21ai_1 _30613_ (.B1(_04888_),
    .Y(_04891_),
    .A1(_04887_),
    .A2(_04889_));
 sg13g2_nand2b_1 _30614_ (.Y(_04892_),
    .B(_04890_),
    .A_N(_04887_));
 sg13g2_nor2b_1 _30615_ (.A(\u_inv.d_reg[130] ),
    .B_N(\u_inv.d_next[130] ),
    .Y(_04893_));
 sg13g2_o21ai_1 _30616_ (.B1(_04893_),
    .Y(_04894_),
    .A1(\u_inv.d_next[131] ),
    .A2(_14678_));
 sg13g2_o21ai_1 _30617_ (.B1(_04894_),
    .Y(_04895_),
    .A1(_14212_),
    .A2(\u_inv.d_reg[131] ));
 sg13g2_a21oi_1 _30618_ (.A1(_04885_),
    .A2(_04891_),
    .Y(_04896_),
    .B1(_04895_));
 sg13g2_nand2b_1 _30619_ (.Y(_04897_),
    .B(\u_inv.d_next[132] ),
    .A_N(\u_inv.d_reg[132] ));
 sg13g2_o21ai_1 _30620_ (.B1(_04897_),
    .Y(_04898_),
    .A1(_14211_),
    .A2(\u_inv.d_reg[133] ));
 sg13g2_o21ai_1 _30621_ (.B1(_04898_),
    .Y(_04899_),
    .A1(\u_inv.d_next[133] ),
    .A2(_14676_));
 sg13g2_nor2_1 _30622_ (.A(_04874_),
    .B(_04899_),
    .Y(_04900_));
 sg13g2_nor2b_2 _30623_ (.A(\u_inv.d_reg[134] ),
    .B_N(\u_inv.d_next[134] ),
    .Y(_04901_));
 sg13g2_a21oi_1 _30624_ (.A1(\u_inv.d_next[135] ),
    .A2(_14674_),
    .Y(_04902_),
    .B1(_04900_));
 sg13g2_o21ai_1 _30625_ (.B1(_04902_),
    .Y(_04903_),
    .A1(_04881_),
    .A2(_04896_));
 sg13g2_a21oi_2 _30626_ (.B1(_04903_),
    .Y(_04904_),
    .A2(_04901_),
    .A1(_04870_));
 sg13g2_inv_1 _30627_ (.Y(_04905_),
    .A(_04904_));
 sg13g2_xnor2_1 _30628_ (.Y(_04906_),
    .A(\u_inv.d_next[137] ),
    .B(\u_inv.d_reg[137] ));
 sg13g2_xor2_1 _30629_ (.B(\u_inv.d_reg[137] ),
    .A(\u_inv.d_next[137] ),
    .X(_04907_));
 sg13g2_nand2_1 _30630_ (.Y(_04908_),
    .A(\u_inv.d_next[136] ),
    .B(\u_inv.d_reg[136] ));
 sg13g2_xor2_1 _30631_ (.B(\u_inv.d_reg[136] ),
    .A(\u_inv.d_next[136] ),
    .X(_04909_));
 sg13g2_inv_1 _30632_ (.Y(_04910_),
    .A(_04909_));
 sg13g2_nor2_1 _30633_ (.A(_04907_),
    .B(_04909_),
    .Y(_04911_));
 sg13g2_nor4_1 _30634_ (.A(_04849_),
    .B(_04853_),
    .C(_04907_),
    .D(_04909_),
    .Y(_04912_));
 sg13g2_nand2_1 _30635_ (.Y(_04913_),
    .A(\u_inv.d_next[152] ),
    .B(_14657_));
 sg13g2_nor2_1 _30636_ (.A(_04806_),
    .B(_04913_),
    .Y(_04914_));
 sg13g2_a21oi_1 _30637_ (.A1(\u_inv.d_next[153] ),
    .A2(_14656_),
    .Y(_04915_),
    .B1(_04914_));
 sg13g2_nor2b_1 _30638_ (.A(\u_inv.d_reg[154] ),
    .B_N(\u_inv.d_next[154] ),
    .Y(_04916_));
 sg13g2_nor2_1 _30639_ (.A(_14201_),
    .B(\u_inv.d_reg[155] ),
    .Y(_04917_));
 sg13g2_a21oi_1 _30640_ (.A1(_04801_),
    .A2(_04916_),
    .Y(_04918_),
    .B1(_04917_));
 sg13g2_o21ai_1 _30641_ (.B1(_04918_),
    .Y(_04919_),
    .A1(_04805_),
    .A2(_04915_));
 sg13g2_nand2_1 _30642_ (.Y(_04920_),
    .A(\u_inv.d_next[156] ),
    .B(_14653_));
 sg13g2_nor2_1 _30643_ (.A(_04796_),
    .B(_04920_),
    .Y(_04921_));
 sg13g2_a21oi_1 _30644_ (.A1(\u_inv.d_next[157] ),
    .A2(_14652_),
    .Y(_04922_),
    .B1(_04921_));
 sg13g2_nor2_1 _30645_ (.A(_04795_),
    .B(_04922_),
    .Y(_04923_));
 sg13g2_nor2b_1 _30646_ (.A(\u_inv.d_reg[158] ),
    .B_N(\u_inv.d_next[158] ),
    .Y(_04924_));
 sg13g2_nor2b_1 _30647_ (.A(\u_inv.d_reg[144] ),
    .B_N(\u_inv.d_next[144] ),
    .Y(_04925_));
 sg13g2_a21oi_1 _30648_ (.A1(net5876),
    .A2(_14664_),
    .Y(_04926_),
    .B1(_04925_));
 sg13g2_a21oi_1 _30649_ (.A1(_14205_),
    .A2(\u_inv.d_reg[145] ),
    .Y(_04927_),
    .B1(_04926_));
 sg13g2_nand2_1 _30650_ (.Y(_04928_),
    .A(\u_inv.d_next[146] ),
    .B(_14663_));
 sg13g2_nor2_1 _30651_ (.A(_04824_),
    .B(_04928_),
    .Y(_04929_));
 sg13g2_a221oi_1 _30652_ (.B2(_04927_),
    .C1(_04929_),
    .B1(_04827_),
    .A1(\u_inv.d_next[147] ),
    .Y(_04930_),
    .A2(_14662_));
 sg13g2_nor2b_1 _30653_ (.A(\u_inv.d_reg[148] ),
    .B_N(\u_inv.d_next[148] ),
    .Y(_04931_));
 sg13g2_nand2_1 _30654_ (.Y(_04932_),
    .A(_04818_),
    .B(_04931_));
 sg13g2_o21ai_1 _30655_ (.B1(_04932_),
    .Y(_04933_),
    .A1(_14203_),
    .A2(\u_inv.d_reg[149] ));
 sg13g2_nand2_1 _30656_ (.Y(_04934_),
    .A(\u_inv.d_next[150] ),
    .B(_14659_));
 sg13g2_nor2_1 _30657_ (.A(_04811_),
    .B(_04934_),
    .Y(_04935_));
 sg13g2_a221oi_1 _30658_ (.B2(_04933_),
    .C1(_04935_),
    .B1(_04816_),
    .A1(\u_inv.d_next[151] ),
    .Y(_04936_),
    .A2(_14658_));
 sg13g2_o21ai_1 _30659_ (.B1(_04936_),
    .Y(_04937_),
    .A1(_04823_),
    .A2(_04930_));
 sg13g2_inv_1 _30660_ (.Y(_04938_),
    .A(_04937_));
 sg13g2_nand2b_1 _30661_ (.Y(_04939_),
    .B(_04912_),
    .A_N(_04904_));
 sg13g2_nand2_2 _30662_ (.Y(_04940_),
    .A(_04868_),
    .B(_04939_));
 sg13g2_a221oi_1 _30663_ (.B2(_04919_),
    .C1(_04923_),
    .B1(_04800_),
    .A1(\u_inv.d_next[159] ),
    .Y(_04941_),
    .A2(_14650_));
 sg13g2_o21ai_1 _30664_ (.B1(_04941_),
    .Y(_04942_),
    .A1(_04809_),
    .A2(_04938_));
 sg13g2_a221oi_1 _30665_ (.B2(_04834_),
    .C1(_04942_),
    .B1(_04940_),
    .A1(_04791_),
    .Y(_04943_),
    .A2(_04924_));
 sg13g2_inv_4 _30666_ (.A(_04943_),
    .Y(_04944_));
 sg13g2_nor2b_1 _30667_ (.A(net5868),
    .B_N(\u_inv.d_next[160] ),
    .Y(_04945_));
 sg13g2_a21oi_1 _30668_ (.A1(_04778_),
    .A2(_04945_),
    .Y(_04946_),
    .B1(_04777_));
 sg13g2_nor2b_1 _30669_ (.A(\u_inv.d_reg[162] ),
    .B_N(\u_inv.d_next[162] ),
    .Y(_04947_));
 sg13g2_nand2_1 _30670_ (.Y(_04948_),
    .A(\u_inv.d_next[162] ),
    .B(_14647_));
 sg13g2_nor2b_1 _30671_ (.A(\u_inv.d_reg[163] ),
    .B_N(\u_inv.d_next[163] ),
    .Y(_04949_));
 sg13g2_a21oi_1 _30672_ (.A1(_04772_),
    .A2(_04947_),
    .Y(_04950_),
    .B1(_04949_));
 sg13g2_o21ai_1 _30673_ (.B1(_04950_),
    .Y(_04951_),
    .A1(_04776_),
    .A2(_04946_));
 sg13g2_inv_1 _30674_ (.Y(_04952_),
    .A(_04951_));
 sg13g2_nand2_1 _30675_ (.Y(_04953_),
    .A(_04769_),
    .B(_04951_));
 sg13g2_nor2b_1 _30676_ (.A(\u_inv.d_reg[165] ),
    .B_N(\u_inv.d_next[165] ),
    .Y(_04954_));
 sg13g2_nor2b_1 _30677_ (.A(net5867),
    .B_N(\u_inv.d_next[164] ),
    .Y(_04955_));
 sg13g2_a21oi_1 _30678_ (.A1(_04759_),
    .A2(_04955_),
    .Y(_04956_),
    .B1(_04954_));
 sg13g2_or3_1 _30679_ (.A(_04764_),
    .B(_04767_),
    .C(_04956_),
    .X(_04957_));
 sg13g2_nor2_1 _30680_ (.A(_14199_),
    .B(\u_inv.d_reg[167] ),
    .Y(_04958_));
 sg13g2_nor2b_1 _30681_ (.A(\u_inv.d_reg[166] ),
    .B_N(\u_inv.d_next[166] ),
    .Y(_04959_));
 sg13g2_a21oi_1 _30682_ (.A1(_04765_),
    .A2(_04959_),
    .Y(_04960_),
    .B1(_04958_));
 sg13g2_nand3_1 _30683_ (.B(_04957_),
    .C(_04960_),
    .A(_04953_),
    .Y(_04961_));
 sg13g2_nor2_1 _30684_ (.A(_14198_),
    .B(\u_inv.d_reg[172] ),
    .Y(_04962_));
 sg13g2_nor3_1 _30685_ (.A(_14198_),
    .B(\u_inv.d_reg[172] ),
    .C(_04740_),
    .Y(_04963_));
 sg13g2_a21o_1 _30686_ (.A2(_14636_),
    .A1(\u_inv.d_next[173] ),
    .B1(_04963_),
    .X(_04964_));
 sg13g2_nor2b_1 _30687_ (.A(\u_inv.d_reg[174] ),
    .B_N(\u_inv.d_next[174] ),
    .Y(_04965_));
 sg13g2_nand2_1 _30688_ (.Y(_04966_),
    .A(\u_inv.d_next[168] ),
    .B(_14641_));
 sg13g2_nor2_1 _30689_ (.A(_04753_),
    .B(_04966_),
    .Y(_04967_));
 sg13g2_a21oi_1 _30690_ (.A1(\u_inv.d_next[169] ),
    .A2(_14640_),
    .Y(_04968_),
    .B1(_04967_));
 sg13g2_nor2b_1 _30691_ (.A(\u_inv.d_reg[170] ),
    .B_N(\u_inv.d_next[170] ),
    .Y(_04969_));
 sg13g2_nand2_1 _30692_ (.Y(_04970_),
    .A(\u_inv.d_next[171] ),
    .B(_14638_));
 sg13g2_o21ai_1 _30693_ (.B1(_04970_),
    .Y(_04971_),
    .A1(_04752_),
    .A2(_04968_));
 sg13g2_a21oi_1 _30694_ (.A1(_04749_),
    .A2(_04969_),
    .Y(_04972_),
    .B1(_04971_));
 sg13g2_a22oi_1 _30695_ (.Y(_04973_),
    .B1(_04965_),
    .B2(_04736_),
    .A2(_04964_),
    .A1(_04739_));
 sg13g2_o21ai_1 _30696_ (.B1(_04973_),
    .Y(_04974_),
    .A1(_04746_),
    .A2(_04972_));
 sg13g2_a21oi_1 _30697_ (.A1(_04757_),
    .A2(_04961_),
    .Y(_04975_),
    .B1(_04974_));
 sg13g2_o21ai_1 _30698_ (.B1(_04975_),
    .Y(_04976_),
    .A1(_14197_),
    .A2(\u_inv.d_reg[175] ));
 sg13g2_nand2_1 _30699_ (.Y(_04977_),
    .A(\u_inv.d_next[177] ),
    .B(_14632_));
 sg13g2_nand2_1 _30700_ (.Y(_04978_),
    .A(\u_inv.d_next[176] ),
    .B(_14633_));
 sg13g2_o21ai_1 _30701_ (.B1(_04977_),
    .Y(_04979_),
    .A1(_04727_),
    .A2(_04978_));
 sg13g2_inv_1 _30702_ (.Y(_04980_),
    .A(_04979_));
 sg13g2_nor2_1 _30703_ (.A(_14195_),
    .B(\u_inv.d_reg[179] ),
    .Y(_04981_));
 sg13g2_nor2b_1 _30704_ (.A(\u_inv.d_reg[178] ),
    .B_N(\u_inv.d_next[178] ),
    .Y(_04982_));
 sg13g2_a221oi_1 _30705_ (.B2(_04723_),
    .C1(_04981_),
    .B1(_04982_),
    .A1(_04726_),
    .Y(_04983_),
    .A2(_04979_));
 sg13g2_nor2b_1 _30706_ (.A(_04983_),
    .B_N(_04722_),
    .Y(_04984_));
 sg13g2_nor2_1 _30707_ (.A(_14194_),
    .B(\u_inv.d_reg[181] ),
    .Y(_04985_));
 sg13g2_nor2b_1 _30708_ (.A(\u_inv.d_reg[180] ),
    .B_N(\u_inv.d_next[180] ),
    .Y(_04986_));
 sg13g2_nand2_1 _30709_ (.Y(_04987_),
    .A(\u_inv.d_next[180] ),
    .B(_14629_));
 sg13g2_a21oi_1 _30710_ (.A1(_04713_),
    .A2(_04986_),
    .Y(_04988_),
    .B1(_04985_));
 sg13g2_nor2_1 _30711_ (.A(_14193_),
    .B(\u_inv.d_reg[183] ),
    .Y(_04989_));
 sg13g2_nand2_1 _30712_ (.Y(_04990_),
    .A(\u_inv.d_next[182] ),
    .B(_14627_));
 sg13g2_o21ai_1 _30713_ (.B1(_04990_),
    .Y(_04991_),
    .A1(_04721_),
    .A2(_04988_));
 sg13g2_a21oi_1 _30714_ (.A1(_04719_),
    .A2(_04991_),
    .Y(_04992_),
    .B1(_04989_));
 sg13g2_nor2b_1 _30715_ (.A(_04984_),
    .B_N(_04992_),
    .Y(_04993_));
 sg13g2_nor2b_1 _30716_ (.A(\u_inv.d_reg[185] ),
    .B_N(\u_inv.d_next[185] ),
    .Y(_04994_));
 sg13g2_nor2b_1 _30717_ (.A(net5866),
    .B_N(\u_inv.d_next[184] ),
    .Y(_04995_));
 sg13g2_a21o_1 _30718_ (.A2(_04995_),
    .A1(_04706_),
    .B1(_04994_),
    .X(_04996_));
 sg13g2_nand2_1 _30719_ (.Y(_04997_),
    .A(\u_inv.d_next[186] ),
    .B(_14623_));
 sg13g2_a22oi_1 _30720_ (.Y(_04998_),
    .B1(_04702_),
    .B2(_04996_),
    .A2(_14622_),
    .A1(\u_inv.d_next[187] ));
 sg13g2_o21ai_1 _30721_ (.B1(_04998_),
    .Y(_04999_),
    .A1(_04698_),
    .A2(_04997_));
 sg13g2_nor2_1 _30722_ (.A(_14192_),
    .B(\u_inv.d_reg[189] ),
    .Y(_05000_));
 sg13g2_nor2b_1 _30723_ (.A(\u_inv.d_reg[188] ),
    .B_N(\u_inv.d_next[188] ),
    .Y(_05001_));
 sg13g2_a21oi_1 _30724_ (.A1(_04691_),
    .A2(_05001_),
    .Y(_05002_),
    .B1(_05000_));
 sg13g2_nor2_1 _30725_ (.A(_14191_),
    .B(\u_inv.d_reg[190] ),
    .Y(_05003_));
 sg13g2_nor2b_1 _30726_ (.A(\u_inv.d_reg[191] ),
    .B_N(\u_inv.d_next[191] ),
    .Y(_05004_));
 sg13g2_a21oi_1 _30727_ (.A1(_04687_),
    .A2(_05003_),
    .Y(_05005_),
    .B1(_05004_));
 sg13g2_o21ai_1 _30728_ (.B1(_05005_),
    .Y(_05006_),
    .A1(_04690_),
    .A2(_05002_));
 sg13g2_a21oi_1 _30729_ (.A1(_04696_),
    .A2(_04999_),
    .Y(_05007_),
    .B1(_05006_));
 sg13g2_o21ai_1 _30730_ (.B1(_05007_),
    .Y(_05008_),
    .A1(_04712_),
    .A2(_04993_));
 sg13g2_a221oi_1 _30731_ (.B2(_04733_),
    .C1(_05008_),
    .B1(_04976_),
    .A1(_04788_),
    .Y(_05009_),
    .A2(_04944_));
 sg13g2_nand2_1 _30732_ (.Y(_05010_),
    .A(\u_inv.d_next[25] ),
    .B(_14784_));
 sg13g2_or2_1 _30733_ (.X(_05011_),
    .B(\u_inv.d_reg[25] ),
    .A(\u_inv.d_next[25] ));
 sg13g2_nand2_1 _30734_ (.Y(_05012_),
    .A(\u_inv.d_next[25] ),
    .B(\u_inv.d_reg[25] ));
 sg13g2_and2_1 _30735_ (.A(_05011_),
    .B(_05012_),
    .X(_05013_));
 sg13g2_nand2_1 _30736_ (.Y(_05014_),
    .A(\u_inv.d_next[24] ),
    .B(_14785_));
 sg13g2_o21ai_1 _30737_ (.B1(_05010_),
    .Y(_05015_),
    .A1(_05013_),
    .A2(_05014_));
 sg13g2_nor2b_1 _30738_ (.A(\u_inv.d_reg[31] ),
    .B_N(\u_inv.d_next[31] ),
    .Y(_05016_));
 sg13g2_nand2b_1 _30739_ (.Y(_05017_),
    .B(\u_inv.d_reg[31] ),
    .A_N(\u_inv.d_next[31] ));
 sg13g2_nor2b_2 _30740_ (.A(_05016_),
    .B_N(_05017_),
    .Y(_05018_));
 sg13g2_nand2_1 _30741_ (.Y(_05019_),
    .A(\u_inv.d_next[30] ),
    .B(\u_inv.d_reg[30] ));
 sg13g2_xnor2_1 _30742_ (.Y(_05020_),
    .A(\u_inv.d_next[30] ),
    .B(\u_inv.d_reg[30] ));
 sg13g2_nor2_1 _30743_ (.A(\u_inv.d_next[29] ),
    .B(\u_inv.d_reg[29] ),
    .Y(_05021_));
 sg13g2_nand2_1 _30744_ (.Y(_05022_),
    .A(\u_inv.d_next[29] ),
    .B(\u_inv.d_reg[29] ));
 sg13g2_nand2b_2 _30745_ (.Y(_05023_),
    .B(_05022_),
    .A_N(_05021_));
 sg13g2_nand2_1 _30746_ (.Y(_05024_),
    .A(\u_inv.d_next[28] ),
    .B(\u_inv.d_reg[28] ));
 sg13g2_xnor2_1 _30747_ (.Y(_05025_),
    .A(\u_inv.d_next[28] ),
    .B(\u_inv.d_reg[28] ));
 sg13g2_and2_1 _30748_ (.A(_05023_),
    .B(_05025_),
    .X(_05026_));
 sg13g2_nand3_1 _30749_ (.B(_05020_),
    .C(_05026_),
    .A(_05018_),
    .Y(_05027_));
 sg13g2_nand2_1 _30750_ (.Y(_05028_),
    .A(\u_inv.d_next[26] ),
    .B(\u_inv.d_reg[26] ));
 sg13g2_xnor2_1 _30751_ (.Y(_05029_),
    .A(\u_inv.d_next[26] ),
    .B(\u_inv.d_reg[26] ));
 sg13g2_nor2_1 _30752_ (.A(\u_inv.d_next[27] ),
    .B(_14782_),
    .Y(_05030_));
 sg13g2_xnor2_1 _30753_ (.Y(_05031_),
    .A(\u_inv.d_next[27] ),
    .B(\u_inv.d_reg[27] ));
 sg13g2_xor2_1 _30754_ (.B(\u_inv.d_reg[27] ),
    .A(\u_inv.d_next[27] ),
    .X(_05032_));
 sg13g2_nand2_1 _30755_ (.Y(_05033_),
    .A(_05029_),
    .B(_05031_));
 sg13g2_nor2b_1 _30756_ (.A(\u_inv.d_reg[29] ),
    .B_N(\u_inv.d_next[29] ),
    .Y(_05034_));
 sg13g2_nor2b_1 _30757_ (.A(\u_inv.d_reg[28] ),
    .B_N(\u_inv.d_next[28] ),
    .Y(_05035_));
 sg13g2_a21o_1 _30758_ (.A2(_05035_),
    .A1(_05023_),
    .B1(_05034_),
    .X(_05036_));
 sg13g2_and3_1 _30759_ (.X(_05037_),
    .A(_05018_),
    .B(_05020_),
    .C(_05036_));
 sg13g2_nor2b_1 _30760_ (.A(\u_inv.d_reg[30] ),
    .B_N(\u_inv.d_next[30] ),
    .Y(_05038_));
 sg13g2_a21o_1 _30761_ (.A2(_05038_),
    .A1(_05017_),
    .B1(_05016_),
    .X(_05039_));
 sg13g2_nor2b_1 _30762_ (.A(\u_inv.d_reg[26] ),
    .B_N(\u_inv.d_next[26] ),
    .Y(_05040_));
 sg13g2_a21oi_1 _30763_ (.A1(\u_inv.d_next[27] ),
    .A2(_14782_),
    .Y(_05041_),
    .B1(_05040_));
 sg13g2_or2_1 _30764_ (.X(_05042_),
    .B(_05041_),
    .A(_05030_));
 sg13g2_nand2b_1 _30765_ (.Y(_05043_),
    .B(_05015_),
    .A_N(_05033_));
 sg13g2_a21oi_1 _30766_ (.A1(_05042_),
    .A2(_05043_),
    .Y(_05044_),
    .B1(_05027_));
 sg13g2_xor2_1 _30767_ (.B(\u_inv.d_reg[24] ),
    .A(\u_inv.d_next[24] ),
    .X(_05045_));
 sg13g2_nor4_1 _30768_ (.A(_05013_),
    .B(_05027_),
    .C(_05033_),
    .D(_05045_),
    .Y(_05046_));
 sg13g2_xnor2_1 _30769_ (.Y(_05047_),
    .A(\u_inv.d_next[23] ),
    .B(\u_inv.d_reg[23] ));
 sg13g2_xor2_1 _30770_ (.B(\u_inv.d_reg[23] ),
    .A(\u_inv.d_next[23] ),
    .X(_05048_));
 sg13g2_nand2_2 _30771_ (.Y(_05049_),
    .A(\u_inv.d_next[22] ),
    .B(\u_inv.d_reg[22] ));
 sg13g2_or2_1 _30772_ (.X(_05050_),
    .B(\u_inv.d_reg[22] ),
    .A(\u_inv.d_next[22] ));
 sg13g2_nand2_2 _30773_ (.Y(_05051_),
    .A(_05049_),
    .B(_05050_));
 sg13g2_nand2_1 _30774_ (.Y(_05052_),
    .A(_05047_),
    .B(_05051_));
 sg13g2_xnor2_1 _30775_ (.Y(_05053_),
    .A(\u_inv.d_next[21] ),
    .B(\u_inv.d_reg[21] ));
 sg13g2_inv_1 _30776_ (.Y(_05054_),
    .A(_05053_));
 sg13g2_and2_1 _30777_ (.A(\u_inv.d_next[20] ),
    .B(\u_inv.d_reg[20] ),
    .X(_05055_));
 sg13g2_xor2_1 _30778_ (.B(\u_inv.d_reg[20] ),
    .A(\u_inv.d_next[20] ),
    .X(_05056_));
 sg13g2_or2_1 _30779_ (.X(_05057_),
    .B(_05056_),
    .A(_05054_));
 sg13g2_or2_1 _30780_ (.X(_05058_),
    .B(_05057_),
    .A(_05052_));
 sg13g2_nor2_1 _30781_ (.A(\u_inv.d_next[19] ),
    .B(_14790_),
    .Y(_05059_));
 sg13g2_nand2_1 _30782_ (.Y(_05060_),
    .A(\u_inv.d_next[19] ),
    .B(_14790_));
 sg13g2_xor2_1 _30783_ (.B(\u_inv.d_reg[19] ),
    .A(\u_inv.d_next[19] ),
    .X(_05061_));
 sg13g2_xnor2_1 _30784_ (.Y(_05062_),
    .A(\u_inv.d_next[18] ),
    .B(\u_inv.d_reg[18] ));
 sg13g2_nor2b_1 _30785_ (.A(_05061_),
    .B_N(_05062_),
    .Y(_05063_));
 sg13g2_inv_1 _30786_ (.Y(_05064_),
    .A(_05063_));
 sg13g2_nor2b_1 _30787_ (.A(net5873),
    .B_N(\u_inv.d_next[16] ),
    .Y(_05065_));
 sg13g2_a21oi_1 _30788_ (.A1(\u_inv.d_next[17] ),
    .A2(_14792_),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_a21oi_1 _30789_ (.A1(_14238_),
    .A2(\u_inv.d_reg[17] ),
    .Y(_05067_),
    .B1(_05066_));
 sg13g2_nand2_1 _30790_ (.Y(_05068_),
    .A(\u_inv.d_next[18] ),
    .B(_14791_));
 sg13g2_a21oi_1 _30791_ (.A1(_05060_),
    .A2(_05068_),
    .Y(_05069_),
    .B1(_05059_));
 sg13g2_a21oi_1 _30792_ (.A1(_05063_),
    .A2(_05067_),
    .Y(_05070_),
    .B1(_05069_));
 sg13g2_nand2_1 _30793_ (.Y(_05071_),
    .A(\u_inv.d_next[22] ),
    .B(_14787_));
 sg13g2_a21oi_1 _30794_ (.A1(_14236_),
    .A2(\u_inv.d_reg[23] ),
    .Y(_05072_),
    .B1(_05071_));
 sg13g2_a21oi_1 _30795_ (.A1(\u_inv.d_next[23] ),
    .A2(_14786_),
    .Y(_05073_),
    .B1(_05072_));
 sg13g2_nor2_1 _30796_ (.A(_14237_),
    .B(\u_inv.d_reg[21] ),
    .Y(_05074_));
 sg13g2_nor2b_1 _30797_ (.A(\u_inv.d_reg[20] ),
    .B_N(\u_inv.d_next[20] ),
    .Y(_05075_));
 sg13g2_a21oi_1 _30798_ (.A1(_05053_),
    .A2(_05075_),
    .Y(_05076_),
    .B1(_05074_));
 sg13g2_nor2_1 _30799_ (.A(_05052_),
    .B(_05076_),
    .Y(_05077_));
 sg13g2_o21ai_1 _30800_ (.B1(_05073_),
    .Y(_05078_),
    .A1(_05058_),
    .A2(_05070_));
 sg13g2_nor2_1 _30801_ (.A(_05077_),
    .B(_05078_),
    .Y(_05079_));
 sg13g2_nand2_1 _30802_ (.Y(_05080_),
    .A(\u_inv.d_next[14] ),
    .B(_14795_));
 sg13g2_a21oi_1 _30803_ (.A1(_14239_),
    .A2(\u_inv.d_reg[15] ),
    .Y(_05081_),
    .B1(_05080_));
 sg13g2_xnor2_1 _30804_ (.Y(_05082_),
    .A(\u_inv.d_next[15] ),
    .B(\u_inv.d_reg[15] ));
 sg13g2_nand2_2 _30805_ (.Y(_05083_),
    .A(\u_inv.d_next[14] ),
    .B(\u_inv.d_reg[14] ));
 sg13g2_or2_1 _30806_ (.X(_05084_),
    .B(\u_inv.d_reg[14] ),
    .A(\u_inv.d_next[14] ));
 sg13g2_and2_1 _30807_ (.A(_05083_),
    .B(_05084_),
    .X(_05085_));
 sg13g2_nand2_2 _30808_ (.Y(_05086_),
    .A(_05083_),
    .B(_05084_));
 sg13g2_and2_1 _30809_ (.A(_05082_),
    .B(_05086_),
    .X(_05087_));
 sg13g2_xor2_1 _30810_ (.B(\u_inv.d_reg[13] ),
    .A(\u_inv.d_next[13] ),
    .X(_05088_));
 sg13g2_nand2_1 _30811_ (.Y(_05089_),
    .A(\u_inv.d_next[12] ),
    .B(_14797_));
 sg13g2_nor2_1 _30812_ (.A(_05088_),
    .B(_05089_),
    .Y(_05090_));
 sg13g2_nor2_1 _30813_ (.A(_14240_),
    .B(\u_inv.d_reg[13] ),
    .Y(_05091_));
 sg13g2_nand2_1 _30814_ (.Y(_05092_),
    .A(\u_inv.d_next[12] ),
    .B(\u_inv.d_reg[12] ));
 sg13g2_or2_1 _30815_ (.X(_05093_),
    .B(\u_inv.d_reg[12] ),
    .A(\u_inv.d_next[12] ));
 sg13g2_xnor2_1 _30816_ (.Y(_05094_),
    .A(\u_inv.d_next[12] ),
    .B(\u_inv.d_reg[12] ));
 sg13g2_nor2b_1 _30817_ (.A(_05088_),
    .B_N(_05094_),
    .Y(_05095_));
 sg13g2_nand2b_1 _30818_ (.Y(_05096_),
    .B(\u_inv.d_next[11] ),
    .A_N(\u_inv.d_reg[11] ));
 sg13g2_nor2b_1 _30819_ (.A(\u_inv.d_next[11] ),
    .B_N(\u_inv.d_reg[11] ),
    .Y(_05097_));
 sg13g2_nand2b_1 _30820_ (.Y(_05098_),
    .B(\u_inv.d_next[10] ),
    .A_N(\u_inv.d_reg[10] ));
 sg13g2_a21oi_1 _30821_ (.A1(_05096_),
    .A2(_05098_),
    .Y(_05099_),
    .B1(_05097_));
 sg13g2_and2_1 _30822_ (.A(_05095_),
    .B(_05099_),
    .X(_05100_));
 sg13g2_or3_1 _30823_ (.A(_05090_),
    .B(_05091_),
    .C(_05100_),
    .X(_05101_));
 sg13g2_a221oi_1 _30824_ (.B2(_05101_),
    .C1(_05081_),
    .B1(_05087_),
    .A1(\u_inv.d_next[15] ),
    .Y(_05102_),
    .A2(_14794_));
 sg13g2_xnor2_1 _30825_ (.Y(_05103_),
    .A(\u_inv.d_next[11] ),
    .B(net5874));
 sg13g2_xor2_1 _30826_ (.B(net5874),
    .A(\u_inv.d_next[11] ),
    .X(_05104_));
 sg13g2_or2_1 _30827_ (.X(_05105_),
    .B(\u_inv.d_reg[10] ),
    .A(\u_inv.d_next[10] ));
 sg13g2_and2_1 _30828_ (.A(\u_inv.d_next[10] ),
    .B(\u_inv.d_reg[10] ),
    .X(_05106_));
 sg13g2_xor2_1 _30829_ (.B(\u_inv.d_reg[10] ),
    .A(\u_inv.d_next[10] ),
    .X(_05107_));
 sg13g2_nor2_1 _30830_ (.A(_05104_),
    .B(_05107_),
    .Y(_05108_));
 sg13g2_nand3_1 _30831_ (.B(_05095_),
    .C(_05108_),
    .A(_05087_),
    .Y(_05109_));
 sg13g2_nor2b_1 _30832_ (.A(\u_inv.d_reg[9] ),
    .B_N(\u_inv.d_next[9] ),
    .Y(_05110_));
 sg13g2_nand2b_1 _30833_ (.Y(_05111_),
    .B(\u_inv.d_reg[9] ),
    .A_N(\u_inv.d_next[9] ));
 sg13g2_nor2b_1 _30834_ (.A(\u_inv.d_reg[8] ),
    .B_N(\u_inv.d_next[8] ),
    .Y(_05112_));
 sg13g2_a21oi_1 _30835_ (.A1(_05111_),
    .A2(_05112_),
    .Y(_05113_),
    .B1(_05110_));
 sg13g2_inv_1 _30836_ (.Y(_05114_),
    .A(_05113_));
 sg13g2_nor2_1 _30837_ (.A(\u_inv.d_next[7] ),
    .B(_14802_),
    .Y(_05115_));
 sg13g2_nor2b_1 _30838_ (.A(\u_inv.d_reg[7] ),
    .B_N(\u_inv.d_next[7] ),
    .Y(_05116_));
 sg13g2_nor2b_1 _30839_ (.A(\u_inv.d_reg[6] ),
    .B_N(\u_inv.d_next[6] ),
    .Y(_05117_));
 sg13g2_nor2_1 _30840_ (.A(_05116_),
    .B(_05117_),
    .Y(_05118_));
 sg13g2_nand2_1 _30841_ (.Y(_05119_),
    .A(\u_inv.d_next[6] ),
    .B(\u_inv.d_reg[6] ));
 sg13g2_xor2_1 _30842_ (.B(\u_inv.d_reg[6] ),
    .A(\u_inv.d_next[6] ),
    .X(_05120_));
 sg13g2_a21oi_1 _30843_ (.A1(_05118_),
    .A2(_05120_),
    .Y(_05121_),
    .B1(_05115_));
 sg13g2_a21o_1 _30844_ (.A2(_05120_),
    .A1(_05118_),
    .B1(_05115_),
    .X(_05122_));
 sg13g2_nand2_1 _30845_ (.Y(_05123_),
    .A(\u_inv.d_next[4] ),
    .B(_14805_));
 sg13g2_nor2b_1 _30846_ (.A(\u_inv.d_reg[3] ),
    .B_N(\u_inv.d_next[3] ),
    .Y(_05124_));
 sg13g2_xnor2_1 _30847_ (.Y(_05125_),
    .A(\u_inv.d_next[3] ),
    .B(\u_inv.d_reg[3] ));
 sg13g2_and2_1 _30848_ (.A(\u_inv.d_next[2] ),
    .B(\u_inv.d_reg[2] ),
    .X(_05126_));
 sg13g2_xor2_1 _30849_ (.B(\u_inv.d_reg[2] ),
    .A(\u_inv.d_next[2] ),
    .X(_05127_));
 sg13g2_nor2b_1 _30850_ (.A(\u_inv.d_reg[1] ),
    .B_N(\u_inv.d_next[1] ),
    .Y(_05128_));
 sg13g2_nand2_1 _30851_ (.Y(_05129_),
    .A(\u_inv.d_next[1] ),
    .B(\u_inv.d_reg[1] ));
 sg13g2_xnor2_1 _30852_ (.Y(_05130_),
    .A(\u_inv.d_next[1] ),
    .B(\u_inv.d_reg[1] ));
 sg13g2_nand2b_1 _30853_ (.Y(_05131_),
    .B(\u_inv.d_reg[0] ),
    .A_N(\u_inv.d_next[0] ));
 sg13g2_a21oi_1 _30854_ (.A1(_05130_),
    .A2(_05131_),
    .Y(_05132_),
    .B1(_05128_));
 sg13g2_nand2_1 _30855_ (.Y(_05133_),
    .A(\u_inv.d_next[2] ),
    .B(_14807_));
 sg13g2_o21ai_1 _30856_ (.B1(_05133_),
    .Y(_05134_),
    .A1(_05127_),
    .A2(_05132_));
 sg13g2_a21oi_1 _30857_ (.A1(_05125_),
    .A2(_05134_),
    .Y(_05135_),
    .B1(_05124_));
 sg13g2_nand2_1 _30858_ (.Y(_05136_),
    .A(\u_inv.d_next[4] ),
    .B(\u_inv.d_reg[4] ));
 sg13g2_xor2_1 _30859_ (.B(\u_inv.d_reg[4] ),
    .A(\u_inv.d_next[4] ),
    .X(_05137_));
 sg13g2_xnor2_1 _30860_ (.Y(_05138_),
    .A(\u_inv.d_next[4] ),
    .B(\u_inv.d_reg[4] ));
 sg13g2_o21ai_1 _30861_ (.B1(_05123_),
    .Y(_05139_),
    .A1(_05135_),
    .A2(_05137_));
 sg13g2_a21oi_1 _30862_ (.A1(_14241_),
    .A2(\u_inv.d_reg[5] ),
    .Y(_05140_),
    .B1(_05123_));
 sg13g2_a21oi_1 _30863_ (.A1(\u_inv.d_next[5] ),
    .A2(_14804_),
    .Y(_05141_),
    .B1(_05140_));
 sg13g2_xnor2_1 _30864_ (.Y(_05142_),
    .A(\u_inv.d_next[5] ),
    .B(\u_inv.d_reg[5] ));
 sg13g2_nand3b_1 _30865_ (.B(_05138_),
    .C(_05142_),
    .Y(_05143_),
    .A_N(_05135_));
 sg13g2_and2_1 _30866_ (.A(_05141_),
    .B(_05143_),
    .X(_05144_));
 sg13g2_and2_1 _30867_ (.A(_05118_),
    .B(_05144_),
    .X(_05145_));
 sg13g2_nand3_1 _30868_ (.B(_05141_),
    .C(_05143_),
    .A(_05118_),
    .Y(_05146_));
 sg13g2_nor2_2 _30869_ (.A(_05122_),
    .B(_05145_),
    .Y(_05147_));
 sg13g2_xnor2_1 _30870_ (.Y(_05148_),
    .A(\u_inv.d_next[9] ),
    .B(\u_inv.d_reg[9] ));
 sg13g2_nand2b_1 _30871_ (.Y(_05149_),
    .B(_05111_),
    .A_N(_05110_));
 sg13g2_nand2_1 _30872_ (.Y(_05150_),
    .A(\u_inv.d_next[8] ),
    .B(\u_inv.d_reg[8] ));
 sg13g2_xor2_1 _30873_ (.B(\u_inv.d_reg[8] ),
    .A(\u_inv.d_next[8] ),
    .X(_05151_));
 sg13g2_nor2_1 _30874_ (.A(_05149_),
    .B(_05151_),
    .Y(_05152_));
 sg13g2_a21oi_1 _30875_ (.A1(_05147_),
    .A2(_05152_),
    .Y(_05153_),
    .B1(_05114_));
 sg13g2_a21o_1 _30876_ (.A2(_05152_),
    .A1(_05147_),
    .B1(_05114_),
    .X(_05154_));
 sg13g2_nor2b_1 _30877_ (.A(_05109_),
    .B_N(_05152_),
    .Y(_05155_));
 sg13g2_and3_2 _30878_ (.X(_05156_),
    .A(_05121_),
    .B(_05146_),
    .C(_05155_));
 sg13g2_nand3_1 _30879_ (.B(_05146_),
    .C(_05155_),
    .A(_05121_),
    .Y(_05157_));
 sg13g2_o21ai_1 _30880_ (.B1(_05102_),
    .Y(_05158_),
    .A1(_05109_),
    .A2(_05113_));
 sg13g2_inv_1 _30881_ (.Y(_05159_),
    .A(_05158_));
 sg13g2_nor2_1 _30882_ (.A(_05156_),
    .B(_05158_),
    .Y(_05160_));
 sg13g2_xnor2_1 _30883_ (.Y(_05161_),
    .A(\u_inv.d_next[17] ),
    .B(\u_inv.d_reg[17] ));
 sg13g2_nand2_1 _30884_ (.Y(_05162_),
    .A(\u_inv.d_next[16] ),
    .B(net5873));
 sg13g2_xor2_1 _30885_ (.B(net5873),
    .A(\u_inv.d_next[16] ),
    .X(_05163_));
 sg13g2_xnor2_1 _30886_ (.Y(_05164_),
    .A(\u_inv.d_next[16] ),
    .B(net5873));
 sg13g2_nand2_1 _30887_ (.Y(_05165_),
    .A(_05161_),
    .B(_05164_));
 sg13g2_nor3_1 _30888_ (.A(_05058_),
    .B(_05064_),
    .C(_05165_),
    .Y(_05166_));
 sg13g2_o21ai_1 _30889_ (.B1(_05166_),
    .Y(_05167_),
    .A1(_05156_),
    .A2(_05158_));
 sg13g2_nor2b_1 _30890_ (.A(_05079_),
    .B_N(_05046_),
    .Y(_05168_));
 sg13g2_nor4_1 _30891_ (.A(_05037_),
    .B(_05039_),
    .C(_05044_),
    .D(_05168_),
    .Y(_05169_));
 sg13g2_nand2_1 _30892_ (.Y(_05170_),
    .A(_05046_),
    .B(_05166_));
 sg13g2_a21o_2 _30893_ (.A2(_05159_),
    .A1(_05157_),
    .B1(_05170_),
    .X(_05171_));
 sg13g2_nand2_2 _30894_ (.Y(_05172_),
    .A(_05169_),
    .B(_05171_));
 sg13g2_nor2b_1 _30895_ (.A(\u_inv.d_reg[47] ),
    .B_N(\u_inv.d_next[47] ),
    .Y(_05173_));
 sg13g2_nand2b_1 _30896_ (.Y(_05174_),
    .B(\u_inv.d_reg[47] ),
    .A_N(\u_inv.d_next[47] ));
 sg13g2_nor2b_2 _30897_ (.A(_05173_),
    .B_N(_05174_),
    .Y(_05175_));
 sg13g2_nand2_1 _30898_ (.Y(_05176_),
    .A(\u_inv.d_next[46] ),
    .B(\u_inv.d_reg[46] ));
 sg13g2_xnor2_1 _30899_ (.Y(_05177_),
    .A(\u_inv.d_next[46] ),
    .B(\u_inv.d_reg[46] ));
 sg13g2_nand2_2 _30900_ (.Y(_05178_),
    .A(_05175_),
    .B(_05177_));
 sg13g2_nor2_1 _30901_ (.A(\u_inv.d_next[45] ),
    .B(\u_inv.d_reg[45] ),
    .Y(_05179_));
 sg13g2_nand2_1 _30902_ (.Y(_05180_),
    .A(\u_inv.d_next[45] ),
    .B(\u_inv.d_reg[45] ));
 sg13g2_nor2b_1 _30903_ (.A(_05179_),
    .B_N(_05180_),
    .Y(_05181_));
 sg13g2_nand2b_2 _30904_ (.Y(_05182_),
    .B(_05180_),
    .A_N(_05179_));
 sg13g2_nand2_1 _30905_ (.Y(_05183_),
    .A(\u_inv.d_next[44] ),
    .B(\u_inv.d_reg[44] ));
 sg13g2_xnor2_1 _30906_ (.Y(_05184_),
    .A(\u_inv.d_next[44] ),
    .B(\u_inv.d_reg[44] ));
 sg13g2_nand2_2 _30907_ (.Y(_05185_),
    .A(_05182_),
    .B(_05184_));
 sg13g2_nor2_1 _30908_ (.A(_05178_),
    .B(_05185_),
    .Y(_05186_));
 sg13g2_xnor2_1 _30909_ (.Y(_05187_),
    .A(\u_inv.d_next[41] ),
    .B(\u_inv.d_reg[41] ));
 sg13g2_inv_2 _30910_ (.Y(_05188_),
    .A(_05187_));
 sg13g2_nand2_1 _30911_ (.Y(_05189_),
    .A(\u_inv.d_next[40] ),
    .B(\u_inv.d_reg[40] ));
 sg13g2_xor2_1 _30912_ (.B(\u_inv.d_reg[40] ),
    .A(\u_inv.d_next[40] ),
    .X(_05190_));
 sg13g2_xnor2_1 _30913_ (.Y(_05191_),
    .A(\u_inv.d_next[40] ),
    .B(\u_inv.d_reg[40] ));
 sg13g2_nand2_1 _30914_ (.Y(_05192_),
    .A(_05187_),
    .B(_05191_));
 sg13g2_nor2b_1 _30915_ (.A(\u_inv.d_next[43] ),
    .B_N(\u_inv.d_reg[43] ),
    .Y(_05193_));
 sg13g2_nand2b_1 _30916_ (.Y(_05194_),
    .B(\u_inv.d_next[43] ),
    .A_N(\u_inv.d_reg[43] ));
 sg13g2_nand2b_2 _30917_ (.Y(_05195_),
    .B(_05194_),
    .A_N(_05193_));
 sg13g2_nor2_1 _30918_ (.A(_14231_),
    .B(_14767_),
    .Y(_05196_));
 sg13g2_nand2_1 _30919_ (.Y(_05197_),
    .A(\u_inv.d_next[42] ),
    .B(\u_inv.d_reg[42] ));
 sg13g2_nand2_2 _30920_ (.Y(_05198_),
    .A(_14231_),
    .B(_14767_));
 sg13g2_nand2_2 _30921_ (.Y(_05199_),
    .A(_05197_),
    .B(_05198_));
 sg13g2_a21oi_1 _30922_ (.A1(_05197_),
    .A2(_05198_),
    .Y(_05200_),
    .B1(_05195_));
 sg13g2_nand2b_1 _30923_ (.Y(_05201_),
    .B(_05199_),
    .A_N(_05195_));
 sg13g2_nor4_2 _30924_ (.A(_05178_),
    .B(_05185_),
    .C(_05192_),
    .Y(_05202_),
    .D(_05201_));
 sg13g2_nor2b_1 _30925_ (.A(\u_inv.d_reg[39] ),
    .B_N(\u_inv.d_next[39] ),
    .Y(_05203_));
 sg13g2_nand2b_1 _30926_ (.Y(_05204_),
    .B(\u_inv.d_reg[39] ),
    .A_N(\u_inv.d_next[39] ));
 sg13g2_nor2b_2 _30927_ (.A(_05203_),
    .B_N(_05204_),
    .Y(_05205_));
 sg13g2_nand2_1 _30928_ (.Y(_05206_),
    .A(\u_inv.d_next[38] ),
    .B(\u_inv.d_reg[38] ));
 sg13g2_or2_1 _30929_ (.X(_05207_),
    .B(\u_inv.d_reg[38] ),
    .A(\u_inv.d_next[38] ));
 sg13g2_nand2_2 _30930_ (.Y(_05208_),
    .A(_05206_),
    .B(_05207_));
 sg13g2_and2_1 _30931_ (.A(_05205_),
    .B(_05208_),
    .X(_05209_));
 sg13g2_nor2_1 _30932_ (.A(\u_inv.d_next[37] ),
    .B(\u_inv.d_reg[37] ),
    .Y(_05210_));
 sg13g2_xor2_1 _30933_ (.B(\u_inv.d_reg[37] ),
    .A(\u_inv.d_next[37] ),
    .X(_05211_));
 sg13g2_nand2_1 _30934_ (.Y(_05212_),
    .A(\u_inv.d_next[36] ),
    .B(\u_inv.d_reg[36] ));
 sg13g2_xor2_1 _30935_ (.B(\u_inv.d_reg[36] ),
    .A(\u_inv.d_next[36] ),
    .X(_05213_));
 sg13g2_xnor2_1 _30936_ (.Y(_05214_),
    .A(\u_inv.d_next[36] ),
    .B(\u_inv.d_reg[36] ));
 sg13g2_nor2_1 _30937_ (.A(_05211_),
    .B(_05213_),
    .Y(_05215_));
 sg13g2_nand2_1 _30938_ (.Y(_05216_),
    .A(_05209_),
    .B(_05215_));
 sg13g2_xnor2_1 _30939_ (.Y(_05217_),
    .A(\u_inv.d_next[34] ),
    .B(\u_inv.d_reg[34] ));
 sg13g2_xnor2_1 _30940_ (.Y(_05218_),
    .A(\u_inv.d_next[35] ),
    .B(\u_inv.d_reg[35] ));
 sg13g2_nand2_1 _30941_ (.Y(_05219_),
    .A(_05217_),
    .B(_05218_));
 sg13g2_nor2b_1 _30942_ (.A(\u_inv.d_reg[33] ),
    .B_N(\u_inv.d_next[33] ),
    .Y(_05220_));
 sg13g2_nand2b_1 _30943_ (.Y(_05221_),
    .B(\u_inv.d_reg[33] ),
    .A_N(\u_inv.d_next[33] ));
 sg13g2_xor2_1 _30944_ (.B(\u_inv.d_reg[33] ),
    .A(\u_inv.d_next[33] ),
    .X(_05222_));
 sg13g2_and2_1 _30945_ (.A(\u_inv.d_next[32] ),
    .B(\u_inv.d_reg[32] ),
    .X(_05223_));
 sg13g2_xor2_1 _30946_ (.B(\u_inv.d_reg[32] ),
    .A(\u_inv.d_next[32] ),
    .X(_05224_));
 sg13g2_inv_1 _30947_ (.Y(_05225_),
    .A(_05224_));
 sg13g2_nor2_1 _30948_ (.A(net5618),
    .B(_05224_),
    .Y(_05226_));
 sg13g2_nor4_1 _30949_ (.A(_05216_),
    .B(_05219_),
    .C(net5618),
    .D(_05224_),
    .Y(_05227_));
 sg13g2_and2_1 _30950_ (.A(_05202_),
    .B(_05227_),
    .X(_05228_));
 sg13g2_inv_1 _30951_ (.Y(_05229_),
    .A(_05228_));
 sg13g2_a21o_2 _30952_ (.A2(_05171_),
    .A1(_05169_),
    .B1(_05229_),
    .X(_05230_));
 sg13g2_nor2b_1 _30953_ (.A(\u_inv.d_reg[32] ),
    .B_N(\u_inv.d_next[32] ),
    .Y(_05231_));
 sg13g2_a21oi_1 _30954_ (.A1(_05221_),
    .A2(_05231_),
    .Y(_05232_),
    .B1(_05220_));
 sg13g2_nor2_1 _30955_ (.A(_05219_),
    .B(_05232_),
    .Y(_05233_));
 sg13g2_nor2_1 _30956_ (.A(_14235_),
    .B(\u_inv.d_reg[34] ),
    .Y(_05234_));
 sg13g2_a21oi_1 _30957_ (.A1(\u_inv.d_next[35] ),
    .A2(_14774_),
    .Y(_05235_),
    .B1(_05234_));
 sg13g2_a21oi_1 _30958_ (.A1(_14234_),
    .A2(\u_inv.d_reg[35] ),
    .Y(_05236_),
    .B1(_05235_));
 sg13g2_inv_1 _30959_ (.Y(_05237_),
    .A(_05236_));
 sg13g2_nor2_1 _30960_ (.A(_05233_),
    .B(_05236_),
    .Y(_05238_));
 sg13g2_nor2b_1 _30961_ (.A(\u_inv.d_reg[36] ),
    .B_N(\u_inv.d_next[36] ),
    .Y(_05239_));
 sg13g2_nand2b_1 _30962_ (.Y(_05240_),
    .B(_05239_),
    .A_N(_05211_));
 sg13g2_o21ai_1 _30963_ (.B1(_05240_),
    .Y(_05241_),
    .A1(_14233_),
    .A2(\u_inv.d_reg[37] ));
 sg13g2_nor2b_1 _30964_ (.A(\u_inv.d_reg[38] ),
    .B_N(\u_inv.d_next[38] ),
    .Y(_05242_));
 sg13g2_a221oi_1 _30965_ (.B2(_05204_),
    .C1(_05203_),
    .B1(_05242_),
    .A1(_05209_),
    .Y(_05243_),
    .A2(_05241_));
 sg13g2_o21ai_1 _30966_ (.B1(_05243_),
    .Y(_05244_),
    .A1(_05216_),
    .A2(_05238_));
 sg13g2_nor2b_1 _30967_ (.A(\u_inv.d_reg[45] ),
    .B_N(\u_inv.d_next[45] ),
    .Y(_05245_));
 sg13g2_nor2b_1 _30968_ (.A(\u_inv.d_reg[44] ),
    .B_N(\u_inv.d_next[44] ),
    .Y(_05246_));
 sg13g2_a21oi_1 _30969_ (.A1(_05182_),
    .A2(_05246_),
    .Y(_05247_),
    .B1(_05245_));
 sg13g2_nor2b_1 _30970_ (.A(\u_inv.d_reg[46] ),
    .B_N(\u_inv.d_next[46] ),
    .Y(_05248_));
 sg13g2_a21oi_1 _30971_ (.A1(_05174_),
    .A2(_05248_),
    .Y(_05249_),
    .B1(_05173_));
 sg13g2_o21ai_1 _30972_ (.B1(_05249_),
    .Y(_05250_),
    .A1(_05178_),
    .A2(_05247_));
 sg13g2_nor2_1 _30973_ (.A(_14232_),
    .B(\u_inv.d_reg[41] ),
    .Y(_05251_));
 sg13g2_nor2b_1 _30974_ (.A(\u_inv.d_reg[40] ),
    .B_N(\u_inv.d_next[40] ),
    .Y(_05252_));
 sg13g2_a21oi_1 _30975_ (.A1(_05187_),
    .A2(_05252_),
    .Y(_05253_),
    .B1(_05251_));
 sg13g2_nand2_1 _30976_ (.Y(_05254_),
    .A(\u_inv.d_next[42] ),
    .B(_14767_));
 sg13g2_a21oi_1 _30977_ (.A1(_05194_),
    .A2(_05254_),
    .Y(_05255_),
    .B1(_05193_));
 sg13g2_inv_1 _30978_ (.Y(_05256_),
    .A(_05255_));
 sg13g2_o21ai_1 _30979_ (.B1(_05256_),
    .Y(_05257_),
    .A1(_05201_),
    .A2(_05253_));
 sg13g2_a221oi_1 _30980_ (.B2(_05186_),
    .C1(_05250_),
    .B1(_05257_),
    .A1(_05202_),
    .Y(_05258_),
    .A2(_05244_));
 sg13g2_and2_1 _30981_ (.A(_05230_),
    .B(_05258_),
    .X(_05259_));
 sg13g2_and2_1 _30982_ (.A(\u_inv.d_next[48] ),
    .B(\u_inv.d_reg[48] ),
    .X(_05260_));
 sg13g2_nand2_1 _30983_ (.Y(_05261_),
    .A(\u_inv.d_next[48] ),
    .B(\u_inv.d_reg[48] ));
 sg13g2_or2_1 _30984_ (.X(_05262_),
    .B(\u_inv.d_reg[48] ),
    .A(\u_inv.d_next[48] ));
 sg13g2_and2_1 _30985_ (.A(_05261_),
    .B(_05262_),
    .X(_05263_));
 sg13g2_nor2_1 _30986_ (.A(\u_inv.d_next[49] ),
    .B(_14760_),
    .Y(_05264_));
 sg13g2_nand2_1 _30987_ (.Y(_05265_),
    .A(\u_inv.d_next[49] ),
    .B(_14760_));
 sg13g2_xor2_1 _30988_ (.B(\u_inv.d_reg[49] ),
    .A(\u_inv.d_next[49] ),
    .X(_05266_));
 sg13g2_xor2_1 _30989_ (.B(\u_inv.d_reg[63] ),
    .A(\u_inv.d_next[63] ),
    .X(_05267_));
 sg13g2_xnor2_1 _30990_ (.Y(_05268_),
    .A(\u_inv.d_next[63] ),
    .B(\u_inv.d_reg[63] ));
 sg13g2_nand2_1 _30991_ (.Y(_05269_),
    .A(\u_inv.d_next[62] ),
    .B(\u_inv.d_reg[62] ));
 sg13g2_xor2_1 _30992_ (.B(\u_inv.d_reg[62] ),
    .A(\u_inv.d_next[62] ),
    .X(_05270_));
 sg13g2_nor2_1 _30993_ (.A(_05267_),
    .B(_05270_),
    .Y(_05271_));
 sg13g2_nand2_1 _30994_ (.Y(_05272_),
    .A(\u_inv.d_next[61] ),
    .B(_14748_));
 sg13g2_nor2_1 _30995_ (.A(\u_inv.d_next[61] ),
    .B(_14748_),
    .Y(_05273_));
 sg13g2_xnor2_1 _30996_ (.Y(_05274_),
    .A(\u_inv.d_next[61] ),
    .B(\u_inv.d_reg[61] ));
 sg13g2_nand2_2 _30997_ (.Y(_05275_),
    .A(\u_inv.d_next[60] ),
    .B(\u_inv.d_reg[60] ));
 sg13g2_or2_1 _30998_ (.X(_05276_),
    .B(\u_inv.d_reg[60] ),
    .A(\u_inv.d_next[60] ));
 sg13g2_nand2_2 _30999_ (.Y(_05277_),
    .A(_05275_),
    .B(_05276_));
 sg13g2_and2_1 _31000_ (.A(_05274_),
    .B(_05277_),
    .X(_05278_));
 sg13g2_nand2_1 _31001_ (.Y(_05279_),
    .A(_05271_),
    .B(_05278_));
 sg13g2_xnor2_1 _31002_ (.Y(_05280_),
    .A(\u_inv.d_next[57] ),
    .B(\u_inv.d_reg[57] ));
 sg13g2_nand2_1 _31003_ (.Y(_05281_),
    .A(\u_inv.d_next[56] ),
    .B(\u_inv.d_reg[56] ));
 sg13g2_xor2_1 _31004_ (.B(\u_inv.d_reg[56] ),
    .A(\u_inv.d_next[56] ),
    .X(_05282_));
 sg13g2_nand2b_1 _31005_ (.Y(_05283_),
    .B(_05280_),
    .A_N(_05282_));
 sg13g2_nor2_2 _31006_ (.A(\u_inv.d_next[59] ),
    .B(_14750_),
    .Y(_05284_));
 sg13g2_nor2b_1 _31007_ (.A(\u_inv.d_reg[59] ),
    .B_N(\u_inv.d_next[59] ),
    .Y(_05285_));
 sg13g2_nor2_2 _31008_ (.A(_05284_),
    .B(_05285_),
    .Y(_05286_));
 sg13g2_nand2_1 _31009_ (.Y(_05287_),
    .A(\u_inv.d_next[58] ),
    .B(\u_inv.d_reg[58] ));
 sg13g2_xnor2_1 _31010_ (.Y(_05288_),
    .A(\u_inv.d_next[58] ),
    .B(\u_inv.d_reg[58] ));
 sg13g2_and2_1 _31011_ (.A(_05286_),
    .B(_05288_),
    .X(_05289_));
 sg13g2_nand2_1 _31012_ (.Y(_05290_),
    .A(_05286_),
    .B(_05288_));
 sg13g2_or3_1 _31013_ (.A(_05279_),
    .B(_05283_),
    .C(_05290_),
    .X(_05291_));
 sg13g2_xnor2_1 _31014_ (.Y(_05292_),
    .A(\u_inv.d_next[55] ),
    .B(\u_inv.d_reg[55] ));
 sg13g2_inv_2 _31015_ (.Y(_05293_),
    .A(_05292_));
 sg13g2_nand2_1 _31016_ (.Y(_05294_),
    .A(\u_inv.d_next[54] ),
    .B(\u_inv.d_reg[54] ));
 sg13g2_or2_1 _31017_ (.X(_05295_),
    .B(\u_inv.d_reg[54] ),
    .A(\u_inv.d_next[54] ));
 sg13g2_and2_1 _31018_ (.A(_05294_),
    .B(_05295_),
    .X(_05296_));
 sg13g2_nand2_1 _31019_ (.Y(_05297_),
    .A(_05294_),
    .B(_05295_));
 sg13g2_nand2_1 _31020_ (.Y(_05298_),
    .A(_05292_),
    .B(_05297_));
 sg13g2_xor2_1 _31021_ (.B(\u_inv.d_reg[53] ),
    .A(\u_inv.d_next[53] ),
    .X(_05299_));
 sg13g2_xnor2_1 _31022_ (.Y(_05300_),
    .A(\u_inv.d_next[53] ),
    .B(\u_inv.d_reg[53] ));
 sg13g2_and2_1 _31023_ (.A(\u_inv.d_next[52] ),
    .B(\u_inv.d_reg[52] ),
    .X(_05301_));
 sg13g2_xor2_1 _31024_ (.B(\u_inv.d_reg[52] ),
    .A(\u_inv.d_next[52] ),
    .X(_05302_));
 sg13g2_or3_1 _31025_ (.A(_05298_),
    .B(_05299_),
    .C(_05302_),
    .X(_05303_));
 sg13g2_nand2_1 _31026_ (.Y(_05304_),
    .A(\u_inv.d_next[50] ),
    .B(\u_inv.d_reg[50] ));
 sg13g2_xor2_1 _31027_ (.B(\u_inv.d_reg[50] ),
    .A(\u_inv.d_next[50] ),
    .X(_05305_));
 sg13g2_xnor2_1 _31028_ (.Y(_05306_),
    .A(\u_inv.d_next[50] ),
    .B(\u_inv.d_reg[50] ));
 sg13g2_nand2b_1 _31029_ (.Y(_05307_),
    .B(\u_inv.d_reg[51] ),
    .A_N(\u_inv.d_next[51] ));
 sg13g2_nor2b_1 _31030_ (.A(\u_inv.d_reg[51] ),
    .B_N(\u_inv.d_next[51] ),
    .Y(_05308_));
 sg13g2_xor2_1 _31031_ (.B(\u_inv.d_reg[51] ),
    .A(\u_inv.d_next[51] ),
    .X(_05309_));
 sg13g2_nor2_1 _31032_ (.A(_05305_),
    .B(_05309_),
    .Y(_05310_));
 sg13g2_nor2b_1 _31033_ (.A(_05303_),
    .B_N(_05310_),
    .Y(_05311_));
 sg13g2_nor3_1 _31034_ (.A(_05263_),
    .B(net5617),
    .C(_05291_),
    .Y(_05312_));
 sg13g2_nand2_1 _31035_ (.Y(_05313_),
    .A(_05311_),
    .B(_05312_));
 sg13g2_a21oi_2 _31036_ (.B1(_05313_),
    .Y(_05314_),
    .A2(_05258_),
    .A1(_05230_));
 sg13g2_a21o_2 _31037_ (.A2(_05258_),
    .A1(_05230_),
    .B1(_05313_),
    .X(_05315_));
 sg13g2_nor2b_2 _31038_ (.A(\u_inv.d_reg[50] ),
    .B_N(\u_inv.d_next[50] ),
    .Y(_05316_));
 sg13g2_a21oi_2 _31039_ (.B1(_05308_),
    .Y(_05317_),
    .A2(_05316_),
    .A1(_05307_));
 sg13g2_nor2b_1 _31040_ (.A(\u_inv.d_reg[52] ),
    .B_N(\u_inv.d_next[52] ),
    .Y(_05318_));
 sg13g2_nand2_1 _31041_ (.Y(_05319_),
    .A(_05300_),
    .B(_05318_));
 sg13g2_o21ai_1 _31042_ (.B1(_05319_),
    .Y(_05320_),
    .A1(_14230_),
    .A2(\u_inv.d_reg[53] ));
 sg13g2_nor2b_1 _31043_ (.A(_05298_),
    .B_N(_05320_),
    .Y(_05321_));
 sg13g2_nand2_1 _31044_ (.Y(_05322_),
    .A(\u_inv.d_next[54] ),
    .B(_14755_));
 sg13g2_a21oi_1 _31045_ (.A1(_14229_),
    .A2(\u_inv.d_reg[55] ),
    .Y(_05323_),
    .B1(_05322_));
 sg13g2_a21oi_1 _31046_ (.A1(\u_inv.d_next[55] ),
    .A2(_14754_),
    .Y(_05324_),
    .B1(_05323_));
 sg13g2_o21ai_1 _31047_ (.B1(_05324_),
    .Y(_05325_),
    .A1(_05303_),
    .A2(_05317_));
 sg13g2_nor2_2 _31048_ (.A(_05321_),
    .B(_05325_),
    .Y(_05326_));
 sg13g2_nand2_1 _31049_ (.Y(_05327_),
    .A(\u_inv.d_next[48] ),
    .B(_14761_));
 sg13g2_a21oi_2 _31050_ (.B1(_05264_),
    .Y(_05328_),
    .A2(_05327_),
    .A1(_05265_));
 sg13g2_nand2_1 _31051_ (.Y(_05329_),
    .A(\u_inv.d_next[60] ),
    .B(_14749_));
 sg13g2_o21ai_1 _31052_ (.B1(_05272_),
    .Y(_05330_),
    .A1(_05273_),
    .A2(_05329_));
 sg13g2_inv_1 _31053_ (.Y(_05331_),
    .A(_05330_));
 sg13g2_nor2_1 _31054_ (.A(_14226_),
    .B(\u_inv.d_reg[63] ),
    .Y(_05332_));
 sg13g2_nor2b_1 _31055_ (.A(\u_inv.d_reg[62] ),
    .B_N(\u_inv.d_next[62] ),
    .Y(_05333_));
 sg13g2_nor2b_1 _31056_ (.A(\u_inv.d_reg[56] ),
    .B_N(\u_inv.d_next[56] ),
    .Y(_05334_));
 sg13g2_o21ai_1 _31057_ (.B1(_05334_),
    .Y(_05335_),
    .A1(\u_inv.d_next[57] ),
    .A2(_14752_));
 sg13g2_o21ai_1 _31058_ (.B1(_05335_),
    .Y(_05336_),
    .A1(_14228_),
    .A2(\u_inv.d_reg[57] ));
 sg13g2_inv_1 _31059_ (.Y(_05337_),
    .A(_05336_));
 sg13g2_nand2_1 _31060_ (.Y(_05338_),
    .A(\u_inv.d_next[58] ),
    .B(_14751_));
 sg13g2_a21oi_1 _31061_ (.A1(\u_inv.d_next[58] ),
    .A2(_14751_),
    .Y(_05339_),
    .B1(_05285_));
 sg13g2_nor2_2 _31062_ (.A(_05284_),
    .B(_05339_),
    .Y(_05340_));
 sg13g2_a21oi_1 _31063_ (.A1(_05289_),
    .A2(_05336_),
    .Y(_05341_),
    .B1(_05340_));
 sg13g2_nand2_1 _31064_ (.Y(_05342_),
    .A(_05311_),
    .B(_05328_));
 sg13g2_a21oi_2 _31065_ (.B1(_05291_),
    .Y(_05343_),
    .A2(_05342_),
    .A1(_05326_));
 sg13g2_a22oi_1 _31066_ (.Y(_05344_),
    .B1(_05333_),
    .B2(_05268_),
    .A2(_05330_),
    .A1(_05271_));
 sg13g2_o21ai_1 _31067_ (.B1(_05344_),
    .Y(_05345_),
    .A1(_05279_),
    .A2(_05341_));
 sg13g2_nor3_2 _31068_ (.A(_05332_),
    .B(_05343_),
    .C(_05345_),
    .Y(_05346_));
 sg13g2_inv_1 _31069_ (.Y(_05347_),
    .A(_05346_));
 sg13g2_nand2_2 _31070_ (.Y(_05348_),
    .A(_05315_),
    .B(_05346_));
 sg13g2_xnor2_1 _31071_ (.Y(_05349_),
    .A(\u_inv.d_next[79] ),
    .B(\u_inv.d_reg[79] ));
 sg13g2_xor2_1 _31072_ (.B(\u_inv.d_reg[79] ),
    .A(\u_inv.d_next[79] ),
    .X(_05350_));
 sg13g2_nand2_1 _31073_ (.Y(_05351_),
    .A(\u_inv.d_next[78] ),
    .B(\u_inv.d_reg[78] ));
 sg13g2_xnor2_1 _31074_ (.Y(_05352_),
    .A(\u_inv.d_next[78] ),
    .B(\u_inv.d_reg[78] ));
 sg13g2_inv_1 _31075_ (.Y(_05353_),
    .A(_05352_));
 sg13g2_nand2_2 _31076_ (.Y(_05354_),
    .A(_05349_),
    .B(_05352_));
 sg13g2_xor2_1 _31077_ (.B(net5872),
    .A(\u_inv.d_next[77] ),
    .X(_05355_));
 sg13g2_xnor2_1 _31078_ (.Y(_05356_),
    .A(\u_inv.d_next[77] ),
    .B(net5872));
 sg13g2_and2_1 _31079_ (.A(\u_inv.d_next[76] ),
    .B(\u_inv.d_reg[76] ),
    .X(_05357_));
 sg13g2_xor2_1 _31080_ (.B(\u_inv.d_reg[76] ),
    .A(\u_inv.d_next[76] ),
    .X(_05358_));
 sg13g2_xnor2_1 _31081_ (.Y(_05359_),
    .A(\u_inv.d_next[76] ),
    .B(\u_inv.d_reg[76] ));
 sg13g2_nand2_1 _31082_ (.Y(_05360_),
    .A(_05356_),
    .B(_05359_));
 sg13g2_nor2_1 _31083_ (.A(_05354_),
    .B(_05360_),
    .Y(_05361_));
 sg13g2_nor2_1 _31084_ (.A(\u_inv.d_next[75] ),
    .B(_14734_),
    .Y(_05362_));
 sg13g2_nand2_1 _31085_ (.Y(_05363_),
    .A(\u_inv.d_next[75] ),
    .B(_14734_));
 sg13g2_nor2b_2 _31086_ (.A(_05362_),
    .B_N(_05363_),
    .Y(_05364_));
 sg13g2_nand2b_2 _31087_ (.Y(_05365_),
    .B(_05363_),
    .A_N(_05362_));
 sg13g2_xor2_1 _31088_ (.B(\u_inv.d_reg[74] ),
    .A(net5877),
    .X(_05366_));
 sg13g2_xnor2_1 _31089_ (.Y(_05367_),
    .A(net5877),
    .B(\u_inv.d_reg[74] ));
 sg13g2_nand2_2 _31090_ (.Y(_05368_),
    .A(_05364_),
    .B(_05367_));
 sg13g2_nor2_1 _31091_ (.A(\u_inv.d_next[73] ),
    .B(\u_inv.d_reg[73] ),
    .Y(_05369_));
 sg13g2_xnor2_1 _31092_ (.Y(_05370_),
    .A(\u_inv.d_next[73] ),
    .B(\u_inv.d_reg[73] ));
 sg13g2_and2_1 _31093_ (.A(net5878),
    .B(\u_inv.d_reg[72] ),
    .X(_05371_));
 sg13g2_xor2_1 _31094_ (.B(\u_inv.d_reg[72] ),
    .A(net5878),
    .X(_05372_));
 sg13g2_xnor2_1 _31095_ (.Y(_05373_),
    .A(net5878),
    .B(\u_inv.d_reg[72] ));
 sg13g2_nand2_2 _31096_ (.Y(_05374_),
    .A(_05370_),
    .B(_05373_));
 sg13g2_nor4_2 _31097_ (.A(_05354_),
    .B(_05360_),
    .C(_05368_),
    .Y(_05375_),
    .D(_05374_));
 sg13g2_nand2_1 _31098_ (.Y(_05376_),
    .A(\u_inv.d_next[71] ),
    .B(_14738_));
 sg13g2_xor2_1 _31099_ (.B(\u_inv.d_reg[71] ),
    .A(\u_inv.d_next[71] ),
    .X(_05377_));
 sg13g2_nand2_1 _31100_ (.Y(_05378_),
    .A(net5879),
    .B(\u_inv.d_reg[70] ));
 sg13g2_nor2_1 _31101_ (.A(net5879),
    .B(\u_inv.d_reg[70] ),
    .Y(_05379_));
 sg13g2_xor2_1 _31102_ (.B(\u_inv.d_reg[70] ),
    .A(net5879),
    .X(_05380_));
 sg13g2_nor2_1 _31103_ (.A(_05377_),
    .B(_05380_),
    .Y(_05381_));
 sg13g2_or2_1 _31104_ (.X(_05382_),
    .B(\u_inv.d_reg[69] ),
    .A(\u_inv.d_next[69] ));
 sg13g2_and2_1 _31105_ (.A(\u_inv.d_next[69] ),
    .B(\u_inv.d_reg[69] ),
    .X(_05383_));
 sg13g2_xor2_1 _31106_ (.B(\u_inv.d_reg[69] ),
    .A(\u_inv.d_next[69] ),
    .X(_05384_));
 sg13g2_xnor2_1 _31107_ (.Y(_05385_),
    .A(\u_inv.d_next[69] ),
    .B(\u_inv.d_reg[69] ));
 sg13g2_and2_1 _31108_ (.A(\u_inv.d_next[68] ),
    .B(\u_inv.d_reg[68] ),
    .X(_05386_));
 sg13g2_xor2_1 _31109_ (.B(\u_inv.d_reg[68] ),
    .A(\u_inv.d_next[68] ),
    .X(_05387_));
 sg13g2_xnor2_1 _31110_ (.Y(_05388_),
    .A(\u_inv.d_next[68] ),
    .B(\u_inv.d_reg[68] ));
 sg13g2_nor2_1 _31111_ (.A(_05384_),
    .B(_05387_),
    .Y(_05389_));
 sg13g2_and2_1 _31112_ (.A(_05381_),
    .B(_05389_),
    .X(_05390_));
 sg13g2_nor2_1 _31113_ (.A(\u_inv.d_next[67] ),
    .B(_14742_),
    .Y(_05391_));
 sg13g2_nand2_1 _31114_ (.Y(_05392_),
    .A(\u_inv.d_next[67] ),
    .B(_14742_));
 sg13g2_xnor2_1 _31115_ (.Y(_05393_),
    .A(\u_inv.d_next[67] ),
    .B(\u_inv.d_reg[67] ));
 sg13g2_xor2_1 _31116_ (.B(\u_inv.d_reg[67] ),
    .A(\u_inv.d_next[67] ),
    .X(_05394_));
 sg13g2_xor2_1 _31117_ (.B(\u_inv.d_reg[66] ),
    .A(net5880),
    .X(_05395_));
 sg13g2_xnor2_1 _31118_ (.Y(_05396_),
    .A(net5880),
    .B(\u_inv.d_reg[66] ));
 sg13g2_nand2_1 _31119_ (.Y(_05397_),
    .A(_05393_),
    .B(_05396_));
 sg13g2_nor2b_1 _31120_ (.A(\u_inv.d_reg[65] ),
    .B_N(\u_inv.d_next[65] ),
    .Y(_05398_));
 sg13g2_nand2b_1 _31121_ (.Y(_05399_),
    .B(\u_inv.d_reg[65] ),
    .A_N(\u_inv.d_next[65] ));
 sg13g2_xor2_1 _31122_ (.B(\u_inv.d_reg[65] ),
    .A(\u_inv.d_next[65] ),
    .X(_05400_));
 sg13g2_and2_1 _31123_ (.A(\u_inv.d_next[64] ),
    .B(\u_inv.d_reg[64] ),
    .X(_05401_));
 sg13g2_xor2_1 _31124_ (.B(\u_inv.d_reg[64] ),
    .A(\u_inv.d_next[64] ),
    .X(_05402_));
 sg13g2_xnor2_1 _31125_ (.Y(_05403_),
    .A(\u_inv.d_next[64] ),
    .B(\u_inv.d_reg[64] ));
 sg13g2_nor2_1 _31126_ (.A(_05400_),
    .B(_05402_),
    .Y(_05404_));
 sg13g2_and4_1 _31127_ (.A(_05390_),
    .B(_05393_),
    .C(_05396_),
    .D(_05404_),
    .X(_05405_));
 sg13g2_nand2_2 _31128_ (.Y(_05406_),
    .A(_05375_),
    .B(_05405_));
 sg13g2_xor2_1 _31129_ (.B(\u_inv.d_reg[125] ),
    .A(\u_inv.d_next[125] ),
    .X(_05407_));
 sg13g2_xnor2_1 _31130_ (.Y(_05408_),
    .A(\u_inv.d_next[125] ),
    .B(\u_inv.d_reg[125] ));
 sg13g2_nand2_1 _31131_ (.Y(_05409_),
    .A(\u_inv.d_next[124] ),
    .B(\u_inv.d_reg[124] ));
 sg13g2_xor2_1 _31132_ (.B(\u_inv.d_reg[124] ),
    .A(\u_inv.d_next[124] ),
    .X(_05410_));
 sg13g2_xnor2_1 _31133_ (.Y(_05411_),
    .A(\u_inv.d_next[124] ),
    .B(\u_inv.d_reg[124] ));
 sg13g2_nand2_1 _31134_ (.Y(_05412_),
    .A(_05408_),
    .B(_05411_));
 sg13g2_inv_1 _31135_ (.Y(_05413_),
    .A(_05412_));
 sg13g2_nor2_1 _31136_ (.A(\u_inv.d_next[127] ),
    .B(\u_inv.d_reg[127] ),
    .Y(_05414_));
 sg13g2_nand2_1 _31137_ (.Y(_05415_),
    .A(\u_inv.d_next[127] ),
    .B(\u_inv.d_reg[127] ));
 sg13g2_nand2b_2 _31138_ (.Y(_05416_),
    .B(_05415_),
    .A_N(_05414_));
 sg13g2_nand2_1 _31139_ (.Y(_05417_),
    .A(\u_inv.d_next[126] ),
    .B(\u_inv.d_reg[126] ));
 sg13g2_inv_1 _31140_ (.Y(_05418_),
    .A(_05417_));
 sg13g2_xor2_1 _31141_ (.B(\u_inv.d_reg[126] ),
    .A(\u_inv.d_next[126] ),
    .X(_05419_));
 sg13g2_xnor2_1 _31142_ (.Y(_05420_),
    .A(\u_inv.d_next[126] ),
    .B(\u_inv.d_reg[126] ));
 sg13g2_nand2_1 _31143_ (.Y(_05421_),
    .A(_05416_),
    .B(_05420_));
 sg13g2_nor2_1 _31144_ (.A(_05412_),
    .B(_05421_),
    .Y(_05422_));
 sg13g2_nor2_1 _31145_ (.A(\u_inv.d_next[123] ),
    .B(\u_inv.d_reg[123] ),
    .Y(_05423_));
 sg13g2_xnor2_1 _31146_ (.Y(_05424_),
    .A(\u_inv.d_next[123] ),
    .B(\u_inv.d_reg[123] ));
 sg13g2_inv_1 _31147_ (.Y(_05425_),
    .A(_05424_));
 sg13g2_nand2_1 _31148_ (.Y(_05426_),
    .A(\u_inv.d_next[122] ),
    .B(\u_inv.d_reg[122] ));
 sg13g2_xnor2_1 _31149_ (.Y(_05427_),
    .A(\u_inv.d_next[122] ),
    .B(\u_inv.d_reg[122] ));
 sg13g2_nand2_1 _31150_ (.Y(_05428_),
    .A(_05424_),
    .B(_05427_));
 sg13g2_nand2_1 _31151_ (.Y(_05429_),
    .A(\u_inv.d_next[121] ),
    .B(_14688_));
 sg13g2_nor2_1 _31152_ (.A(\u_inv.d_next[121] ),
    .B(_14688_),
    .Y(_05430_));
 sg13g2_xnor2_1 _31153_ (.Y(_05431_),
    .A(\u_inv.d_next[121] ),
    .B(\u_inv.d_reg[121] ));
 sg13g2_xor2_1 _31154_ (.B(\u_inv.d_reg[121] ),
    .A(\u_inv.d_next[121] ),
    .X(_05432_));
 sg13g2_nand2_1 _31155_ (.Y(_05433_),
    .A(\u_inv.d_next[120] ),
    .B(\u_inv.d_reg[120] ));
 sg13g2_xor2_1 _31156_ (.B(\u_inv.d_reg[120] ),
    .A(\u_inv.d_next[120] ),
    .X(_05434_));
 sg13g2_xnor2_1 _31157_ (.Y(_05435_),
    .A(\u_inv.d_next[120] ),
    .B(\u_inv.d_reg[120] ));
 sg13g2_nand2_1 _31158_ (.Y(_05436_),
    .A(_05431_),
    .B(_05435_));
 sg13g2_nor4_1 _31159_ (.A(_05412_),
    .B(_05421_),
    .C(_05428_),
    .D(_05436_),
    .Y(_05437_));
 sg13g2_xnor2_1 _31160_ (.Y(_05438_),
    .A(\u_inv.d_next[117] ),
    .B(\u_inv.d_reg[117] ));
 sg13g2_xor2_1 _31161_ (.B(\u_inv.d_reg[117] ),
    .A(\u_inv.d_next[117] ),
    .X(_05439_));
 sg13g2_xnor2_1 _31162_ (.Y(_05440_),
    .A(\u_inv.d_next[116] ),
    .B(\u_inv.d_reg[116] ));
 sg13g2_and2_1 _31163_ (.A(_05438_),
    .B(_05440_),
    .X(_05441_));
 sg13g2_nand2_1 _31164_ (.Y(_05442_),
    .A(\u_inv.d_next[118] ),
    .B(\u_inv.d_reg[118] ));
 sg13g2_xor2_1 _31165_ (.B(\u_inv.d_reg[118] ),
    .A(\u_inv.d_next[118] ),
    .X(_05443_));
 sg13g2_nand2_1 _31166_ (.Y(_05444_),
    .A(\u_inv.d_next[119] ),
    .B(\u_inv.d_reg[119] ));
 sg13g2_nor2_1 _31167_ (.A(\u_inv.d_next[119] ),
    .B(\u_inv.d_reg[119] ),
    .Y(_05445_));
 sg13g2_xnor2_1 _31168_ (.Y(_05446_),
    .A(\u_inv.d_next[119] ),
    .B(\u_inv.d_reg[119] ));
 sg13g2_nand2_1 _31169_ (.Y(_05447_),
    .A(_05441_),
    .B(_05446_));
 sg13g2_nor2_1 _31170_ (.A(_05443_),
    .B(_05447_),
    .Y(_05448_));
 sg13g2_xnor2_1 _31171_ (.Y(_05449_),
    .A(\u_inv.d_next[115] ),
    .B(\u_inv.d_reg[115] ));
 sg13g2_xnor2_1 _31172_ (.Y(_05450_),
    .A(\u_inv.d_next[114] ),
    .B(\u_inv.d_reg[114] ));
 sg13g2_nand2_1 _31173_ (.Y(_05451_),
    .A(_05449_),
    .B(_05450_));
 sg13g2_nor2b_1 _31174_ (.A(\u_inv.d_reg[113] ),
    .B_N(\u_inv.d_next[113] ),
    .Y(_05452_));
 sg13g2_nand2b_1 _31175_ (.Y(_05453_),
    .B(\u_inv.d_reg[113] ),
    .A_N(\u_inv.d_next[113] ));
 sg13g2_nor2b_2 _31176_ (.A(_05452_),
    .B_N(_05453_),
    .Y(_05454_));
 sg13g2_xor2_1 _31177_ (.B(\u_inv.d_reg[113] ),
    .A(\u_inv.d_next[113] ),
    .X(_05455_));
 sg13g2_and2_1 _31178_ (.A(\u_inv.d_next[112] ),
    .B(\u_inv.d_reg[112] ),
    .X(_05456_));
 sg13g2_xnor2_1 _31179_ (.Y(_05457_),
    .A(\u_inv.d_next[112] ),
    .B(\u_inv.d_reg[112] ));
 sg13g2_nand2_1 _31180_ (.Y(_05458_),
    .A(_05454_),
    .B(_05457_));
 sg13g2_nor4_1 _31181_ (.A(_05443_),
    .B(_05447_),
    .C(_05451_),
    .D(_05458_),
    .Y(_05459_));
 sg13g2_and2_1 _31182_ (.A(_05437_),
    .B(_05459_),
    .X(_05460_));
 sg13g2_nand2_1 _31183_ (.Y(_05461_),
    .A(\u_inv.d_next[111] ),
    .B(\u_inv.d_reg[111] ));
 sg13g2_xor2_1 _31184_ (.B(\u_inv.d_reg[111] ),
    .A(\u_inv.d_next[111] ),
    .X(_05462_));
 sg13g2_xnor2_1 _31185_ (.Y(_05463_),
    .A(\u_inv.d_next[111] ),
    .B(\u_inv.d_reg[111] ));
 sg13g2_and2_1 _31186_ (.A(\u_inv.d_next[110] ),
    .B(\u_inv.d_reg[110] ),
    .X(_05464_));
 sg13g2_xnor2_1 _31187_ (.Y(_05465_),
    .A(\u_inv.d_next[110] ),
    .B(\u_inv.d_reg[110] ));
 sg13g2_nand2_1 _31188_ (.Y(_05466_),
    .A(_05463_),
    .B(_05465_));
 sg13g2_nor2b_1 _31189_ (.A(\u_inv.d_reg[109] ),
    .B_N(\u_inv.d_next[109] ),
    .Y(_05467_));
 sg13g2_nand2b_1 _31190_ (.Y(_05468_),
    .B(\u_inv.d_reg[109] ),
    .A_N(\u_inv.d_next[109] ));
 sg13g2_nand2b_2 _31191_ (.Y(_05469_),
    .B(_05468_),
    .A_N(_05467_));
 sg13g2_xor2_1 _31192_ (.B(\u_inv.d_reg[108] ),
    .A(\u_inv.d_next[108] ),
    .X(_05470_));
 sg13g2_or2_1 _31193_ (.X(_05471_),
    .B(_05470_),
    .A(_05469_));
 sg13g2_or2_1 _31194_ (.X(_05472_),
    .B(_05471_),
    .A(_05466_));
 sg13g2_nor2_1 _31195_ (.A(\u_inv.d_next[107] ),
    .B(_14702_),
    .Y(_05473_));
 sg13g2_xnor2_1 _31196_ (.Y(_05474_),
    .A(\u_inv.d_next[107] ),
    .B(\u_inv.d_reg[107] ));
 sg13g2_xor2_1 _31197_ (.B(\u_inv.d_reg[107] ),
    .A(\u_inv.d_next[107] ),
    .X(_05475_));
 sg13g2_nand2_1 _31198_ (.Y(_05476_),
    .A(\u_inv.d_next[106] ),
    .B(\u_inv.d_reg[106] ));
 sg13g2_xor2_1 _31199_ (.B(\u_inv.d_reg[106] ),
    .A(\u_inv.d_next[106] ),
    .X(_05477_));
 sg13g2_xnor2_1 _31200_ (.Y(_05478_),
    .A(\u_inv.d_next[106] ),
    .B(\u_inv.d_reg[106] ));
 sg13g2_nor2_1 _31201_ (.A(_05475_),
    .B(_05477_),
    .Y(_05479_));
 sg13g2_xor2_1 _31202_ (.B(\u_inv.d_reg[105] ),
    .A(\u_inv.d_next[105] ),
    .X(_05480_));
 sg13g2_and2_1 _31203_ (.A(\u_inv.d_next[104] ),
    .B(\u_inv.d_reg[104] ),
    .X(_05481_));
 sg13g2_xnor2_1 _31204_ (.Y(_05482_),
    .A(\u_inv.d_next[104] ),
    .B(\u_inv.d_reg[104] ));
 sg13g2_nor2b_1 _31205_ (.A(_05480_),
    .B_N(_05482_),
    .Y(_05483_));
 sg13g2_and2_1 _31206_ (.A(_05479_),
    .B(_05483_),
    .X(_05484_));
 sg13g2_nand2b_1 _31207_ (.Y(_05485_),
    .B(_05484_),
    .A_N(_05472_));
 sg13g2_nor2_1 _31208_ (.A(_14218_),
    .B(\u_inv.d_reg[103] ),
    .Y(_05486_));
 sg13g2_xnor2_1 _31209_ (.Y(_05487_),
    .A(\u_inv.d_next[103] ),
    .B(\u_inv.d_reg[103] ));
 sg13g2_nand2_1 _31210_ (.Y(_05488_),
    .A(\u_inv.d_next[102] ),
    .B(\u_inv.d_reg[102] ));
 sg13g2_xnor2_1 _31211_ (.Y(_05489_),
    .A(\u_inv.d_next[102] ),
    .B(\u_inv.d_reg[102] ));
 sg13g2_nand2_1 _31212_ (.Y(_05490_),
    .A(_05487_),
    .B(_05489_));
 sg13g2_xor2_1 _31213_ (.B(\u_inv.d_reg[101] ),
    .A(\u_inv.d_next[101] ),
    .X(_05491_));
 sg13g2_xor2_1 _31214_ (.B(\u_inv.d_reg[100] ),
    .A(\u_inv.d_next[100] ),
    .X(_05492_));
 sg13g2_or2_1 _31215_ (.X(_05493_),
    .B(_05492_),
    .A(_05491_));
 sg13g2_or2_1 _31216_ (.X(_05494_),
    .B(_05493_),
    .A(_05490_));
 sg13g2_nor2b_1 _31217_ (.A(\u_inv.d_reg[99] ),
    .B_N(\u_inv.d_next[99] ),
    .Y(_05495_));
 sg13g2_nand2b_1 _31218_ (.Y(_05496_),
    .B(\u_inv.d_reg[99] ),
    .A_N(\u_inv.d_next[99] ));
 sg13g2_nor2b_2 _31219_ (.A(_05495_),
    .B_N(_05496_),
    .Y(_05497_));
 sg13g2_xor2_1 _31220_ (.B(\u_inv.d_reg[99] ),
    .A(\u_inv.d_next[99] ),
    .X(_05498_));
 sg13g2_nand2_1 _31221_ (.Y(_05499_),
    .A(\u_inv.d_next[98] ),
    .B(net5870));
 sg13g2_xnor2_1 _31222_ (.Y(_05500_),
    .A(\u_inv.d_next[98] ),
    .B(net5870));
 sg13g2_nor2b_1 _31223_ (.A(_05498_),
    .B_N(_05500_),
    .Y(_05501_));
 sg13g2_nand2_1 _31224_ (.Y(_05502_),
    .A(\u_inv.d_next[97] ),
    .B(_14712_));
 sg13g2_nor2_1 _31225_ (.A(\u_inv.d_next[97] ),
    .B(_14712_),
    .Y(_05503_));
 sg13g2_xnor2_1 _31226_ (.Y(_05504_),
    .A(\u_inv.d_next[97] ),
    .B(\u_inv.d_reg[97] ));
 sg13g2_xor2_1 _31227_ (.B(\u_inv.d_reg[97] ),
    .A(\u_inv.d_next[97] ),
    .X(_05505_));
 sg13g2_and2_1 _31228_ (.A(\u_inv.d_next[96] ),
    .B(\u_inv.d_reg[96] ),
    .X(_05506_));
 sg13g2_xor2_1 _31229_ (.B(\u_inv.d_reg[96] ),
    .A(\u_inv.d_next[96] ),
    .X(_05507_));
 sg13g2_xnor2_1 _31230_ (.Y(_05508_),
    .A(\u_inv.d_next[96] ),
    .B(\u_inv.d_reg[96] ));
 sg13g2_nor2_1 _31231_ (.A(_05505_),
    .B(_05507_),
    .Y(_05509_));
 sg13g2_and2_1 _31232_ (.A(_05501_),
    .B(_05509_),
    .X(_05510_));
 sg13g2_nand2b_2 _31233_ (.Y(_05511_),
    .B(_05510_),
    .A_N(_05494_));
 sg13g2_nor2_1 _31234_ (.A(_05485_),
    .B(_05511_),
    .Y(_05512_));
 sg13g2_and2_1 _31235_ (.A(_05460_),
    .B(_05512_),
    .X(_05513_));
 sg13g2_nor2_1 _31236_ (.A(\u_inv.d_next[95] ),
    .B(\u_inv.d_reg[95] ),
    .Y(_05514_));
 sg13g2_xnor2_1 _31237_ (.Y(_05515_),
    .A(\u_inv.d_next[95] ),
    .B(\u_inv.d_reg[95] ));
 sg13g2_nand2_1 _31238_ (.Y(_05516_),
    .A(\u_inv.d_next[94] ),
    .B(\u_inv.d_reg[94] ));
 sg13g2_xnor2_1 _31239_ (.Y(_05517_),
    .A(\u_inv.d_next[94] ),
    .B(\u_inv.d_reg[94] ));
 sg13g2_nand2_1 _31240_ (.Y(_05518_),
    .A(_05515_),
    .B(_05517_));
 sg13g2_xnor2_1 _31241_ (.Y(_05519_),
    .A(\u_inv.d_next[93] ),
    .B(\u_inv.d_reg[93] ));
 sg13g2_xor2_1 _31242_ (.B(\u_inv.d_reg[93] ),
    .A(\u_inv.d_next[93] ),
    .X(_05520_));
 sg13g2_nand2_1 _31243_ (.Y(_05521_),
    .A(\u_inv.d_next[92] ),
    .B(\u_inv.d_reg[92] ));
 sg13g2_xor2_1 _31244_ (.B(\u_inv.d_reg[92] ),
    .A(\u_inv.d_next[92] ),
    .X(_05522_));
 sg13g2_nand2b_1 _31245_ (.Y(_05523_),
    .B(_05519_),
    .A_N(_05522_));
 sg13g2_nor2_1 _31246_ (.A(_05518_),
    .B(_05523_),
    .Y(_05524_));
 sg13g2_nor2_1 _31247_ (.A(\u_inv.d_next[91] ),
    .B(_14718_),
    .Y(_05525_));
 sg13g2_xnor2_1 _31248_ (.Y(_05526_),
    .A(\u_inv.d_next[91] ),
    .B(\u_inv.d_reg[91] ));
 sg13g2_inv_1 _31249_ (.Y(_05527_),
    .A(_05526_));
 sg13g2_nand2_1 _31250_ (.Y(_05528_),
    .A(\u_inv.d_next[90] ),
    .B(net5871));
 sg13g2_xnor2_1 _31251_ (.Y(_05529_),
    .A(\u_inv.d_next[90] ),
    .B(net5871));
 sg13g2_and2_1 _31252_ (.A(_05526_),
    .B(_05529_),
    .X(_05530_));
 sg13g2_xnor2_1 _31253_ (.Y(_05531_),
    .A(\u_inv.d_next[89] ),
    .B(\u_inv.d_reg[89] ));
 sg13g2_nand2_1 _31254_ (.Y(_05532_),
    .A(\u_inv.d_next[88] ),
    .B(\u_inv.d_reg[88] ));
 sg13g2_xor2_1 _31255_ (.B(\u_inv.d_reg[88] ),
    .A(\u_inv.d_next[88] ),
    .X(_05533_));
 sg13g2_xnor2_1 _31256_ (.Y(_05534_),
    .A(\u_inv.d_next[88] ),
    .B(\u_inv.d_reg[88] ));
 sg13g2_and2_1 _31257_ (.A(_05531_),
    .B(_05534_),
    .X(_05535_));
 sg13g2_inv_1 _31258_ (.Y(_05536_),
    .A(_05535_));
 sg13g2_nand3_1 _31259_ (.B(_05530_),
    .C(_05535_),
    .A(_05524_),
    .Y(_05537_));
 sg13g2_nor2b_1 _31260_ (.A(\u_inv.d_reg[87] ),
    .B_N(\u_inv.d_next[87] ),
    .Y(_05538_));
 sg13g2_nand2b_1 _31261_ (.Y(_05539_),
    .B(\u_inv.d_reg[87] ),
    .A_N(\u_inv.d_next[87] ));
 sg13g2_nor2b_1 _31262_ (.A(_05538_),
    .B_N(_05539_),
    .Y(_05540_));
 sg13g2_nand2b_2 _31263_ (.Y(_05541_),
    .B(_05539_),
    .A_N(_05538_));
 sg13g2_and2_1 _31264_ (.A(\u_inv.d_next[86] ),
    .B(\u_inv.d_reg[86] ),
    .X(_05542_));
 sg13g2_xor2_1 _31265_ (.B(\u_inv.d_reg[86] ),
    .A(\u_inv.d_next[86] ),
    .X(_05543_));
 sg13g2_inv_1 _31266_ (.Y(_05544_),
    .A(_05543_));
 sg13g2_nor2_1 _31267_ (.A(_05541_),
    .B(_05543_),
    .Y(_05545_));
 sg13g2_xor2_1 _31268_ (.B(\u_inv.d_reg[85] ),
    .A(\u_inv.d_next[85] ),
    .X(_05546_));
 sg13g2_xor2_1 _31269_ (.B(\u_inv.d_reg[84] ),
    .A(\u_inv.d_next[84] ),
    .X(_05547_));
 sg13g2_xnor2_1 _31270_ (.Y(_05548_),
    .A(\u_inv.d_next[84] ),
    .B(\u_inv.d_reg[84] ));
 sg13g2_nor2_1 _31271_ (.A(_05546_),
    .B(_05547_),
    .Y(_05549_));
 sg13g2_nand2_1 _31272_ (.Y(_05550_),
    .A(_05545_),
    .B(_05549_));
 sg13g2_xnor2_1 _31273_ (.Y(_05551_),
    .A(\u_inv.d_next[83] ),
    .B(\u_inv.d_reg[83] ));
 sg13g2_nor2_1 _31274_ (.A(\u_inv.d_next[82] ),
    .B(\u_inv.d_reg[82] ),
    .Y(_05552_));
 sg13g2_nand2_1 _31275_ (.Y(_05553_),
    .A(\u_inv.d_next[82] ),
    .B(\u_inv.d_reg[82] ));
 sg13g2_nand2b_2 _31276_ (.Y(_05554_),
    .B(_05553_),
    .A_N(_05552_));
 sg13g2_and2_1 _31277_ (.A(_05551_),
    .B(_05554_),
    .X(_05555_));
 sg13g2_nor2b_1 _31278_ (.A(\u_inv.d_reg[81] ),
    .B_N(\u_inv.d_next[81] ),
    .Y(_05556_));
 sg13g2_nand2_1 _31279_ (.Y(_05557_),
    .A(\u_inv.d_next[81] ),
    .B(_14728_));
 sg13g2_nand2b_1 _31280_ (.Y(_05558_),
    .B(\u_inv.d_reg[81] ),
    .A_N(\u_inv.d_next[81] ));
 sg13g2_xor2_1 _31281_ (.B(\u_inv.d_reg[81] ),
    .A(\u_inv.d_next[81] ),
    .X(_05559_));
 sg13g2_and2_1 _31282_ (.A(\u_inv.d_next[80] ),
    .B(\u_inv.d_reg[80] ),
    .X(_05560_));
 sg13g2_xor2_1 _31283_ (.B(\u_inv.d_reg[80] ),
    .A(\u_inv.d_next[80] ),
    .X(_05561_));
 sg13g2_xnor2_1 _31284_ (.Y(_05562_),
    .A(\u_inv.d_next[80] ),
    .B(\u_inv.d_reg[80] ));
 sg13g2_nand2b_1 _31285_ (.Y(_05563_),
    .B(_05562_),
    .A_N(_05559_));
 sg13g2_nand4_1 _31286_ (.B(_05557_),
    .C(_05558_),
    .A(_05555_),
    .Y(_05564_),
    .D(_05562_));
 sg13g2_or2_1 _31287_ (.X(_05565_),
    .B(_05564_),
    .A(_05550_));
 sg13g2_nor2_2 _31288_ (.A(_05537_),
    .B(_05565_),
    .Y(_05566_));
 sg13g2_nor2b_2 _31289_ (.A(_05406_),
    .B_N(_05566_),
    .Y(_05567_));
 sg13g2_and2_1 _31290_ (.A(_05513_),
    .B(_05567_),
    .X(_05568_));
 sg13g2_o21ai_1 _31291_ (.B1(_05568_),
    .Y(_05569_),
    .A1(_05314_),
    .A2(_05347_));
 sg13g2_nand2_1 _31292_ (.Y(_05570_),
    .A(\u_inv.d_next[123] ),
    .B(_14686_));
 sg13g2_nor2b_1 _31293_ (.A(\u_inv.d_reg[122] ),
    .B_N(\u_inv.d_next[122] ),
    .Y(_05571_));
 sg13g2_nand2_1 _31294_ (.Y(_05572_),
    .A(\u_inv.d_next[120] ),
    .B(_14689_));
 sg13g2_o21ai_1 _31295_ (.B1(_05429_),
    .Y(_05573_),
    .A1(_05430_),
    .A2(_05572_));
 sg13g2_inv_1 _31296_ (.Y(_05574_),
    .A(_05573_));
 sg13g2_a21oi_1 _31297_ (.A1(_05427_),
    .A2(_05573_),
    .Y(_05575_),
    .B1(_05571_));
 sg13g2_o21ai_1 _31298_ (.B1(_05570_),
    .Y(_05576_),
    .A1(_05425_),
    .A2(_05575_));
 sg13g2_nor2b_1 _31299_ (.A(\u_inv.d_reg[127] ),
    .B_N(\u_inv.d_next[127] ),
    .Y(_05577_));
 sg13g2_nand2_1 _31300_ (.Y(_05578_),
    .A(\u_inv.d_next[126] ),
    .B(_14683_));
 sg13g2_nand2_1 _31301_ (.Y(_05579_),
    .A(\u_inv.d_next[124] ),
    .B(_14685_));
 sg13g2_nor2_1 _31302_ (.A(_05407_),
    .B(_05579_),
    .Y(_05580_));
 sg13g2_a21oi_1 _31303_ (.A1(\u_inv.d_next[125] ),
    .A2(_14684_),
    .Y(_05581_),
    .B1(_05580_));
 sg13g2_o21ai_1 _31304_ (.B1(_05578_),
    .Y(_05582_),
    .A1(_05419_),
    .A2(_05581_));
 sg13g2_a21oi_1 _31305_ (.A1(_05416_),
    .A2(_05582_),
    .Y(_05583_),
    .B1(_05577_));
 sg13g2_nor2b_1 _31306_ (.A(\u_inv.d_reg[112] ),
    .B_N(\u_inv.d_next[112] ),
    .Y(_05584_));
 sg13g2_a21oi_1 _31307_ (.A1(_05453_),
    .A2(_05584_),
    .Y(_05585_),
    .B1(_05452_));
 sg13g2_nor2_1 _31308_ (.A(_05451_),
    .B(_05585_),
    .Y(_05586_));
 sg13g2_nor2_1 _31309_ (.A(_14216_),
    .B(\u_inv.d_reg[114] ),
    .Y(_05587_));
 sg13g2_o21ai_1 _31310_ (.B1(_05587_),
    .Y(_05588_),
    .A1(\u_inv.d_next[115] ),
    .A2(_14694_));
 sg13g2_a21oi_1 _31311_ (.A1(\u_inv.d_next[115] ),
    .A2(_14694_),
    .Y(_05589_),
    .B1(_05586_));
 sg13g2_nand2_1 _31312_ (.Y(_05590_),
    .A(_05588_),
    .B(_05589_));
 sg13g2_nor2b_1 _31313_ (.A(\u_inv.d_reg[116] ),
    .B_N(\u_inv.d_next[116] ),
    .Y(_05591_));
 sg13g2_a21oi_1 _31314_ (.A1(\u_inv.d_next[117] ),
    .A2(_14692_),
    .Y(_05592_),
    .B1(_05591_));
 sg13g2_a21o_1 _31315_ (.A2(\u_inv.d_reg[117] ),
    .A1(_14215_),
    .B1(_05592_),
    .X(_05593_));
 sg13g2_nand2_1 _31316_ (.Y(_05594_),
    .A(\u_inv.d_next[118] ),
    .B(_14691_));
 sg13g2_o21ai_1 _31317_ (.B1(_05594_),
    .Y(_05595_),
    .A1(_05443_),
    .A2(_05593_));
 sg13g2_a22oi_1 _31318_ (.Y(_05596_),
    .B1(_05595_),
    .B2(_05446_),
    .A2(_05590_),
    .A1(_05448_));
 sg13g2_o21ai_1 _31319_ (.B1(_05596_),
    .Y(_05597_),
    .A1(_14214_),
    .A2(\u_inv.d_reg[119] ));
 sg13g2_a22oi_1 _31320_ (.Y(_05598_),
    .B1(_05597_),
    .B2(_05437_),
    .A2(_05576_),
    .A1(_05422_));
 sg13g2_nor2b_1 _31321_ (.A(\u_inv.d_reg[80] ),
    .B_N(\u_inv.d_next[80] ),
    .Y(_05599_));
 sg13g2_a21oi_1 _31322_ (.A1(_05558_),
    .A2(_05599_),
    .Y(_05600_),
    .B1(_05556_));
 sg13g2_inv_1 _31323_ (.Y(_05601_),
    .A(_05600_));
 sg13g2_nand2_1 _31324_ (.Y(_05602_),
    .A(\u_inv.d_next[82] ),
    .B(_14727_));
 sg13g2_a21oi_1 _31325_ (.A1(_14223_),
    .A2(\u_inv.d_reg[83] ),
    .Y(_05603_),
    .B1(_05602_));
 sg13g2_a221oi_1 _31326_ (.B2(_05601_),
    .C1(_05603_),
    .B1(_05555_),
    .A1(\u_inv.d_next[83] ),
    .Y(_05604_),
    .A2(_14726_));
 sg13g2_inv_1 _31327_ (.Y(_05605_),
    .A(_05604_));
 sg13g2_nor2b_2 _31328_ (.A(\u_inv.d_reg[86] ),
    .B_N(\u_inv.d_next[86] ),
    .Y(_05606_));
 sg13g2_a21oi_1 _31329_ (.A1(_05539_),
    .A2(_05606_),
    .Y(_05607_),
    .B1(_05538_));
 sg13g2_nand2_1 _31330_ (.Y(_05608_),
    .A(\u_inv.d_next[85] ),
    .B(_14724_));
 sg13g2_nor2b_1 _31331_ (.A(\u_inv.d_reg[84] ),
    .B_N(\u_inv.d_next[84] ),
    .Y(_05609_));
 sg13g2_nand2b_1 _31332_ (.Y(_05610_),
    .B(_05609_),
    .A_N(_05546_));
 sg13g2_and2_1 _31333_ (.A(_05608_),
    .B(_05610_),
    .X(_05611_));
 sg13g2_nand2_1 _31334_ (.Y(_05612_),
    .A(_05608_),
    .B(_05610_));
 sg13g2_o21ai_1 _31335_ (.B1(_05607_),
    .Y(_05613_),
    .A1(_05550_),
    .A2(_05604_));
 sg13g2_a21oi_2 _31336_ (.B1(_05613_),
    .Y(_05614_),
    .A2(_05612_),
    .A1(_05545_));
 sg13g2_a22oi_1 _31337_ (.Y(_05615_),
    .B1(_14721_),
    .B2(\u_inv.d_next[88] ),
    .A2(_14720_),
    .A1(\u_inv.d_next[89] ));
 sg13g2_a21oi_1 _31338_ (.A1(_14221_),
    .A2(\u_inv.d_reg[89] ),
    .Y(_05616_),
    .B1(_05615_));
 sg13g2_nor2_1 _31339_ (.A(_14220_),
    .B(net5871),
    .Y(_05617_));
 sg13g2_nor3_1 _31340_ (.A(_14220_),
    .B(net5871),
    .C(_05525_),
    .Y(_05618_));
 sg13g2_a221oi_1 _31341_ (.B2(_05616_),
    .C1(_05618_),
    .B1(_05530_),
    .A1(\u_inv.d_next[91] ),
    .Y(_05619_),
    .A2(_14718_));
 sg13g2_inv_1 _31342_ (.Y(_05620_),
    .A(_05619_));
 sg13g2_nor2b_1 _31343_ (.A(\u_inv.d_reg[94] ),
    .B_N(\u_inv.d_next[94] ),
    .Y(_05621_));
 sg13g2_nand2_1 _31344_ (.Y(_05622_),
    .A(_05515_),
    .B(_05621_));
 sg13g2_nand2_1 _31345_ (.Y(_05623_),
    .A(\u_inv.d_next[92] ),
    .B(_14717_));
 sg13g2_o21ai_1 _31346_ (.B1(_05623_),
    .Y(_05624_),
    .A1(_14219_),
    .A2(\u_inv.d_reg[93] ));
 sg13g2_o21ai_1 _31347_ (.B1(_05624_),
    .Y(_05625_),
    .A1(\u_inv.d_next[93] ),
    .A2(_14716_));
 sg13g2_nor2_1 _31348_ (.A(_05518_),
    .B(_05625_),
    .Y(_05626_));
 sg13g2_nand2_1 _31349_ (.Y(_05627_),
    .A(\u_inv.d_next[96] ),
    .B(_14713_));
 sg13g2_o21ai_1 _31350_ (.B1(_05502_),
    .Y(_05628_),
    .A1(_05503_),
    .A2(_05627_));
 sg13g2_nor2b_1 _31351_ (.A(net5870),
    .B_N(\u_inv.d_next[98] ),
    .Y(_05629_));
 sg13g2_a221oi_1 _31352_ (.B2(_05496_),
    .C1(_05495_),
    .B1(_05629_),
    .A1(_05501_),
    .Y(_05630_),
    .A2(_05628_));
 sg13g2_inv_1 _31353_ (.Y(_05631_),
    .A(_05630_));
 sg13g2_nor2_1 _31354_ (.A(_05494_),
    .B(_05630_),
    .Y(_05632_));
 sg13g2_nand2_1 _31355_ (.Y(_05633_),
    .A(\u_inv.d_next[102] ),
    .B(_14707_));
 sg13g2_a21oi_1 _31356_ (.A1(_14218_),
    .A2(\u_inv.d_reg[103] ),
    .Y(_05634_),
    .B1(_05633_));
 sg13g2_nand2_1 _31357_ (.Y(_05635_),
    .A(\u_inv.d_next[100] ),
    .B(_14709_));
 sg13g2_nor2_1 _31358_ (.A(_05491_),
    .B(_05635_),
    .Y(_05636_));
 sg13g2_a21oi_1 _31359_ (.A1(\u_inv.d_next[101] ),
    .A2(_14708_),
    .Y(_05637_),
    .B1(_05636_));
 sg13g2_nor2_1 _31360_ (.A(_05490_),
    .B(_05637_),
    .Y(_05638_));
 sg13g2_nor4_1 _31361_ (.A(_05486_),
    .B(_05632_),
    .C(_05634_),
    .D(_05638_),
    .Y(_05639_));
 sg13g2_nor2_1 _31362_ (.A(_05485_),
    .B(_05639_),
    .Y(_05640_));
 sg13g2_nor2b_1 _31363_ (.A(\u_inv.d_reg[104] ),
    .B_N(\u_inv.d_next[104] ),
    .Y(_05641_));
 sg13g2_a21oi_1 _31364_ (.A1(\u_inv.d_next[105] ),
    .A2(_14704_),
    .Y(_05642_),
    .B1(_05641_));
 sg13g2_a21oi_1 _31365_ (.A1(_14217_),
    .A2(\u_inv.d_reg[105] ),
    .Y(_05643_),
    .B1(_05642_));
 sg13g2_nand2_1 _31366_ (.Y(_05644_),
    .A(\u_inv.d_next[106] ),
    .B(_14703_));
 sg13g2_a22oi_1 _31367_ (.Y(_05645_),
    .B1(_05479_),
    .B2(_05643_),
    .A2(_14702_),
    .A1(\u_inv.d_next[107] ));
 sg13g2_o21ai_1 _31368_ (.B1(_05645_),
    .Y(_05646_),
    .A1(_05473_),
    .A2(_05644_));
 sg13g2_nor2b_1 _31369_ (.A(_05472_),
    .B_N(_05646_),
    .Y(_05647_));
 sg13g2_nor2b_1 _31370_ (.A(\u_inv.d_reg[108] ),
    .B_N(\u_inv.d_next[108] ),
    .Y(_05648_));
 sg13g2_a21oi_1 _31371_ (.A1(_05468_),
    .A2(_05648_),
    .Y(_05649_),
    .B1(_05467_));
 sg13g2_nand2_1 _31372_ (.Y(_05650_),
    .A(\u_inv.d_next[110] ),
    .B(_14699_));
 sg13g2_nand2_1 _31373_ (.Y(_05651_),
    .A(\u_inv.d_next[111] ),
    .B(_14698_));
 sg13g2_o21ai_1 _31374_ (.B1(_05651_),
    .Y(_05652_),
    .A1(_05466_),
    .A2(_05649_));
 sg13g2_nor3_1 _31375_ (.A(_05640_),
    .B(_05647_),
    .C(_05652_),
    .Y(_05653_));
 sg13g2_o21ai_1 _31376_ (.B1(_05653_),
    .Y(_05654_),
    .A1(_05462_),
    .A2(_05650_));
 sg13g2_nor2b_1 _31377_ (.A(\u_inv.d_reg[64] ),
    .B_N(\u_inv.d_next[64] ),
    .Y(_05655_));
 sg13g2_a21oi_1 _31378_ (.A1(_05399_),
    .A2(_05655_),
    .Y(_05656_),
    .B1(_05398_));
 sg13g2_nor2_1 _31379_ (.A(_05397_),
    .B(_05656_),
    .Y(_05657_));
 sg13g2_nand2_1 _31380_ (.Y(_05658_),
    .A(net5880),
    .B(_14743_));
 sg13g2_a21oi_1 _31381_ (.A1(_05392_),
    .A2(_05658_),
    .Y(_05659_),
    .B1(_05391_));
 sg13g2_o21ai_1 _31382_ (.B1(_05390_),
    .Y(_05660_),
    .A1(_05657_),
    .A2(_05659_));
 sg13g2_nand2b_1 _31383_ (.Y(_05661_),
    .B(\u_inv.d_next[68] ),
    .A_N(\u_inv.d_reg[68] ));
 sg13g2_nor2_1 _31384_ (.A(_05384_),
    .B(_05661_),
    .Y(_05662_));
 sg13g2_a21oi_1 _31385_ (.A1(\u_inv.d_next[69] ),
    .A2(_14740_),
    .Y(_05663_),
    .B1(_05662_));
 sg13g2_nand2b_1 _31386_ (.Y(_05664_),
    .B(_05381_),
    .A_N(_05663_));
 sg13g2_nor2b_1 _31387_ (.A(\u_inv.d_reg[70] ),
    .B_N(net5879),
    .Y(_05665_));
 sg13g2_o21ai_1 _31388_ (.B1(_05665_),
    .Y(_05666_),
    .A1(\u_inv.d_next[71] ),
    .A2(_14738_));
 sg13g2_nand4_1 _31389_ (.B(_05660_),
    .C(_05664_),
    .A(_05376_),
    .Y(_05667_),
    .D(_05666_));
 sg13g2_inv_1 _31390_ (.Y(_05668_),
    .A(_05667_));
 sg13g2_nor2b_1 _31391_ (.A(net5872),
    .B_N(\u_inv.d_next[77] ),
    .Y(_05669_));
 sg13g2_nor2b_1 _31392_ (.A(\u_inv.d_reg[76] ),
    .B_N(\u_inv.d_next[76] ),
    .Y(_05670_));
 sg13g2_a21oi_1 _31393_ (.A1(_05356_),
    .A2(_05670_),
    .Y(_05671_),
    .B1(_05669_));
 sg13g2_nor2b_1 _31394_ (.A(\u_inv.d_reg[78] ),
    .B_N(\u_inv.d_next[78] ),
    .Y(_05672_));
 sg13g2_a21o_1 _31395_ (.A2(_14730_),
    .A1(\u_inv.d_next[79] ),
    .B1(_05672_),
    .X(_05673_));
 sg13g2_o21ai_1 _31396_ (.B1(_05673_),
    .Y(_05674_),
    .A1(\u_inv.d_next[79] ),
    .A2(_14730_));
 sg13g2_o21ai_1 _31397_ (.B1(_05674_),
    .Y(_05675_),
    .A1(_05354_),
    .A2(_05671_));
 sg13g2_and3_1 _31398_ (.X(_05676_),
    .A(net5878),
    .B(_14737_),
    .C(_05370_));
 sg13g2_a21oi_2 _31399_ (.B1(_05676_),
    .Y(_05677_),
    .A2(_14736_),
    .A1(\u_inv.d_next[73] ));
 sg13g2_nand2_1 _31400_ (.Y(_05678_),
    .A(net5877),
    .B(_14735_));
 sg13g2_o21ai_1 _31401_ (.B1(_05363_),
    .Y(_05679_),
    .A1(_05362_),
    .A2(_05678_));
 sg13g2_inv_1 _31402_ (.Y(_05680_),
    .A(_05679_));
 sg13g2_o21ai_1 _31403_ (.B1(_05680_),
    .Y(_05681_),
    .A1(_05368_),
    .A2(_05677_));
 sg13g2_a22oi_1 _31404_ (.Y(_05682_),
    .B1(_05681_),
    .B2(_05361_),
    .A2(_05667_),
    .A1(_05375_));
 sg13g2_nand2b_2 _31405_ (.Y(_05683_),
    .B(_05682_),
    .A_N(_05675_));
 sg13g2_inv_2 _31406_ (.Y(_05684_),
    .A(_05683_));
 sg13g2_a221oi_1 _31407_ (.B2(_05620_),
    .C1(_05626_),
    .B1(_05524_),
    .A1(\u_inv.d_next[95] ),
    .Y(_05685_),
    .A2(_14714_));
 sg13g2_o21ai_1 _31408_ (.B1(_05685_),
    .Y(_05686_),
    .A1(_05537_),
    .A2(_05614_));
 sg13g2_a21oi_1 _31409_ (.A1(_05566_),
    .A2(_05683_),
    .Y(_05687_),
    .B1(_05686_));
 sg13g2_nand2_2 _31410_ (.Y(_05688_),
    .A(_05622_),
    .B(_05687_));
 sg13g2_a22oi_1 _31411_ (.Y(_05689_),
    .B1(_05688_),
    .B2(_05513_),
    .A2(_05654_),
    .A1(_05460_));
 sg13g2_and3_2 _31412_ (.X(_05690_),
    .A(_05583_),
    .B(_05598_),
    .C(_05689_));
 sg13g2_and2_1 _31413_ (.A(_05569_),
    .B(_05690_),
    .X(_05691_));
 sg13g2_nor2b_2 _31414_ (.A(_04887_),
    .B_N(_04888_),
    .Y(_05692_));
 sg13g2_inv_2 _31415_ (.Y(_05693_),
    .A(_05692_));
 sg13g2_nand2_1 _31416_ (.Y(_05694_),
    .A(\u_inv.d_next[128] ),
    .B(\u_inv.d_reg[128] ));
 sg13g2_xor2_1 _31417_ (.B(\u_inv.d_reg[128] ),
    .A(\u_inv.d_next[128] ),
    .X(_05695_));
 sg13g2_xnor2_1 _31418_ (.Y(_05696_),
    .A(\u_inv.d_next[128] ),
    .B(\u_inv.d_reg[128] ));
 sg13g2_nand2_1 _31419_ (.Y(_05697_),
    .A(_05692_),
    .B(_05696_));
 sg13g2_nor2_1 _31420_ (.A(_04881_),
    .B(_05697_),
    .Y(_05698_));
 sg13g2_nand2_1 _31421_ (.Y(_05699_),
    .A(_04885_),
    .B(_05698_));
 sg13g2_nand4_1 _31422_ (.B(_04885_),
    .C(_04912_),
    .A(_04834_),
    .Y(_05700_),
    .D(_05698_));
 sg13g2_or2_1 _31423_ (.X(_05701_),
    .B(_05700_),
    .A(_04789_));
 sg13g2_a21o_2 _31424_ (.A2(_05690_),
    .A1(_05569_),
    .B1(_05701_),
    .X(_05702_));
 sg13g2_nand2_2 _31425_ (.Y(_05703_),
    .A(_05009_),
    .B(_05702_));
 sg13g2_a21oi_2 _31426_ (.B1(_04684_),
    .Y(_05704_),
    .A2(_05702_),
    .A1(_05009_));
 sg13g2_nor2b_1 _31427_ (.A(\u_inv.d_reg[226] ),
    .B_N(\u_inv.d_next[226] ),
    .Y(_05705_));
 sg13g2_nand2_1 _31428_ (.Y(_05706_),
    .A(\u_inv.d_next[224] ),
    .B(_14585_));
 sg13g2_nor2_1 _31429_ (.A(_04566_),
    .B(_05706_),
    .Y(_05707_));
 sg13g2_a21oi_1 _31430_ (.A1(net5875),
    .A2(_14584_),
    .Y(_05708_),
    .B1(_05707_));
 sg13g2_a21o_1 _31431_ (.A2(_14584_),
    .A1(net5875),
    .B1(_05707_),
    .X(_05709_));
 sg13g2_a21oi_1 _31432_ (.A1(_04562_),
    .A2(_05709_),
    .Y(_05710_),
    .B1(_05705_));
 sg13g2_nor2_1 _31433_ (.A(_04559_),
    .B(_05710_),
    .Y(_05711_));
 sg13g2_a21oi_2 _31434_ (.B1(_05711_),
    .Y(_05712_),
    .A2(_14582_),
    .A1(\u_inv.d_next[227] ));
 sg13g2_nor2b_1 _31435_ (.A(\u_inv.d_reg[231] ),
    .B_N(\u_inv.d_next[231] ),
    .Y(_05713_));
 sg13g2_nor2b_1 _31436_ (.A(\u_inv.d_reg[230] ),
    .B_N(\u_inv.d_next[230] ),
    .Y(_05714_));
 sg13g2_nand2_1 _31437_ (.Y(_05715_),
    .A(\u_inv.d_next[230] ),
    .B(_14579_));
 sg13g2_nand2_1 _31438_ (.Y(_05716_),
    .A(\u_inv.d_next[229] ),
    .B(_14580_));
 sg13g2_nor2b_1 _31439_ (.A(\u_inv.d_reg[228] ),
    .B_N(\u_inv.d_next[228] ),
    .Y(_05717_));
 sg13g2_nand2_1 _31440_ (.Y(_05718_),
    .A(\u_inv.d_next[228] ),
    .B(_14581_));
 sg13g2_o21ai_1 _31441_ (.B1(_05716_),
    .Y(_05719_),
    .A1(_04548_),
    .A2(_05718_));
 sg13g2_a21oi_1 _31442_ (.A1(_04556_),
    .A2(_05714_),
    .Y(_05720_),
    .B1(_05713_));
 sg13g2_o21ai_1 _31443_ (.B1(_05720_),
    .Y(_05721_),
    .A1(_04558_),
    .A2(_05712_));
 sg13g2_a21oi_2 _31444_ (.B1(_05721_),
    .Y(_05722_),
    .A2(_05719_),
    .A1(_04557_));
 sg13g2_inv_1 _31445_ (.Y(_05723_),
    .A(_05722_));
 sg13g2_nor2b_1 _31446_ (.A(\u_inv.d_reg[237] ),
    .B_N(\u_inv.d_next[237] ),
    .Y(_05724_));
 sg13g2_nor2b_1 _31447_ (.A(\u_inv.d_reg[236] ),
    .B_N(\u_inv.d_next[236] ),
    .Y(_05725_));
 sg13g2_nand2_1 _31448_ (.Y(_05726_),
    .A(\u_inv.d_next[236] ),
    .B(_14573_));
 sg13g2_a21oi_1 _31449_ (.A1(_04523_),
    .A2(_05725_),
    .Y(_05727_),
    .B1(_05724_));
 sg13g2_nor2b_1 _31450_ (.A(\u_inv.d_reg[238] ),
    .B_N(\u_inv.d_next[238] ),
    .Y(_05728_));
 sg13g2_nor2_1 _31451_ (.A(_14175_),
    .B(\u_inv.d_reg[239] ),
    .Y(_05729_));
 sg13g2_a21oi_1 _31452_ (.A1(_04516_),
    .A2(_05728_),
    .Y(_05730_),
    .B1(_05729_));
 sg13g2_o21ai_1 _31453_ (.B1(_05730_),
    .Y(_05731_),
    .A1(_04520_),
    .A2(_05727_));
 sg13g2_nor2_1 _31454_ (.A(_14177_),
    .B(\u_inv.d_reg[232] ),
    .Y(_05732_));
 sg13g2_nand2_1 _31455_ (.Y(_05733_),
    .A(_04540_),
    .B(_05732_));
 sg13g2_o21ai_1 _31456_ (.B1(_05733_),
    .Y(_05734_),
    .A1(_14176_),
    .A2(\u_inv.d_reg[233] ));
 sg13g2_nand2_1 _31457_ (.Y(_05735_),
    .A(\u_inv.d_next[234] ),
    .B(_14575_));
 sg13g2_a22oi_1 _31458_ (.Y(_05736_),
    .B1(_04538_),
    .B2(_05734_),
    .A2(_14574_),
    .A1(\u_inv.d_next[235] ));
 sg13g2_o21ai_1 _31459_ (.B1(_05736_),
    .Y(_05737_),
    .A1(_04532_),
    .A2(_05735_));
 sg13g2_a221oi_1 _31460_ (.B2(_04529_),
    .C1(_05731_),
    .B1(_05737_),
    .A1(_04547_),
    .Y(_05738_),
    .A2(_05723_));
 sg13g2_nand2b_1 _31461_ (.Y(_05739_),
    .B(_04514_),
    .A_N(_05738_));
 sg13g2_nor2b_1 _31462_ (.A(\u_inv.d_reg[192] ),
    .B_N(\u_inv.d_next[192] ),
    .Y(_05740_));
 sg13g2_a21oi_1 _31463_ (.A1(\u_inv.d_next[193] ),
    .A2(_14616_),
    .Y(_05741_),
    .B1(_05740_));
 sg13g2_a21oi_1 _31464_ (.A1(_14190_),
    .A2(\u_inv.d_reg[193] ),
    .Y(_05742_),
    .B1(_05741_));
 sg13g2_nand2_1 _31465_ (.Y(_05743_),
    .A(\u_inv.d_next[194] ),
    .B(_14615_));
 sg13g2_nor2b_1 _31466_ (.A(_05743_),
    .B_N(_04675_),
    .Y(_05744_));
 sg13g2_a22oi_1 _31467_ (.Y(_05745_),
    .B1(_04678_),
    .B2(_05742_),
    .A2(_14614_),
    .A1(\u_inv.d_next[195] ));
 sg13g2_nand2b_2 _31468_ (.Y(_05746_),
    .B(_05745_),
    .A_N(_05744_));
 sg13g2_nand2_1 _31469_ (.Y(_05747_),
    .A(_04670_),
    .B(_05746_));
 sg13g2_nor2b_1 _31470_ (.A(\u_inv.d_reg[197] ),
    .B_N(\u_inv.d_next[197] ),
    .Y(_05748_));
 sg13g2_nor2b_1 _31471_ (.A(\u_inv.d_reg[196] ),
    .B_N(\u_inv.d_next[196] ),
    .Y(_05749_));
 sg13g2_nand2_1 _31472_ (.Y(_05750_),
    .A(\u_inv.d_next[196] ),
    .B(_14613_));
 sg13g2_a21oi_1 _31473_ (.A1(_04661_),
    .A2(_05749_),
    .Y(_05751_),
    .B1(_05748_));
 sg13g2_nor2_1 _31474_ (.A(_14188_),
    .B(\u_inv.d_reg[199] ),
    .Y(_05752_));
 sg13g2_nand2_1 _31475_ (.Y(_05753_),
    .A(\u_inv.d_next[198] ),
    .B(_14611_));
 sg13g2_o21ai_1 _31476_ (.B1(_05753_),
    .Y(_05754_),
    .A1(_04669_),
    .A2(_05751_));
 sg13g2_a21oi_1 _31477_ (.A1(_04667_),
    .A2(_05754_),
    .Y(_05755_),
    .B1(_05752_));
 sg13g2_nand2_2 _31478_ (.Y(_05756_),
    .A(_05747_),
    .B(_05755_));
 sg13g2_nor2_1 _31479_ (.A(_14186_),
    .B(\u_inv.d_reg[205] ),
    .Y(_05757_));
 sg13g2_nor2b_1 _31480_ (.A(\u_inv.d_reg[204] ),
    .B_N(\u_inv.d_next[204] ),
    .Y(_05758_));
 sg13g2_a21o_1 _31481_ (.A2(_05758_),
    .A1(_04640_),
    .B1(_05757_),
    .X(_05759_));
 sg13g2_nand2_1 _31482_ (.Y(_05760_),
    .A(\u_inv.d_next[206] ),
    .B(_14603_));
 sg13g2_nor2_1 _31483_ (.A(_04633_),
    .B(_05760_),
    .Y(_05761_));
 sg13g2_nand2_1 _31484_ (.Y(_05762_),
    .A(\u_inv.d_next[200] ),
    .B(_14609_));
 sg13g2_nor2_1 _31485_ (.A(_04652_),
    .B(_05762_),
    .Y(_05763_));
 sg13g2_a21oi_1 _31486_ (.A1(\u_inv.d_next[201] ),
    .A2(_14608_),
    .Y(_05764_),
    .B1(_05763_));
 sg13g2_nor2b_1 _31487_ (.A(\u_inv.d_reg[202] ),
    .B_N(\u_inv.d_next[202] ),
    .Y(_05765_));
 sg13g2_nand2_1 _31488_ (.Y(_05766_),
    .A(\u_inv.d_next[203] ),
    .B(_14606_));
 sg13g2_o21ai_1 _31489_ (.B1(_05766_),
    .Y(_05767_),
    .A1(_04649_),
    .A2(_05764_));
 sg13g2_a21oi_1 _31490_ (.A1(_04646_),
    .A2(_05765_),
    .Y(_05768_),
    .B1(_05767_));
 sg13g2_a21oi_1 _31491_ (.A1(_04637_),
    .A2(_05759_),
    .Y(_05769_),
    .B1(_05761_));
 sg13g2_o21ai_1 _31492_ (.B1(_05769_),
    .Y(_05770_),
    .A1(_04645_),
    .A2(_05768_));
 sg13g2_a21oi_1 _31493_ (.A1(_04658_),
    .A2(_05756_),
    .Y(_05771_),
    .B1(_05770_));
 sg13g2_o21ai_1 _31494_ (.B1(_05771_),
    .Y(_05772_),
    .A1(_14185_),
    .A2(\u_inv.d_reg[207] ));
 sg13g2_nor2b_1 _31495_ (.A(\u_inv.d_reg[216] ),
    .B_N(\u_inv.d_next[216] ),
    .Y(_05773_));
 sg13g2_nand2b_1 _31496_ (.Y(_05774_),
    .B(_05773_),
    .A_N(_04599_));
 sg13g2_o21ai_1 _31497_ (.B1(_05774_),
    .Y(_05775_),
    .A1(_14182_),
    .A2(\u_inv.d_reg[217] ));
 sg13g2_nand2_1 _31498_ (.Y(_05776_),
    .A(\u_inv.d_next[218] ),
    .B(_14591_));
 sg13g2_inv_1 _31499_ (.Y(_05777_),
    .A(_05776_));
 sg13g2_a22oi_1 _31500_ (.Y(_05778_),
    .B1(_04596_),
    .B2(_05775_),
    .A2(_14590_),
    .A1(\u_inv.d_next[219] ));
 sg13g2_o21ai_1 _31501_ (.B1(_05778_),
    .Y(_05779_),
    .A1(_04591_),
    .A2(_05776_));
 sg13g2_nand2_1 _31502_ (.Y(_05780_),
    .A(\u_inv.d_next[220] ),
    .B(_14589_));
 sg13g2_nor2_1 _31503_ (.A(_04583_),
    .B(_05780_),
    .Y(_05781_));
 sg13g2_a21oi_1 _31504_ (.A1(\u_inv.d_next[221] ),
    .A2(_14588_),
    .Y(_05782_),
    .B1(_05781_));
 sg13g2_nor2_1 _31505_ (.A(_14180_),
    .B(\u_inv.d_reg[222] ),
    .Y(_05783_));
 sg13g2_nand2_1 _31506_ (.Y(_05784_),
    .A(_04578_),
    .B(_05783_));
 sg13g2_o21ai_1 _31507_ (.B1(_05784_),
    .Y(_05785_),
    .A1(_04582_),
    .A2(_05782_));
 sg13g2_a221oi_1 _31508_ (.B2(_05779_),
    .C1(_05785_),
    .B1(_04589_),
    .A1(\u_inv.d_next[223] ),
    .Y(_05786_),
    .A2(_14586_));
 sg13g2_nor2b_1 _31509_ (.A(\u_inv.d_reg[208] ),
    .B_N(\u_inv.d_next[208] ),
    .Y(_05787_));
 sg13g2_nand2_1 _31510_ (.Y(_05788_),
    .A(_04627_),
    .B(_05787_));
 sg13g2_o21ai_1 _31511_ (.B1(_05788_),
    .Y(_05789_),
    .A1(_14184_),
    .A2(\u_inv.d_reg[209] ));
 sg13g2_nor2b_1 _31512_ (.A(\u_inv.d_reg[211] ),
    .B_N(\u_inv.d_next[211] ),
    .Y(_05790_));
 sg13g2_nor2b_1 _31513_ (.A(\u_inv.d_reg[210] ),
    .B_N(\u_inv.d_next[210] ),
    .Y(_05791_));
 sg13g2_a221oi_1 _31514_ (.B2(_04622_),
    .C1(_05790_),
    .B1(_05791_),
    .A1(_04625_),
    .Y(_05792_),
    .A2(_05789_));
 sg13g2_nand2_1 _31515_ (.Y(_05793_),
    .A(\u_inv.d_next[213] ),
    .B(_14596_));
 sg13g2_nand2_1 _31516_ (.Y(_05794_),
    .A(\u_inv.d_next[212] ),
    .B(_14597_));
 sg13g2_o21ai_1 _31517_ (.B1(_05793_),
    .Y(_05795_),
    .A1(_04606_),
    .A2(_05794_));
 sg13g2_nand2_1 _31518_ (.Y(_05796_),
    .A(\u_inv.d_next[214] ),
    .B(_14595_));
 sg13g2_nor2_1 _31519_ (.A(_04616_),
    .B(_05796_),
    .Y(_05797_));
 sg13g2_a21oi_1 _31520_ (.A1(\u_inv.d_next[215] ),
    .A2(_14594_),
    .Y(_05798_),
    .B1(_05797_));
 sg13g2_o21ai_1 _31521_ (.B1(_05798_),
    .Y(_05799_),
    .A1(_04619_),
    .A2(_05792_));
 sg13g2_a21oi_1 _31522_ (.A1(_04618_),
    .A2(_05795_),
    .Y(_05800_),
    .B1(_05799_));
 sg13g2_o21ai_1 _31523_ (.B1(_05786_),
    .Y(_05801_),
    .A1(_04605_),
    .A2(_05800_));
 sg13g2_a21o_2 _31524_ (.A2(_05772_),
    .A1(_04632_),
    .B1(_05801_),
    .X(_05802_));
 sg13g2_nand2b_1 _31525_ (.Y(_05803_),
    .B(_05802_),
    .A_N(_04576_));
 sg13g2_nand2_1 _31526_ (.Y(_05804_),
    .A(\u_inv.d_next[242] ),
    .B(_14567_));
 sg13g2_nor2b_1 _31527_ (.A(net5865),
    .B_N(\u_inv.d_next[240] ),
    .Y(_05805_));
 sg13g2_nand2_1 _31528_ (.Y(_05806_),
    .A(_04504_),
    .B(_05805_));
 sg13g2_o21ai_1 _31529_ (.B1(_05806_),
    .Y(_05807_),
    .A1(_14174_),
    .A2(\u_inv.d_reg[241] ));
 sg13g2_a22oi_1 _31530_ (.Y(_05808_),
    .B1(_04503_),
    .B2(_05807_),
    .A2(_14566_),
    .A1(\u_inv.d_next[243] ));
 sg13g2_o21ai_1 _31531_ (.B1(_05808_),
    .Y(_05809_),
    .A1(_04498_),
    .A2(_05804_));
 sg13g2_nand2_1 _31532_ (.Y(_05810_),
    .A(\u_inv.d_next[244] ),
    .B(_14565_));
 sg13g2_nor2b_1 _31533_ (.A(_05810_),
    .B_N(_04485_),
    .Y(_05811_));
 sg13g2_a21oi_1 _31534_ (.A1(\u_inv.d_next[245] ),
    .A2(_14564_),
    .Y(_05812_),
    .B1(_05811_));
 sg13g2_nor2_1 _31535_ (.A(_14173_),
    .B(\u_inv.d_reg[246] ),
    .Y(_05813_));
 sg13g2_nor2_1 _31536_ (.A(_04492_),
    .B(_05812_),
    .Y(_05814_));
 sg13g2_o21ai_1 _31537_ (.B1(_04494_),
    .Y(_05815_),
    .A1(_05813_),
    .A2(_05814_));
 sg13g2_a22oi_1 _31538_ (.Y(_05816_),
    .B1(_04495_),
    .B2(_05809_),
    .A2(_14562_),
    .A1(\u_inv.d_next[247] ));
 sg13g2_nand2_2 _31539_ (.Y(_05817_),
    .A(_05815_),
    .B(_05816_));
 sg13g2_nor2b_1 _31540_ (.A(\u_inv.d_reg[250] ),
    .B_N(\u_inv.d_next[250] ),
    .Y(_05818_));
 sg13g2_nand2_1 _31541_ (.Y(_05819_),
    .A(\u_inv.d_next[248] ),
    .B(_14561_));
 sg13g2_nor2_1 _31542_ (.A(_04474_),
    .B(_05819_),
    .Y(_05820_));
 sg13g2_a21oi_1 _31543_ (.A1(\u_inv.d_next[249] ),
    .A2(_14560_),
    .Y(_05821_),
    .B1(_05820_));
 sg13g2_inv_1 _31544_ (.Y(_05822_),
    .A(_05821_));
 sg13g2_nor2b_1 _31545_ (.A(_04470_),
    .B_N(_05818_),
    .Y(_05823_));
 sg13g2_a221oi_1 _31546_ (.B2(_05822_),
    .C1(_05823_),
    .B1(_04471_),
    .A1(\u_inv.d_next[251] ),
    .Y(_05824_),
    .A2(_14558_));
 sg13g2_nand2_1 _31547_ (.Y(_05825_),
    .A(\u_inv.d_next[253] ),
    .B(_14556_));
 sg13g2_nand2_1 _31548_ (.Y(_05826_),
    .A(\u_inv.d_next[252] ),
    .B(_14557_));
 sg13g2_o21ai_1 _31549_ (.B1(_05825_),
    .Y(_05827_),
    .A1(_04460_),
    .A2(_05826_));
 sg13g2_nand2_1 _31550_ (.Y(_05828_),
    .A(\u_inv.d_next[254] ),
    .B(_14555_));
 sg13g2_nor2_1 _31551_ (.A(_04452_),
    .B(_05828_),
    .Y(_05829_));
 sg13g2_a221oi_1 _31552_ (.B2(_05827_),
    .C1(_05829_),
    .B1(_04457_),
    .A1(\u_inv.d_next[255] ),
    .Y(_05830_),
    .A2(_14554_));
 sg13g2_o21ai_1 _31553_ (.B1(_05830_),
    .Y(_05831_),
    .A1(_04466_),
    .A2(_05824_));
 sg13g2_a21oi_1 _31554_ (.A1(_04482_),
    .A2(_05817_),
    .Y(_05832_),
    .B1(_05831_));
 sg13g2_nand3_1 _31555_ (.B(_05803_),
    .C(_05832_),
    .A(_05739_),
    .Y(_05833_));
 sg13g2_o21ai_1 _31556_ (.B1(_04448_),
    .Y(_05834_),
    .A1(_05704_),
    .A2(_05833_));
 sg13g2_a21oi_2 _31557_ (.B1(net5020),
    .Y(_05835_),
    .A2(\u_inv.d_reg[256] ),
    .A1(_14172_));
 sg13g2_nor2_1 _31558_ (.A(_04453_),
    .B(_04456_),
    .Y(_05836_));
 sg13g2_nand2_1 _31559_ (.Y(_05837_),
    .A(_04460_),
    .B(_04463_));
 sg13g2_nor3_1 _31560_ (.A(_04453_),
    .B(_04456_),
    .C(_05837_),
    .Y(_05838_));
 sg13g2_and2_1 _31561_ (.A(_04468_),
    .B(_04470_),
    .X(_05839_));
 sg13g2_nand2_1 _31562_ (.Y(_05840_),
    .A(_04474_),
    .B(_04477_));
 sg13g2_nand4_1 _31563_ (.B(_04477_),
    .C(_05838_),
    .A(_04474_),
    .Y(_05841_),
    .D(_05839_));
 sg13g2_and2_1 _31564_ (.A(_04492_),
    .B(_04493_),
    .X(_05842_));
 sg13g2_nor2_1 _31565_ (.A(_04485_),
    .B(_04489_),
    .Y(_05843_));
 sg13g2_nand2_1 _31566_ (.Y(_05844_),
    .A(_05842_),
    .B(_05843_));
 sg13g2_nand2_1 _31567_ (.Y(_05845_),
    .A(_04498_),
    .B(_04501_));
 sg13g2_nor2b_1 _31568_ (.A(_04504_),
    .B_N(_04507_),
    .Y(_05846_));
 sg13g2_nand3_1 _31569_ (.B(_05843_),
    .C(_05846_),
    .A(_05842_),
    .Y(_05847_));
 sg13g2_or2_1 _31570_ (.X(_05848_),
    .B(_05847_),
    .A(_05845_));
 sg13g2_inv_1 _31571_ (.Y(_05849_),
    .A(_05848_));
 sg13g2_nor2_1 _31572_ (.A(_05841_),
    .B(_05848_),
    .Y(_05850_));
 sg13g2_nor2_1 _31573_ (.A(_04516_),
    .B(_04518_),
    .Y(_05851_));
 sg13g2_nor2_1 _31574_ (.A(_04523_),
    .B(_04526_),
    .Y(_05852_));
 sg13g2_nand2_1 _31575_ (.Y(_05853_),
    .A(_05851_),
    .B(_05852_));
 sg13g2_nand2_1 _31576_ (.Y(_05854_),
    .A(_04532_),
    .B(_04536_));
 sg13g2_nand2_1 _31577_ (.Y(_05855_),
    .A(_04539_),
    .B(_04541_));
 sg13g2_inv_1 _31578_ (.Y(_05856_),
    .A(_05855_));
 sg13g2_nor3_1 _31579_ (.A(_05853_),
    .B(_05854_),
    .C(_05855_),
    .Y(_05857_));
 sg13g2_nor2_1 _31580_ (.A(_04554_),
    .B(_04556_),
    .Y(_05858_));
 sg13g2_nor2_1 _31581_ (.A(_04560_),
    .B(_04562_),
    .Y(_05859_));
 sg13g2_inv_1 _31582_ (.Y(_05860_),
    .A(_05859_));
 sg13g2_and2_1 _31583_ (.A(_04548_),
    .B(_04550_),
    .X(_05861_));
 sg13g2_and2_1 _31584_ (.A(_05858_),
    .B(_05861_),
    .X(_05862_));
 sg13g2_and4_1 _31585_ (.A(_04566_),
    .B(_04569_),
    .C(_05859_),
    .D(_05862_),
    .X(_05863_));
 sg13g2_inv_1 _31586_ (.Y(_05864_),
    .A(_05863_));
 sg13g2_and2_1 _31587_ (.A(_05857_),
    .B(_05863_),
    .X(_05865_));
 sg13g2_inv_1 _31588_ (.Y(_05866_),
    .A(_05865_));
 sg13g2_nand2_1 _31589_ (.Y(_05867_),
    .A(_05850_),
    .B(_05865_));
 sg13g2_a22oi_1 _31590_ (.Y(_05868_),
    .B1(net5865),
    .B2(\u_inv.d_next[240] ),
    .A2(\u_inv.d_reg[241] ),
    .A1(\u_inv.d_next[241] ));
 sg13g2_a21o_1 _31591_ (.A2(_14568_),
    .A1(_14174_),
    .B1(_05868_),
    .X(_05869_));
 sg13g2_nor2_1 _31592_ (.A(_05845_),
    .B(_05869_),
    .Y(_05870_));
 sg13g2_o21ai_1 _31593_ (.B1(_04497_),
    .Y(_05871_),
    .A1(_04496_),
    .A2(_04500_));
 sg13g2_nor2_1 _31594_ (.A(_05870_),
    .B(_05871_),
    .Y(_05872_));
 sg13g2_a22oi_1 _31595_ (.Y(_05873_),
    .B1(\u_inv.d_reg[246] ),
    .B2(\u_inv.d_next[246] ),
    .A2(\u_inv.d_reg[247] ),
    .A1(\u_inv.d_next[247] ));
 sg13g2_inv_1 _31596_ (.Y(_05874_),
    .A(_05873_));
 sg13g2_o21ai_1 _31597_ (.B1(_05874_),
    .Y(_05875_),
    .A1(\u_inv.d_next[247] ),
    .A2(\u_inv.d_reg[247] ));
 sg13g2_o21ai_1 _31598_ (.B1(_04484_),
    .Y(_05876_),
    .A1(_04483_),
    .A2(_04486_));
 sg13g2_o21ai_1 _31599_ (.B1(_05875_),
    .Y(_05877_),
    .A1(_05844_),
    .A2(_05872_));
 sg13g2_a21oi_2 _31600_ (.B1(_05877_),
    .Y(_05878_),
    .A2(_05876_),
    .A1(_05842_));
 sg13g2_o21ai_1 _31601_ (.B1(_04473_),
    .Y(_05879_),
    .A1(_04472_),
    .A2(_04476_));
 sg13g2_a22oi_1 _31602_ (.Y(_05880_),
    .B1(_05839_),
    .B2(_05879_),
    .A2(\u_inv.d_reg[251] ),
    .A1(\u_inv.d_next[251] ));
 sg13g2_o21ai_1 _31603_ (.B1(_05880_),
    .Y(_05881_),
    .A1(_04467_),
    .A2(_04469_));
 sg13g2_o21ai_1 _31604_ (.B1(_04459_),
    .Y(_05882_),
    .A1(_04458_),
    .A2(_04461_));
 sg13g2_o21ai_1 _31605_ (.B1(_04451_),
    .Y(_05883_),
    .A1(_04450_),
    .A2(_04454_));
 sg13g2_a221oi_1 _31606_ (.B2(_05836_),
    .C1(_05883_),
    .B1(_05882_),
    .A1(_05838_),
    .Y(_05884_),
    .A2(_05881_));
 sg13g2_o21ai_1 _31607_ (.B1(_05884_),
    .Y(_05885_),
    .A1(_05841_),
    .A2(_05878_));
 sg13g2_a22oi_1 _31608_ (.Y(_05886_),
    .B1(\u_inv.d_reg[230] ),
    .B2(\u_inv.d_next[230] ),
    .A2(\u_inv.d_reg[231] ),
    .A1(\u_inv.d_next[231] ));
 sg13g2_a21oi_1 _31609_ (.A1(\u_inv.d_next[229] ),
    .A2(\u_inv.d_reg[229] ),
    .Y(_05887_),
    .B1(_04549_));
 sg13g2_a21oi_1 _31610_ (.A1(_14178_),
    .A2(_14580_),
    .Y(_05888_),
    .B1(_05887_));
 sg13g2_a21oi_1 _31611_ (.A1(_04564_),
    .A2(_04568_),
    .Y(_05889_),
    .B1(_04565_));
 sg13g2_inv_1 _31612_ (.Y(_05890_),
    .A(_05889_));
 sg13g2_a21oi_1 _31613_ (.A1(_14179_),
    .A2(_14582_),
    .Y(_05891_),
    .B1(_04561_));
 sg13g2_a21oi_1 _31614_ (.A1(\u_inv.d_next[227] ),
    .A2(\u_inv.d_reg[227] ),
    .Y(_05892_),
    .B1(_05891_));
 sg13g2_o21ai_1 _31615_ (.B1(_05892_),
    .Y(_05893_),
    .A1(_05860_),
    .A2(_05890_));
 sg13g2_a22oi_1 _31616_ (.Y(_05894_),
    .B1(_05893_),
    .B2(_05862_),
    .A2(_05888_),
    .A1(_05858_));
 sg13g2_o21ai_1 _31617_ (.B1(_05894_),
    .Y(_05895_),
    .A1(_04555_),
    .A2(_05886_));
 sg13g2_a22oi_1 _31618_ (.Y(_05896_),
    .B1(\u_inv.d_reg[232] ),
    .B2(\u_inv.d_next[232] ),
    .A2(\u_inv.d_reg[233] ),
    .A1(\u_inv.d_next[233] ));
 sg13g2_a21o_1 _31619_ (.A2(_14576_),
    .A1(_14176_),
    .B1(_05896_),
    .X(_05897_));
 sg13g2_o21ai_1 _31620_ (.B1(_04531_),
    .Y(_05898_),
    .A1(_05854_),
    .A2(_05897_));
 sg13g2_a21oi_1 _31621_ (.A1(_04530_),
    .A2(_04535_),
    .Y(_05899_),
    .B1(_05898_));
 sg13g2_o21ai_1 _31622_ (.B1(_04522_),
    .Y(_05900_),
    .A1(_04521_),
    .A2(_04524_));
 sg13g2_a21oi_1 _31623_ (.A1(_14175_),
    .A2(_14570_),
    .Y(_05901_),
    .B1(_04517_));
 sg13g2_a221oi_1 _31624_ (.B2(_05900_),
    .C1(_05901_),
    .B1(_05851_),
    .A1(\u_inv.d_next[239] ),
    .Y(_05902_),
    .A2(\u_inv.d_reg[239] ));
 sg13g2_o21ai_1 _31625_ (.B1(_05902_),
    .Y(_05903_),
    .A1(_05853_),
    .A2(_05899_));
 sg13g2_a21o_2 _31626_ (.A2(_05895_),
    .A1(_05857_),
    .B1(_05903_),
    .X(_05904_));
 sg13g2_a21oi_1 _31627_ (.A1(_05850_),
    .A2(_05904_),
    .Y(_05905_),
    .B1(_05885_));
 sg13g2_nor2_1 _31628_ (.A(_04741_),
    .B(_04743_),
    .Y(_05906_));
 sg13g2_or4_1 _31629_ (.A(_04736_),
    .B(_04738_),
    .C(_04741_),
    .D(_04743_),
    .X(_05907_));
 sg13g2_or2_1 _31630_ (.X(_05908_),
    .B(_04751_),
    .A(_04749_));
 sg13g2_nand2_1 _31631_ (.Y(_05909_),
    .A(_04753_),
    .B(_04754_));
 sg13g2_or3_1 _31632_ (.A(_05907_),
    .B(_05908_),
    .C(_05909_),
    .X(_05910_));
 sg13g2_nand2_1 _31633_ (.Y(_05911_),
    .A(_04764_),
    .B(_04767_));
 sg13g2_nor3_2 _31634_ (.A(_04759_),
    .B(_04762_),
    .C(_05911_),
    .Y(_05912_));
 sg13g2_nand2b_2 _31635_ (.Y(_05913_),
    .B(_05912_),
    .A_N(_05910_));
 sg13g2_nor2_1 _31636_ (.A(_04691_),
    .B(_04694_),
    .Y(_05914_));
 sg13g2_nor4_1 _31637_ (.A(_04687_),
    .B(_04689_),
    .C(_04691_),
    .D(_04694_),
    .Y(_05915_));
 sg13g2_inv_1 _31638_ (.Y(_05916_),
    .A(_05915_));
 sg13g2_nand2_1 _31639_ (.Y(_05917_),
    .A(_04705_),
    .B(_04708_));
 sg13g2_nand2_1 _31640_ (.Y(_05918_),
    .A(_04698_),
    .B(_04701_));
 sg13g2_nor3_2 _31641_ (.A(_05916_),
    .B(_05917_),
    .C(_05918_),
    .Y(_05919_));
 sg13g2_and2_1 _31642_ (.A(_04718_),
    .B(_04721_),
    .X(_05920_));
 sg13g2_nor2_1 _31643_ (.A(_04713_),
    .B(_04716_),
    .Y(_05921_));
 sg13g2_nand2_1 _31644_ (.Y(_05922_),
    .A(_05920_),
    .B(_05921_));
 sg13g2_nor2_1 _31645_ (.A(_04723_),
    .B(_04725_),
    .Y(_05923_));
 sg13g2_and2_1 _31646_ (.A(_04727_),
    .B(_04729_),
    .X(_05924_));
 sg13g2_and4_1 _31647_ (.A(_05920_),
    .B(_05921_),
    .C(_05923_),
    .D(_05924_),
    .X(_05925_));
 sg13g2_nand2_2 _31648_ (.Y(_05926_),
    .A(_05919_),
    .B(_05925_));
 sg13g2_nor2_1 _31649_ (.A(_04772_),
    .B(_04775_),
    .Y(_05927_));
 sg13g2_nand3_1 _31650_ (.B(_04782_),
    .C(_05927_),
    .A(_04780_),
    .Y(_05928_));
 sg13g2_nor3_2 _31651_ (.A(_05913_),
    .B(_05926_),
    .C(_05928_),
    .Y(_05929_));
 sg13g2_a21oi_1 _31652_ (.A1(\u_inv.d_next[177] ),
    .A2(\u_inv.d_reg[177] ),
    .Y(_05930_),
    .B1(_04728_));
 sg13g2_a21oi_1 _31653_ (.A1(_14196_),
    .A2(_14632_),
    .Y(_05931_),
    .B1(_05930_));
 sg13g2_a21oi_1 _31654_ (.A1(_14195_),
    .A2(_14630_),
    .Y(_05932_),
    .B1(_04724_));
 sg13g2_a221oi_1 _31655_ (.B2(_05931_),
    .C1(_05932_),
    .B1(_05923_),
    .A1(\u_inv.d_next[179] ),
    .Y(_05933_),
    .A2(\u_inv.d_reg[179] ));
 sg13g2_a21oi_1 _31656_ (.A1(_14193_),
    .A2(_14626_),
    .Y(_05934_),
    .B1(_04720_));
 sg13g2_a21oi_1 _31657_ (.A1(\u_inv.d_next[181] ),
    .A2(\u_inv.d_reg[181] ),
    .Y(_05935_),
    .B1(_04714_));
 sg13g2_a21oi_1 _31658_ (.A1(_14194_),
    .A2(_14628_),
    .Y(_05936_),
    .B1(_05935_));
 sg13g2_a221oi_1 _31659_ (.B2(_05936_),
    .C1(_05934_),
    .B1(_05920_),
    .A1(\u_inv.d_next[183] ),
    .Y(_05937_),
    .A2(\u_inv.d_reg[183] ));
 sg13g2_o21ai_1 _31660_ (.B1(_05937_),
    .Y(_05938_),
    .A1(_05922_),
    .A2(_05933_));
 sg13g2_o21ai_1 _31661_ (.B1(_04704_),
    .Y(_05939_),
    .A1(_04703_),
    .A2(_04707_));
 sg13g2_nor2b_1 _31662_ (.A(_05918_),
    .B_N(_05939_),
    .Y(_05940_));
 sg13g2_a21oi_1 _31663_ (.A1(\u_inv.d_next[187] ),
    .A2(\u_inv.d_reg[187] ),
    .Y(_05941_),
    .B1(_05940_));
 sg13g2_o21ai_1 _31664_ (.B1(_05941_),
    .Y(_05942_),
    .A1(_04697_),
    .A2(_04700_));
 sg13g2_a21oi_1 _31665_ (.A1(_14192_),
    .A2(_14620_),
    .Y(_05943_),
    .B1(_04693_));
 sg13g2_a21oi_1 _31666_ (.A1(\u_inv.d_next[189] ),
    .A2(\u_inv.d_reg[189] ),
    .Y(_05944_),
    .B1(_05943_));
 sg13g2_nor3_1 _31667_ (.A(_04687_),
    .B(_04689_),
    .C(_05944_),
    .Y(_05945_));
 sg13g2_o21ai_1 _31668_ (.B1(_04686_),
    .Y(_05946_),
    .A1(_04685_),
    .A2(_04688_));
 sg13g2_or2_1 _31669_ (.X(_05947_),
    .B(_05946_),
    .A(_05945_));
 sg13g2_a221oi_1 _31670_ (.B2(_05915_),
    .C1(_05947_),
    .B1(_05942_),
    .A1(_05919_),
    .Y(_05948_),
    .A2(_05938_));
 sg13g2_nand2_1 _31671_ (.Y(_05949_),
    .A(\u_inv.d_next[161] ),
    .B(\u_inv.d_reg[161] ));
 sg13g2_o21ai_1 _31672_ (.B1(_05949_),
    .Y(_05950_),
    .A1(_04779_),
    .A2(_04781_));
 sg13g2_o21ai_1 _31673_ (.B1(_04771_),
    .Y(_05951_),
    .A1(_04770_),
    .A2(_04773_));
 sg13g2_a21o_1 _31674_ (.A2(_05950_),
    .A1(_05927_),
    .B1(_05951_),
    .X(_05952_));
 sg13g2_a21oi_1 _31675_ (.A1(_14199_),
    .A2(_14642_),
    .Y(_05953_),
    .B1(_04766_));
 sg13g2_a22oi_1 _31676_ (.Y(_05954_),
    .B1(net5867),
    .B2(\u_inv.d_next[164] ),
    .A2(\u_inv.d_reg[165] ),
    .A1(\u_inv.d_next[165] ));
 sg13g2_inv_1 _31677_ (.Y(_05955_),
    .A(_05954_));
 sg13g2_o21ai_1 _31678_ (.B1(_05955_),
    .Y(_05956_),
    .A1(\u_inv.d_next[165] ),
    .A2(\u_inv.d_reg[165] ));
 sg13g2_nor2_1 _31679_ (.A(_05911_),
    .B(_05956_),
    .Y(_05957_));
 sg13g2_a221oi_1 _31680_ (.B2(_05952_),
    .C1(_05953_),
    .B1(_05912_),
    .A1(\u_inv.d_next[167] ),
    .Y(_05958_),
    .A2(\u_inv.d_reg[167] ));
 sg13g2_nor2b_1 _31681_ (.A(_05957_),
    .B_N(_05958_),
    .Y(_05959_));
 sg13g2_inv_1 _31682_ (.Y(_05960_),
    .A(_05959_));
 sg13g2_nor2_1 _31683_ (.A(_05910_),
    .B(_05959_),
    .Y(_05961_));
 sg13g2_a22oi_1 _31684_ (.Y(_05962_),
    .B1(\u_inv.d_reg[168] ),
    .B2(\u_inv.d_next[168] ),
    .A2(\u_inv.d_reg[169] ),
    .A1(\u_inv.d_next[169] ));
 sg13g2_inv_1 _31685_ (.Y(_05963_),
    .A(_05962_));
 sg13g2_o21ai_1 _31686_ (.B1(_05963_),
    .Y(_05964_),
    .A1(\u_inv.d_next[169] ),
    .A2(\u_inv.d_reg[169] ));
 sg13g2_nor2_1 _31687_ (.A(_04747_),
    .B(_04750_),
    .Y(_05965_));
 sg13g2_o21ai_1 _31688_ (.B1(_04748_),
    .Y(_05966_),
    .A1(_05908_),
    .A2(_05964_));
 sg13g2_nor2_1 _31689_ (.A(_05965_),
    .B(_05966_),
    .Y(_05967_));
 sg13g2_inv_1 _31690_ (.Y(_05968_),
    .A(_05967_));
 sg13g2_nor2_1 _31691_ (.A(_05907_),
    .B(_05967_),
    .Y(_05969_));
 sg13g2_a21oi_1 _31692_ (.A1(\u_inv.d_next[173] ),
    .A2(\u_inv.d_reg[173] ),
    .Y(_05970_),
    .B1(_04742_));
 sg13g2_inv_1 _31693_ (.Y(_05971_),
    .A(_05970_));
 sg13g2_o21ai_1 _31694_ (.B1(_05971_),
    .Y(_05972_),
    .A1(\u_inv.d_next[173] ),
    .A2(\u_inv.d_reg[173] ));
 sg13g2_nor3_1 _31695_ (.A(_04736_),
    .B(_04738_),
    .C(_05972_),
    .Y(_05973_));
 sg13g2_o21ai_1 _31696_ (.B1(_04735_),
    .Y(_05974_),
    .A1(_04734_),
    .A2(_04737_));
 sg13g2_nor4_1 _31697_ (.A(_05961_),
    .B(_05969_),
    .C(_05973_),
    .D(_05974_),
    .Y(_05975_));
 sg13g2_nor2_1 _31698_ (.A(_05926_),
    .B(_05975_),
    .Y(_05976_));
 sg13g2_nand2_1 _31699_ (.Y(_05977_),
    .A(_05407_),
    .B(_05410_));
 sg13g2_nor3_1 _31700_ (.A(_05416_),
    .B(_05420_),
    .C(_05977_),
    .Y(_05978_));
 sg13g2_nor2_2 _31701_ (.A(_05424_),
    .B(_05427_),
    .Y(_05979_));
 sg13g2_nand4_1 _31702_ (.B(_05434_),
    .C(_05978_),
    .A(_05432_),
    .Y(_05980_),
    .D(_05979_));
 sg13g2_nand3b_1 _31703_ (.B(_05443_),
    .C(_05444_),
    .Y(_05981_),
    .A_N(_05445_));
 sg13g2_nor3_1 _31704_ (.A(_05438_),
    .B(_05440_),
    .C(_05981_),
    .Y(_05982_));
 sg13g2_a21oi_1 _31705_ (.A1(_14216_),
    .A2(_14695_),
    .Y(_05983_),
    .B1(_05449_));
 sg13g2_nor4_1 _31706_ (.A(_05449_),
    .B(_05450_),
    .C(_05454_),
    .D(_05457_),
    .Y(_05984_));
 sg13g2_nand2_1 _31707_ (.Y(_05985_),
    .A(_05982_),
    .B(_05984_));
 sg13g2_inv_1 _31708_ (.Y(_05986_),
    .A(_05985_));
 sg13g2_nor2_1 _31709_ (.A(_05980_),
    .B(_05985_),
    .Y(_05987_));
 sg13g2_nor2_1 _31710_ (.A(_05463_),
    .B(_05465_),
    .Y(_05988_));
 sg13g2_and2_1 _31711_ (.A(_05469_),
    .B(_05470_),
    .X(_05989_));
 sg13g2_nand2_1 _31712_ (.Y(_05990_),
    .A(_05988_),
    .B(_05989_));
 sg13g2_nand2_1 _31713_ (.Y(_05991_),
    .A(_05475_),
    .B(_05477_));
 sg13g2_nand2b_1 _31714_ (.Y(_05992_),
    .B(_05480_),
    .A_N(_05482_));
 sg13g2_nor3_1 _31715_ (.A(_05990_),
    .B(_05991_),
    .C(_05992_),
    .Y(_05993_));
 sg13g2_nand2_1 _31716_ (.Y(_05994_),
    .A(_05491_),
    .B(_05492_));
 sg13g2_nor3_2 _31717_ (.A(_05487_),
    .B(_05489_),
    .C(_05994_),
    .Y(_05995_));
 sg13g2_nor4_2 _31718_ (.A(_05497_),
    .B(_05500_),
    .C(_05504_),
    .Y(_05996_),
    .D(_05508_));
 sg13g2_inv_1 _31719_ (.Y(_05997_),
    .A(_05996_));
 sg13g2_and4_1 _31720_ (.A(_05987_),
    .B(_05993_),
    .C(_05995_),
    .D(_05996_),
    .X(_05998_));
 sg13g2_and2_1 _31721_ (.A(\u_inv.d_next[113] ),
    .B(\u_inv.d_reg[113] ),
    .X(_05999_));
 sg13g2_a21oi_1 _31722_ (.A1(_05455_),
    .A2(_05456_),
    .Y(_06000_),
    .B1(_05999_));
 sg13g2_o21ai_1 _31723_ (.B1(_06000_),
    .Y(_06001_),
    .A1(_14216_),
    .A2(_14695_));
 sg13g2_a22oi_1 _31724_ (.Y(_06002_),
    .B1(_05983_),
    .B2(_06001_),
    .A2(\u_inv.d_reg[115] ),
    .A1(\u_inv.d_next[115] ));
 sg13g2_nor2b_1 _31725_ (.A(_06002_),
    .B_N(_05982_),
    .Y(_06003_));
 sg13g2_nand3_1 _31726_ (.B(\u_inv.d_reg[116] ),
    .C(_05439_),
    .A(\u_inv.d_next[116] ),
    .Y(_06004_));
 sg13g2_o21ai_1 _31727_ (.B1(_06004_),
    .Y(_06005_),
    .A1(_14215_),
    .A2(_14692_));
 sg13g2_nor2b_1 _31728_ (.A(_05981_),
    .B_N(_06005_),
    .Y(_06006_));
 sg13g2_o21ai_1 _31729_ (.B1(_05444_),
    .Y(_06007_),
    .A1(_05442_),
    .A2(_05445_));
 sg13g2_nor3_1 _31730_ (.A(_06003_),
    .B(_06006_),
    .C(_06007_),
    .Y(_06008_));
 sg13g2_nor2_1 _31731_ (.A(_05980_),
    .B(_06008_),
    .Y(_06009_));
 sg13g2_nand2_1 _31732_ (.Y(_06010_),
    .A(\u_inv.d_next[121] ),
    .B(\u_inv.d_reg[121] ));
 sg13g2_o21ai_1 _31733_ (.B1(_06010_),
    .Y(_06011_),
    .A1(_05431_),
    .A2(_05433_));
 sg13g2_a22oi_1 _31734_ (.Y(_06012_),
    .B1(_05979_),
    .B2(_06011_),
    .A2(\u_inv.d_reg[123] ),
    .A1(\u_inv.d_next[123] ));
 sg13g2_o21ai_1 _31735_ (.B1(_06012_),
    .Y(_06013_),
    .A1(_05423_),
    .A2(_05426_));
 sg13g2_and2_1 _31736_ (.A(_05978_),
    .B(_06013_),
    .X(_06014_));
 sg13g2_o21ai_1 _31737_ (.B1(_05415_),
    .Y(_06015_),
    .A1(_05414_),
    .A2(_05417_));
 sg13g2_o21ai_1 _31738_ (.B1(_05409_),
    .Y(_06016_),
    .A1(_14213_),
    .A2(_14684_));
 sg13g2_o21ai_1 _31739_ (.B1(_06016_),
    .Y(_06017_),
    .A1(\u_inv.d_next[125] ),
    .A2(\u_inv.d_reg[125] ));
 sg13g2_nor3_1 _31740_ (.A(_05416_),
    .B(_05420_),
    .C(_06017_),
    .Y(_06018_));
 sg13g2_nor4_1 _31741_ (.A(_06009_),
    .B(_06014_),
    .C(_06015_),
    .D(_06018_),
    .Y(_06019_));
 sg13g2_and2_1 _31742_ (.A(\u_inv.d_next[97] ),
    .B(\u_inv.d_reg[97] ),
    .X(_06020_));
 sg13g2_a21oi_1 _31743_ (.A1(_05505_),
    .A2(_05506_),
    .Y(_06021_),
    .B1(_06020_));
 sg13g2_o21ai_1 _31744_ (.B1(_05498_),
    .Y(_06022_),
    .A1(\u_inv.d_next[98] ),
    .A2(net5870));
 sg13g2_a21oi_1 _31745_ (.A1(_05499_),
    .A2(_06021_),
    .Y(_06023_),
    .B1(_06022_));
 sg13g2_a21o_1 _31746_ (.A2(\u_inv.d_reg[99] ),
    .A1(\u_inv.d_next[99] ),
    .B1(_06023_),
    .X(_06024_));
 sg13g2_a22oi_1 _31747_ (.Y(_06025_),
    .B1(\u_inv.d_reg[100] ),
    .B2(\u_inv.d_next[100] ),
    .A2(\u_inv.d_reg[101] ),
    .A1(\u_inv.d_next[101] ));
 sg13g2_inv_1 _31748_ (.Y(_06026_),
    .A(_06025_));
 sg13g2_o21ai_1 _31749_ (.B1(_06026_),
    .Y(_06027_),
    .A1(\u_inv.d_next[101] ),
    .A2(\u_inv.d_reg[101] ));
 sg13g2_nand2_1 _31750_ (.Y(_06028_),
    .A(_05488_),
    .B(_06027_));
 sg13g2_o21ai_1 _31751_ (.B1(_06028_),
    .Y(_06029_),
    .A1(\u_inv.d_next[102] ),
    .A2(\u_inv.d_reg[102] ));
 sg13g2_a22oi_1 _31752_ (.Y(_06030_),
    .B1(_05995_),
    .B2(_06024_),
    .A2(\u_inv.d_reg[103] ),
    .A1(\u_inv.d_next[103] ));
 sg13g2_o21ai_1 _31753_ (.B1(_06030_),
    .Y(_06031_),
    .A1(_05487_),
    .A2(_06029_));
 sg13g2_nand2_1 _31754_ (.Y(_06032_),
    .A(_05480_),
    .B(_05481_));
 sg13g2_and2_1 _31755_ (.A(\u_inv.d_next[105] ),
    .B(\u_inv.d_reg[105] ),
    .X(_06033_));
 sg13g2_a21oi_1 _31756_ (.A1(_05480_),
    .A2(_05481_),
    .Y(_06034_),
    .B1(_06033_));
 sg13g2_o21ai_1 _31757_ (.B1(_05475_),
    .Y(_06035_),
    .A1(\u_inv.d_next[106] ),
    .A2(\u_inv.d_reg[106] ));
 sg13g2_a21oi_1 _31758_ (.A1(_05476_),
    .A2(_06034_),
    .Y(_06036_),
    .B1(_06035_));
 sg13g2_a21o_2 _31759_ (.A2(\u_inv.d_reg[107] ),
    .A1(\u_inv.d_next[107] ),
    .B1(_06036_),
    .X(_06037_));
 sg13g2_nand2b_1 _31760_ (.Y(_06038_),
    .B(_06037_),
    .A_N(_05990_));
 sg13g2_o21ai_1 _31761_ (.B1(_05464_),
    .Y(_06039_),
    .A1(\u_inv.d_next[111] ),
    .A2(\u_inv.d_reg[111] ));
 sg13g2_and3_1 _31762_ (.X(_06040_),
    .A(\u_inv.d_next[108] ),
    .B(\u_inv.d_reg[108] ),
    .C(_05469_));
 sg13g2_a21oi_1 _31763_ (.A1(\u_inv.d_next[109] ),
    .A2(\u_inv.d_reg[109] ),
    .Y(_06041_),
    .B1(_06040_));
 sg13g2_nand2b_1 _31764_ (.Y(_06042_),
    .B(_05988_),
    .A_N(_06041_));
 sg13g2_nand4_1 _31765_ (.B(_06038_),
    .C(_06039_),
    .A(_05461_),
    .Y(_06043_),
    .D(_06042_));
 sg13g2_a21o_2 _31766_ (.A2(_06031_),
    .A1(_05993_),
    .B1(_06043_),
    .X(_06044_));
 sg13g2_nand2_1 _31767_ (.Y(_06045_),
    .A(_05987_),
    .B(_06044_));
 sg13g2_nand3_1 _31768_ (.B(_05995_),
    .C(_05996_),
    .A(_05993_),
    .Y(_06046_));
 sg13g2_nand2_1 _31769_ (.Y(_06047_),
    .A(_05520_),
    .B(_05522_));
 sg13g2_nor3_1 _31770_ (.A(_05515_),
    .B(_05517_),
    .C(_06047_),
    .Y(_06048_));
 sg13g2_nor4_1 _31771_ (.A(_05526_),
    .B(_05529_),
    .C(_05531_),
    .D(_05534_),
    .Y(_06049_));
 sg13g2_nand2_1 _31772_ (.Y(_06050_),
    .A(_06048_),
    .B(_06049_));
 sg13g2_nand2_1 _31773_ (.Y(_06051_),
    .A(_05546_),
    .B(_05547_));
 sg13g2_nor3_1 _31774_ (.A(_05540_),
    .B(_05544_),
    .C(_06051_),
    .Y(_06052_));
 sg13g2_nor2_1 _31775_ (.A(_05551_),
    .B(_05554_),
    .Y(_06053_));
 sg13g2_nand4_1 _31776_ (.B(_05561_),
    .C(_06052_),
    .A(net5616),
    .Y(_06054_),
    .D(_06053_));
 sg13g2_or2_1 _31777_ (.X(_06055_),
    .B(_06054_),
    .A(_06050_));
 sg13g2_nand2b_1 _31778_ (.Y(_06056_),
    .B(_05350_),
    .A_N(_05352_));
 sg13g2_nor3_1 _31779_ (.A(_05356_),
    .B(_05359_),
    .C(_06056_),
    .Y(_06057_));
 sg13g2_nor2_1 _31780_ (.A(_05370_),
    .B(_05373_),
    .Y(_06058_));
 sg13g2_and4_1 _31781_ (.A(_05365_),
    .B(_05366_),
    .C(_06057_),
    .D(_06058_),
    .X(_06059_));
 sg13g2_nor2_1 _31782_ (.A(_05385_),
    .B(_05388_),
    .Y(_06060_));
 sg13g2_and3_2 _31783_ (.X(_06061_),
    .A(_05377_),
    .B(_05380_),
    .C(_06060_));
 sg13g2_inv_1 _31784_ (.Y(_06062_),
    .A(_06061_));
 sg13g2_nand2_1 _31785_ (.Y(_06063_),
    .A(\u_inv.d_next[67] ),
    .B(\u_inv.d_reg[67] ));
 sg13g2_and2_1 _31786_ (.A(_05400_),
    .B(_05401_),
    .X(_06064_));
 sg13g2_and2_1 _31787_ (.A(\u_inv.d_next[65] ),
    .B(\u_inv.d_reg[65] ),
    .X(_06065_));
 sg13g2_nor2_1 _31788_ (.A(_06064_),
    .B(_06065_),
    .Y(_06066_));
 sg13g2_a221oi_1 _31789_ (.B2(_05401_),
    .C1(_06065_),
    .B1(_05400_),
    .A1(net5880),
    .Y(_06067_),
    .A2(\u_inv.d_reg[66] ));
 sg13g2_o21ai_1 _31790_ (.B1(_05394_),
    .Y(_06068_),
    .A1(net5880),
    .A2(\u_inv.d_reg[66] ));
 sg13g2_o21ai_1 _31791_ (.B1(_06063_),
    .Y(_06069_),
    .A1(_06067_),
    .A2(_06068_));
 sg13g2_a221oi_1 _31792_ (.B2(_05386_),
    .C1(_05383_),
    .B1(_05382_),
    .A1(net5879),
    .Y(_06070_),
    .A2(\u_inv.d_reg[70] ));
 sg13g2_o21ai_1 _31793_ (.B1(_05377_),
    .Y(_06071_),
    .A1(net5879),
    .A2(\u_inv.d_reg[70] ));
 sg13g2_nand2_1 _31794_ (.Y(_06072_),
    .A(\u_inv.d_next[71] ),
    .B(\u_inv.d_reg[71] ));
 sg13g2_o21ai_1 _31795_ (.B1(_06072_),
    .Y(_06073_),
    .A1(_06070_),
    .A2(_06071_));
 sg13g2_a21oi_1 _31796_ (.A1(_06061_),
    .A2(_06069_),
    .Y(_06074_),
    .B1(_06073_));
 sg13g2_a21o_1 _31797_ (.A2(_06069_),
    .A1(_06061_),
    .B1(_06073_),
    .X(_06075_));
 sg13g2_a22oi_1 _31798_ (.Y(_06076_),
    .B1(\u_inv.d_reg[76] ),
    .B2(\u_inv.d_next[76] ),
    .A2(net5872),
    .A1(\u_inv.d_next[77] ));
 sg13g2_inv_1 _31799_ (.Y(_06077_),
    .A(_06076_));
 sg13g2_o21ai_1 _31800_ (.B1(_06077_),
    .Y(_06078_),
    .A1(\u_inv.d_next[77] ),
    .A2(net5872));
 sg13g2_nor2_1 _31801_ (.A(_05349_),
    .B(_05351_),
    .Y(_06079_));
 sg13g2_a21oi_1 _31802_ (.A1(\u_inv.d_next[79] ),
    .A2(\u_inv.d_reg[79] ),
    .Y(_06080_),
    .B1(_06079_));
 sg13g2_o21ai_1 _31803_ (.B1(_06080_),
    .Y(_06081_),
    .A1(_06056_),
    .A2(_06078_));
 sg13g2_nand2_1 _31804_ (.Y(_06082_),
    .A(\u_inv.d_next[75] ),
    .B(\u_inv.d_reg[75] ));
 sg13g2_a22oi_1 _31805_ (.Y(_06083_),
    .B1(\u_inv.d_reg[72] ),
    .B2(net5878),
    .A2(\u_inv.d_reg[73] ),
    .A1(\u_inv.d_next[73] ));
 sg13g2_or2_1 _31806_ (.X(_06084_),
    .B(_06083_),
    .A(_05369_));
 sg13g2_nor3_1 _31807_ (.A(_05367_),
    .B(_05369_),
    .C(_06083_),
    .Y(_06085_));
 sg13g2_a21oi_1 _31808_ (.A1(net5877),
    .A2(\u_inv.d_reg[74] ),
    .Y(_06086_),
    .B1(_06085_));
 sg13g2_o21ai_1 _31809_ (.B1(_06082_),
    .Y(_06087_),
    .A1(_05364_),
    .A2(_06086_));
 sg13g2_a221oi_1 _31810_ (.B2(_06057_),
    .C1(_06081_),
    .B1(_06087_),
    .A1(_06059_),
    .Y(_06088_),
    .A2(_06075_));
 sg13g2_nor2_1 _31811_ (.A(_06055_),
    .B(_06088_),
    .Y(_06089_));
 sg13g2_nand2_1 _31812_ (.Y(_06090_),
    .A(\u_inv.d_next[91] ),
    .B(\u_inv.d_reg[91] ));
 sg13g2_nor2_1 _31813_ (.A(_05531_),
    .B(_05532_),
    .Y(_06091_));
 sg13g2_a21oi_1 _31814_ (.A1(\u_inv.d_next[89] ),
    .A2(\u_inv.d_reg[89] ),
    .Y(_06092_),
    .B1(_06091_));
 sg13g2_a221oi_1 _31815_ (.B2(\u_inv.d_next[89] ),
    .C1(_06091_),
    .B1(\u_inv.d_reg[89] ),
    .A1(\u_inv.d_next[90] ),
    .Y(_06093_),
    .A2(net5871));
 sg13g2_o21ai_1 _31816_ (.B1(_05527_),
    .Y(_06094_),
    .A1(\u_inv.d_next[90] ),
    .A2(\u_inv.d_reg[90] ));
 sg13g2_o21ai_1 _31817_ (.B1(_06090_),
    .Y(_06095_),
    .A1(_06093_),
    .A2(_06094_));
 sg13g2_nand2b_1 _31818_ (.Y(_06096_),
    .B(_05520_),
    .A_N(_05521_));
 sg13g2_nand2_1 _31819_ (.Y(_06097_),
    .A(\u_inv.d_next[93] ),
    .B(\u_inv.d_reg[93] ));
 sg13g2_and2_1 _31820_ (.A(_06096_),
    .B(_06097_),
    .X(_06098_));
 sg13g2_nor3_1 _31821_ (.A(_05515_),
    .B(_05517_),
    .C(_06098_),
    .Y(_06099_));
 sg13g2_a221oi_1 _31822_ (.B2(_06095_),
    .C1(_06099_),
    .B1(_06048_),
    .A1(\u_inv.d_next[95] ),
    .Y(_06100_),
    .A2(\u_inv.d_reg[95] ));
 sg13g2_o21ai_1 _31823_ (.B1(_06100_),
    .Y(_06101_),
    .A1(_05514_),
    .A2(_05516_));
 sg13g2_nand2_1 _31824_ (.Y(_06102_),
    .A(\u_inv.d_next[83] ),
    .B(\u_inv.d_reg[83] ));
 sg13g2_nand2_1 _31825_ (.Y(_06103_),
    .A(net5616),
    .B(_05560_));
 sg13g2_and2_1 _31826_ (.A(\u_inv.d_next[81] ),
    .B(\u_inv.d_reg[81] ),
    .X(_06104_));
 sg13g2_a21oi_1 _31827_ (.A1(net5616),
    .A2(_05560_),
    .Y(_06105_),
    .B1(_06104_));
 sg13g2_a221oi_1 _31828_ (.B2(_05560_),
    .C1(_06104_),
    .B1(net5616),
    .A1(\u_inv.d_next[82] ),
    .Y(_06106_),
    .A2(\u_inv.d_reg[82] ));
 sg13g2_or2_1 _31829_ (.X(_06107_),
    .B(_05552_),
    .A(_05551_));
 sg13g2_o21ai_1 _31830_ (.B1(_06102_),
    .Y(_06108_),
    .A1(_06106_),
    .A2(_06107_));
 sg13g2_a22oi_1 _31831_ (.Y(_06109_),
    .B1(\u_inv.d_reg[84] ),
    .B2(\u_inv.d_next[84] ),
    .A2(\u_inv.d_reg[85] ),
    .A1(\u_inv.d_next[85] ));
 sg13g2_a21oi_1 _31832_ (.A1(_14222_),
    .A2(_14724_),
    .Y(_06110_),
    .B1(_06109_));
 sg13g2_a21oi_1 _31833_ (.A1(_05543_),
    .A2(_06110_),
    .Y(_06111_),
    .B1(_05542_));
 sg13g2_a22oi_1 _31834_ (.Y(_06112_),
    .B1(_06052_),
    .B2(_06108_),
    .A2(\u_inv.d_reg[87] ),
    .A1(\u_inv.d_next[87] ));
 sg13g2_o21ai_1 _31835_ (.B1(_06112_),
    .Y(_06113_),
    .A1(_05540_),
    .A2(_06111_));
 sg13g2_nor2b_1 _31836_ (.A(_06050_),
    .B_N(_06113_),
    .Y(_06114_));
 sg13g2_nor3_2 _31837_ (.A(_06089_),
    .B(_06101_),
    .C(_06114_),
    .Y(_06115_));
 sg13g2_nand2_1 _31838_ (.Y(_06116_),
    .A(_05267_),
    .B(_05270_));
 sg13g2_nor3_1 _31839_ (.A(_05274_),
    .B(_05277_),
    .C(_06116_),
    .Y(_06117_));
 sg13g2_nor2_1 _31840_ (.A(_05286_),
    .B(_05288_),
    .Y(_06118_));
 sg13g2_nor2b_1 _31841_ (.A(_05280_),
    .B_N(_05282_),
    .Y(_06119_));
 sg13g2_nand3_1 _31842_ (.B(_06118_),
    .C(_06119_),
    .A(_06117_),
    .Y(_06120_));
 sg13g2_nand2_1 _31843_ (.Y(_06121_),
    .A(_05299_),
    .B(_05302_));
 sg13g2_nor3_1 _31844_ (.A(_05292_),
    .B(_05297_),
    .C(_06121_),
    .Y(_06122_));
 sg13g2_nand4_1 _31845_ (.B(_05296_),
    .C(_05299_),
    .A(_05293_),
    .Y(_06123_),
    .D(_05302_));
 sg13g2_and2_1 _31846_ (.A(\u_inv.d_next[49] ),
    .B(\u_inv.d_reg[49] ),
    .X(_06124_));
 sg13g2_a21oi_1 _31847_ (.A1(_05260_),
    .A2(net5617),
    .Y(_06125_),
    .B1(_06124_));
 sg13g2_o21ai_1 _31848_ (.B1(_05309_),
    .Y(_06126_),
    .A1(\u_inv.d_next[50] ),
    .A2(\u_inv.d_reg[50] ));
 sg13g2_a21oi_1 _31849_ (.A1(_05304_),
    .A2(_06125_),
    .Y(_06127_),
    .B1(_06126_));
 sg13g2_and2_1 _31850_ (.A(\u_inv.d_next[51] ),
    .B(\u_inv.d_reg[51] ),
    .X(_06128_));
 sg13g2_nor2_1 _31851_ (.A(_06127_),
    .B(_06128_),
    .Y(_06129_));
 sg13g2_o21ai_1 _31852_ (.B1(_06122_),
    .Y(_06130_),
    .A1(_06127_),
    .A2(_06128_));
 sg13g2_a22oi_1 _31853_ (.Y(_06131_),
    .B1(\u_inv.d_reg[52] ),
    .B2(\u_inv.d_next[52] ),
    .A2(\u_inv.d_reg[53] ),
    .A1(\u_inv.d_next[53] ));
 sg13g2_a21o_1 _31854_ (.A2(_14756_),
    .A1(_14230_),
    .B1(_06131_),
    .X(_06132_));
 sg13g2_nand2_1 _31855_ (.Y(_06133_),
    .A(_05294_),
    .B(_06132_));
 sg13g2_nor2b_1 _31856_ (.A(_05292_),
    .B_N(_05295_),
    .Y(_06134_));
 sg13g2_a22oi_1 _31857_ (.Y(_06135_),
    .B1(_06133_),
    .B2(_06134_),
    .A2(\u_inv.d_reg[55] ),
    .A1(\u_inv.d_next[55] ));
 sg13g2_and2_1 _31858_ (.A(_06130_),
    .B(_06135_),
    .X(_06136_));
 sg13g2_or2_1 _31859_ (.X(_06137_),
    .B(_06136_),
    .A(_06120_));
 sg13g2_nor2_1 _31860_ (.A(_05280_),
    .B(_05281_),
    .Y(_06138_));
 sg13g2_a21oi_1 _31861_ (.A1(\u_inv.d_next[57] ),
    .A2(\u_inv.d_reg[57] ),
    .Y(_06139_),
    .B1(_06138_));
 sg13g2_nand2_1 _31862_ (.Y(_06140_),
    .A(_05287_),
    .B(_06139_));
 sg13g2_a21oi_1 _31863_ (.A1(_14227_),
    .A2(_14751_),
    .Y(_06141_),
    .B1(_05286_));
 sg13g2_a22oi_1 _31864_ (.Y(_06142_),
    .B1(_06140_),
    .B2(_06141_),
    .A2(\u_inv.d_reg[59] ),
    .A1(\u_inv.d_next[59] ));
 sg13g2_nand2b_1 _31865_ (.Y(_06143_),
    .B(_06117_),
    .A_N(_06142_));
 sg13g2_a21oi_1 _31866_ (.A1(_14226_),
    .A2(_14746_),
    .Y(_06144_),
    .B1(_05269_));
 sg13g2_a21oi_1 _31867_ (.A1(\u_inv.d_next[63] ),
    .A2(\u_inv.d_reg[63] ),
    .Y(_06145_),
    .B1(_06144_));
 sg13g2_nand2_1 _31868_ (.Y(_06146_),
    .A(\u_inv.d_next[61] ),
    .B(\u_inv.d_reg[61] ));
 sg13g2_o21ai_1 _31869_ (.B1(_06146_),
    .Y(_06147_),
    .A1(_05274_),
    .A2(_05275_));
 sg13g2_nand2b_1 _31870_ (.Y(_06148_),
    .B(_06147_),
    .A_N(_06116_));
 sg13g2_nand4_1 _31871_ (.B(_06143_),
    .C(_06145_),
    .A(_06137_),
    .Y(_06149_),
    .D(_06148_));
 sg13g2_nand4_1 _31872_ (.B(_05266_),
    .C(_05305_),
    .A(_05263_),
    .Y(_06150_),
    .D(_05309_));
 sg13g2_inv_1 _31873_ (.Y(_06151_),
    .A(_06150_));
 sg13g2_nor3_2 _31874_ (.A(_06120_),
    .B(_06123_),
    .C(_06150_),
    .Y(_06152_));
 sg13g2_nor2_1 _31875_ (.A(_05175_),
    .B(_05177_),
    .Y(_06153_));
 sg13g2_nor2_1 _31876_ (.A(_05182_),
    .B(_05184_),
    .Y(_06154_));
 sg13g2_and2_1 _31877_ (.A(_06153_),
    .B(_06154_),
    .X(_06155_));
 sg13g2_nand2_1 _31878_ (.Y(_06156_),
    .A(_05188_),
    .B(_05190_));
 sg13g2_nor2b_1 _31879_ (.A(_05199_),
    .B_N(_05195_),
    .Y(_06157_));
 sg13g2_and4_1 _31880_ (.A(_05188_),
    .B(_05190_),
    .C(_06155_),
    .D(_06157_),
    .X(_06158_));
 sg13g2_nand2_1 _31881_ (.Y(_06159_),
    .A(_05211_),
    .B(_05213_));
 sg13g2_nor3_1 _31882_ (.A(_05205_),
    .B(_05208_),
    .C(_06159_),
    .Y(_06160_));
 sg13g2_nand2_1 _31883_ (.Y(_06161_),
    .A(\u_inv.d_next[35] ),
    .B(\u_inv.d_reg[35] ));
 sg13g2_and2_1 _31884_ (.A(net5618),
    .B(_05223_),
    .X(_06162_));
 sg13g2_and2_1 _31885_ (.A(\u_inv.d_next[33] ),
    .B(\u_inv.d_reg[33] ),
    .X(_06163_));
 sg13g2_nor2_1 _31886_ (.A(_06162_),
    .B(_06163_),
    .Y(_06164_));
 sg13g2_a221oi_1 _31887_ (.B2(_05223_),
    .C1(_06163_),
    .B1(net5618),
    .A1(\u_inv.d_next[34] ),
    .Y(_06165_),
    .A2(\u_inv.d_reg[34] ));
 sg13g2_a21o_1 _31888_ (.A2(_14775_),
    .A1(_14235_),
    .B1(_05218_),
    .X(_06166_));
 sg13g2_o21ai_1 _31889_ (.B1(_06161_),
    .Y(_06167_),
    .A1(_06165_),
    .A2(_06166_));
 sg13g2_a22oi_1 _31890_ (.Y(_06168_),
    .B1(\u_inv.d_reg[36] ),
    .B2(\u_inv.d_next[36] ),
    .A2(\u_inv.d_reg[37] ),
    .A1(\u_inv.d_next[37] ));
 sg13g2_nor2_1 _31891_ (.A(_05210_),
    .B(_06168_),
    .Y(_06169_));
 sg13g2_o21ai_1 _31892_ (.B1(_05206_),
    .Y(_06170_),
    .A1(_05210_),
    .A2(_06168_));
 sg13g2_nand2_1 _31893_ (.Y(_06171_),
    .A(_05207_),
    .B(_06170_));
 sg13g2_a22oi_1 _31894_ (.Y(_06172_),
    .B1(_06160_),
    .B2(_06167_),
    .A2(\u_inv.d_reg[39] ),
    .A1(\u_inv.d_next[39] ));
 sg13g2_o21ai_1 _31895_ (.B1(_06172_),
    .Y(_06173_),
    .A1(_05205_),
    .A2(_06171_));
 sg13g2_nor2_1 _31896_ (.A(_05018_),
    .B(_05020_),
    .Y(_06174_));
 sg13g2_or4_1 _31897_ (.A(_05018_),
    .B(_05020_),
    .C(_05023_),
    .D(_05025_),
    .X(_06175_));
 sg13g2_o21ai_1 _31898_ (.B1(_05032_),
    .Y(_06176_),
    .A1(\u_inv.d_next[26] ),
    .A2(\u_inv.d_reg[26] ));
 sg13g2_nand2_1 _31899_ (.Y(_06177_),
    .A(_05013_),
    .B(_05045_));
 sg13g2_nor3_1 _31900_ (.A(_05029_),
    .B(_05031_),
    .C(_06177_),
    .Y(_06178_));
 sg13g2_nand2b_2 _31901_ (.Y(_06179_),
    .B(_06178_),
    .A_N(_06175_));
 sg13g2_nor2b_1 _31902_ (.A(_05053_),
    .B_N(_05056_),
    .Y(_06180_));
 sg13g2_nand4_1 _31903_ (.B(_05049_),
    .C(_05050_),
    .A(_05048_),
    .Y(_06181_),
    .D(_06180_));
 sg13g2_nor2_1 _31904_ (.A(_05161_),
    .B(_05162_),
    .Y(_06182_));
 sg13g2_nand2_1 _31905_ (.Y(_06183_),
    .A(\u_inv.d_next[17] ),
    .B(\u_inv.d_reg[17] ));
 sg13g2_nor2b_1 _31906_ (.A(_06182_),
    .B_N(_06183_),
    .Y(_06184_));
 sg13g2_o21ai_1 _31907_ (.B1(_06183_),
    .Y(_06185_),
    .A1(_05161_),
    .A2(_05162_));
 sg13g2_and3_1 _31908_ (.X(_06186_),
    .A(\u_inv.d_next[18] ),
    .B(\u_inv.d_reg[18] ),
    .C(_05061_));
 sg13g2_nor2b_1 _31909_ (.A(_05062_),
    .B_N(_05061_),
    .Y(_06187_));
 sg13g2_a221oi_1 _31910_ (.B2(_06187_),
    .C1(_06186_),
    .B1(_06185_),
    .A1(\u_inv.d_next[19] ),
    .Y(_06188_),
    .A2(\u_inv.d_reg[19] ));
 sg13g2_a22oi_1 _31911_ (.Y(_06189_),
    .B1(\u_inv.d_reg[20] ),
    .B2(\u_inv.d_next[20] ),
    .A2(\u_inv.d_reg[21] ),
    .A1(\u_inv.d_next[21] ));
 sg13g2_a21oi_1 _31912_ (.A1(_14237_),
    .A2(_14788_),
    .Y(_06190_),
    .B1(_06189_));
 sg13g2_nand2b_1 _31913_ (.Y(_06191_),
    .B(_06190_),
    .A_N(_05051_));
 sg13g2_a21oi_1 _31914_ (.A1(_05049_),
    .A2(_06191_),
    .Y(_06192_),
    .B1(_05047_));
 sg13g2_nand2_1 _31915_ (.Y(_06193_),
    .A(\u_inv.d_next[23] ),
    .B(\u_inv.d_reg[23] ));
 sg13g2_o21ai_1 _31916_ (.B1(_06193_),
    .Y(_06194_),
    .A1(_06181_),
    .A2(_06188_));
 sg13g2_nor2_1 _31917_ (.A(_06192_),
    .B(_06194_),
    .Y(_06195_));
 sg13g2_nor2_2 _31918_ (.A(_06179_),
    .B(_06195_),
    .Y(_06196_));
 sg13g2_o21ai_1 _31919_ (.B1(_05022_),
    .Y(_06197_),
    .A1(_05021_),
    .A2(_05024_));
 sg13g2_nor2_1 _31920_ (.A(_05018_),
    .B(_05019_),
    .Y(_06198_));
 sg13g2_nand3_1 _31921_ (.B(\u_inv.d_reg[24] ),
    .C(_05011_),
    .A(\u_inv.d_next[24] ),
    .Y(_06199_));
 sg13g2_and2_1 _31922_ (.A(_05012_),
    .B(_06199_),
    .X(_06200_));
 sg13g2_a21oi_1 _31923_ (.A1(_05028_),
    .A2(_06200_),
    .Y(_06201_),
    .B1(_06176_));
 sg13g2_a21oi_1 _31924_ (.A1(\u_inv.d_next[27] ),
    .A2(\u_inv.d_reg[27] ),
    .Y(_06202_),
    .B1(_06201_));
 sg13g2_inv_1 _31925_ (.Y(_06203_),
    .A(_06202_));
 sg13g2_a22oi_1 _31926_ (.Y(_06204_),
    .B1(_06174_),
    .B2(_06197_),
    .A2(\u_inv.d_reg[31] ),
    .A1(\u_inv.d_next[31] ));
 sg13g2_o21ai_1 _31927_ (.B1(_06204_),
    .Y(_06205_),
    .A1(_06175_),
    .A2(_06202_));
 sg13g2_nor3_2 _31928_ (.A(_06196_),
    .B(_06198_),
    .C(_06205_),
    .Y(_06206_));
 sg13g2_nand2_1 _31929_ (.Y(_06207_),
    .A(\u_inv.d_next[3] ),
    .B(\u_inv.d_reg[3] ));
 sg13g2_nand2_1 _31930_ (.Y(_06208_),
    .A(\u_inv.d_next[0] ),
    .B(\u_inv.d_reg[0] ));
 sg13g2_o21ai_1 _31931_ (.B1(_05129_),
    .Y(_06209_),
    .A1(_05130_),
    .A2(_06208_));
 sg13g2_a21oi_1 _31932_ (.A1(_05127_),
    .A2(_06209_),
    .Y(_06210_),
    .B1(_05126_));
 sg13g2_o21ai_1 _31933_ (.B1(_06207_),
    .Y(_06211_),
    .A1(_05125_),
    .A2(_06210_));
 sg13g2_nand2_1 _31934_ (.Y(_06212_),
    .A(_05137_),
    .B(_06211_));
 sg13g2_nor2_1 _31935_ (.A(_05138_),
    .B(_05142_),
    .Y(_06213_));
 sg13g2_nor2_1 _31936_ (.A(_05142_),
    .B(_06212_),
    .Y(_06214_));
 sg13g2_nor2_1 _31937_ (.A(_05115_),
    .B(_05116_),
    .Y(_06215_));
 sg13g2_or2_1 _31938_ (.X(_06216_),
    .B(_05116_),
    .A(_05115_));
 sg13g2_nand4_1 _31939_ (.B(_06211_),
    .C(_06213_),
    .A(_05120_),
    .Y(_06217_),
    .D(_06216_));
 sg13g2_nand2_1 _31940_ (.Y(_06218_),
    .A(\u_inv.d_next[5] ),
    .B(\u_inv.d_reg[5] ));
 sg13g2_o21ai_1 _31941_ (.B1(_06218_),
    .Y(_06219_),
    .A1(_05136_),
    .A2(_05142_));
 sg13g2_nand2_1 _31942_ (.Y(_06220_),
    .A(_05120_),
    .B(_06219_));
 sg13g2_a21oi_1 _31943_ (.A1(_05119_),
    .A2(_06220_),
    .Y(_06221_),
    .B1(_06215_));
 sg13g2_a21oi_1 _31944_ (.A1(\u_inv.d_next[7] ),
    .A2(\u_inv.d_reg[7] ),
    .Y(_06222_),
    .B1(_06221_));
 sg13g2_nand2_1 _31945_ (.Y(_06223_),
    .A(_06217_),
    .B(_06222_));
 sg13g2_nand3_1 _31946_ (.B(_05092_),
    .C(_05093_),
    .A(_05088_),
    .Y(_06224_));
 sg13g2_nor3_1 _31947_ (.A(_05082_),
    .B(_05086_),
    .C(_06224_),
    .Y(_06225_));
 sg13g2_and2_1 _31948_ (.A(_05104_),
    .B(_05107_),
    .X(_06226_));
 sg13g2_and4_1 _31949_ (.A(_05149_),
    .B(_05151_),
    .C(_06225_),
    .D(_06226_),
    .X(_06227_));
 sg13g2_inv_1 _31950_ (.Y(_06228_),
    .A(_06227_));
 sg13g2_a21oi_2 _31951_ (.B1(_06228_),
    .Y(_06229_),
    .A2(_06222_),
    .A1(_06217_));
 sg13g2_nand2_1 _31952_ (.Y(_06230_),
    .A(\u_inv.d_next[11] ),
    .B(net5874));
 sg13g2_nand2_1 _31953_ (.Y(_06231_),
    .A(\u_inv.d_next[9] ),
    .B(\u_inv.d_reg[9] ));
 sg13g2_o21ai_1 _31954_ (.B1(_06231_),
    .Y(_06232_),
    .A1(_05148_),
    .A2(_05150_));
 sg13g2_a21oi_1 _31955_ (.A1(_05105_),
    .A2(_06232_),
    .Y(_06233_),
    .B1(_05106_));
 sg13g2_o21ai_1 _31956_ (.B1(_06230_),
    .Y(_06234_),
    .A1(_05103_),
    .A2(_06233_));
 sg13g2_nand2_1 _31957_ (.Y(_06235_),
    .A(_06225_),
    .B(_06234_));
 sg13g2_a21oi_1 _31958_ (.A1(_14240_),
    .A2(_14796_),
    .Y(_06236_),
    .B1(_05092_));
 sg13g2_a21oi_1 _31959_ (.A1(\u_inv.d_next[13] ),
    .A2(\u_inv.d_reg[13] ),
    .Y(_06237_),
    .B1(_06236_));
 sg13g2_o21ai_1 _31960_ (.B1(_05083_),
    .Y(_06238_),
    .A1(_05086_),
    .A2(_06237_));
 sg13g2_nand2b_1 _31961_ (.Y(_06239_),
    .B(_06238_),
    .A_N(_05082_));
 sg13g2_nand2_1 _31962_ (.Y(_06240_),
    .A(\u_inv.d_next[15] ),
    .B(\u_inv.d_reg[15] ));
 sg13g2_nand3_1 _31963_ (.B(_06239_),
    .C(_06240_),
    .A(_06235_),
    .Y(_06241_));
 sg13g2_nor2_1 _31964_ (.A(_06229_),
    .B(_06241_),
    .Y(_06242_));
 sg13g2_nor2_1 _31965_ (.A(_05161_),
    .B(_05164_),
    .Y(_06243_));
 sg13g2_and2_1 _31966_ (.A(_06187_),
    .B(_06243_),
    .X(_06244_));
 sg13g2_inv_1 _31967_ (.Y(_06245_),
    .A(_06244_));
 sg13g2_nor3_1 _31968_ (.A(_06179_),
    .B(_06181_),
    .C(_06245_),
    .Y(_06246_));
 sg13g2_o21ai_1 _31969_ (.B1(_06246_),
    .Y(_06247_),
    .A1(_06241_),
    .A2(_06229_));
 sg13g2_nand2_2 _31970_ (.Y(_06248_),
    .A(_06206_),
    .B(net1070));
 sg13g2_nor2_1 _31971_ (.A(_05217_),
    .B(_05218_),
    .Y(_06249_));
 sg13g2_and4_1 _31972_ (.A(_05222_),
    .B(_05224_),
    .C(_06160_),
    .D(_06249_),
    .X(_06250_));
 sg13g2_a21oi_2 _31973_ (.B1(_06173_),
    .Y(_06251_),
    .A2(_06250_),
    .A1(_06248_));
 sg13g2_o21ai_1 _31974_ (.B1(_05180_),
    .Y(_06252_),
    .A1(_05179_),
    .A2(_05183_));
 sg13g2_nor2_1 _31975_ (.A(_05175_),
    .B(_05176_),
    .Y(_06253_));
 sg13g2_a221oi_1 _31976_ (.B2(_06252_),
    .C1(_06253_),
    .B1(_06153_),
    .A1(\u_inv.d_next[47] ),
    .Y(_06254_),
    .A2(\u_inv.d_reg[47] ));
 sg13g2_a21oi_1 _31977_ (.A1(_14232_),
    .A2(_14768_),
    .Y(_06255_),
    .B1(_05189_));
 sg13g2_a21oi_1 _31978_ (.A1(\u_inv.d_next[41] ),
    .A2(\u_inv.d_reg[41] ),
    .Y(_06256_),
    .B1(_06255_));
 sg13g2_nand2_1 _31979_ (.Y(_06257_),
    .A(_05195_),
    .B(_05198_));
 sg13g2_a21oi_1 _31980_ (.A1(_05197_),
    .A2(_06256_),
    .Y(_06258_),
    .B1(_06257_));
 sg13g2_a21o_1 _31981_ (.A2(\u_inv.d_reg[43] ),
    .A1(\u_inv.d_next[43] ),
    .B1(_06258_),
    .X(_06259_));
 sg13g2_a22oi_1 _31982_ (.Y(_06260_),
    .B1(_06259_),
    .B2(_06155_),
    .A2(_06173_),
    .A1(_06158_));
 sg13g2_nand2_2 _31983_ (.Y(_06261_),
    .A(_06254_),
    .B(_06260_));
 sg13g2_and2_1 _31984_ (.A(_06158_),
    .B(_06250_),
    .X(_06262_));
 sg13g2_inv_1 _31985_ (.Y(_06263_),
    .A(_06262_));
 sg13g2_a21oi_2 _31986_ (.B1(_06263_),
    .Y(_06264_),
    .A2(net1070),
    .A1(_06206_));
 sg13g2_a21o_2 _31987_ (.A2(_06261_),
    .A1(_06152_),
    .B1(_06149_),
    .X(_06265_));
 sg13g2_nand2_1 _31988_ (.Y(_06266_),
    .A(_06152_),
    .B(_06262_));
 sg13g2_a21oi_2 _31989_ (.B1(_06266_),
    .Y(_06267_),
    .A2(net1070),
    .A1(_06206_));
 sg13g2_or2_1 _31990_ (.X(_06268_),
    .B(_06267_),
    .A(_06265_));
 sg13g2_and4_1 _31991_ (.A(_05394_),
    .B(_05395_),
    .C(_05400_),
    .D(_05402_),
    .X(_06269_));
 sg13g2_nand3_1 _31992_ (.B(_06061_),
    .C(_06269_),
    .A(_06059_),
    .Y(_06270_));
 sg13g2_nor2_1 _31993_ (.A(_06055_),
    .B(_06270_),
    .Y(_06271_));
 sg13g2_o21ai_1 _31994_ (.B1(_06271_),
    .Y(_06272_),
    .A1(_06265_),
    .A2(_06267_));
 sg13g2_and3_1 _31995_ (.X(_06273_),
    .A(_06059_),
    .B(_06061_),
    .C(_06269_));
 sg13g2_nand2b_2 _31996_ (.Y(_06274_),
    .B(_05998_),
    .A_N(_06115_));
 sg13g2_and3_2 _31997_ (.X(_06275_),
    .A(_06019_),
    .B(_06045_),
    .C(_06274_));
 sg13g2_and2_1 _31998_ (.A(_05998_),
    .B(_06271_),
    .X(_06276_));
 sg13g2_o21ai_1 _31999_ (.B1(_06276_),
    .Y(_06277_),
    .A1(_06265_),
    .A2(_06267_));
 sg13g2_nand2_1 _32000_ (.Y(_06278_),
    .A(_06275_),
    .B(_06277_));
 sg13g2_nand2_1 _32001_ (.Y(_06279_),
    .A(_04790_),
    .B(_04793_));
 sg13g2_nand2_1 _32002_ (.Y(_06280_),
    .A(_04796_),
    .B(_04797_));
 sg13g2_nor2_1 _32003_ (.A(_06279_),
    .B(_06280_),
    .Y(_06281_));
 sg13g2_nor2_1 _32004_ (.A(_04801_),
    .B(_04803_),
    .Y(_06282_));
 sg13g2_nand2_1 _32005_ (.Y(_06283_),
    .A(_04806_),
    .B(_04807_));
 sg13g2_and4_1 _32006_ (.A(_04806_),
    .B(_04807_),
    .C(_06281_),
    .D(_06282_),
    .X(_06284_));
 sg13g2_and2_1 _32007_ (.A(_04817_),
    .B(_04820_),
    .X(_06285_));
 sg13g2_and2_1 _32008_ (.A(_04829_),
    .B(_04831_),
    .X(_06286_));
 sg13g2_nand2_1 _32009_ (.Y(_06287_),
    .A(_04824_),
    .B(_04826_));
 sg13g2_nand3_1 _32010_ (.B(_04826_),
    .C(_06285_),
    .A(_04824_),
    .Y(_06288_));
 sg13g2_nand3_1 _32011_ (.B(_04814_),
    .C(_06286_),
    .A(_04811_),
    .Y(_06289_));
 sg13g2_nor2_1 _32012_ (.A(_06288_),
    .B(_06289_),
    .Y(_06290_));
 sg13g2_nand2_2 _32013_ (.Y(_06291_),
    .A(_06284_),
    .B(_06290_));
 sg13g2_nand2_1 _32014_ (.Y(_06292_),
    .A(_04845_),
    .B(_04848_));
 sg13g2_or2_1 _32015_ (.X(_06293_),
    .B(_04841_),
    .A(_04839_));
 sg13g2_nor2_1 _32016_ (.A(_06292_),
    .B(_06293_),
    .Y(_06294_));
 sg13g2_nor2_1 _32017_ (.A(_04906_),
    .B(_04910_),
    .Y(_06295_));
 sg13g2_and2_1 _32018_ (.A(_04850_),
    .B(_04852_),
    .X(_06296_));
 sg13g2_nand3_1 _32019_ (.B(_06295_),
    .C(_06296_),
    .A(_06294_),
    .Y(_06297_));
 sg13g2_nor2_1 _32020_ (.A(_04870_),
    .B(_04873_),
    .Y(_06298_));
 sg13g2_nand3_1 _32021_ (.B(_04878_),
    .C(_06298_),
    .A(_04876_),
    .Y(_06299_));
 sg13g2_nor2_1 _32022_ (.A(net5619),
    .B(_04884_),
    .Y(_06300_));
 sg13g2_nor4_1 _32023_ (.A(_04882_),
    .B(_04884_),
    .C(_05692_),
    .D(_05696_),
    .Y(_06301_));
 sg13g2_nand2b_2 _32024_ (.Y(_06302_),
    .B(_06301_),
    .A_N(_06299_));
 sg13g2_nor3_1 _32025_ (.A(_06291_),
    .B(_06297_),
    .C(_06302_),
    .Y(_06303_));
 sg13g2_inv_1 _32026_ (.Y(_06304_),
    .A(_06303_));
 sg13g2_a21o_2 _32027_ (.A2(_06277_),
    .A1(_06275_),
    .B1(_06304_),
    .X(_06305_));
 sg13g2_nor2_1 _32028_ (.A(_05692_),
    .B(_05694_),
    .Y(_06306_));
 sg13g2_nand2_1 _32029_ (.Y(_06307_),
    .A(\u_inv.d_next[129] ),
    .B(\u_inv.d_reg[129] ));
 sg13g2_nor2b_1 _32030_ (.A(_06306_),
    .B_N(_06307_),
    .Y(_06308_));
 sg13g2_o21ai_1 _32031_ (.B1(_06307_),
    .Y(_06309_),
    .A1(_05692_),
    .A2(_05694_));
 sg13g2_nor2_1 _32032_ (.A(net5619),
    .B(_04883_),
    .Y(_06310_));
 sg13g2_a221oi_1 _32033_ (.B2(_06309_),
    .C1(_06310_),
    .B1(_06300_),
    .A1(\u_inv.d_next[131] ),
    .Y(_06311_),
    .A2(\u_inv.d_reg[131] ));
 sg13g2_nor2_1 _32034_ (.A(_04875_),
    .B(_04877_),
    .Y(_06312_));
 sg13g2_a21oi_1 _32035_ (.A1(\u_inv.d_next[133] ),
    .A2(\u_inv.d_reg[133] ),
    .Y(_06313_),
    .B1(_06312_));
 sg13g2_a21o_1 _32036_ (.A2(\u_inv.d_reg[133] ),
    .A1(\u_inv.d_next[133] ),
    .B1(_06312_),
    .X(_06314_));
 sg13g2_a21oi_1 _32037_ (.A1(_14210_),
    .A2(_14674_),
    .Y(_06315_),
    .B1(_04871_));
 sg13g2_a221oi_1 _32038_ (.B2(_06314_),
    .C1(_06315_),
    .B1(_06298_),
    .A1(\u_inv.d_next[135] ),
    .Y(_06316_),
    .A2(\u_inv.d_reg[135] ));
 sg13g2_o21ai_1 _32039_ (.B1(_06316_),
    .Y(_06317_),
    .A1(_06299_),
    .A2(_06311_));
 sg13g2_nor2b_1 _32040_ (.A(_06297_),
    .B_N(_06317_),
    .Y(_06318_));
 sg13g2_a22oi_1 _32041_ (.Y(_06319_),
    .B1(net5869),
    .B2(\u_inv.d_next[140] ),
    .A2(\u_inv.d_reg[141] ),
    .A1(\u_inv.d_next[141] ));
 sg13g2_a21oi_1 _32042_ (.A1(_14207_),
    .A2(_14668_),
    .Y(_06320_),
    .B1(_06319_));
 sg13g2_nor2b_1 _32043_ (.A(_06292_),
    .B_N(_06320_),
    .Y(_06321_));
 sg13g2_o21ai_1 _32044_ (.B1(_04844_),
    .Y(_06322_),
    .A1(_04843_),
    .A2(_04847_));
 sg13g2_nand2_1 _32045_ (.Y(_06323_),
    .A(\u_inv.d_next[137] ),
    .B(\u_inv.d_reg[137] ));
 sg13g2_o21ai_1 _32046_ (.B1(_06323_),
    .Y(_06324_),
    .A1(_04906_),
    .A2(_04908_));
 sg13g2_o21ai_1 _32047_ (.B1(_04851_),
    .Y(_06325_),
    .A1(\u_inv.d_next[139] ),
    .A2(\u_inv.d_reg[139] ));
 sg13g2_o21ai_1 _32048_ (.B1(_06325_),
    .Y(_06326_),
    .A1(_14208_),
    .A2(_14670_));
 sg13g2_a21oi_1 _32049_ (.A1(_06296_),
    .A2(_06324_),
    .Y(_06327_),
    .B1(_06326_));
 sg13g2_nor2b_1 _32050_ (.A(_06327_),
    .B_N(_06294_),
    .Y(_06328_));
 sg13g2_nor4_2 _32051_ (.A(_06318_),
    .B(_06321_),
    .C(_06322_),
    .Y(_06329_),
    .D(_06328_));
 sg13g2_a22oi_1 _32052_ (.Y(_06330_),
    .B1(\u_inv.d_reg[148] ),
    .B2(\u_inv.d_next[148] ),
    .A2(\u_inv.d_reg[149] ),
    .A1(\u_inv.d_next[149] ));
 sg13g2_a21oi_1 _32053_ (.A1(_14203_),
    .A2(_14660_),
    .Y(_06331_),
    .B1(_06330_));
 sg13g2_a22oi_1 _32054_ (.Y(_06332_),
    .B1(\u_inv.d_reg[146] ),
    .B2(\u_inv.d_next[146] ),
    .A2(\u_inv.d_reg[147] ),
    .A1(\u_inv.d_next[147] ));
 sg13g2_a21oi_1 _32055_ (.A1(_14204_),
    .A2(_14662_),
    .Y(_06333_),
    .B1(_06332_));
 sg13g2_inv_1 _32056_ (.Y(_06334_),
    .A(_06333_));
 sg13g2_nor2_1 _32057_ (.A(_04828_),
    .B(_04830_),
    .Y(_06335_));
 sg13g2_a21oi_1 _32058_ (.A1(net5876),
    .A2(\u_inv.d_reg[145] ),
    .Y(_06336_),
    .B1(_06335_));
 sg13g2_a21oi_1 _32059_ (.A1(_06285_),
    .A2(_06333_),
    .Y(_06337_),
    .B1(_06331_));
 sg13g2_o21ai_1 _32060_ (.B1(_06337_),
    .Y(_06338_),
    .A1(_06288_),
    .A2(_06336_));
 sg13g2_nand3_1 _32061_ (.B(_04814_),
    .C(_06338_),
    .A(_04811_),
    .Y(_06339_));
 sg13g2_a22oi_1 _32062_ (.Y(_06340_),
    .B1(\u_inv.d_reg[150] ),
    .B2(\u_inv.d_next[150] ),
    .A2(\u_inv.d_reg[151] ),
    .A1(\u_inv.d_next[151] ));
 sg13g2_o21ai_1 _32063_ (.B1(_06339_),
    .Y(_06341_),
    .A1(_04810_),
    .A2(_06340_));
 sg13g2_a22oi_1 _32064_ (.Y(_06342_),
    .B1(\u_inv.d_reg[152] ),
    .B2(\u_inv.d_next[152] ),
    .A2(\u_inv.d_reg[153] ),
    .A1(\u_inv.d_next[153] ));
 sg13g2_a21oi_1 _32065_ (.A1(_14202_),
    .A2(_14656_),
    .Y(_06343_),
    .B1(_06342_));
 sg13g2_inv_1 _32066_ (.Y(_06344_),
    .A(_06343_));
 sg13g2_o21ai_1 _32067_ (.B1(_04802_),
    .Y(_06345_),
    .A1(\u_inv.d_next[155] ),
    .A2(\u_inv.d_reg[155] ));
 sg13g2_o21ai_1 _32068_ (.B1(_06345_),
    .Y(_06346_),
    .A1(_14201_),
    .A2(_14654_));
 sg13g2_a21o_1 _32069_ (.A2(_06343_),
    .A1(_06282_),
    .B1(_06346_),
    .X(_06347_));
 sg13g2_a21oi_1 _32070_ (.A1(_14200_),
    .A2(_14650_),
    .Y(_06348_),
    .B1(_04792_));
 sg13g2_a21oi_1 _32071_ (.A1(\u_inv.d_next[159] ),
    .A2(\u_inv.d_reg[159] ),
    .Y(_06349_),
    .B1(_06348_));
 sg13g2_a22oi_1 _32072_ (.Y(_06350_),
    .B1(\u_inv.d_reg[156] ),
    .B2(\u_inv.d_next[156] ),
    .A2(\u_inv.d_reg[157] ),
    .A1(\u_inv.d_next[157] ));
 sg13g2_inv_1 _32073_ (.Y(_06351_),
    .A(_06350_));
 sg13g2_o21ai_1 _32074_ (.B1(_06351_),
    .Y(_06352_),
    .A1(\u_inv.d_next[157] ),
    .A2(\u_inv.d_reg[157] ));
 sg13g2_o21ai_1 _32075_ (.B1(_06349_),
    .Y(_06353_),
    .A1(_06279_),
    .A2(_06352_));
 sg13g2_a221oi_1 _32076_ (.B2(_06281_),
    .C1(_06353_),
    .B1(_06347_),
    .A1(_06284_),
    .Y(_06354_),
    .A2(_06341_));
 sg13g2_o21ai_1 _32077_ (.B1(_06354_),
    .Y(_06355_),
    .A1(_06291_),
    .A2(_06329_));
 sg13g2_inv_1 _32078_ (.Y(_06356_),
    .A(_06355_));
 sg13g2_a21oi_2 _32079_ (.B1(_05976_),
    .Y(_06357_),
    .A2(_06355_),
    .A1(_05929_));
 sg13g2_nand2_2 _32080_ (.Y(_06358_),
    .A(_05948_),
    .B(_06357_));
 sg13g2_and2_1 _32081_ (.A(_05929_),
    .B(_06303_),
    .X(_06359_));
 sg13g2_inv_1 _32082_ (.Y(_06360_),
    .A(_06359_));
 sg13g2_a21oi_2 _32083_ (.B1(_06360_),
    .Y(_06361_),
    .A2(_06277_),
    .A1(_06275_));
 sg13g2_nor2_2 _32084_ (.A(_06358_),
    .B(_06361_),
    .Y(_06362_));
 sg13g2_nor2_1 _32085_ (.A(_04584_),
    .B(_04587_),
    .Y(_06363_));
 sg13g2_inv_1 _32086_ (.Y(_06364_),
    .A(_06363_));
 sg13g2_nand3b_1 _32087_ (.B(_04580_),
    .C(_06363_),
    .Y(_06365_),
    .A_N(_04578_));
 sg13g2_nor2_1 _32088_ (.A(_04592_),
    .B(_04595_),
    .Y(_06366_));
 sg13g2_nand2_1 _32089_ (.Y(_06367_),
    .A(_04599_),
    .B(_04601_));
 sg13g2_nor4_2 _32090_ (.A(_04592_),
    .B(_04595_),
    .C(_06365_),
    .Y(_06368_),
    .D(_06367_));
 sg13g2_nor2_1 _32091_ (.A(_04614_),
    .B(_04617_),
    .Y(_06369_));
 sg13g2_nor2_1 _32092_ (.A(_04622_),
    .B(_04624_),
    .Y(_06370_));
 sg13g2_or2_1 _32093_ (.X(_06371_),
    .B(_04624_),
    .A(_04622_));
 sg13g2_nor2_1 _32094_ (.A(_04607_),
    .B(_04610_),
    .Y(_06372_));
 sg13g2_nand2_1 _32095_ (.Y(_06373_),
    .A(_06369_),
    .B(_06372_));
 sg13g2_nor3_1 _32096_ (.A(_04627_),
    .B(_06371_),
    .C(_06373_),
    .Y(_06374_));
 sg13g2_nand3_1 _32097_ (.B(_06368_),
    .C(_06374_),
    .A(_04628_),
    .Y(_06375_));
 sg13g2_and2_1 _32098_ (.A(_04633_),
    .B(_04636_),
    .X(_06376_));
 sg13g2_nor2_1 _32099_ (.A(_04640_),
    .B(_04642_),
    .Y(_06377_));
 sg13g2_and2_1 _32100_ (.A(_06376_),
    .B(_06377_),
    .X(_06378_));
 sg13g2_nor2_2 _32101_ (.A(_04646_),
    .B(_04648_),
    .Y(_06379_));
 sg13g2_inv_1 _32102_ (.Y(_06380_),
    .A(_06379_));
 sg13g2_and2_1 _32103_ (.A(_04652_),
    .B(_04655_),
    .X(_06381_));
 sg13g2_nand3_1 _32104_ (.B(_06379_),
    .C(_06381_),
    .A(_06378_),
    .Y(_06382_));
 sg13g2_and2_1 _32105_ (.A(_04666_),
    .B(_04669_),
    .X(_06383_));
 sg13g2_nor2_1 _32106_ (.A(_04661_),
    .B(_04663_),
    .Y(_06384_));
 sg13g2_nand2_2 _32107_ (.Y(_06385_),
    .A(_06383_),
    .B(_06384_));
 sg13g2_nor2_1 _32108_ (.A(_04675_),
    .B(_04677_),
    .Y(_06386_));
 sg13g2_nor2_1 _32109_ (.A(_04671_),
    .B(_04673_),
    .Y(_06387_));
 sg13g2_nand2_2 _32110_ (.Y(_06388_),
    .A(_06386_),
    .B(_06387_));
 sg13g2_nor3_1 _32111_ (.A(_06382_),
    .B(_06385_),
    .C(_06388_),
    .Y(_06389_));
 sg13g2_nor2b_1 _32112_ (.A(_06375_),
    .B_N(_06389_),
    .Y(_06390_));
 sg13g2_o21ai_1 _32113_ (.B1(_06390_),
    .Y(_06391_),
    .A1(_06361_),
    .A2(_06358_));
 sg13g2_a22oi_1 _32114_ (.Y(_06392_),
    .B1(\u_inv.d_reg[214] ),
    .B2(\u_inv.d_next[214] ),
    .A2(\u_inv.d_reg[215] ),
    .A1(\u_inv.d_next[215] ));
 sg13g2_a21oi_1 _32115_ (.A1(\u_inv.d_next[213] ),
    .A2(\u_inv.d_reg[213] ),
    .Y(_06393_),
    .B1(_04608_));
 sg13g2_a21oi_1 _32116_ (.A1(_14183_),
    .A2(_14596_),
    .Y(_06394_),
    .B1(_06393_));
 sg13g2_a22oi_1 _32117_ (.Y(_06395_),
    .B1(\u_inv.d_reg[208] ),
    .B2(\u_inv.d_next[208] ),
    .A2(\u_inv.d_reg[209] ),
    .A1(\u_inv.d_next[209] ));
 sg13g2_a21oi_1 _32118_ (.A1(_14184_),
    .A2(_14600_),
    .Y(_06396_),
    .B1(_06395_));
 sg13g2_a21oi_1 _32119_ (.A1(_04620_),
    .A2(_04623_),
    .Y(_06397_),
    .B1(_04621_));
 sg13g2_inv_1 _32120_ (.Y(_06398_),
    .A(_06397_));
 sg13g2_a21oi_1 _32121_ (.A1(_06370_),
    .A2(_06396_),
    .Y(_06399_),
    .B1(_06397_));
 sg13g2_nor2_1 _32122_ (.A(_06373_),
    .B(_06399_),
    .Y(_06400_));
 sg13g2_a21oi_1 _32123_ (.A1(_06369_),
    .A2(_06394_),
    .Y(_06401_),
    .B1(_06400_));
 sg13g2_o21ai_1 _32124_ (.B1(_06401_),
    .Y(_06402_),
    .A1(_04615_),
    .A2(_06392_));
 sg13g2_nand2_1 _32125_ (.Y(_06403_),
    .A(_06368_),
    .B(_06402_));
 sg13g2_o21ai_1 _32126_ (.B1(_04598_),
    .Y(_06404_),
    .A1(_04597_),
    .A2(_04600_));
 sg13g2_a22oi_1 _32127_ (.Y(_06405_),
    .B1(_06366_),
    .B2(_06404_),
    .A2(\u_inv.d_reg[219] ),
    .A1(\u_inv.d_next[219] ));
 sg13g2_o21ai_1 _32128_ (.B1(_06405_),
    .Y(_06406_),
    .A1(_04590_),
    .A2(_04593_));
 sg13g2_nand2b_1 _32129_ (.Y(_06407_),
    .B(_06406_),
    .A_N(_06365_));
 sg13g2_o21ai_1 _32130_ (.B1(_04579_),
    .Y(_06408_),
    .A1(\u_inv.d_next[223] ),
    .A2(\u_inv.d_reg[223] ));
 sg13g2_a21oi_1 _32131_ (.A1(_14181_),
    .A2(_14588_),
    .Y(_06409_),
    .B1(_04585_));
 sg13g2_a21oi_1 _32132_ (.A1(\u_inv.d_next[221] ),
    .A2(\u_inv.d_reg[221] ),
    .Y(_06410_),
    .B1(_06409_));
 sg13g2_nor3_1 _32133_ (.A(_04578_),
    .B(_04581_),
    .C(_06410_),
    .Y(_06411_));
 sg13g2_or2_1 _32134_ (.X(_06412_),
    .B(_04672_),
    .A(_04671_));
 sg13g2_nand2_1 _32135_ (.Y(_06413_),
    .A(\u_inv.d_next[193] ),
    .B(\u_inv.d_reg[193] ));
 sg13g2_and2_1 _32136_ (.A(_06412_),
    .B(_06413_),
    .X(_06414_));
 sg13g2_nand2_1 _32137_ (.Y(_06415_),
    .A(_06412_),
    .B(_06413_));
 sg13g2_a21oi_1 _32138_ (.A1(_14189_),
    .A2(_14614_),
    .Y(_06416_),
    .B1(_04676_));
 sg13g2_a221oi_1 _32139_ (.B2(_06415_),
    .C1(_06416_),
    .B1(_06386_),
    .A1(\u_inv.d_next[195] ),
    .Y(_06417_),
    .A2(\u_inv.d_reg[195] ));
 sg13g2_o21ai_1 _32140_ (.B1(_04660_),
    .Y(_06418_),
    .A1(_04659_),
    .A2(_04662_));
 sg13g2_a21oi_1 _32141_ (.A1(_14188_),
    .A2(_14610_),
    .Y(_06419_),
    .B1(_04668_));
 sg13g2_a221oi_1 _32142_ (.B2(_06418_),
    .C1(_06419_),
    .B1(_06383_),
    .A1(\u_inv.d_next[199] ),
    .Y(_06420_),
    .A2(\u_inv.d_reg[199] ));
 sg13g2_o21ai_1 _32143_ (.B1(_06420_),
    .Y(_06421_),
    .A1(_06385_),
    .A2(_06417_));
 sg13g2_o21ai_1 _32144_ (.B1(_04651_),
    .Y(_06422_),
    .A1(_04650_),
    .A2(_04654_));
 sg13g2_a21oi_1 _32145_ (.A1(_14187_),
    .A2(_14606_),
    .Y(_06423_),
    .B1(_04647_));
 sg13g2_a221oi_1 _32146_ (.B2(_06422_),
    .C1(_06423_),
    .B1(_06379_),
    .A1(\u_inv.d_next[203] ),
    .Y(_06424_),
    .A2(\u_inv.d_reg[203] ));
 sg13g2_nand2b_1 _32147_ (.Y(_06425_),
    .B(_06378_),
    .A_N(_06424_));
 sg13g2_nand2_1 _32148_ (.Y(_06426_),
    .A(_04638_),
    .B(_04641_));
 sg13g2_nand2_1 _32149_ (.Y(_06427_),
    .A(_04639_),
    .B(_06426_));
 sg13g2_a21oi_1 _32150_ (.A1(_14185_),
    .A2(_14602_),
    .Y(_06428_),
    .B1(_04635_));
 sg13g2_a21oi_1 _32151_ (.A1(\u_inv.d_next[207] ),
    .A2(\u_inv.d_reg[207] ),
    .Y(_06429_),
    .B1(_06428_));
 sg13g2_nand4_1 _32152_ (.B(_06379_),
    .C(_06381_),
    .A(_06378_),
    .Y(_06430_),
    .D(_06421_));
 sg13g2_nand3_1 _32153_ (.B(_06429_),
    .C(_06430_),
    .A(_06425_),
    .Y(_06431_));
 sg13g2_a21oi_2 _32154_ (.B1(_06431_),
    .Y(_06432_),
    .A2(_06427_),
    .A1(_06376_));
 sg13g2_nor2_2 _32155_ (.A(_06375_),
    .B(_06432_),
    .Y(_06433_));
 sg13g2_nand4_1 _32156_ (.B(_06403_),
    .C(_06407_),
    .A(_04577_),
    .Y(_06434_),
    .D(_06408_));
 sg13g2_nor3_2 _32157_ (.A(_06411_),
    .B(_06433_),
    .C(_06434_),
    .Y(_06435_));
 sg13g2_and2_1 _32158_ (.A(_05905_),
    .B(_06435_),
    .X(_06436_));
 sg13g2_a22oi_1 _32159_ (.Y(_06437_),
    .B1(_06391_),
    .B2(_06436_),
    .A2(_05905_),
    .A1(_05867_));
 sg13g2_nand3_1 _32160_ (.B(_04449_),
    .C(_06437_),
    .A(net5720),
    .Y(_06438_));
 sg13g2_o21ai_1 _32161_ (.B1(net5020),
    .Y(_06439_),
    .A1(net5720),
    .A2(\u_inv.d_next[256] ));
 sg13g2_a21oi_1 _32162_ (.A1(_14172_),
    .A2(_14553_),
    .Y(_06440_),
    .B1(_06439_));
 sg13g2_and2_1 _32163_ (.A(_06438_),
    .B(_06440_),
    .X(_06441_));
 sg13g2_a21oi_1 _32164_ (.A1(_05834_),
    .A2(_05835_),
    .Y(_06442_),
    .B1(_06441_));
 sg13g2_a21o_2 _32165_ (.A2(_05835_),
    .A1(_05834_),
    .B1(_06441_),
    .X(_06443_));
 sg13g2_nand2_1 _32166_ (.Y(_06444_),
    .A(\u_inv.d_reg[0] ),
    .B(net4924));
 sg13g2_xnor2_1 _32167_ (.Y(_06445_),
    .A(_05130_),
    .B(_06208_));
 sg13g2_nand2_1 _32168_ (.Y(_06446_),
    .A(net5720),
    .B(_06445_));
 sg13g2_o21ai_1 _32169_ (.B1(_06446_),
    .Y(_06447_),
    .A1(net5721),
    .A2(\u_inv.d_next[1] ));
 sg13g2_xnor2_1 _32170_ (.Y(_06448_),
    .A(_06444_),
    .B(_06447_));
 sg13g2_nand2_1 _32171_ (.Y(_06449_),
    .A(net5720),
    .B(\u_inv.d_reg[0] ));
 sg13g2_xnor2_1 _32172_ (.Y(_06450_),
    .A(\u_inv.d_next[0] ),
    .B(_06449_));
 sg13g2_xnor2_1 _32173_ (.Y(_06451_),
    .A(_14242_),
    .B(_06449_));
 sg13g2_nor2_1 _32174_ (.A(_06448_),
    .B(net5349),
    .Y(_06452_));
 sg13g2_nand2_1 _32175_ (.Y(_06453_),
    .A(net4791),
    .B(net5391));
 sg13g2_nand2_1 _32176_ (.Y(_06454_),
    .A(net4791),
    .B(_06452_));
 sg13g2_xor2_1 _32177_ (.B(_06453_),
    .A(_06448_),
    .X(_06455_));
 sg13g2_xnor2_1 _32178_ (.Y(_06456_),
    .A(_06448_),
    .B(_06453_));
 sg13g2_xnor2_1 _32179_ (.Y(_06457_),
    .A(_05127_),
    .B(_06209_));
 sg13g2_nand2_1 _32180_ (.Y(_06458_),
    .A(net5721),
    .B(_06457_));
 sg13g2_o21ai_1 _32181_ (.B1(_06458_),
    .Y(_06459_),
    .A1(net5720),
    .A2(\u_inv.d_next[2] ));
 sg13g2_xnor2_1 _32182_ (.Y(_06460_),
    .A(_05127_),
    .B(_05132_));
 sg13g2_mux2_1 _32183_ (.A0(_06460_),
    .A1(_06459_),
    .S(net5020),
    .X(_06461_));
 sg13g2_inv_1 _32184_ (.Y(_06462_),
    .A(_06461_));
 sg13g2_xnor2_1 _32185_ (.Y(_06463_),
    .A(_06454_),
    .B(_06462_));
 sg13g2_inv_1 _32186_ (.Y(_06464_),
    .A(_06463_));
 sg13g2_a21oi_1 _32187_ (.A1(_19007_),
    .A2(_06463_),
    .Y(_06465_),
    .B1(net4691));
 sg13g2_a221oi_1 _32188_ (.B2(net4691),
    .C1(_06465_),
    .B1(_19007_),
    .A1(_18919_),
    .Y(_06466_),
    .A2(_19003_));
 sg13g2_a21oi_2 _32189_ (.B1(_04682_),
    .Y(_06467_),
    .A2(_05702_),
    .A1(_05009_));
 sg13g2_nor2_1 _32190_ (.A(_05802_),
    .B(_06467_),
    .Y(_06468_));
 sg13g2_o21ai_1 _32191_ (.B1(_04575_),
    .Y(_06469_),
    .A1(_05802_),
    .A2(_06467_));
 sg13g2_a21oi_2 _32192_ (.B1(_04513_),
    .Y(_06470_),
    .A2(_06469_),
    .A1(_05738_));
 sg13g2_o21ai_1 _32193_ (.B1(_04478_),
    .Y(_06471_),
    .A1(_05817_),
    .A2(_06470_));
 sg13g2_o21ai_1 _32194_ (.B1(_04479_),
    .Y(_06472_),
    .A1(_05817_),
    .A2(_06470_));
 sg13g2_o21ai_1 _32195_ (.B1(_04481_),
    .Y(_06473_),
    .A1(_05817_),
    .A2(_06470_));
 sg13g2_nand2_1 _32196_ (.Y(_06474_),
    .A(_05824_),
    .B(_06473_));
 sg13g2_a21oi_1 _32197_ (.A1(_05824_),
    .A2(_06473_),
    .Y(_06475_),
    .B1(_04465_));
 sg13g2_nor3_1 _32198_ (.A(_04456_),
    .B(_05827_),
    .C(_06475_),
    .Y(_06476_));
 sg13g2_o21ai_1 _32199_ (.B1(_04456_),
    .Y(_06477_),
    .A1(_05827_),
    .A2(_06475_));
 sg13g2_nor2b_1 _32200_ (.A(_06476_),
    .B_N(_06477_),
    .Y(_06478_));
 sg13g2_nand2_1 _32201_ (.Y(_06479_),
    .A(_06391_),
    .B(_06435_));
 sg13g2_a21oi_2 _32202_ (.B1(_05866_),
    .Y(_06480_),
    .A2(_06435_),
    .A1(_06391_));
 sg13g2_o21ai_1 _32203_ (.B1(_05849_),
    .Y(_06481_),
    .A1(_05904_),
    .A2(_06480_));
 sg13g2_nand2_1 _32204_ (.Y(_06482_),
    .A(_05878_),
    .B(_06481_));
 sg13g2_a21oi_1 _32205_ (.A1(_05878_),
    .A2(_06481_),
    .Y(_06483_),
    .B1(_05840_));
 sg13g2_nor2_1 _32206_ (.A(_05879_),
    .B(_06483_),
    .Y(_06484_));
 sg13g2_a21oi_1 _32207_ (.A1(_05839_),
    .A2(_06483_),
    .Y(_06485_),
    .B1(_05881_));
 sg13g2_nor2_1 _32208_ (.A(_05837_),
    .B(_06485_),
    .Y(_06486_));
 sg13g2_nor3_1 _32209_ (.A(_04455_),
    .B(_05882_),
    .C(_06486_),
    .Y(_06487_));
 sg13g2_o21ai_1 _32210_ (.B1(_04455_),
    .Y(_06488_),
    .A1(_05882_),
    .A2(_06486_));
 sg13g2_nand2_1 _32211_ (.Y(_06489_),
    .A(net5720),
    .B(_06488_));
 sg13g2_a21oi_1 _32212_ (.A1(net5654),
    .A2(\u_inv.d_next[254] ),
    .Y(_06490_),
    .B1(net4924));
 sg13g2_o21ai_1 _32213_ (.B1(_06490_),
    .Y(_06491_),
    .A1(_06487_),
    .A2(_06489_));
 sg13g2_o21ai_1 _32214_ (.B1(_06491_),
    .Y(_06492_),
    .A1(net5018),
    .A2(_06478_));
 sg13g2_nor2_1 _32215_ (.A(net4788),
    .B(_06492_),
    .Y(_06493_));
 sg13g2_xnor2_1 _32216_ (.Y(_06494_),
    .A(net4788),
    .B(_06492_));
 sg13g2_inv_1 _32217_ (.Y(_06495_),
    .A(_06494_));
 sg13g2_a21o_1 _32218_ (.A2(_06488_),
    .A1(_04454_),
    .B1(_04453_),
    .X(_06496_));
 sg13g2_nand3_1 _32219_ (.B(_04454_),
    .C(_06488_),
    .A(_04453_),
    .Y(_06497_));
 sg13g2_nand3_1 _32220_ (.B(_06496_),
    .C(_06497_),
    .A(net5720),
    .Y(_06498_));
 sg13g2_a21oi_1 _32221_ (.A1(net5654),
    .A2(\u_inv.d_next[255] ),
    .Y(_06499_),
    .B1(net4924));
 sg13g2_nand3_1 _32222_ (.B(_05828_),
    .C(_06477_),
    .A(_04453_),
    .Y(_06500_));
 sg13g2_a21oi_1 _32223_ (.A1(_05828_),
    .A2(_06477_),
    .Y(_06501_),
    .B1(_04453_));
 sg13g2_nor2_1 _32224_ (.A(net5020),
    .B(_06501_),
    .Y(_06502_));
 sg13g2_a22oi_1 _32225_ (.Y(_06503_),
    .B1(_06500_),
    .B2(_06502_),
    .A2(_06499_),
    .A1(_06498_));
 sg13g2_xnor2_1 _32226_ (.Y(_06504_),
    .A(net4788),
    .B(_06503_));
 sg13g2_nand2_1 _32227_ (.Y(_06505_),
    .A(_06495_),
    .B(_06504_));
 sg13g2_nand2b_1 _32228_ (.Y(_06506_),
    .B(_04463_),
    .A_N(_06485_));
 sg13g2_nand2_1 _32229_ (.Y(_06507_),
    .A(_04461_),
    .B(_06506_));
 sg13g2_a21oi_1 _32230_ (.A1(_04460_),
    .A2(_06507_),
    .Y(_06508_),
    .B1(net5650));
 sg13g2_o21ai_1 _32231_ (.B1(_06508_),
    .Y(_06509_),
    .A1(_04460_),
    .A2(_06507_));
 sg13g2_a21oi_1 _32232_ (.A1(net5654),
    .A2(\u_inv.d_next[253] ),
    .Y(_06510_),
    .B1(net4920));
 sg13g2_a21oi_1 _32233_ (.A1(_05824_),
    .A2(_06473_),
    .Y(_06511_),
    .B1(_04463_));
 sg13g2_a21o_1 _32234_ (.A2(_14557_),
    .A1(\u_inv.d_next[252] ),
    .B1(_06511_),
    .X(_06512_));
 sg13g2_or2_1 _32235_ (.X(_06513_),
    .B(_06512_),
    .A(_04460_));
 sg13g2_a21oi_1 _32236_ (.A1(_04460_),
    .A2(_06512_),
    .Y(_06514_),
    .B1(net5018));
 sg13g2_a22oi_1 _32237_ (.Y(_06515_),
    .B1(_06513_),
    .B2(_06514_),
    .A2(_06510_),
    .A1(_06509_));
 sg13g2_nor2_1 _32238_ (.A(net4731),
    .B(_06515_),
    .Y(_06516_));
 sg13g2_xnor2_1 _32239_ (.Y(_06517_),
    .A(net4788),
    .B(_06515_));
 sg13g2_xnor2_1 _32240_ (.Y(_06518_),
    .A(_04462_),
    .B(_06474_));
 sg13g2_nand2_1 _32241_ (.Y(_06519_),
    .A(_04462_),
    .B(_06485_));
 sg13g2_nand3_1 _32242_ (.B(_06506_),
    .C(_06519_),
    .A(net5718),
    .Y(_06520_));
 sg13g2_a21oi_1 _32243_ (.A1(net5650),
    .A2(\u_inv.d_next[252] ),
    .Y(_06521_),
    .B1(net4920));
 sg13g2_a22oi_1 _32244_ (.Y(_06522_),
    .B1(_06520_),
    .B2(_06521_),
    .A2(_06518_),
    .A1(net4921));
 sg13g2_nand2_1 _32245_ (.Y(_06523_),
    .A(net4731),
    .B(_06522_));
 sg13g2_xnor2_1 _32246_ (.Y(_06524_),
    .A(net4788),
    .B(_06522_));
 sg13g2_and2_1 _32247_ (.A(_06517_),
    .B(_06524_),
    .X(_06525_));
 sg13g2_inv_1 _32248_ (.Y(_06526_),
    .A(_06525_));
 sg13g2_a21oi_1 _32249_ (.A1(_05821_),
    .A2(_06472_),
    .Y(_06527_),
    .B1(_04468_));
 sg13g2_o21ai_1 _32250_ (.B1(_04470_),
    .Y(_06528_),
    .A1(_05818_),
    .A2(_06527_));
 sg13g2_or3_1 _32251_ (.A(_04470_),
    .B(_05818_),
    .C(_06527_),
    .X(_06529_));
 sg13g2_nand3_1 _32252_ (.B(_06528_),
    .C(_06529_),
    .A(net4920),
    .Y(_06530_));
 sg13g2_o21ai_1 _32253_ (.B1(_04468_),
    .Y(_06531_),
    .A1(_05879_),
    .A2(_06483_));
 sg13g2_nand2_1 _32254_ (.Y(_06532_),
    .A(_04467_),
    .B(_06531_));
 sg13g2_xnor2_1 _32255_ (.Y(_06533_),
    .A(_04470_),
    .B(_06532_));
 sg13g2_nor2b_1 _32256_ (.A(net5718),
    .B_N(\u_inv.d_next[251] ),
    .Y(_06534_));
 sg13g2_o21ai_1 _32257_ (.B1(net5018),
    .Y(_06535_),
    .A1(net5650),
    .A2(_06533_));
 sg13g2_o21ai_1 _32258_ (.B1(_06530_),
    .Y(_06536_),
    .A1(_06534_),
    .A2(_06535_));
 sg13g2_xnor2_1 _32259_ (.Y(_06537_),
    .A(net4787),
    .B(_06536_));
 sg13g2_nand3_1 _32260_ (.B(_05821_),
    .C(_06472_),
    .A(_04468_),
    .Y(_06538_));
 sg13g2_nand2b_1 _32261_ (.Y(_06539_),
    .B(_06538_),
    .A_N(_06527_));
 sg13g2_xnor2_1 _32262_ (.Y(_06540_),
    .A(_04468_),
    .B(_06484_));
 sg13g2_nand2_1 _32263_ (.Y(_06541_),
    .A(net5650),
    .B(\u_inv.d_next[250] ));
 sg13g2_a21oi_1 _32264_ (.A1(net5718),
    .A2(_06540_),
    .Y(_06542_),
    .B1(net4920));
 sg13g2_a22oi_1 _32265_ (.Y(_06543_),
    .B1(_06541_),
    .B2(_06542_),
    .A2(_06539_),
    .A1(net4920));
 sg13g2_nand2_1 _32266_ (.Y(_06544_),
    .A(net4730),
    .B(_06543_));
 sg13g2_xnor2_1 _32267_ (.Y(_06545_),
    .A(net4730),
    .B(_06543_));
 sg13g2_nor2_1 _32268_ (.A(_06537_),
    .B(_06545_),
    .Y(_06546_));
 sg13g2_nand2_1 _32269_ (.Y(_06547_),
    .A(_04477_),
    .B(_06482_));
 sg13g2_xnor2_1 _32270_ (.Y(_06548_),
    .A(_04477_),
    .B(_06482_));
 sg13g2_o21ai_1 _32271_ (.B1(net5018),
    .Y(_06549_),
    .A1(net5718),
    .A2(\u_inv.d_next[248] ));
 sg13g2_a21o_1 _32272_ (.A2(_06548_),
    .A1(net5719),
    .B1(_06549_),
    .X(_06550_));
 sg13g2_nor3_1 _32273_ (.A(_04478_),
    .B(_05817_),
    .C(_06470_),
    .Y(_06551_));
 sg13g2_nand2_1 _32274_ (.Y(_06552_),
    .A(net4920),
    .B(_06471_));
 sg13g2_o21ai_1 _32275_ (.B1(_06550_),
    .Y(_06553_),
    .A1(_06551_),
    .A2(_06552_));
 sg13g2_nand2_1 _32276_ (.Y(_06554_),
    .A(net4730),
    .B(_06553_));
 sg13g2_xnor2_1 _32277_ (.Y(_06555_),
    .A(net4730),
    .B(_06553_));
 sg13g2_and2_1 _32278_ (.A(_04476_),
    .B(_06547_),
    .X(_06556_));
 sg13g2_a21oi_1 _32279_ (.A1(_04475_),
    .A2(_06556_),
    .Y(_06557_),
    .B1(net5650));
 sg13g2_o21ai_1 _32280_ (.B1(_06557_),
    .Y(_06558_),
    .A1(_04475_),
    .A2(_06556_));
 sg13g2_a21oi_1 _32281_ (.A1(net5650),
    .A2(\u_inv.d_next[249] ),
    .Y(_06559_),
    .B1(net4920));
 sg13g2_and2_1 _32282_ (.A(_05819_),
    .B(_06471_),
    .X(_06560_));
 sg13g2_o21ai_1 _32283_ (.B1(net4920),
    .Y(_06561_),
    .A1(_04475_),
    .A2(_06560_));
 sg13g2_a21oi_1 _32284_ (.A1(_04475_),
    .A2(_06560_),
    .Y(_06562_),
    .B1(_06561_));
 sg13g2_a21o_2 _32285_ (.A2(_06559_),
    .A1(_06558_),
    .B1(_06562_),
    .X(_06563_));
 sg13g2_nand2_1 _32286_ (.Y(_06564_),
    .A(net4787),
    .B(_06563_));
 sg13g2_xnor2_1 _32287_ (.Y(_06565_),
    .A(net4787),
    .B(_06563_));
 sg13g2_nor4_1 _32288_ (.A(_06537_),
    .B(_06545_),
    .C(_06555_),
    .D(_06565_),
    .Y(_06566_));
 sg13g2_inv_1 _32289_ (.Y(_06567_),
    .A(_06566_));
 sg13g2_and4_1 _32290_ (.A(_06495_),
    .B(_06504_),
    .C(_06525_),
    .D(_06566_),
    .X(_06568_));
 sg13g2_o21ai_1 _32291_ (.B1(_05846_),
    .Y(_06569_),
    .A1(_05904_),
    .A2(_06480_));
 sg13g2_nand2_1 _32292_ (.Y(_06570_),
    .A(_05869_),
    .B(_06569_));
 sg13g2_o21ai_1 _32293_ (.B1(_05872_),
    .Y(_06571_),
    .A1(_05845_),
    .A2(_06569_));
 sg13g2_a21oi_1 _32294_ (.A1(_05843_),
    .A2(_06571_),
    .Y(_06572_),
    .B1(_05876_));
 sg13g2_nand2b_1 _32295_ (.Y(_06573_),
    .B(_04492_),
    .A_N(_06572_));
 sg13g2_o21ai_1 _32296_ (.B1(_06573_),
    .Y(_06574_),
    .A1(_14173_),
    .A2(_14563_));
 sg13g2_xnor2_1 _32297_ (.Y(_06575_),
    .A(_04494_),
    .B(_06574_));
 sg13g2_nand2_1 _32298_ (.Y(_06576_),
    .A(net5718),
    .B(_06575_));
 sg13g2_a21oi_1 _32299_ (.A1(net5649),
    .A2(\u_inv.d_next[247] ),
    .Y(_06577_),
    .B1(net4921));
 sg13g2_a21oi_1 _32300_ (.A1(_05738_),
    .A2(_06469_),
    .Y(_06578_),
    .B1(_04507_));
 sg13g2_a21oi_1 _32301_ (.A1(_05738_),
    .A2(_06469_),
    .Y(_06579_),
    .B1(_04509_));
 sg13g2_a21oi_1 _32302_ (.A1(_05738_),
    .A2(_06469_),
    .Y(_06580_),
    .B1(_04511_));
 sg13g2_nor2_1 _32303_ (.A(_05809_),
    .B(_06580_),
    .Y(_06581_));
 sg13g2_o21ai_1 _32304_ (.B1(_04491_),
    .Y(_06582_),
    .A1(_05809_),
    .A2(_06580_));
 sg13g2_a21oi_1 _32305_ (.A1(_05812_),
    .A2(_06582_),
    .Y(_06583_),
    .B1(_04492_));
 sg13g2_nor3_1 _32306_ (.A(_04493_),
    .B(_05813_),
    .C(_06583_),
    .Y(_06584_));
 sg13g2_o21ai_1 _32307_ (.B1(_04493_),
    .Y(_06585_),
    .A1(_05813_),
    .A2(_06583_));
 sg13g2_nor2_1 _32308_ (.A(net5018),
    .B(_06584_),
    .Y(_06586_));
 sg13g2_a22oi_1 _32309_ (.Y(_06587_),
    .B1(_06585_),
    .B2(_06586_),
    .A2(_06577_),
    .A1(_06576_));
 sg13g2_and2_1 _32310_ (.A(net4730),
    .B(_06587_),
    .X(_06588_));
 sg13g2_xnor2_1 _32311_ (.Y(_06589_),
    .A(net4730),
    .B(_06587_));
 sg13g2_nand3_1 _32312_ (.B(_05812_),
    .C(_06582_),
    .A(_04492_),
    .Y(_06590_));
 sg13g2_nand2b_1 _32313_ (.Y(_06591_),
    .B(_06590_),
    .A_N(_06583_));
 sg13g2_xnor2_1 _32314_ (.Y(_06592_),
    .A(_04492_),
    .B(_06572_));
 sg13g2_nand2_1 _32315_ (.Y(_06593_),
    .A(net5649),
    .B(\u_inv.d_next[246] ));
 sg13g2_a21oi_1 _32316_ (.A1(net5718),
    .A2(_06592_),
    .Y(_06594_),
    .B1(net4919));
 sg13g2_a22oi_1 _32317_ (.Y(_06595_),
    .B1(_06593_),
    .B2(_06594_),
    .A2(_06591_),
    .A1(net4921));
 sg13g2_and2_1 _32318_ (.A(net4730),
    .B(_06595_),
    .X(_06596_));
 sg13g2_xnor2_1 _32319_ (.Y(_06597_),
    .A(net4730),
    .B(_06595_));
 sg13g2_o21ai_1 _32320_ (.B1(_04489_),
    .Y(_06598_),
    .A1(_05809_),
    .A2(_06580_));
 sg13g2_xnor2_1 _32321_ (.Y(_06599_),
    .A(_04489_),
    .B(_06581_));
 sg13g2_xor2_1 _32322_ (.B(_06571_),
    .A(_04489_),
    .X(_06600_));
 sg13g2_a21oi_1 _32323_ (.A1(net5649),
    .A2(\u_inv.d_next[244] ),
    .Y(_06601_),
    .B1(net4919));
 sg13g2_o21ai_1 _32324_ (.B1(_06601_),
    .Y(_06602_),
    .A1(net5649),
    .A2(_06600_));
 sg13g2_o21ai_1 _32325_ (.B1(_06602_),
    .Y(_06603_),
    .A1(net5018),
    .A2(_06599_));
 sg13g2_nor2_1 _32326_ (.A(net4787),
    .B(_06603_),
    .Y(_06604_));
 sg13g2_nand2b_1 _32327_ (.Y(_06605_),
    .B(net4731),
    .A_N(_06603_));
 sg13g2_xnor2_1 _32328_ (.Y(_06606_),
    .A(net4787),
    .B(_06603_));
 sg13g2_a21oi_1 _32329_ (.A1(_04488_),
    .A2(_06571_),
    .Y(_06607_),
    .B1(_04487_));
 sg13g2_nand2_1 _32330_ (.Y(_06608_),
    .A(_04485_),
    .B(_06607_));
 sg13g2_nor2_1 _32331_ (.A(_04485_),
    .B(_06607_),
    .Y(_06609_));
 sg13g2_nor2_1 _32332_ (.A(net5650),
    .B(_06609_),
    .Y(_06610_));
 sg13g2_a221oi_1 _32333_ (.B2(_06610_),
    .C1(net4921),
    .B1(_06608_),
    .A1(net5650),
    .Y(_06611_),
    .A2(\u_inv.d_next[245] ));
 sg13g2_a21oi_1 _32334_ (.A1(_05810_),
    .A2(_06598_),
    .Y(_06612_),
    .B1(_04485_));
 sg13g2_nand3_1 _32335_ (.B(_05810_),
    .C(_06598_),
    .A(_04485_),
    .Y(_06613_));
 sg13g2_nor2_1 _32336_ (.A(net5018),
    .B(_06612_),
    .Y(_06614_));
 sg13g2_a21oi_2 _32337_ (.B1(_06611_),
    .Y(_06615_),
    .A2(_06614_),
    .A1(_06613_));
 sg13g2_and2_1 _32338_ (.A(net4731),
    .B(_06615_),
    .X(_06616_));
 sg13g2_nand2b_1 _32339_ (.Y(_06617_),
    .B(net4787),
    .A_N(_06615_));
 sg13g2_xnor2_1 _32340_ (.Y(_06618_),
    .A(net4731),
    .B(_06615_));
 sg13g2_or2_1 _32341_ (.X(_06619_),
    .B(_06618_),
    .A(_06606_));
 sg13g2_nor2_1 _32342_ (.A(_05807_),
    .B(_06579_),
    .Y(_06620_));
 sg13g2_o21ai_1 _32343_ (.B1(_04502_),
    .Y(_06621_),
    .A1(_05807_),
    .A2(_06579_));
 sg13g2_xnor2_1 _32344_ (.Y(_06622_),
    .A(_04501_),
    .B(_06620_));
 sg13g2_nand2_1 _32345_ (.Y(_06623_),
    .A(_04501_),
    .B(_06570_));
 sg13g2_nor2_1 _32346_ (.A(_04501_),
    .B(_06570_),
    .Y(_06624_));
 sg13g2_nor2_1 _32347_ (.A(net5649),
    .B(_06624_),
    .Y(_06625_));
 sg13g2_a221oi_1 _32348_ (.B2(_06625_),
    .C1(net4919),
    .B1(_06623_),
    .A1(net5649),
    .Y(_06626_),
    .A2(\u_inv.d_next[242] ));
 sg13g2_a21o_2 _32349_ (.A2(_06622_),
    .A1(net4919),
    .B1(_06626_),
    .X(_06627_));
 sg13g2_nand2b_1 _32350_ (.Y(_06628_),
    .B(net4732),
    .A_N(_06627_));
 sg13g2_inv_1 _32351_ (.Y(_06629_),
    .A(_06628_));
 sg13g2_xnor2_1 _32352_ (.Y(_06630_),
    .A(net4789),
    .B(_06627_));
 sg13g2_a21o_1 _32353_ (.A2(_06621_),
    .A1(_05804_),
    .B1(_04499_),
    .X(_06631_));
 sg13g2_nand3_1 _32354_ (.B(_05804_),
    .C(_06621_),
    .A(_04499_),
    .Y(_06632_));
 sg13g2_nand3_1 _32355_ (.B(_06631_),
    .C(_06632_),
    .A(net4919),
    .Y(_06633_));
 sg13g2_nand3_1 _32356_ (.B(_04500_),
    .C(_06623_),
    .A(_04499_),
    .Y(_06634_));
 sg13g2_a21o_1 _32357_ (.A2(_06623_),
    .A1(_04500_),
    .B1(_04499_),
    .X(_06635_));
 sg13g2_nand3_1 _32358_ (.B(_06634_),
    .C(_06635_),
    .A(net5718),
    .Y(_06636_));
 sg13g2_nand2_1 _32359_ (.Y(_06637_),
    .A(net5649),
    .B(\u_inv.d_next[243] ));
 sg13g2_nand3_1 _32360_ (.B(_06636_),
    .C(_06637_),
    .A(net5018),
    .Y(_06638_));
 sg13g2_and3_2 _32361_ (.X(_06639_),
    .A(net4732),
    .B(_06633_),
    .C(_06638_));
 sg13g2_a21oi_1 _32362_ (.A1(_06633_),
    .A2(_06638_),
    .Y(_06640_),
    .B1(net4732));
 sg13g2_nor2_1 _32363_ (.A(_06639_),
    .B(_06640_),
    .Y(_06641_));
 sg13g2_nor3_1 _32364_ (.A(_06630_),
    .B(_06639_),
    .C(_06640_),
    .Y(_06642_));
 sg13g2_o21ai_1 _32365_ (.B1(_04507_),
    .Y(_06643_),
    .A1(_05904_),
    .A2(_06480_));
 sg13g2_nor3_1 _32366_ (.A(_04507_),
    .B(_05904_),
    .C(_06480_),
    .Y(_06644_));
 sg13g2_nor2_1 _32367_ (.A(net5651),
    .B(_06644_),
    .Y(_06645_));
 sg13g2_nand3_1 _32368_ (.B(_05738_),
    .C(_06469_),
    .A(_04507_),
    .Y(_06646_));
 sg13g2_nand2b_1 _32369_ (.Y(_06647_),
    .B(_06646_),
    .A_N(_06578_));
 sg13g2_a221oi_1 _32370_ (.B2(_06645_),
    .C1(net4922),
    .B1(_06643_),
    .A1(net5651),
    .Y(_06648_),
    .A2(\u_inv.d_next[240] ));
 sg13g2_a21oi_2 _32371_ (.B1(_06648_),
    .Y(_06649_),
    .A2(_06647_),
    .A1(net4919));
 sg13g2_inv_1 _32372_ (.Y(_06650_),
    .A(_06649_));
 sg13g2_xnor2_1 _32373_ (.Y(_06651_),
    .A(net4789),
    .B(_06649_));
 sg13g2_o21ai_1 _32374_ (.B1(_04505_),
    .Y(_06652_),
    .A1(_05805_),
    .A2(_06578_));
 sg13g2_or3_1 _32375_ (.A(_04505_),
    .B(_05805_),
    .C(_06578_),
    .X(_06653_));
 sg13g2_nand3_1 _32376_ (.B(_06652_),
    .C(_06653_),
    .A(net4919),
    .Y(_06654_));
 sg13g2_nand3_1 _32377_ (.B(_04506_),
    .C(_06643_),
    .A(_04504_),
    .Y(_06655_));
 sg13g2_a21o_1 _32378_ (.A2(_06643_),
    .A1(_04506_),
    .B1(_04504_),
    .X(_06656_));
 sg13g2_nand3_1 _32379_ (.B(_06655_),
    .C(_06656_),
    .A(net5718),
    .Y(_06657_));
 sg13g2_a21oi_1 _32380_ (.A1(net5649),
    .A2(\u_inv.d_next[241] ),
    .Y(_06658_),
    .B1(net4919));
 sg13g2_nand2_1 _32381_ (.Y(_06659_),
    .A(_06657_),
    .B(_06658_));
 sg13g2_nand2_2 _32382_ (.Y(_06660_),
    .A(_06654_),
    .B(_06659_));
 sg13g2_and2_1 _32383_ (.A(net4789),
    .B(_06660_),
    .X(_06661_));
 sg13g2_xnor2_1 _32384_ (.Y(_06662_),
    .A(net4732),
    .B(_06660_));
 sg13g2_nand3_1 _32385_ (.B(_06651_),
    .C(_06662_),
    .A(_06642_),
    .Y(_06663_));
 sg13g2_nor4_2 _32386_ (.A(_06589_),
    .B(_06597_),
    .C(_06619_),
    .Y(_06664_),
    .D(_06663_));
 sg13g2_o21ai_1 _32387_ (.B1(_04574_),
    .Y(_06665_),
    .A1(_05802_),
    .A2(_06467_));
 sg13g2_nand2_1 _32388_ (.Y(_06666_),
    .A(_05722_),
    .B(_06665_));
 sg13g2_a21oi_1 _32389_ (.A1(_05722_),
    .A2(_06665_),
    .Y(_06667_),
    .B1(_04544_));
 sg13g2_a21oi_1 _32390_ (.A1(_05722_),
    .A2(_06665_),
    .Y(_06668_),
    .B1(_04546_));
 sg13g2_nor2_1 _32391_ (.A(_05737_),
    .B(_06668_),
    .Y(_06669_));
 sg13g2_o21ai_1 _32392_ (.B1(_04528_),
    .Y(_06670_),
    .A1(_05737_),
    .A2(_06668_));
 sg13g2_nand2_1 _32393_ (.Y(_06671_),
    .A(_05727_),
    .B(_06670_));
 sg13g2_a21oi_1 _32394_ (.A1(_05727_),
    .A2(_06670_),
    .Y(_06672_),
    .B1(_04519_));
 sg13g2_xnor2_1 _32395_ (.Y(_06673_),
    .A(_04518_),
    .B(_06671_));
 sg13g2_a21oi_2 _32396_ (.B1(_05864_),
    .Y(_06674_),
    .A2(_06435_),
    .A1(_06391_));
 sg13g2_nor2_1 _32397_ (.A(_05895_),
    .B(_06674_),
    .Y(_06675_));
 sg13g2_o21ai_1 _32398_ (.B1(_05856_),
    .Y(_06676_),
    .A1(_05895_),
    .A2(_06674_));
 sg13g2_nand2_1 _32399_ (.Y(_06677_),
    .A(_05897_),
    .B(_06676_));
 sg13g2_o21ai_1 _32400_ (.B1(_05899_),
    .Y(_06678_),
    .A1(_05854_),
    .A2(_06676_));
 sg13g2_a21oi_1 _32401_ (.A1(_05852_),
    .A2(_06678_),
    .Y(_06679_),
    .B1(_05900_));
 sg13g2_xnor2_1 _32402_ (.Y(_06680_),
    .A(_04519_),
    .B(_06679_));
 sg13g2_nand2_1 _32403_ (.Y(_06681_),
    .A(net5651),
    .B(\u_inv.d_next[238] ));
 sg13g2_a21oi_1 _32404_ (.A1(net5719),
    .A2(_06680_),
    .Y(_06682_),
    .B1(net4922));
 sg13g2_a22oi_1 _32405_ (.Y(_06683_),
    .B1(_06681_),
    .B2(_06682_),
    .A2(_06673_),
    .A1(net4922));
 sg13g2_and2_1 _32406_ (.A(net4732),
    .B(_06683_),
    .X(_06684_));
 sg13g2_xnor2_1 _32407_ (.Y(_06685_),
    .A(net4789),
    .B(_06683_));
 sg13g2_inv_1 _32408_ (.Y(_06686_),
    .A(_06685_));
 sg13g2_o21ai_1 _32409_ (.B1(_04517_),
    .Y(_06687_),
    .A1(_04518_),
    .A2(_06679_));
 sg13g2_o21ai_1 _32410_ (.B1(net5719),
    .Y(_06688_),
    .A1(_04515_),
    .A2(_06687_));
 sg13g2_a21oi_1 _32411_ (.A1(_04515_),
    .A2(_06687_),
    .Y(_06689_),
    .B1(_06688_));
 sg13g2_a21oi_1 _32412_ (.A1(net5651),
    .A2(\u_inv.d_next[239] ),
    .Y(_06690_),
    .B1(net4922));
 sg13g2_nand2b_1 _32413_ (.Y(_06691_),
    .B(_06690_),
    .A_N(_06689_));
 sg13g2_o21ai_1 _32414_ (.B1(_04515_),
    .Y(_06692_),
    .A1(_05728_),
    .A2(_06672_));
 sg13g2_or3_1 _32415_ (.A(_04515_),
    .B(_05728_),
    .C(_06672_),
    .X(_06693_));
 sg13g2_nand3_1 _32416_ (.B(_06692_),
    .C(_06693_),
    .A(net4922),
    .Y(_06694_));
 sg13g2_and2_1 _32417_ (.A(_06691_),
    .B(_06694_),
    .X(_06695_));
 sg13g2_nand3_1 _32418_ (.B(_06691_),
    .C(_06694_),
    .A(net4732),
    .Y(_06696_));
 sg13g2_a21o_1 _32419_ (.A2(_06694_),
    .A1(_06691_),
    .B1(net4733),
    .X(_06697_));
 sg13g2_nand2_1 _32420_ (.Y(_06698_),
    .A(_06696_),
    .B(_06697_));
 sg13g2_nand2_1 _32421_ (.Y(_06699_),
    .A(_04525_),
    .B(_06678_));
 sg13g2_nand3_1 _32422_ (.B(_04524_),
    .C(_06699_),
    .A(_04523_),
    .Y(_06700_));
 sg13g2_a21o_1 _32423_ (.A2(_06699_),
    .A1(_04524_),
    .B1(_04523_),
    .X(_06701_));
 sg13g2_nand3_1 _32424_ (.B(_06700_),
    .C(_06701_),
    .A(net5719),
    .Y(_06702_));
 sg13g2_nand2_1 _32425_ (.Y(_06703_),
    .A(net5651),
    .B(\u_inv.d_next[237] ));
 sg13g2_nand3_1 _32426_ (.B(_06702_),
    .C(_06703_),
    .A(net5019),
    .Y(_06704_));
 sg13g2_o21ai_1 _32427_ (.B1(_04526_),
    .Y(_06705_),
    .A1(_05737_),
    .A2(_06668_));
 sg13g2_a21o_1 _32428_ (.A2(_06705_),
    .A1(_05726_),
    .B1(_04523_),
    .X(_06706_));
 sg13g2_nand3_1 _32429_ (.B(_05726_),
    .C(_06705_),
    .A(_04523_),
    .Y(_06707_));
 sg13g2_nand3_1 _32430_ (.B(_06706_),
    .C(_06707_),
    .A(net4922),
    .Y(_06708_));
 sg13g2_and3_1 _32431_ (.X(_06709_),
    .A(net4733),
    .B(_06704_),
    .C(_06708_));
 sg13g2_a21oi_1 _32432_ (.A1(_06704_),
    .A2(_06708_),
    .Y(_06710_),
    .B1(net4733));
 sg13g2_or2_1 _32433_ (.X(_06711_),
    .B(_06710_),
    .A(_06709_));
 sg13g2_xnor2_1 _32434_ (.Y(_06712_),
    .A(_04525_),
    .B(_06669_));
 sg13g2_nand2b_1 _32435_ (.Y(_06713_),
    .B(_04526_),
    .A_N(_06678_));
 sg13g2_nand3_1 _32436_ (.B(_06699_),
    .C(_06713_),
    .A(net5719),
    .Y(_06714_));
 sg13g2_a21oi_1 _32437_ (.A1(net5651),
    .A2(\u_inv.d_next[236] ),
    .Y(_06715_),
    .B1(net4922));
 sg13g2_a22oi_1 _32438_ (.Y(_06716_),
    .B1(_06714_),
    .B2(_06715_),
    .A2(_06712_),
    .A1(net4922));
 sg13g2_and2_1 _32439_ (.A(net4732),
    .B(_06716_),
    .X(_06717_));
 sg13g2_xnor2_1 _32440_ (.Y(_06718_),
    .A(net4732),
    .B(_06716_));
 sg13g2_nor3_1 _32441_ (.A(_06709_),
    .B(_06710_),
    .C(_06718_),
    .Y(_06719_));
 sg13g2_nand4_1 _32442_ (.B(_06696_),
    .C(_06697_),
    .A(_06685_),
    .Y(_06720_),
    .D(_06719_));
 sg13g2_nor2_1 _32443_ (.A(_05734_),
    .B(_06667_),
    .Y(_06721_));
 sg13g2_o21ai_1 _32444_ (.B1(_04537_),
    .Y(_06722_),
    .A1(_05734_),
    .A2(_06667_));
 sg13g2_nand3_1 _32445_ (.B(_05735_),
    .C(_06722_),
    .A(_04533_),
    .Y(_06723_));
 sg13g2_a21o_1 _32446_ (.A2(_06722_),
    .A1(_05735_),
    .B1(_04533_),
    .X(_06724_));
 sg13g2_nand3_1 _32447_ (.B(_06723_),
    .C(_06724_),
    .A(net4923),
    .Y(_06725_));
 sg13g2_a21oi_1 _32448_ (.A1(_04536_),
    .A2(_06677_),
    .Y(_06726_),
    .B1(_04535_));
 sg13g2_xnor2_1 _32449_ (.Y(_06727_),
    .A(_04533_),
    .B(_06726_));
 sg13g2_o21ai_1 _32450_ (.B1(net5019),
    .Y(_06728_),
    .A1(net5652),
    .A2(_06727_));
 sg13g2_a21o_1 _32451_ (.A2(\u_inv.d_next[235] ),
    .A1(net5652),
    .B1(_06728_),
    .X(_06729_));
 sg13g2_and3_1 _32452_ (.X(_06730_),
    .A(net4734),
    .B(_06725_),
    .C(_06729_));
 sg13g2_a21oi_1 _32453_ (.A1(_06725_),
    .A2(_06729_),
    .Y(_06731_),
    .B1(net4734));
 sg13g2_nor2_1 _32454_ (.A(_06730_),
    .B(_06731_),
    .Y(_06732_));
 sg13g2_xnor2_1 _32455_ (.Y(_06733_),
    .A(_04537_),
    .B(_06721_));
 sg13g2_xnor2_1 _32456_ (.Y(_06734_),
    .A(_04536_),
    .B(_06677_));
 sg13g2_a21oi_1 _32457_ (.A1(net5652),
    .A2(\u_inv.d_next[234] ),
    .Y(_06735_),
    .B1(net4923));
 sg13g2_o21ai_1 _32458_ (.B1(_06735_),
    .Y(_06736_),
    .A1(net5652),
    .A2(_06734_));
 sg13g2_o21ai_1 _32459_ (.B1(_06736_),
    .Y(_06737_),
    .A1(net5019),
    .A2(_06733_));
 sg13g2_nand2b_1 _32460_ (.Y(_06738_),
    .B(net4734),
    .A_N(_06737_));
 sg13g2_xnor2_1 _32461_ (.Y(_06739_),
    .A(net4789),
    .B(_06737_));
 sg13g2_nor3_1 _32462_ (.A(_06730_),
    .B(_06731_),
    .C(_06739_),
    .Y(_06740_));
 sg13g2_a21oi_1 _32463_ (.A1(_04542_),
    .A2(_06666_),
    .Y(_06741_),
    .B1(_05732_));
 sg13g2_a21oi_1 _32464_ (.A1(_04540_),
    .A2(_06741_),
    .Y(_06742_),
    .B1(net5019));
 sg13g2_o21ai_1 _32465_ (.B1(_06742_),
    .Y(_06743_),
    .A1(_04540_),
    .A2(_06741_));
 sg13g2_o21ai_1 _32466_ (.B1(_04541_),
    .Y(_06744_),
    .A1(_05895_),
    .A2(_06674_));
 sg13g2_o21ai_1 _32467_ (.B1(_06744_),
    .Y(_06745_),
    .A1(_14177_),
    .A2(_14577_));
 sg13g2_xnor2_1 _32468_ (.Y(_06746_),
    .A(_04539_),
    .B(_06745_));
 sg13g2_nor2_1 _32469_ (.A(net5652),
    .B(_06746_),
    .Y(_06747_));
 sg13g2_o21ai_1 _32470_ (.B1(net5019),
    .Y(_06748_),
    .A1(net5719),
    .A2(_14176_));
 sg13g2_o21ai_1 _32471_ (.B1(_06743_),
    .Y(_06749_),
    .A1(_06747_),
    .A2(_06748_));
 sg13g2_nand2_1 _32472_ (.Y(_06750_),
    .A(net4789),
    .B(_06749_));
 sg13g2_xnor2_1 _32473_ (.Y(_06751_),
    .A(net4733),
    .B(_06749_));
 sg13g2_xnor2_1 _32474_ (.Y(_06752_),
    .A(_04542_),
    .B(_06666_));
 sg13g2_a21oi_1 _32475_ (.A1(_04542_),
    .A2(_06675_),
    .Y(_06753_),
    .B1(net5651));
 sg13g2_nand2_1 _32476_ (.Y(_06754_),
    .A(_06744_),
    .B(_06753_));
 sg13g2_a21oi_1 _32477_ (.A1(net5651),
    .A2(\u_inv.d_next[232] ),
    .Y(_06755_),
    .B1(net4923));
 sg13g2_a22oi_1 _32478_ (.Y(_06756_),
    .B1(_06754_),
    .B2(_06755_),
    .A2(_06752_),
    .A1(net4923));
 sg13g2_nand2_1 _32479_ (.Y(_06757_),
    .A(net4733),
    .B(_06756_));
 sg13g2_xnor2_1 _32480_ (.Y(_06758_),
    .A(net4733),
    .B(_06756_));
 sg13g2_inv_1 _32481_ (.Y(_06759_),
    .A(_06758_));
 sg13g2_nand3_1 _32482_ (.B(_06751_),
    .C(_06759_),
    .A(_06740_),
    .Y(_06760_));
 sg13g2_nor2_1 _32483_ (.A(_06720_),
    .B(_06760_),
    .Y(_06761_));
 sg13g2_a21oi_1 _32484_ (.A1(_06391_),
    .A2(_06435_),
    .Y(_06762_),
    .B1(_04570_));
 sg13g2_nand2_1 _32485_ (.Y(_06763_),
    .A(_04569_),
    .B(_06479_));
 sg13g2_a21oi_2 _32486_ (.B1(_05889_),
    .Y(_06764_),
    .A2(_06762_),
    .A1(_04566_));
 sg13g2_o21ai_1 _32487_ (.B1(_05892_),
    .Y(_06765_),
    .A1(_05860_),
    .A2(_06764_));
 sg13g2_a21oi_1 _32488_ (.A1(_05861_),
    .A2(_06765_),
    .Y(_06766_),
    .B1(_05888_));
 sg13g2_o21ai_1 _32489_ (.B1(_04553_),
    .Y(_06767_),
    .A1(_04554_),
    .A2(_06766_));
 sg13g2_xnor2_1 _32490_ (.Y(_06768_),
    .A(_04556_),
    .B(_06767_));
 sg13g2_a21o_1 _32491_ (.A2(\u_inv.d_next[231] ),
    .A1(net5654),
    .B1(net4925),
    .X(_06769_));
 sg13g2_a21o_1 _32492_ (.A2(_06768_),
    .A1(net5722),
    .B1(_06769_),
    .X(_06770_));
 sg13g2_o21ai_1 _32493_ (.B1(_04571_),
    .Y(_06771_),
    .A1(_05802_),
    .A2(_06467_));
 sg13g2_o21ai_1 _32494_ (.B1(_04573_),
    .Y(_06772_),
    .A1(_05802_),
    .A2(_06467_));
 sg13g2_nand2_1 _32495_ (.Y(_06773_),
    .A(_05712_),
    .B(_06772_));
 sg13g2_a21oi_1 _32496_ (.A1(_05712_),
    .A2(_06772_),
    .Y(_06774_),
    .B1(_04552_));
 sg13g2_o21ai_1 _32497_ (.B1(_04554_),
    .Y(_06775_),
    .A1(_05719_),
    .A2(_06774_));
 sg13g2_nand3_1 _32498_ (.B(_05715_),
    .C(_06775_),
    .A(_04556_),
    .Y(_06776_));
 sg13g2_a21o_1 _32499_ (.A2(_06775_),
    .A1(_05715_),
    .B1(_04556_),
    .X(_06777_));
 sg13g2_nand3_1 _32500_ (.B(_06776_),
    .C(_06777_),
    .A(net4925),
    .Y(_06778_));
 sg13g2_and3_2 _32501_ (.X(_06779_),
    .A(net4735),
    .B(_06770_),
    .C(_06778_));
 sg13g2_a21oi_1 _32502_ (.A1(_06770_),
    .A2(_06778_),
    .Y(_06780_),
    .B1(net4735));
 sg13g2_nor2_1 _32503_ (.A(_06779_),
    .B(_06780_),
    .Y(_06781_));
 sg13g2_or3_1 _32504_ (.A(_04554_),
    .B(_05719_),
    .C(_06774_),
    .X(_06782_));
 sg13g2_nand2_1 _32505_ (.Y(_06783_),
    .A(_06775_),
    .B(_06782_));
 sg13g2_xor2_1 _32506_ (.B(_06766_),
    .A(_04554_),
    .X(_06784_));
 sg13g2_nand2_1 _32507_ (.Y(_06785_),
    .A(net5654),
    .B(\u_inv.d_next[230] ));
 sg13g2_a21oi_1 _32508_ (.A1(net5722),
    .A2(_06784_),
    .Y(_06786_),
    .B1(net4925));
 sg13g2_a22oi_1 _32509_ (.Y(_06787_),
    .B1(_06785_),
    .B2(_06786_),
    .A2(_06783_),
    .A1(net4925));
 sg13g2_nand2_1 _32510_ (.Y(_06788_),
    .A(net4735),
    .B(_06787_));
 sg13g2_xnor2_1 _32511_ (.Y(_06789_),
    .A(net4735),
    .B(_06787_));
 sg13g2_nor3_1 _32512_ (.A(_06779_),
    .B(_06780_),
    .C(_06789_),
    .Y(_06790_));
 sg13g2_a21oi_1 _32513_ (.A1(_05712_),
    .A2(_06772_),
    .Y(_06791_),
    .B1(_04550_));
 sg13g2_xor2_1 _32514_ (.B(_06773_),
    .A(_04550_),
    .X(_06792_));
 sg13g2_xnor2_1 _32515_ (.Y(_06793_),
    .A(_04550_),
    .B(_06765_));
 sg13g2_o21ai_1 _32516_ (.B1(net5021),
    .Y(_06794_),
    .A1(net5722),
    .A2(\u_inv.d_next[228] ));
 sg13g2_a21o_1 _32517_ (.A2(_06793_),
    .A1(net5722),
    .B1(_06794_),
    .X(_06795_));
 sg13g2_o21ai_1 _32518_ (.B1(_06795_),
    .Y(_06796_),
    .A1(net5021),
    .A2(_06792_));
 sg13g2_nand2_1 _32519_ (.Y(_06797_),
    .A(net4735),
    .B(_06796_));
 sg13g2_xnor2_1 _32520_ (.Y(_06798_),
    .A(net4792),
    .B(_06796_));
 sg13g2_inv_2 _32521_ (.Y(_06799_),
    .A(_06798_));
 sg13g2_a21oi_1 _32522_ (.A1(_04550_),
    .A2(_06765_),
    .Y(_06800_),
    .B1(_04549_));
 sg13g2_xnor2_1 _32523_ (.Y(_06801_),
    .A(_04548_),
    .B(_06800_));
 sg13g2_o21ai_1 _32524_ (.B1(net5021),
    .Y(_06802_),
    .A1(net5723),
    .A2(_14178_));
 sg13g2_a21o_1 _32525_ (.A2(_06801_),
    .A1(net5723),
    .B1(_06802_),
    .X(_06803_));
 sg13g2_or3_1 _32526_ (.A(_04548_),
    .B(_05717_),
    .C(_06791_),
    .X(_06804_));
 sg13g2_o21ai_1 _32527_ (.B1(_04548_),
    .Y(_06805_),
    .A1(_05717_),
    .A2(_06791_));
 sg13g2_nand3_1 _32528_ (.B(_06804_),
    .C(_06805_),
    .A(net4925),
    .Y(_06806_));
 sg13g2_nand3_1 _32529_ (.B(_06803_),
    .C(_06806_),
    .A(net4735),
    .Y(_06807_));
 sg13g2_a21o_1 _32530_ (.A2(_06806_),
    .A1(_06803_),
    .B1(net4736),
    .X(_06808_));
 sg13g2_and2_1 _32531_ (.A(_06807_),
    .B(_06808_),
    .X(_06809_));
 sg13g2_nand3_1 _32532_ (.B(_06807_),
    .C(_06808_),
    .A(_06798_),
    .Y(_06810_));
 sg13g2_nor4_1 _32533_ (.A(_06779_),
    .B(_06780_),
    .C(_06789_),
    .D(_06810_),
    .Y(_06811_));
 sg13g2_o21ai_1 _32534_ (.B1(_04561_),
    .Y(_06812_),
    .A1(_04562_),
    .A2(_06764_));
 sg13g2_xnor2_1 _32535_ (.Y(_06813_),
    .A(_04559_),
    .B(_06812_));
 sg13g2_a21oi_1 _32536_ (.A1(net5654),
    .A2(\u_inv.d_next[227] ),
    .Y(_06814_),
    .B1(net4925));
 sg13g2_o21ai_1 _32537_ (.B1(_06814_),
    .Y(_06815_),
    .A1(net5654),
    .A2(_06813_));
 sg13g2_a21oi_1 _32538_ (.A1(_05708_),
    .A2(_06771_),
    .Y(_06816_),
    .B1(_04563_));
 sg13g2_a21o_1 _32539_ (.A2(_06771_),
    .A1(_05708_),
    .B1(_04563_),
    .X(_06817_));
 sg13g2_o21ai_1 _32540_ (.B1(_04559_),
    .Y(_06818_),
    .A1(_05705_),
    .A2(_06816_));
 sg13g2_or3_1 _32541_ (.A(_04559_),
    .B(_05705_),
    .C(_06816_),
    .X(_06819_));
 sg13g2_nand3_1 _32542_ (.B(_06818_),
    .C(_06819_),
    .A(net4925),
    .Y(_06820_));
 sg13g2_nand3_1 _32543_ (.B(_06815_),
    .C(_06820_),
    .A(net4736),
    .Y(_06821_));
 sg13g2_a21o_1 _32544_ (.A2(_06820_),
    .A1(_06815_),
    .B1(net4736),
    .X(_06822_));
 sg13g2_nand2_1 _32545_ (.Y(_06823_),
    .A(_06821_),
    .B(_06822_));
 sg13g2_nand3_1 _32546_ (.B(_05708_),
    .C(_06771_),
    .A(_04563_),
    .Y(_06824_));
 sg13g2_a21oi_1 _32547_ (.A1(_06817_),
    .A2(_06824_),
    .Y(_06825_),
    .B1(net5021));
 sg13g2_xnor2_1 _32548_ (.Y(_06826_),
    .A(_04562_),
    .B(_06764_));
 sg13g2_o21ai_1 _32549_ (.B1(net5020),
    .Y(_06827_),
    .A1(net5655),
    .A2(_06826_));
 sg13g2_a21oi_1 _32550_ (.A1(net5655),
    .A2(\u_inv.d_next[226] ),
    .Y(_06828_),
    .B1(_06827_));
 sg13g2_nor2_2 _32551_ (.A(_06825_),
    .B(_06828_),
    .Y(_06829_));
 sg13g2_nor3_1 _32552_ (.A(net4792),
    .B(_06825_),
    .C(_06828_),
    .Y(_06830_));
 sg13g2_inv_1 _32553_ (.Y(_06831_),
    .A(_06830_));
 sg13g2_xnor2_1 _32554_ (.Y(_06832_),
    .A(net4792),
    .B(_06829_));
 sg13g2_xnor2_1 _32555_ (.Y(_06833_),
    .A(net4736),
    .B(_06829_));
 sg13g2_nor2_1 _32556_ (.A(_04569_),
    .B(_06479_),
    .Y(_06834_));
 sg13g2_nor2_1 _32557_ (.A(net5662),
    .B(_06834_),
    .Y(_06835_));
 sg13g2_xnor2_1 _32558_ (.Y(_06836_),
    .A(_04569_),
    .B(_06468_));
 sg13g2_a221oi_1 _32559_ (.B2(_06835_),
    .C1(net4932),
    .B1(_06763_),
    .A1(net5658),
    .Y(_06837_),
    .A2(\u_inv.d_next[224] ));
 sg13g2_a21oi_2 _32560_ (.B1(_06837_),
    .Y(_06838_),
    .A2(_06836_),
    .A1(net4937));
 sg13g2_nand2_1 _32561_ (.Y(_06839_),
    .A(net4735),
    .B(_06838_));
 sg13g2_inv_1 _32562_ (.Y(_06840_),
    .A(_06839_));
 sg13g2_xnor2_1 _32563_ (.Y(_06841_),
    .A(net4791),
    .B(_06838_));
 sg13g2_o21ai_1 _32564_ (.B1(_05706_),
    .Y(_06842_),
    .A1(_04569_),
    .A2(_06468_));
 sg13g2_and2_1 _32565_ (.A(_04566_),
    .B(_06842_),
    .X(_06843_));
 sg13g2_o21ai_1 _32566_ (.B1(net4937),
    .Y(_06844_),
    .A1(_04566_),
    .A2(_06842_));
 sg13g2_a21o_1 _32567_ (.A2(_06763_),
    .A1(_04568_),
    .B1(_04567_),
    .X(_06845_));
 sg13g2_nand3_1 _32568_ (.B(_04568_),
    .C(_06763_),
    .A(_04567_),
    .Y(_06846_));
 sg13g2_nand3_1 _32569_ (.B(_06845_),
    .C(_06846_),
    .A(net5733),
    .Y(_06847_));
 sg13g2_a21oi_1 _32570_ (.A1(net5662),
    .A2(net5875),
    .Y(_06848_),
    .B1(net4925));
 sg13g2_nand2_1 _32571_ (.Y(_06849_),
    .A(_06847_),
    .B(_06848_));
 sg13g2_o21ai_1 _32572_ (.B1(_06849_),
    .Y(_06850_),
    .A1(_06843_),
    .A2(_06844_));
 sg13g2_and2_1 _32573_ (.A(net4792),
    .B(_06850_),
    .X(_06851_));
 sg13g2_xnor2_1 _32574_ (.Y(_06852_),
    .A(net4735),
    .B(_06850_));
 sg13g2_nand2_1 _32575_ (.Y(_06853_),
    .A(_06841_),
    .B(_06852_));
 sg13g2_nor3_1 _32576_ (.A(_06823_),
    .B(_06833_),
    .C(_06853_),
    .Y(_06854_));
 sg13g2_and2_1 _32577_ (.A(_06811_),
    .B(_06854_),
    .X(_06855_));
 sg13g2_and2_1 _32578_ (.A(_06761_),
    .B(_06855_),
    .X(_06856_));
 sg13g2_nand3_1 _32579_ (.B(_06664_),
    .C(_06856_),
    .A(_06568_),
    .Y(_06857_));
 sg13g2_a21oi_1 _32580_ (.A1(_05009_),
    .A2(_05702_),
    .Y(_06858_),
    .B1(_04674_));
 sg13g2_a21oi_2 _32581_ (.B1(_04680_),
    .Y(_06859_),
    .A2(_05702_),
    .A1(_05009_));
 sg13g2_a21oi_2 _32582_ (.B1(_05756_),
    .Y(_06860_),
    .A2(_06859_),
    .A1(_04670_));
 sg13g2_a21oi_2 _32583_ (.B1(_05772_),
    .Y(_06861_),
    .A2(_05703_),
    .A1(_04681_));
 sg13g2_o21ai_1 _32584_ (.B1(_05800_),
    .Y(_06862_),
    .A1(_04631_),
    .A2(_06861_));
 sg13g2_a21oi_2 _32585_ (.B1(_05779_),
    .Y(_06863_),
    .A2(_06862_),
    .A1(_04604_));
 sg13g2_o21ai_1 _32586_ (.B1(_05782_),
    .Y(_06864_),
    .A1(_04588_),
    .A2(_06863_));
 sg13g2_xnor2_1 _32587_ (.Y(_06865_),
    .A(_04580_),
    .B(_06864_));
 sg13g2_or2_1 _32588_ (.X(_06866_),
    .B(_06362_),
    .A(_04673_));
 sg13g2_o21ai_1 _32589_ (.B1(_06387_),
    .Y(_06867_),
    .A1(_06358_),
    .A2(_06361_));
 sg13g2_nor3_2 _32590_ (.A(_06362_),
    .B(_06385_),
    .C(_06388_),
    .Y(_06868_));
 sg13g2_o21ai_1 _32591_ (.B1(_06389_),
    .Y(_06869_),
    .A1(_06358_),
    .A2(_06361_));
 sg13g2_a21oi_2 _32592_ (.B1(_04629_),
    .Y(_06870_),
    .A2(_06869_),
    .A1(_06432_));
 sg13g2_a21oi_2 _32593_ (.B1(_06402_),
    .Y(_06871_),
    .A2(_06870_),
    .A1(_06374_));
 sg13g2_nor2_1 _32594_ (.A(_06367_),
    .B(_06871_),
    .Y(_06872_));
 sg13g2_or2_1 _32595_ (.X(_06873_),
    .B(_06872_),
    .A(_06404_));
 sg13g2_a21oi_2 _32596_ (.B1(_06406_),
    .Y(_06874_),
    .A2(_06872_),
    .A1(_06366_));
 sg13g2_o21ai_1 _32597_ (.B1(_06410_),
    .Y(_06875_),
    .A1(_06364_),
    .A2(_06874_));
 sg13g2_xnor2_1 _32598_ (.Y(_06876_),
    .A(_04580_),
    .B(_06875_));
 sg13g2_a21oi_1 _32599_ (.A1(net5658),
    .A2(\u_inv.d_next[222] ),
    .Y(_06877_),
    .B1(net4932));
 sg13g2_o21ai_1 _32600_ (.B1(_06877_),
    .Y(_06878_),
    .A1(net5658),
    .A2(_06876_));
 sg13g2_o21ai_1 _32601_ (.B1(_06878_),
    .Y(_06879_),
    .A1(net5030),
    .A2(_06865_));
 sg13g2_nand2b_1 _32602_ (.Y(_06880_),
    .B(net4738),
    .A_N(_06879_));
 sg13g2_xnor2_1 _32603_ (.Y(_06881_),
    .A(net4738),
    .B(_06879_));
 sg13g2_a21oi_1 _32604_ (.A1(_04580_),
    .A2(_06875_),
    .Y(_06882_),
    .B1(_04579_));
 sg13g2_xnor2_1 _32605_ (.Y(_06883_),
    .A(_04578_),
    .B(_06882_));
 sg13g2_a21oi_1 _32606_ (.A1(net5658),
    .A2(\u_inv.d_next[223] ),
    .Y(_06884_),
    .B1(net4932));
 sg13g2_o21ai_1 _32607_ (.B1(_06884_),
    .Y(_06885_),
    .A1(net5658),
    .A2(_06883_));
 sg13g2_a21oi_1 _32608_ (.A1(_04581_),
    .A2(_06864_),
    .Y(_06886_),
    .B1(_05783_));
 sg13g2_and2_1 _32609_ (.A(_04578_),
    .B(_06886_),
    .X(_06887_));
 sg13g2_o21ai_1 _32610_ (.B1(net4932),
    .Y(_06888_),
    .A1(_04578_),
    .A2(_06886_));
 sg13g2_o21ai_1 _32611_ (.B1(_06885_),
    .Y(_06889_),
    .A1(_06887_),
    .A2(_06888_));
 sg13g2_inv_1 _32612_ (.Y(_06890_),
    .A(_06889_));
 sg13g2_nand2_1 _32613_ (.Y(_06891_),
    .A(net4738),
    .B(_06890_));
 sg13g2_xnor2_1 _32614_ (.Y(_06892_),
    .A(net4738),
    .B(_06889_));
 sg13g2_o21ai_1 _32615_ (.B1(_04585_),
    .Y(_06893_),
    .A1(_04587_),
    .A2(_06874_));
 sg13g2_a21oi_1 _32616_ (.A1(_04583_),
    .A2(_06893_),
    .Y(_06894_),
    .B1(net5659));
 sg13g2_o21ai_1 _32617_ (.B1(_06894_),
    .Y(_06895_),
    .A1(_04583_),
    .A2(_06893_));
 sg13g2_a21oi_1 _32618_ (.A1(net5659),
    .A2(\u_inv.d_next[221] ),
    .Y(_06896_),
    .B1(net4932));
 sg13g2_o21ai_1 _32619_ (.B1(_05780_),
    .Y(_06897_),
    .A1(_04586_),
    .A2(_06863_));
 sg13g2_o21ai_1 _32620_ (.B1(net4932),
    .Y(_06898_),
    .A1(_04583_),
    .A2(_06897_));
 sg13g2_a21oi_1 _32621_ (.A1(_04583_),
    .A2(_06897_),
    .Y(_06899_),
    .B1(_06898_));
 sg13g2_a21o_2 _32622_ (.A2(_06896_),
    .A1(_06895_),
    .B1(_06899_),
    .X(_06900_));
 sg13g2_nand2_1 _32623_ (.Y(_06901_),
    .A(net4797),
    .B(_06900_));
 sg13g2_xnor2_1 _32624_ (.Y(_06902_),
    .A(net4738),
    .B(_06900_));
 sg13g2_xnor2_1 _32625_ (.Y(_06903_),
    .A(_04587_),
    .B(_06863_));
 sg13g2_xnor2_1 _32626_ (.Y(_06904_),
    .A(_04587_),
    .B(_06874_));
 sg13g2_a21oi_1 _32627_ (.A1(net5659),
    .A2(\u_inv.d_next[220] ),
    .Y(_06905_),
    .B1(net4935));
 sg13g2_o21ai_1 _32628_ (.B1(_06905_),
    .Y(_06906_),
    .A1(net5659),
    .A2(_06904_));
 sg13g2_o21ai_1 _32629_ (.B1(_06906_),
    .Y(_06907_),
    .A1(net5028),
    .A2(_06903_));
 sg13g2_nand2b_1 _32630_ (.Y(_06908_),
    .B(net4738),
    .A_N(_06907_));
 sg13g2_xnor2_1 _32631_ (.Y(_06909_),
    .A(net4738),
    .B(_06907_));
 sg13g2_inv_1 _32632_ (.Y(_06910_),
    .A(_06909_));
 sg13g2_and4_1 _32633_ (.A(_06881_),
    .B(_06892_),
    .C(_06902_),
    .D(_06909_),
    .X(_06911_));
 sg13g2_a21o_1 _32634_ (.A2(_06862_),
    .A1(_04603_),
    .B1(_05775_),
    .X(_06912_));
 sg13g2_xnor2_1 _32635_ (.Y(_06913_),
    .A(_04595_),
    .B(_06912_));
 sg13g2_nand2_1 _32636_ (.Y(_06914_),
    .A(_04594_),
    .B(_06873_));
 sg13g2_xnor2_1 _32637_ (.Y(_06915_),
    .A(_04595_),
    .B(_06873_));
 sg13g2_nand2_1 _32638_ (.Y(_06916_),
    .A(net5659),
    .B(\u_inv.d_next[218] ));
 sg13g2_a21oi_1 _32639_ (.A1(net5732),
    .A2(_06915_),
    .Y(_06917_),
    .B1(net4935));
 sg13g2_a22oi_1 _32640_ (.Y(_06918_),
    .B1(_06916_),
    .B2(_06917_),
    .A2(_06913_),
    .A1(net4935));
 sg13g2_xnor2_1 _32641_ (.Y(_06919_),
    .A(net4796),
    .B(_06918_));
 sg13g2_inv_1 _32642_ (.Y(_06920_),
    .A(_06919_));
 sg13g2_nand3_1 _32643_ (.B(_04593_),
    .C(_06914_),
    .A(_04592_),
    .Y(_06921_));
 sg13g2_a21o_1 _32644_ (.A2(_06914_),
    .A1(_04593_),
    .B1(_04592_),
    .X(_06922_));
 sg13g2_nand3_1 _32645_ (.B(_06921_),
    .C(_06922_),
    .A(net5732),
    .Y(_06923_));
 sg13g2_a21oi_1 _32646_ (.A1(net5659),
    .A2(\u_inv.d_next[219] ),
    .Y(_06924_),
    .B1(net4935));
 sg13g2_a21oi_1 _32647_ (.A1(_04595_),
    .A2(_06912_),
    .Y(_06925_),
    .B1(_05777_));
 sg13g2_nand2b_1 _32648_ (.Y(_06926_),
    .B(_04591_),
    .A_N(_06925_));
 sg13g2_a21oi_1 _32649_ (.A1(_04592_),
    .A2(_06925_),
    .Y(_06927_),
    .B1(net5028));
 sg13g2_a22oi_1 _32650_ (.Y(_06928_),
    .B1(_06926_),
    .B2(_06927_),
    .A2(_06924_),
    .A1(_06923_));
 sg13g2_xnor2_1 _32651_ (.Y(_06929_),
    .A(net4796),
    .B(_06928_));
 sg13g2_o21ai_1 _32652_ (.B1(_04600_),
    .Y(_06930_),
    .A1(_04602_),
    .A2(_06871_));
 sg13g2_a21oi_1 _32653_ (.A1(_04599_),
    .A2(_06930_),
    .Y(_06931_),
    .B1(net5659));
 sg13g2_o21ai_1 _32654_ (.B1(_06931_),
    .Y(_06932_),
    .A1(_04599_),
    .A2(_06930_));
 sg13g2_a21oi_1 _32655_ (.A1(net5659),
    .A2(\u_inv.d_next[217] ),
    .Y(_06933_),
    .B1(net4935));
 sg13g2_a21o_1 _32656_ (.A2(_06862_),
    .A1(_04602_),
    .B1(_05773_),
    .X(_06934_));
 sg13g2_or2_1 _32657_ (.X(_06935_),
    .B(_06934_),
    .A(_04599_));
 sg13g2_a21oi_1 _32658_ (.A1(_04599_),
    .A2(_06934_),
    .Y(_06936_),
    .B1(net5028));
 sg13g2_a22oi_1 _32659_ (.Y(_06937_),
    .B1(_06935_),
    .B2(_06936_),
    .A2(_06933_),
    .A1(_06932_));
 sg13g2_nand2_1 _32660_ (.Y(_06938_),
    .A(net4739),
    .B(_06937_));
 sg13g2_nor2_1 _32661_ (.A(net4739),
    .B(_06937_),
    .Y(_06939_));
 sg13g2_xnor2_1 _32662_ (.Y(_06940_),
    .A(net4796),
    .B(_06937_));
 sg13g2_xnor2_1 _32663_ (.Y(_06941_),
    .A(_04602_),
    .B(_06862_));
 sg13g2_xnor2_1 _32664_ (.Y(_06942_),
    .A(_04602_),
    .B(_06871_));
 sg13g2_o21ai_1 _32665_ (.B1(net5028),
    .Y(_06943_),
    .A1(net5732),
    .A2(\u_inv.d_next[216] ));
 sg13g2_a21o_1 _32666_ (.A2(_06942_),
    .A1(net5732),
    .B1(_06943_),
    .X(_06944_));
 sg13g2_o21ai_1 _32667_ (.B1(_06944_),
    .Y(_06945_),
    .A1(net5028),
    .A2(_06941_));
 sg13g2_nand2_1 _32668_ (.Y(_06946_),
    .A(net4739),
    .B(_06945_));
 sg13g2_xnor2_1 _32669_ (.Y(_06947_),
    .A(net4739),
    .B(_06945_));
 sg13g2_inv_2 _32670_ (.Y(_06948_),
    .A(_06947_));
 sg13g2_and4_1 _32671_ (.A(_06919_),
    .B(_06929_),
    .C(_06940_),
    .D(_06948_),
    .X(_06949_));
 sg13g2_nand2_1 _32672_ (.Y(_06950_),
    .A(_06911_),
    .B(_06949_));
 sg13g2_nor2_1 _32673_ (.A(_04628_),
    .B(_06861_),
    .Y(_06951_));
 sg13g2_o21ai_1 _32674_ (.B1(_05792_),
    .Y(_06952_),
    .A1(_04630_),
    .A2(_06861_));
 sg13g2_a21oi_1 _32675_ (.A1(_04611_),
    .A2(_06952_),
    .Y(_06953_),
    .B1(_05795_));
 sg13g2_xnor2_1 _32676_ (.Y(_06954_),
    .A(_04613_),
    .B(_06953_));
 sg13g2_a21oi_1 _32677_ (.A1(\u_inv.d_next[208] ),
    .A2(\u_inv.d_reg[208] ),
    .Y(_06955_),
    .B1(_06870_));
 sg13g2_a21oi_2 _32678_ (.B1(_06396_),
    .Y(_06956_),
    .A2(_06870_),
    .A1(_04626_));
 sg13g2_o21ai_1 _32679_ (.B1(_06398_),
    .Y(_06957_),
    .A1(_06371_),
    .A2(_06956_));
 sg13g2_a21oi_1 _32680_ (.A1(_06372_),
    .A2(_06957_),
    .Y(_06958_),
    .B1(_06394_));
 sg13g2_xnor2_1 _32681_ (.Y(_06959_),
    .A(_04613_),
    .B(_06958_));
 sg13g2_nand2_1 _32682_ (.Y(_06960_),
    .A(net5660),
    .B(\u_inv.d_next[214] ));
 sg13g2_a21oi_1 _32683_ (.A1(net5732),
    .A2(_06959_),
    .Y(_06961_),
    .B1(net4935));
 sg13g2_a22oi_1 _32684_ (.Y(_06962_),
    .B1(_06960_),
    .B2(_06961_),
    .A2(_06954_),
    .A1(net4935));
 sg13g2_nand2_1 _32685_ (.Y(_06963_),
    .A(net4739),
    .B(_06962_));
 sg13g2_xnor2_1 _32686_ (.Y(_06964_),
    .A(net4796),
    .B(_06962_));
 sg13g2_o21ai_1 _32687_ (.B1(_04612_),
    .Y(_06965_),
    .A1(_04614_),
    .A2(_06958_));
 sg13g2_o21ai_1 _32688_ (.B1(net5731),
    .Y(_06966_),
    .A1(_04616_),
    .A2(_06965_));
 sg13g2_a21o_1 _32689_ (.A2(_06965_),
    .A1(_04616_),
    .B1(_06966_),
    .X(_06967_));
 sg13g2_a21oi_1 _32690_ (.A1(net5660),
    .A2(\u_inv.d_next[215] ),
    .Y(_06968_),
    .B1(net4935));
 sg13g2_o21ai_1 _32691_ (.B1(_05796_),
    .Y(_06969_),
    .A1(_04613_),
    .A2(_06953_));
 sg13g2_nand2b_1 _32692_ (.Y(_06970_),
    .B(_04617_),
    .A_N(_06969_));
 sg13g2_a21oi_1 _32693_ (.A1(_04616_),
    .A2(_06969_),
    .Y(_06971_),
    .B1(net5028));
 sg13g2_a22oi_1 _32694_ (.Y(_06972_),
    .B1(_06970_),
    .B2(_06971_),
    .A2(_06968_),
    .A1(_06967_));
 sg13g2_xnor2_1 _32695_ (.Y(_06973_),
    .A(net4796),
    .B(_06972_));
 sg13g2_nand2_1 _32696_ (.Y(_06974_),
    .A(_06964_),
    .B(_06973_));
 sg13g2_a21o_1 _32697_ (.A2(_06957_),
    .A1(_04609_),
    .B1(_04608_),
    .X(_06975_));
 sg13g2_a21oi_1 _32698_ (.A1(_04606_),
    .A2(_06975_),
    .Y(_06976_),
    .B1(net5660));
 sg13g2_o21ai_1 _32699_ (.B1(_06976_),
    .Y(_06977_),
    .A1(_04606_),
    .A2(_06975_));
 sg13g2_a21oi_1 _32700_ (.A1(net5660),
    .A2(\u_inv.d_next[213] ),
    .Y(_06978_),
    .B1(net4936));
 sg13g2_nand2_1 _32701_ (.Y(_06979_),
    .A(_04610_),
    .B(_06952_));
 sg13g2_nand3_1 _32702_ (.B(_05794_),
    .C(_06979_),
    .A(_04607_),
    .Y(_06980_));
 sg13g2_a21oi_1 _32703_ (.A1(_05794_),
    .A2(_06979_),
    .Y(_06981_),
    .B1(_04607_));
 sg13g2_nor2_1 _32704_ (.A(net5029),
    .B(_06981_),
    .Y(_06982_));
 sg13g2_a22oi_1 _32705_ (.Y(_06983_),
    .B1(_06980_),
    .B2(_06982_),
    .A2(_06978_),
    .A1(_06977_));
 sg13g2_nand2b_1 _32706_ (.Y(_06984_),
    .B(net4796),
    .A_N(_06983_));
 sg13g2_xnor2_1 _32707_ (.Y(_06985_),
    .A(net4742),
    .B(_06983_));
 sg13g2_xnor2_1 _32708_ (.Y(_06986_),
    .A(_04610_),
    .B(_06952_));
 sg13g2_xor2_1 _32709_ (.B(_06957_),
    .A(_04610_),
    .X(_06987_));
 sg13g2_o21ai_1 _32710_ (.B1(net5028),
    .Y(_06988_),
    .A1(net5745),
    .A2(\u_inv.d_next[212] ));
 sg13g2_a21o_1 _32711_ (.A2(_06987_),
    .A1(net5745),
    .B1(_06988_),
    .X(_06989_));
 sg13g2_o21ai_1 _32712_ (.B1(_06989_),
    .Y(_06990_),
    .A1(net5028),
    .A2(_06986_));
 sg13g2_nand2_1 _32713_ (.Y(_06991_),
    .A(net4742),
    .B(_06990_));
 sg13g2_xnor2_1 _32714_ (.Y(_06992_),
    .A(net4742),
    .B(_06990_));
 sg13g2_nor3_1 _32715_ (.A(_06974_),
    .B(_06985_),
    .C(_06992_),
    .Y(_06993_));
 sg13g2_o21ai_1 _32716_ (.B1(_04623_),
    .Y(_06994_),
    .A1(_04624_),
    .A2(_06956_));
 sg13g2_xnor2_1 _32717_ (.Y(_06995_),
    .A(_04622_),
    .B(_06994_));
 sg13g2_nand2_1 _32718_ (.Y(_06996_),
    .A(net5748),
    .B(_06995_));
 sg13g2_a21oi_1 _32719_ (.A1(net5668),
    .A2(\u_inv.d_next[211] ),
    .Y(_06997_),
    .B1(net4945));
 sg13g2_a21o_1 _32720_ (.A2(_06951_),
    .A1(_04627_),
    .B1(_05789_),
    .X(_06998_));
 sg13g2_a21oi_1 _32721_ (.A1(_04624_),
    .A2(_06998_),
    .Y(_06999_),
    .B1(_05791_));
 sg13g2_xor2_1 _32722_ (.B(_06999_),
    .A(_04622_),
    .X(_07000_));
 sg13g2_a22oi_1 _32723_ (.Y(_07001_),
    .B1(_07000_),
    .B2(net4945),
    .A2(_06997_),
    .A1(_06996_));
 sg13g2_xnor2_1 _32724_ (.Y(_07002_),
    .A(net4802),
    .B(_07001_));
 sg13g2_xnor2_1 _32725_ (.Y(_07003_),
    .A(_04624_),
    .B(_06998_));
 sg13g2_xor2_1 _32726_ (.B(_06956_),
    .A(_04624_),
    .X(_07004_));
 sg13g2_nand2_1 _32727_ (.Y(_07005_),
    .A(net5671),
    .B(\u_inv.d_next[210] ));
 sg13g2_a21oi_1 _32728_ (.A1(net5745),
    .A2(_07004_),
    .Y(_07006_),
    .B1(net4945));
 sg13g2_a22oi_1 _32729_ (.Y(_07007_),
    .B1(_07005_),
    .B2(_07006_),
    .A2(_07003_),
    .A1(net4945));
 sg13g2_and2_1 _32730_ (.A(net4742),
    .B(_07007_),
    .X(_07008_));
 sg13g2_xnor2_1 _32731_ (.Y(_07009_),
    .A(net4802),
    .B(_07007_));
 sg13g2_nand2_1 _32732_ (.Y(_07010_),
    .A(_07002_),
    .B(_07009_));
 sg13g2_or3_1 _32733_ (.A(_04626_),
    .B(_05787_),
    .C(_06951_),
    .X(_07011_));
 sg13g2_o21ai_1 _32734_ (.B1(_04626_),
    .Y(_07012_),
    .A1(_05787_),
    .A2(_06951_));
 sg13g2_nand3_1 _32735_ (.B(_07011_),
    .C(_07012_),
    .A(net4945),
    .Y(_07013_));
 sg13g2_xnor2_1 _32736_ (.Y(_07014_),
    .A(_04627_),
    .B(_06955_));
 sg13g2_a21oi_1 _32737_ (.A1(net5671),
    .A2(\u_inv.d_next[209] ),
    .Y(_07015_),
    .B1(net4945));
 sg13g2_o21ai_1 _32738_ (.B1(_07015_),
    .Y(_07016_),
    .A1(net5671),
    .A2(_07014_));
 sg13g2_nand2_1 _32739_ (.Y(_07017_),
    .A(_07013_),
    .B(_07016_));
 sg13g2_nand3_1 _32740_ (.B(_07013_),
    .C(_07016_),
    .A(net4742),
    .Y(_07018_));
 sg13g2_nand2_1 _32741_ (.Y(_07019_),
    .A(net4802),
    .B(_07017_));
 sg13g2_and2_1 _32742_ (.A(_07018_),
    .B(_07019_),
    .X(_07020_));
 sg13g2_xnor2_1 _32743_ (.Y(_07021_),
    .A(_04628_),
    .B(_06861_));
 sg13g2_nand3_1 _32744_ (.B(_06432_),
    .C(_06869_),
    .A(_04629_),
    .Y(_07022_));
 sg13g2_nand3b_1 _32745_ (.B(_07022_),
    .C(net5745),
    .Y(_07023_),
    .A_N(_06870_));
 sg13g2_a21oi_1 _32746_ (.A1(net5668),
    .A2(\u_inv.d_next[208] ),
    .Y(_07024_),
    .B1(net4945));
 sg13g2_a22oi_1 _32747_ (.Y(_07025_),
    .B1(_07023_),
    .B2(_07024_),
    .A2(_07021_),
    .A1(net4945));
 sg13g2_nand2_1 _32748_ (.Y(_07026_),
    .A(net4742),
    .B(_07025_));
 sg13g2_xnor2_1 _32749_ (.Y(_07027_),
    .A(net4742),
    .B(_07025_));
 sg13g2_inv_1 _32750_ (.Y(_07028_),
    .A(_07027_));
 sg13g2_nand4_1 _32751_ (.B(_07009_),
    .C(_07020_),
    .A(_07002_),
    .Y(_07029_),
    .D(_07028_));
 sg13g2_inv_1 _32752_ (.Y(_07030_),
    .A(_07029_));
 sg13g2_nor4_1 _32753_ (.A(_06974_),
    .B(_06985_),
    .C(_06992_),
    .D(_07029_),
    .Y(_07031_));
 sg13g2_inv_1 _32754_ (.Y(_07032_),
    .A(_07031_));
 sg13g2_and3_1 _32755_ (.X(_07033_),
    .A(_06911_),
    .B(_06949_),
    .C(_07031_));
 sg13g2_o21ai_1 _32756_ (.B1(_05768_),
    .Y(_07034_),
    .A1(_04657_),
    .A2(_06860_));
 sg13g2_a21oi_1 _32757_ (.A1(_04644_),
    .A2(_07034_),
    .Y(_07035_),
    .B1(_05759_));
 sg13g2_xor2_1 _32758_ (.B(_07035_),
    .A(_04636_),
    .X(_07036_));
 sg13g2_o21ai_1 _32759_ (.B1(_06381_),
    .Y(_07037_),
    .A1(_06421_),
    .A2(_06868_));
 sg13g2_nor2b_1 _32760_ (.A(_06422_),
    .B_N(_07037_),
    .Y(_07038_));
 sg13g2_o21ai_1 _32761_ (.B1(_06424_),
    .Y(_07039_),
    .A1(_06380_),
    .A2(_07037_));
 sg13g2_a21oi_1 _32762_ (.A1(_06377_),
    .A2(_07039_),
    .Y(_07040_),
    .B1(_06427_));
 sg13g2_nand2b_1 _32763_ (.Y(_07041_),
    .B(_04636_),
    .A_N(_07040_));
 sg13g2_xor2_1 _32764_ (.B(_07040_),
    .A(_04636_),
    .X(_07042_));
 sg13g2_a21oi_1 _32765_ (.A1(net5668),
    .A2(\u_inv.d_next[206] ),
    .Y(_07043_),
    .B1(net4950));
 sg13g2_o21ai_1 _32766_ (.B1(_07043_),
    .Y(_07044_),
    .A1(net5668),
    .A2(_07042_));
 sg13g2_o21ai_1 _32767_ (.B1(_07044_),
    .Y(_07045_),
    .A1(net5038),
    .A2(_07036_));
 sg13g2_nor2_1 _32768_ (.A(net4799),
    .B(_07045_),
    .Y(_07046_));
 sg13g2_nand2_1 _32769_ (.Y(_07047_),
    .A(net4800),
    .B(_07045_));
 sg13g2_xnor2_1 _32770_ (.Y(_07048_),
    .A(net4800),
    .B(_07045_));
 sg13g2_nand3_1 _32771_ (.B(_04635_),
    .C(_07041_),
    .A(_04634_),
    .Y(_07049_));
 sg13g2_a21o_1 _32772_ (.A2(_07041_),
    .A1(_04635_),
    .B1(_04634_),
    .X(_07050_));
 sg13g2_nand3_1 _32773_ (.B(_07049_),
    .C(_07050_),
    .A(net5745),
    .Y(_07051_));
 sg13g2_a21oi_1 _32774_ (.A1(net5668),
    .A2(\u_inv.d_next[207] ),
    .Y(_07052_),
    .B1(net4950));
 sg13g2_o21ai_1 _32775_ (.B1(_05760_),
    .Y(_07053_),
    .A1(_04636_),
    .A2(_07035_));
 sg13g2_nand2b_1 _32776_ (.Y(_07054_),
    .B(_04634_),
    .A_N(_07053_));
 sg13g2_a21oi_1 _32777_ (.A1(_04633_),
    .A2(_07053_),
    .Y(_07055_),
    .B1(net5040));
 sg13g2_a22oi_1 _32778_ (.Y(_07056_),
    .B1(_07054_),
    .B2(_07055_),
    .A2(_07052_),
    .A1(_07051_));
 sg13g2_xnor2_1 _32779_ (.Y(_07057_),
    .A(net4745),
    .B(_07056_));
 sg13g2_xnor2_1 _32780_ (.Y(_07058_),
    .A(_04643_),
    .B(_07034_));
 sg13g2_xnor2_1 _32781_ (.Y(_07059_),
    .A(_04643_),
    .B(_07039_));
 sg13g2_a21oi_1 _32782_ (.A1(net5669),
    .A2(\u_inv.d_next[204] ),
    .Y(_07060_),
    .B1(net4946));
 sg13g2_o21ai_1 _32783_ (.B1(_07060_),
    .Y(_07061_),
    .A1(net5669),
    .A2(_07059_));
 sg13g2_o21ai_1 _32784_ (.B1(_07061_),
    .Y(_07062_),
    .A1(net5038),
    .A2(_07058_));
 sg13g2_nand2b_1 _32785_ (.Y(_07063_),
    .B(net4745),
    .A_N(_07062_));
 sg13g2_xnor2_1 _32786_ (.Y(_07064_),
    .A(net4800),
    .B(_07062_));
 sg13g2_a21oi_1 _32787_ (.A1(_04643_),
    .A2(_07039_),
    .Y(_07065_),
    .B1(_04641_));
 sg13g2_xor2_1 _32788_ (.B(_07065_),
    .A(_04640_),
    .X(_07066_));
 sg13g2_o21ai_1 _32789_ (.B1(net5040),
    .Y(_07067_),
    .A1(net5745),
    .A2(_14186_));
 sg13g2_a21oi_1 _32790_ (.A1(net5747),
    .A2(_07066_),
    .Y(_07068_),
    .B1(_07067_));
 sg13g2_a21oi_1 _32791_ (.A1(_04642_),
    .A2(_07034_),
    .Y(_07069_),
    .B1(_05758_));
 sg13g2_or2_1 _32792_ (.X(_07070_),
    .B(_07069_),
    .A(_04640_));
 sg13g2_a21oi_1 _32793_ (.A1(_04640_),
    .A2(_07069_),
    .Y(_07071_),
    .B1(net5040));
 sg13g2_a21o_2 _32794_ (.A2(_07071_),
    .A1(_07070_),
    .B1(_07068_),
    .X(_07072_));
 sg13g2_xnor2_1 _32795_ (.Y(_07073_),
    .A(net4745),
    .B(_07072_));
 sg13g2_nand2b_1 _32796_ (.Y(_07074_),
    .B(_07073_),
    .A_N(_07064_));
 sg13g2_nor3_1 _32797_ (.A(_07048_),
    .B(_07057_),
    .C(_07074_),
    .Y(_07075_));
 sg13g2_o21ai_1 _32798_ (.B1(_05764_),
    .Y(_07076_),
    .A1(_04656_),
    .A2(_06860_));
 sg13g2_xnor2_1 _32799_ (.Y(_07077_),
    .A(_04648_),
    .B(_07076_));
 sg13g2_xor2_1 _32800_ (.B(_07038_),
    .A(_04648_),
    .X(_07078_));
 sg13g2_nand2_1 _32801_ (.Y(_07079_),
    .A(net5669),
    .B(\u_inv.d_next[202] ));
 sg13g2_a21oi_1 _32802_ (.A1(net5747),
    .A2(_07078_),
    .Y(_07080_),
    .B1(net4948));
 sg13g2_a22oi_1 _32803_ (.Y(_07081_),
    .B1(_07079_),
    .B2(_07080_),
    .A2(_07077_),
    .A1(net4948));
 sg13g2_and2_1 _32804_ (.A(net4745),
    .B(_07081_),
    .X(_07082_));
 sg13g2_xnor2_1 _32805_ (.Y(_07083_),
    .A(net4800),
    .B(_07081_));
 sg13g2_o21ai_1 _32806_ (.B1(_04647_),
    .Y(_07084_),
    .A1(_04648_),
    .A2(_07038_));
 sg13g2_xnor2_1 _32807_ (.Y(_07085_),
    .A(_04646_),
    .B(_07084_));
 sg13g2_nand2_1 _32808_ (.Y(_07086_),
    .A(net5747),
    .B(_07085_));
 sg13g2_a21oi_1 _32809_ (.A1(net5669),
    .A2(\u_inv.d_next[203] ),
    .Y(_07087_),
    .B1(net4948));
 sg13g2_a21oi_1 _32810_ (.A1(_04648_),
    .A2(_07076_),
    .Y(_07088_),
    .B1(_05765_));
 sg13g2_or2_1 _32811_ (.X(_07089_),
    .B(_07088_),
    .A(_04646_));
 sg13g2_a21oi_1 _32812_ (.A1(_04646_),
    .A2(_07088_),
    .Y(_07090_),
    .B1(net5040));
 sg13g2_a22oi_1 _32813_ (.Y(_07091_),
    .B1(_07089_),
    .B2(_07090_),
    .A2(_07087_),
    .A1(_07086_));
 sg13g2_xnor2_1 _32814_ (.Y(_07092_),
    .A(net4800),
    .B(_07091_));
 sg13g2_nand2_1 _32815_ (.Y(_07093_),
    .A(_07083_),
    .B(_07092_));
 sg13g2_o21ai_1 _32816_ (.B1(_04655_),
    .Y(_07094_),
    .A1(_06421_),
    .A2(_06868_));
 sg13g2_nand3_1 _32817_ (.B(_04654_),
    .C(_07094_),
    .A(_04653_),
    .Y(_07095_));
 sg13g2_a21o_1 _32818_ (.A2(_07094_),
    .A1(_04654_),
    .B1(_04653_),
    .X(_07096_));
 sg13g2_nand3_1 _32819_ (.B(_07095_),
    .C(_07096_),
    .A(net5747),
    .Y(_07097_));
 sg13g2_a21oi_1 _32820_ (.A1(net5669),
    .A2(\u_inv.d_next[201] ),
    .Y(_07098_),
    .B1(net4948));
 sg13g2_o21ai_1 _32821_ (.B1(_05762_),
    .Y(_07099_),
    .A1(_04655_),
    .A2(_06860_));
 sg13g2_o21ai_1 _32822_ (.B1(net4948),
    .Y(_07100_),
    .A1(_04652_),
    .A2(_07099_));
 sg13g2_a21oi_1 _32823_ (.A1(_04652_),
    .A2(_07099_),
    .Y(_07101_),
    .B1(_07100_));
 sg13g2_a21oi_2 _32824_ (.B1(_07101_),
    .Y(_07102_),
    .A2(_07098_),
    .A1(_07097_));
 sg13g2_inv_1 _32825_ (.Y(_07103_),
    .A(_07102_));
 sg13g2_xnor2_1 _32826_ (.Y(_07104_),
    .A(net4745),
    .B(_07102_));
 sg13g2_xnor2_1 _32827_ (.Y(_07105_),
    .A(_04655_),
    .B(_06860_));
 sg13g2_nor3_1 _32828_ (.A(_04655_),
    .B(_06421_),
    .C(_06868_),
    .Y(_07106_));
 sg13g2_nor2_1 _32829_ (.A(net5669),
    .B(_07106_),
    .Y(_07107_));
 sg13g2_a221oi_1 _32830_ (.B2(_07107_),
    .C1(net4948),
    .B1(_07094_),
    .A1(net5669),
    .Y(_07108_),
    .A2(\u_inv.d_next[200] ));
 sg13g2_a21oi_2 _32831_ (.B1(_07108_),
    .Y(_07109_),
    .A2(_07105_),
    .A1(net4948));
 sg13g2_nand2_1 _32832_ (.Y(_07110_),
    .A(net4746),
    .B(_07109_));
 sg13g2_xnor2_1 _32833_ (.Y(_07111_),
    .A(net4746),
    .B(_07109_));
 sg13g2_nor3_1 _32834_ (.A(_07093_),
    .B(_07104_),
    .C(_07111_),
    .Y(_07112_));
 sg13g2_nand2_1 _32835_ (.Y(_07113_),
    .A(_07075_),
    .B(_07112_));
 sg13g2_nor2_1 _32836_ (.A(_05746_),
    .B(_06859_),
    .Y(_07114_));
 sg13g2_o21ai_1 _32837_ (.B1(_04665_),
    .Y(_07115_),
    .A1(_05746_),
    .A2(_06859_));
 sg13g2_nand3_1 _32838_ (.B(_05751_),
    .C(_07115_),
    .A(_04669_),
    .Y(_07116_));
 sg13g2_a21o_1 _32839_ (.A2(_07115_),
    .A1(_05751_),
    .B1(_04669_),
    .X(_07117_));
 sg13g2_a21oi_1 _32840_ (.A1(_07116_),
    .A2(_07117_),
    .Y(_07118_),
    .B1(net5039));
 sg13g2_o21ai_1 _32841_ (.B1(_06417_),
    .Y(_07119_),
    .A1(_06362_),
    .A2(_06388_));
 sg13g2_a21oi_1 _32842_ (.A1(_06384_),
    .A2(_07119_),
    .Y(_07120_),
    .B1(_06418_));
 sg13g2_nand2b_1 _32843_ (.Y(_07121_),
    .B(_04669_),
    .A_N(_07120_));
 sg13g2_xor2_1 _32844_ (.B(_07120_),
    .A(_04669_),
    .X(_07122_));
 sg13g2_a21oi_1 _32845_ (.A1(net5669),
    .A2(\u_inv.d_next[198] ),
    .Y(_07123_),
    .B1(net4949));
 sg13g2_o21ai_1 _32846_ (.B1(_07123_),
    .Y(_07124_),
    .A1(net5671),
    .A2(_07122_));
 sg13g2_nand2b_2 _32847_ (.Y(_07125_),
    .B(_07124_),
    .A_N(_07118_));
 sg13g2_nor2_1 _32848_ (.A(net4802),
    .B(_07125_),
    .Y(_07126_));
 sg13g2_nand2_1 _32849_ (.Y(_07127_),
    .A(net4802),
    .B(_07125_));
 sg13g2_nand2b_1 _32850_ (.Y(_07128_),
    .B(_07127_),
    .A_N(_07126_));
 sg13g2_nand3_1 _32851_ (.B(_04668_),
    .C(_07121_),
    .A(_04667_),
    .Y(_07129_));
 sg13g2_a21o_1 _32852_ (.A2(_07121_),
    .A1(_04668_),
    .B1(_04667_),
    .X(_07130_));
 sg13g2_nand3_1 _32853_ (.B(_07129_),
    .C(_07130_),
    .A(net5746),
    .Y(_07131_));
 sg13g2_nand2_1 _32854_ (.Y(_07132_),
    .A(net5670),
    .B(\u_inv.d_next[199] ));
 sg13g2_nand3_1 _32855_ (.B(_07131_),
    .C(_07132_),
    .A(net5039),
    .Y(_07133_));
 sg13g2_nand3_1 _32856_ (.B(_05753_),
    .C(_07117_),
    .A(_04667_),
    .Y(_07134_));
 sg13g2_a21oi_1 _32857_ (.A1(_05753_),
    .A2(_07117_),
    .Y(_07135_),
    .B1(_04667_));
 sg13g2_nand2_1 _32858_ (.Y(_07136_),
    .A(net4948),
    .B(_07134_));
 sg13g2_o21ai_1 _32859_ (.B1(_07133_),
    .Y(_07137_),
    .A1(_07135_),
    .A2(_07136_));
 sg13g2_xnor2_1 _32860_ (.Y(_07138_),
    .A(net4745),
    .B(_07137_));
 sg13g2_nand2b_1 _32861_ (.Y(_07139_),
    .B(_07138_),
    .A_N(_07128_));
 sg13g2_o21ai_1 _32862_ (.B1(_04663_),
    .Y(_07140_),
    .A1(_05746_),
    .A2(_06859_));
 sg13g2_xor2_1 _32863_ (.B(_07114_),
    .A(_04663_),
    .X(_07141_));
 sg13g2_nand2b_1 _32864_ (.Y(_07142_),
    .B(_07119_),
    .A_N(_04663_));
 sg13g2_xor2_1 _32865_ (.B(_07119_),
    .A(_04663_),
    .X(_07143_));
 sg13g2_o21ai_1 _32866_ (.B1(net5039),
    .Y(_07144_),
    .A1(net5747),
    .A2(\u_inv.d_next[196] ));
 sg13g2_a21o_1 _32867_ (.A2(_07143_),
    .A1(net5747),
    .B1(_07144_),
    .X(_07145_));
 sg13g2_o21ai_1 _32868_ (.B1(_07145_),
    .Y(_07146_),
    .A1(net5039),
    .A2(_07141_));
 sg13g2_and2_1 _32869_ (.A(net4747),
    .B(_07146_),
    .X(_07147_));
 sg13g2_nand3_1 _32870_ (.B(_04662_),
    .C(_07142_),
    .A(_04661_),
    .Y(_07148_));
 sg13g2_a21o_1 _32871_ (.A2(_07142_),
    .A1(_04662_),
    .B1(_04661_),
    .X(_07149_));
 sg13g2_nand3_1 _32872_ (.B(_07148_),
    .C(_07149_),
    .A(net5747),
    .Y(_07150_));
 sg13g2_nand2_1 _32873_ (.Y(_07151_),
    .A(net5670),
    .B(\u_inv.d_next[197] ));
 sg13g2_nand3_1 _32874_ (.B(_07150_),
    .C(_07151_),
    .A(net5039),
    .Y(_07152_));
 sg13g2_nand3_1 _32875_ (.B(_05750_),
    .C(_07140_),
    .A(_04661_),
    .Y(_07153_));
 sg13g2_a21o_1 _32876_ (.A2(_07140_),
    .A1(_05750_),
    .B1(_04661_),
    .X(_07154_));
 sg13g2_nand3_1 _32877_ (.B(_07153_),
    .C(_07154_),
    .A(net4949),
    .Y(_07155_));
 sg13g2_nand2_1 _32878_ (.Y(_07156_),
    .A(_07152_),
    .B(_07155_));
 sg13g2_nand3_1 _32879_ (.B(_07152_),
    .C(_07155_),
    .A(net4747),
    .Y(_07157_));
 sg13g2_nor2b_1 _32880_ (.A(_07147_),
    .B_N(_07157_),
    .Y(_07158_));
 sg13g2_xnor2_1 _32881_ (.Y(_07159_),
    .A(net4804),
    .B(_07146_));
 sg13g2_a21o_1 _32882_ (.A2(_07155_),
    .A1(_07152_),
    .B1(net4748),
    .X(_07160_));
 sg13g2_and2_1 _32883_ (.A(_07157_),
    .B(_07160_),
    .X(_07161_));
 sg13g2_nand3_1 _32884_ (.B(_07159_),
    .C(_07160_),
    .A(_07157_),
    .Y(_07162_));
 sg13g2_nor3_1 _32885_ (.A(_04677_),
    .B(_05742_),
    .C(_06858_),
    .Y(_07163_));
 sg13g2_o21ai_1 _32886_ (.B1(_04677_),
    .Y(_07164_),
    .A1(_05742_),
    .A2(_06858_));
 sg13g2_nor2b_1 _32887_ (.A(_07163_),
    .B_N(_07164_),
    .Y(_07165_));
 sg13g2_nand3_1 _32888_ (.B(_06414_),
    .C(_06867_),
    .A(_04677_),
    .Y(_07166_));
 sg13g2_a21o_1 _32889_ (.A2(_06867_),
    .A1(_06414_),
    .B1(_04677_),
    .X(_07167_));
 sg13g2_nand3_1 _32890_ (.B(_07166_),
    .C(_07167_),
    .A(net5759),
    .Y(_07168_));
 sg13g2_a21oi_1 _32891_ (.A1(net5675),
    .A2(\u_inv.d_next[194] ),
    .Y(_07169_),
    .B1(net4958));
 sg13g2_nand2_1 _32892_ (.Y(_07170_),
    .A(_07168_),
    .B(_07169_));
 sg13g2_o21ai_1 _32893_ (.B1(_07170_),
    .Y(_07171_),
    .A1(net5048),
    .A2(_07165_));
 sg13g2_nand2b_1 _32894_ (.Y(_07172_),
    .B(net4747),
    .A_N(_07171_));
 sg13g2_xnor2_1 _32895_ (.Y(_07173_),
    .A(net4747),
    .B(_07171_));
 sg13g2_nand2_1 _32896_ (.Y(_07174_),
    .A(_04676_),
    .B(_07167_));
 sg13g2_xor2_1 _32897_ (.B(_07174_),
    .A(_04675_),
    .X(_07175_));
 sg13g2_a21oi_1 _32898_ (.A1(net5676),
    .A2(\u_inv.d_next[195] ),
    .Y(_07176_),
    .B1(net4958));
 sg13g2_o21ai_1 _32899_ (.B1(_07176_),
    .Y(_07177_),
    .A1(net5676),
    .A2(_07175_));
 sg13g2_nand3_1 _32900_ (.B(_05743_),
    .C(_07164_),
    .A(_04675_),
    .Y(_07178_));
 sg13g2_a21o_1 _32901_ (.A2(_07164_),
    .A1(_05743_),
    .B1(_04675_),
    .X(_07179_));
 sg13g2_nand3_1 _32902_ (.B(_07178_),
    .C(_07179_),
    .A(net4958),
    .Y(_07180_));
 sg13g2_nand3_1 _32903_ (.B(_07177_),
    .C(_07180_),
    .A(net4747),
    .Y(_07181_));
 sg13g2_a21o_1 _32904_ (.A2(_07180_),
    .A1(_07177_),
    .B1(net4747),
    .X(_07182_));
 sg13g2_and2_1 _32905_ (.A(_07181_),
    .B(_07182_),
    .X(_07183_));
 sg13g2_nand2_1 _32906_ (.Y(_07184_),
    .A(_07173_),
    .B(_07183_));
 sg13g2_nand3_1 _32907_ (.B(_04672_),
    .C(_06866_),
    .A(_04671_),
    .Y(_07185_));
 sg13g2_nand4_1 _32908_ (.B(_06412_),
    .C(_06867_),
    .A(net5759),
    .Y(_07186_),
    .D(_07185_));
 sg13g2_nand2_1 _32909_ (.Y(_07187_),
    .A(net5676),
    .B(\u_inv.d_next[193] ));
 sg13g2_and2_1 _32910_ (.A(net5048),
    .B(_07186_),
    .X(_07188_));
 sg13g2_a21oi_1 _32911_ (.A1(_04673_),
    .A2(_05703_),
    .Y(_07189_),
    .B1(_05740_));
 sg13g2_or2_1 _32912_ (.X(_07190_),
    .B(_07189_),
    .A(_04671_));
 sg13g2_a21oi_1 _32913_ (.A1(_04671_),
    .A2(_07189_),
    .Y(_07191_),
    .B1(net5051));
 sg13g2_a22oi_1 _32914_ (.Y(_07192_),
    .B1(_07190_),
    .B2(_07191_),
    .A2(_07188_),
    .A1(_07187_));
 sg13g2_a221oi_1 _32915_ (.B2(_07191_),
    .C1(net4804),
    .B1(_07190_),
    .A1(_07187_),
    .Y(_07193_),
    .A2(_07188_));
 sg13g2_xnor2_1 _32916_ (.Y(_07194_),
    .A(_04673_),
    .B(_05703_));
 sg13g2_a21oi_1 _32917_ (.A1(_04673_),
    .A2(_06362_),
    .Y(_07195_),
    .B1(net5676));
 sg13g2_nand2_1 _32918_ (.Y(_07196_),
    .A(_06866_),
    .B(_07195_));
 sg13g2_a21oi_1 _32919_ (.A1(net5676),
    .A2(\u_inv.d_next[192] ),
    .Y(_07197_),
    .B1(net4958));
 sg13g2_a22oi_1 _32920_ (.Y(_07198_),
    .B1(_07196_),
    .B2(_07197_),
    .A2(_07194_),
    .A1(net4958));
 sg13g2_nand2_1 _32921_ (.Y(_07199_),
    .A(net4747),
    .B(_07198_));
 sg13g2_nor2b_1 _32922_ (.A(_07193_),
    .B_N(_07199_),
    .Y(_07200_));
 sg13g2_nand2b_1 _32923_ (.Y(_07201_),
    .B(_07199_),
    .A_N(_07193_));
 sg13g2_nand4_1 _32924_ (.B(_07181_),
    .C(_07182_),
    .A(_07173_),
    .Y(_07202_),
    .D(_07201_));
 sg13g2_and2_1 _32925_ (.A(_07172_),
    .B(_07181_),
    .X(_07203_));
 sg13g2_nand2_1 _32926_ (.Y(_07204_),
    .A(_07202_),
    .B(_07203_));
 sg13g2_a21oi_1 _32927_ (.A1(_07202_),
    .A2(_07203_),
    .Y(_07205_),
    .B1(_07162_));
 sg13g2_nor2b_1 _32928_ (.A(_07205_),
    .B_N(_07158_),
    .Y(_07206_));
 sg13g2_nor2_1 _32929_ (.A(_07139_),
    .B(_07206_),
    .Y(_07207_));
 sg13g2_a21o_1 _32930_ (.A2(_07137_),
    .A1(_07125_),
    .B1(net4800),
    .X(_07208_));
 sg13g2_nor2b_1 _32931_ (.A(_07207_),
    .B_N(_07208_),
    .Y(_07209_));
 sg13g2_o21ai_1 _32932_ (.B1(_07208_),
    .Y(_07210_),
    .A1(_07139_),
    .A2(_07206_));
 sg13g2_nand3_1 _32933_ (.B(_07112_),
    .C(_07210_),
    .A(_07075_),
    .Y(_07211_));
 sg13g2_a21o_1 _32934_ (.A2(_07072_),
    .A1(_07062_),
    .B1(net4800),
    .X(_07212_));
 sg13g2_or3_1 _32935_ (.A(_07048_),
    .B(_07057_),
    .C(_07212_),
    .X(_07213_));
 sg13g2_a21oi_1 _32936_ (.A1(net4745),
    .A2(_07056_),
    .Y(_07214_),
    .B1(_07046_));
 sg13g2_o21ai_1 _32937_ (.B1(net4746),
    .Y(_07215_),
    .A1(_07102_),
    .A2(_07109_));
 sg13g2_a21oi_1 _32938_ (.A1(net4745),
    .A2(_07091_),
    .Y(_07216_),
    .B1(_07082_));
 sg13g2_o21ai_1 _32939_ (.B1(_07216_),
    .Y(_07217_),
    .A1(_07093_),
    .A2(_07215_));
 sg13g2_nand2_1 _32940_ (.Y(_07218_),
    .A(_07075_),
    .B(_07217_));
 sg13g2_and4_1 _32941_ (.A(_07211_),
    .B(_07213_),
    .C(_07214_),
    .D(_07218_),
    .X(_07219_));
 sg13g2_inv_1 _32942_ (.Y(_07220_),
    .A(_07219_));
 sg13g2_nor2b_1 _32943_ (.A(_07219_),
    .B_N(_07033_),
    .Y(_07221_));
 sg13g2_nand2_1 _32944_ (.Y(_07222_),
    .A(_06938_),
    .B(_06946_));
 sg13g2_nand3_1 _32945_ (.B(_06929_),
    .C(_07222_),
    .A(_06919_),
    .Y(_07223_));
 sg13g2_o21ai_1 _32946_ (.B1(net4738),
    .Y(_07224_),
    .A1(_06918_),
    .A2(_06928_));
 sg13g2_nand2_1 _32947_ (.Y(_07225_),
    .A(_07223_),
    .B(_07224_));
 sg13g2_nand2_1 _32948_ (.Y(_07226_),
    .A(_06911_),
    .B(_07225_));
 sg13g2_a21o_1 _32949_ (.A2(_06907_),
    .A1(_06900_),
    .B1(net4797),
    .X(_07227_));
 sg13g2_nand3b_1 _32950_ (.B(_06892_),
    .C(_06881_),
    .Y(_07228_),
    .A_N(_07227_));
 sg13g2_nand4_1 _32951_ (.B(_06891_),
    .C(_07226_),
    .A(_06880_),
    .Y(_07229_),
    .D(_07228_));
 sg13g2_and2_1 _32952_ (.A(_07018_),
    .B(_07026_),
    .X(_07230_));
 sg13g2_a21oi_1 _32953_ (.A1(net4743),
    .A2(_07001_),
    .Y(_07231_),
    .B1(_07008_));
 sg13g2_o21ai_1 _32954_ (.B1(_07231_),
    .Y(_07232_),
    .A1(_07010_),
    .A2(_07230_));
 sg13g2_o21ai_1 _32955_ (.B1(net4742),
    .Y(_07233_),
    .A1(_06983_),
    .A2(_06990_));
 sg13g2_o21ai_1 _32956_ (.B1(_06963_),
    .Y(_07234_),
    .A1(_06974_),
    .A2(_07233_));
 sg13g2_a221oi_1 _32957_ (.B2(_07232_),
    .C1(_07234_),
    .B1(_06993_),
    .A1(net4739),
    .Y(_07235_),
    .A2(_06972_));
 sg13g2_nor2_1 _32958_ (.A(_06950_),
    .B(_07235_),
    .Y(_07236_));
 sg13g2_nor3_2 _32959_ (.A(_07221_),
    .B(_07229_),
    .C(_07236_),
    .Y(_07237_));
 sg13g2_o21ai_1 _32960_ (.B1(_06839_),
    .Y(_07238_),
    .A1(net4792),
    .A2(_06850_));
 sg13g2_nand4_1 _32961_ (.B(_06822_),
    .C(_06832_),
    .A(_06821_),
    .Y(_07239_),
    .D(_07238_));
 sg13g2_nand3_1 _32962_ (.B(_06831_),
    .C(_07239_),
    .A(_06821_),
    .Y(_07240_));
 sg13g2_nand2b_1 _32963_ (.Y(_07241_),
    .B(_06788_),
    .A_N(_06779_));
 sg13g2_and2_1 _32964_ (.A(_06797_),
    .B(_06807_),
    .X(_07242_));
 sg13g2_inv_1 _32965_ (.Y(_07243_),
    .A(_07242_));
 sg13g2_a221oi_1 _32966_ (.B2(_06790_),
    .C1(_07241_),
    .B1(_07243_),
    .A1(_06811_),
    .Y(_07244_),
    .A2(_07240_));
 sg13g2_nor3_1 _32967_ (.A(_06720_),
    .B(_06760_),
    .C(_07244_),
    .Y(_07245_));
 sg13g2_o21ai_1 _32968_ (.B1(_06757_),
    .Y(_07246_),
    .A1(net4790),
    .A2(_06749_));
 sg13g2_nand2b_1 _32969_ (.Y(_07247_),
    .B(_06738_),
    .A_N(_06730_));
 sg13g2_a21oi_1 _32970_ (.A1(_06740_),
    .A2(_07246_),
    .Y(_07248_),
    .B1(_07247_));
 sg13g2_nor2_1 _32971_ (.A(_06720_),
    .B(_07248_),
    .Y(_07249_));
 sg13g2_nor2_1 _32972_ (.A(_06709_),
    .B(_06717_),
    .Y(_07250_));
 sg13g2_nor3_1 _32973_ (.A(_06686_),
    .B(_06698_),
    .C(_07250_),
    .Y(_07251_));
 sg13g2_nand2b_1 _32974_ (.Y(_07252_),
    .B(_06696_),
    .A_N(_06684_));
 sg13g2_or4_1 _32975_ (.A(_07245_),
    .B(_07249_),
    .C(_07251_),
    .D(_07252_),
    .X(_07253_));
 sg13g2_and3_1 _32976_ (.X(_07254_),
    .A(_06568_),
    .B(_06664_),
    .C(_07253_));
 sg13g2_a21o_1 _32977_ (.A2(_06660_),
    .A1(_06650_),
    .B1(net4789),
    .X(_07255_));
 sg13g2_nor4_1 _32978_ (.A(_06630_),
    .B(_06639_),
    .C(_06640_),
    .D(_07255_),
    .Y(_07256_));
 sg13g2_nor3_1 _32979_ (.A(_06629_),
    .B(_06639_),
    .C(_07256_),
    .Y(_07257_));
 sg13g2_nor4_1 _32980_ (.A(_06589_),
    .B(_06597_),
    .C(_06619_),
    .D(_07257_),
    .Y(_07258_));
 sg13g2_nor2_1 _32981_ (.A(_06604_),
    .B(_06616_),
    .Y(_07259_));
 sg13g2_nor3_1 _32982_ (.A(_06589_),
    .B(_06597_),
    .C(_07259_),
    .Y(_07260_));
 sg13g2_or4_1 _32983_ (.A(_06588_),
    .B(_06596_),
    .C(_07258_),
    .D(_07260_),
    .X(_07261_));
 sg13g2_and2_1 _32984_ (.A(_06568_),
    .B(_07261_),
    .X(_07262_));
 sg13g2_o21ai_1 _32985_ (.B1(_06554_),
    .Y(_07263_),
    .A1(net4787),
    .A2(_06563_));
 sg13g2_o21ai_1 _32986_ (.B1(_06544_),
    .Y(_07264_),
    .A1(net4787),
    .A2(_06536_));
 sg13g2_a21oi_1 _32987_ (.A1(_06546_),
    .A2(_07263_),
    .Y(_07265_),
    .B1(_07264_));
 sg13g2_nor3_1 _32988_ (.A(_06505_),
    .B(_06526_),
    .C(_07265_),
    .Y(_07266_));
 sg13g2_o21ai_1 _32989_ (.B1(net4731),
    .Y(_07267_),
    .A1(_06515_),
    .A2(_06522_));
 sg13g2_a21oi_1 _32990_ (.A1(net4731),
    .A2(_06503_),
    .Y(_07268_),
    .B1(_06493_));
 sg13g2_o21ai_1 _32991_ (.B1(_07268_),
    .Y(_07269_),
    .A1(_06505_),
    .A2(_07267_));
 sg13g2_nor4_2 _32992_ (.A(_07254_),
    .B(_07262_),
    .C(_07266_),
    .Y(_07270_),
    .D(_07269_));
 sg13g2_o21ai_1 _32993_ (.B1(_07270_),
    .Y(_07271_),
    .A1(_06857_),
    .A2(_07237_));
 sg13g2_nand2b_1 _32994_ (.Y(_07272_),
    .B(net4804),
    .A_N(_07192_));
 sg13g2_nor2b_1 _32995_ (.A(_07193_),
    .B_N(_07272_),
    .Y(_07273_));
 sg13g2_inv_1 _32996_ (.Y(_07274_),
    .A(_07273_));
 sg13g2_xnor2_1 _32997_ (.Y(_07275_),
    .A(net4747),
    .B(_07198_));
 sg13g2_nor3_1 _32998_ (.A(_07184_),
    .B(_07274_),
    .C(_07275_),
    .Y(_07276_));
 sg13g2_nor2_1 _32999_ (.A(_07139_),
    .B(_07162_),
    .Y(_07277_));
 sg13g2_nand2_2 _33000_ (.Y(_07278_),
    .A(_07276_),
    .B(_07277_));
 sg13g2_nor2_2 _33001_ (.A(_07113_),
    .B(_07278_),
    .Y(_07279_));
 sg13g2_nand2_2 _33002_ (.Y(_07280_),
    .A(_07033_),
    .B(_07279_));
 sg13g2_nor2_1 _33003_ (.A(_06857_),
    .B(_07280_),
    .Y(_07281_));
 sg13g2_a21oi_1 _33004_ (.A1(_05569_),
    .A2(_05690_),
    .Y(_07282_),
    .B1(_05699_));
 sg13g2_nand2b_1 _33005_ (.Y(_07283_),
    .B(_04904_),
    .A_N(_07282_));
 sg13g2_a21o_2 _33006_ (.A2(_07282_),
    .A1(_04912_),
    .B1(_04940_),
    .X(_07284_));
 sg13g2_a21oi_2 _33007_ (.B1(_04937_),
    .Y(_07285_),
    .A2(_07284_),
    .A1(_04833_));
 sg13g2_nor3_1 _33008_ (.A(_04805_),
    .B(_04808_),
    .C(_07285_),
    .Y(_07286_));
 sg13g2_nor2_1 _33009_ (.A(_04919_),
    .B(_07286_),
    .Y(_07287_));
 sg13g2_o21ai_1 _33010_ (.B1(_04799_),
    .Y(_07288_),
    .A1(_04919_),
    .A2(_07286_));
 sg13g2_nand2_1 _33011_ (.Y(_07289_),
    .A(_04922_),
    .B(_07288_));
 sg13g2_a21oi_1 _33012_ (.A1(_04922_),
    .A2(_07288_),
    .Y(_07290_),
    .B1(_04793_));
 sg13g2_xnor2_1 _33013_ (.Y(_07291_),
    .A(_04793_),
    .B(_07289_));
 sg13g2_a21o_2 _33014_ (.A2(_06277_),
    .A1(_06275_),
    .B1(_06302_),
    .X(_07292_));
 sg13g2_nand2b_2 _33015_ (.Y(_07293_),
    .B(_07292_),
    .A_N(_06317_));
 sg13g2_o21ai_1 _33016_ (.B1(_06329_),
    .Y(_07294_),
    .A1(_06297_),
    .A2(_07292_));
 sg13g2_a21oi_2 _33017_ (.B1(_06341_),
    .Y(_07295_),
    .A2(_07294_),
    .A1(_06290_));
 sg13g2_o21ai_1 _33018_ (.B1(_06344_),
    .Y(_07296_),
    .A1(_06283_),
    .A2(_07295_));
 sg13g2_a21oi_1 _33019_ (.A1(_06282_),
    .A2(_07296_),
    .Y(_07297_),
    .B1(_06346_));
 sg13g2_or2_1 _33020_ (.X(_07298_),
    .B(_07297_),
    .A(_06280_));
 sg13g2_a21o_1 _33021_ (.A2(_07298_),
    .A1(_06352_),
    .B1(_04794_),
    .X(_07299_));
 sg13g2_nand3_1 _33022_ (.B(_06352_),
    .C(_07298_),
    .A(_04794_),
    .Y(_07300_));
 sg13g2_nand3_1 _33023_ (.B(_07299_),
    .C(_07300_),
    .A(net5775),
    .Y(_07301_));
 sg13g2_a21oi_1 _33024_ (.A1(net5687),
    .A2(\u_inv.d_next[158] ),
    .Y(_07302_),
    .B1(net4972));
 sg13g2_nand2_1 _33025_ (.Y(_07303_),
    .A(_07301_),
    .B(_07302_));
 sg13g2_o21ai_1 _33026_ (.B1(_07303_),
    .Y(_07304_),
    .A1(net5062),
    .A2(_07291_));
 sg13g2_nand2b_1 _33027_ (.Y(_07305_),
    .B(net4760),
    .A_N(_07304_));
 sg13g2_inv_1 _33028_ (.Y(_07306_),
    .A(_07305_));
 sg13g2_xnor2_1 _33029_ (.Y(_07307_),
    .A(net4814),
    .B(_07304_));
 sg13g2_inv_1 _33030_ (.Y(_07308_),
    .A(_07307_));
 sg13g2_o21ai_1 _33031_ (.B1(_04790_),
    .Y(_07309_),
    .A1(_04924_),
    .A2(_07290_));
 sg13g2_or3_1 _33032_ (.A(_04790_),
    .B(_04924_),
    .C(_07290_),
    .X(_07310_));
 sg13g2_nand3_1 _33033_ (.B(_07309_),
    .C(_07310_),
    .A(net4971),
    .Y(_07311_));
 sg13g2_nand3_1 _33034_ (.B(_04792_),
    .C(_07299_),
    .A(_04791_),
    .Y(_07312_));
 sg13g2_a21o_1 _33035_ (.A2(_07299_),
    .A1(_04792_),
    .B1(_04791_),
    .X(_07313_));
 sg13g2_nand3_1 _33036_ (.B(_07312_),
    .C(_07313_),
    .A(net5776),
    .Y(_07314_));
 sg13g2_nand2_1 _33037_ (.Y(_07315_),
    .A(net5688),
    .B(\u_inv.d_next[159] ));
 sg13g2_nand3_1 _33038_ (.B(_07314_),
    .C(_07315_),
    .A(net5063),
    .Y(_07316_));
 sg13g2_and3_1 _33039_ (.X(_07317_),
    .A(net4760),
    .B(_07311_),
    .C(_07316_));
 sg13g2_nand3_1 _33040_ (.B(_07311_),
    .C(_07316_),
    .A(net4760),
    .Y(_07318_));
 sg13g2_a21oi_1 _33041_ (.A1(_07311_),
    .A2(_07316_),
    .Y(_07319_),
    .B1(net4760));
 sg13g2_nor2_1 _33042_ (.A(_07317_),
    .B(_07319_),
    .Y(_07320_));
 sg13g2_nor3_1 _33043_ (.A(_07307_),
    .B(_07317_),
    .C(_07319_),
    .Y(_07321_));
 sg13g2_o21ai_1 _33044_ (.B1(_04920_),
    .Y(_07322_),
    .A1(_04797_),
    .A2(_07287_));
 sg13g2_o21ai_1 _33045_ (.B1(net4972),
    .Y(_07323_),
    .A1(_04796_),
    .A2(_07322_));
 sg13g2_a21oi_1 _33046_ (.A1(_04796_),
    .A2(_07322_),
    .Y(_07324_),
    .B1(_07323_));
 sg13g2_nor2b_1 _33047_ (.A(_07297_),
    .B_N(_04797_),
    .Y(_07325_));
 sg13g2_a21oi_1 _33048_ (.A1(\u_inv.d_next[156] ),
    .A2(\u_inv.d_reg[156] ),
    .Y(_07326_),
    .B1(_07325_));
 sg13g2_xnor2_1 _33049_ (.Y(_07327_),
    .A(_04796_),
    .B(_07326_));
 sg13g2_nand2_1 _33050_ (.Y(_07328_),
    .A(net5687),
    .B(\u_inv.d_next[157] ));
 sg13g2_a21oi_1 _33051_ (.A1(net5775),
    .A2(_07327_),
    .Y(_07329_),
    .B1(net4971));
 sg13g2_a21o_1 _33052_ (.A2(_07329_),
    .A1(_07328_),
    .B1(_07324_),
    .X(_07330_));
 sg13g2_xnor2_1 _33053_ (.Y(_07331_),
    .A(net4760),
    .B(_07330_));
 sg13g2_xnor2_1 _33054_ (.Y(_07332_),
    .A(_04797_),
    .B(_07287_));
 sg13g2_xnor2_1 _33055_ (.Y(_07333_),
    .A(_04797_),
    .B(_07297_));
 sg13g2_nand2_1 _33056_ (.Y(_07334_),
    .A(net5775),
    .B(_07333_));
 sg13g2_a21oi_1 _33057_ (.A1(net5687),
    .A2(\u_inv.d_next[156] ),
    .Y(_07335_),
    .B1(net4971));
 sg13g2_a22oi_1 _33058_ (.Y(_07336_),
    .B1(_07334_),
    .B2(_07335_),
    .A2(_07332_),
    .A1(net4971));
 sg13g2_inv_1 _33059_ (.Y(_07337_),
    .A(_07336_));
 sg13g2_xnor2_1 _33060_ (.Y(_07338_),
    .A(net4814),
    .B(_07336_));
 sg13g2_nand2_1 _33061_ (.Y(_07339_),
    .A(_07331_),
    .B(_07338_));
 sg13g2_o21ai_1 _33062_ (.B1(_04915_),
    .Y(_07340_),
    .A1(_04808_),
    .A2(_07285_));
 sg13g2_xnor2_1 _33063_ (.Y(_07341_),
    .A(_04803_),
    .B(_07340_));
 sg13g2_a21oi_1 _33064_ (.A1(_04804_),
    .A2(_07296_),
    .Y(_07342_),
    .B1(net5687));
 sg13g2_o21ai_1 _33065_ (.B1(_07342_),
    .Y(_07343_),
    .A1(_04804_),
    .A2(_07296_));
 sg13g2_a21oi_1 _33066_ (.A1(net5687),
    .A2(\u_inv.d_next[154] ),
    .Y(_07344_),
    .B1(net4971));
 sg13g2_a22oi_1 _33067_ (.Y(_07345_),
    .B1(_07343_),
    .B2(_07344_),
    .A2(_07341_),
    .A1(net4971));
 sg13g2_and2_1 _33068_ (.A(net4759),
    .B(_07345_),
    .X(_07346_));
 sg13g2_xnor2_1 _33069_ (.Y(_07347_),
    .A(net4812),
    .B(_07345_));
 sg13g2_a21oi_1 _33070_ (.A1(_04803_),
    .A2(_07340_),
    .Y(_07348_),
    .B1(_04916_));
 sg13g2_or2_1 _33071_ (.X(_07349_),
    .B(_07348_),
    .A(_04801_));
 sg13g2_a21oi_1 _33072_ (.A1(_04801_),
    .A2(_07348_),
    .Y(_07350_),
    .B1(net5063));
 sg13g2_a21oi_1 _33073_ (.A1(_04804_),
    .A2(_07296_),
    .Y(_07351_),
    .B1(_04802_));
 sg13g2_o21ai_1 _33074_ (.B1(net5775),
    .Y(_07352_),
    .A1(_04801_),
    .A2(_07351_));
 sg13g2_a21o_1 _33075_ (.A2(_07351_),
    .A1(_04801_),
    .B1(_07352_),
    .X(_07353_));
 sg13g2_a21oi_1 _33076_ (.A1(net5687),
    .A2(\u_inv.d_next[155] ),
    .Y(_07354_),
    .B1(net4971));
 sg13g2_a22oi_1 _33077_ (.Y(_07355_),
    .B1(_07353_),
    .B2(_07354_),
    .A2(_07350_),
    .A1(_07349_));
 sg13g2_xnor2_1 _33078_ (.Y(_07356_),
    .A(net4812),
    .B(_07355_));
 sg13g2_nand2_1 _33079_ (.Y(_07357_),
    .A(_07347_),
    .B(_07356_));
 sg13g2_o21ai_1 _33080_ (.B1(_04913_),
    .Y(_07358_),
    .A1(_04807_),
    .A2(_07285_));
 sg13g2_o21ai_1 _33081_ (.B1(net4971),
    .Y(_07359_),
    .A1(_04806_),
    .A2(_07358_));
 sg13g2_a21oi_1 _33082_ (.A1(_04806_),
    .A2(_07358_),
    .Y(_07360_),
    .B1(_07359_));
 sg13g2_nor2b_1 _33083_ (.A(_07295_),
    .B_N(_04807_),
    .Y(_07361_));
 sg13g2_a21oi_1 _33084_ (.A1(\u_inv.d_next[152] ),
    .A2(\u_inv.d_reg[152] ),
    .Y(_07362_),
    .B1(_07361_));
 sg13g2_xnor2_1 _33085_ (.Y(_07363_),
    .A(_04806_),
    .B(_07362_));
 sg13g2_o21ai_1 _33086_ (.B1(net5063),
    .Y(_07364_),
    .A1(net5775),
    .A2(_14202_));
 sg13g2_a21oi_1 _33087_ (.A1(net5775),
    .A2(_07363_),
    .Y(_07365_),
    .B1(_07364_));
 sg13g2_nor2_2 _33088_ (.A(_07360_),
    .B(_07365_),
    .Y(_07366_));
 sg13g2_inv_1 _33089_ (.Y(_07367_),
    .A(_07366_));
 sg13g2_xor2_1 _33090_ (.B(_07295_),
    .A(_04807_),
    .X(_07368_));
 sg13g2_o21ai_1 _33091_ (.B1(net5063),
    .Y(_07369_),
    .A1(net5775),
    .A2(\u_inv.d_next[152] ));
 sg13g2_a21o_1 _33092_ (.A2(_07368_),
    .A1(net5775),
    .B1(_07369_),
    .X(_07370_));
 sg13g2_xnor2_1 _33093_ (.Y(_07371_),
    .A(_04807_),
    .B(_07285_));
 sg13g2_o21ai_1 _33094_ (.B1(_07370_),
    .Y(_07372_),
    .A1(net5062),
    .A2(_07371_));
 sg13g2_nand2_1 _33095_ (.Y(_07373_),
    .A(net4760),
    .B(_07372_));
 sg13g2_o21ai_1 _33096_ (.B1(net4762),
    .Y(_07374_),
    .A1(_07366_),
    .A2(_07372_));
 sg13g2_a21oi_1 _33097_ (.A1(net4759),
    .A2(_07355_),
    .Y(_07375_),
    .B1(_07346_));
 sg13g2_o21ai_1 _33098_ (.B1(_07375_),
    .Y(_07376_),
    .A1(_07357_),
    .A2(_07374_));
 sg13g2_nand4_1 _33099_ (.B(_07331_),
    .C(_07338_),
    .A(_07321_),
    .Y(_07377_),
    .D(_07376_));
 sg13g2_a21o_1 _33100_ (.A2(_07337_),
    .A1(_07330_),
    .B1(net4814),
    .X(_07378_));
 sg13g2_nand2b_1 _33101_ (.Y(_07379_),
    .B(_07321_),
    .A_N(_07378_));
 sg13g2_nand4_1 _33102_ (.B(_07318_),
    .C(_07377_),
    .A(_07305_),
    .Y(_07380_),
    .D(_07379_));
 sg13g2_xnor2_1 _33103_ (.Y(_07381_),
    .A(net4760),
    .B(_07366_));
 sg13g2_xnor2_1 _33104_ (.Y(_07382_),
    .A(net4762),
    .B(_07372_));
 sg13g2_inv_1 _33105_ (.Y(_07383_),
    .A(_07382_));
 sg13g2_nor3_1 _33106_ (.A(_07357_),
    .B(_07381_),
    .C(_07382_),
    .Y(_07384_));
 sg13g2_and4_1 _33107_ (.A(_07321_),
    .B(_07331_),
    .C(_07338_),
    .D(_07384_),
    .X(_07385_));
 sg13g2_nand4_1 _33108_ (.B(_07331_),
    .C(_07338_),
    .A(_07321_),
    .Y(_07386_),
    .D(_07384_));
 sg13g2_a21oi_1 _33109_ (.A1(_04832_),
    .A2(_07284_),
    .Y(_07387_),
    .B1(_04927_));
 sg13g2_nand3_1 _33110_ (.B(_04832_),
    .C(_07284_),
    .A(_04827_),
    .Y(_07388_));
 sg13g2_a21oi_1 _33111_ (.A1(_04930_),
    .A2(_07388_),
    .Y(_07389_),
    .B1(_04822_));
 sg13g2_nor3_1 _33112_ (.A(_04815_),
    .B(_04933_),
    .C(_07389_),
    .Y(_07390_));
 sg13g2_o21ai_1 _33113_ (.B1(_04815_),
    .Y(_07391_),
    .A1(_04933_),
    .A2(_07389_));
 sg13g2_nand2b_1 _33114_ (.Y(_07392_),
    .B(_07391_),
    .A_N(_07390_));
 sg13g2_and2_1 _33115_ (.A(_06286_),
    .B(_07294_),
    .X(_07393_));
 sg13g2_a221oi_1 _33116_ (.B2(_07294_),
    .C1(_06335_),
    .B1(_06286_),
    .A1(net5876),
    .Y(_07394_),
    .A2(\u_inv.d_reg[145] ));
 sg13g2_o21ai_1 _33117_ (.B1(_06334_),
    .Y(_07395_),
    .A1(_06287_),
    .A2(_07394_));
 sg13g2_a21oi_1 _33118_ (.A1(_06285_),
    .A2(_07395_),
    .Y(_07396_),
    .B1(_06331_));
 sg13g2_xnor2_1 _33119_ (.Y(_07397_),
    .A(_04814_),
    .B(_07396_));
 sg13g2_nand2_1 _33120_ (.Y(_07398_),
    .A(net5694),
    .B(\u_inv.d_next[150] ));
 sg13g2_a21oi_1 _33121_ (.A1(net5786),
    .A2(_07397_),
    .Y(_07399_),
    .B1(net4982));
 sg13g2_a22oi_1 _33122_ (.Y(_07400_),
    .B1(_07398_),
    .B2(_07399_),
    .A2(_07392_),
    .A1(net4982));
 sg13g2_and2_1 _33123_ (.A(net4761),
    .B(_07400_),
    .X(_07401_));
 sg13g2_xnor2_1 _33124_ (.Y(_07402_),
    .A(net4761),
    .B(_07400_));
 sg13g2_inv_2 _33125_ (.Y(_07403_),
    .A(_07402_));
 sg13g2_a21oi_1 _33126_ (.A1(_04934_),
    .A2(_07391_),
    .Y(_07404_),
    .B1(_04812_));
 sg13g2_nand3_1 _33127_ (.B(_04934_),
    .C(_07391_),
    .A(_04812_),
    .Y(_07405_));
 sg13g2_nor2_1 _33128_ (.A(net5070),
    .B(_07404_),
    .Y(_07406_));
 sg13g2_o21ai_1 _33129_ (.B1(_04813_),
    .Y(_07407_),
    .A1(_04815_),
    .A2(_07396_));
 sg13g2_xnor2_1 _33130_ (.Y(_07408_),
    .A(_04812_),
    .B(_07407_));
 sg13g2_nand2_1 _33131_ (.Y(_07409_),
    .A(net5694),
    .B(\u_inv.d_next[151] ));
 sg13g2_a21oi_1 _33132_ (.A1(net5786),
    .A2(_07408_),
    .Y(_07410_),
    .B1(net4982));
 sg13g2_a22oi_1 _33133_ (.Y(_07411_),
    .B1(_07409_),
    .B2(_07410_),
    .A2(_07406_),
    .A1(_07405_));
 sg13g2_xnor2_1 _33134_ (.Y(_07412_),
    .A(net4815),
    .B(_07411_));
 sg13g2_a21oi_1 _33135_ (.A1(_04930_),
    .A2(_07388_),
    .Y(_07413_),
    .B1(_04820_));
 sg13g2_nor2_1 _33136_ (.A(_04931_),
    .B(_07413_),
    .Y(_07414_));
 sg13g2_o21ai_1 _33137_ (.B1(_04817_),
    .Y(_07415_),
    .A1(_04931_),
    .A2(_07413_));
 sg13g2_a21oi_1 _33138_ (.A1(_04818_),
    .A2(_07414_),
    .Y(_07416_),
    .B1(net5070));
 sg13g2_a21oi_1 _33139_ (.A1(_04820_),
    .A2(_07395_),
    .Y(_07417_),
    .B1(_04819_));
 sg13g2_xnor2_1 _33140_ (.Y(_07418_),
    .A(_04817_),
    .B(_07417_));
 sg13g2_nand2_1 _33141_ (.Y(_07419_),
    .A(net5694),
    .B(\u_inv.d_next[149] ));
 sg13g2_a21oi_1 _33142_ (.A1(net5786),
    .A2(_07418_),
    .Y(_07420_),
    .B1(net4982));
 sg13g2_a22oi_1 _33143_ (.Y(_07421_),
    .B1(_07419_),
    .B2(_07420_),
    .A2(_07416_),
    .A1(_07415_));
 sg13g2_inv_1 _33144_ (.Y(_07422_),
    .A(_07421_));
 sg13g2_xnor2_1 _33145_ (.Y(_07423_),
    .A(net4814),
    .B(_07421_));
 sg13g2_xnor2_1 _33146_ (.Y(_07424_),
    .A(_04820_),
    .B(_07395_));
 sg13g2_o21ai_1 _33147_ (.B1(net5070),
    .Y(_07425_),
    .A1(net5786),
    .A2(\u_inv.d_next[148] ));
 sg13g2_a21o_1 _33148_ (.A2(_07424_),
    .A1(net5786),
    .B1(_07425_),
    .X(_07426_));
 sg13g2_nand3_1 _33149_ (.B(_04930_),
    .C(_07388_),
    .A(_04820_),
    .Y(_07427_));
 sg13g2_nand2b_1 _33150_ (.Y(_07428_),
    .B(_07427_),
    .A_N(_07413_));
 sg13g2_o21ai_1 _33151_ (.B1(_07426_),
    .Y(_07429_),
    .A1(net5070),
    .A2(_07428_));
 sg13g2_nand2_1 _33152_ (.Y(_07430_),
    .A(net4761),
    .B(_07429_));
 sg13g2_xnor2_1 _33153_ (.Y(_07431_),
    .A(net4814),
    .B(_07429_));
 sg13g2_and2_1 _33154_ (.A(_07423_),
    .B(_07431_),
    .X(_07432_));
 sg13g2_xnor2_1 _33155_ (.Y(_07433_),
    .A(_04826_),
    .B(_07387_));
 sg13g2_nor2b_1 _33156_ (.A(_07394_),
    .B_N(_04826_),
    .Y(_07434_));
 sg13g2_xnor2_1 _33157_ (.Y(_07435_),
    .A(_04826_),
    .B(_07394_));
 sg13g2_nand2_1 _33158_ (.Y(_07436_),
    .A(net5694),
    .B(\u_inv.d_next[146] ));
 sg13g2_a21oi_1 _33159_ (.A1(net5786),
    .A2(_07435_),
    .Y(_07437_),
    .B1(net4982));
 sg13g2_a22oi_1 _33160_ (.Y(_07438_),
    .B1(_07436_),
    .B2(_07437_),
    .A2(_07433_),
    .A1(net4983));
 sg13g2_and2_1 _33161_ (.A(net4761),
    .B(_07438_),
    .X(_07439_));
 sg13g2_xnor2_1 _33162_ (.Y(_07440_),
    .A(net4814),
    .B(_07438_));
 sg13g2_o21ai_1 _33163_ (.B1(_04928_),
    .Y(_07441_),
    .A1(_04826_),
    .A2(_07387_));
 sg13g2_nand2b_1 _33164_ (.Y(_07442_),
    .B(_04825_),
    .A_N(_07441_));
 sg13g2_a21oi_1 _33165_ (.A1(_04824_),
    .A2(_07441_),
    .Y(_07443_),
    .B1(net5073));
 sg13g2_a21o_1 _33166_ (.A2(\u_inv.d_reg[146] ),
    .A1(\u_inv.d_next[146] ),
    .B1(_07434_),
    .X(_07444_));
 sg13g2_xnor2_1 _33167_ (.Y(_07445_),
    .A(_04825_),
    .B(_07444_));
 sg13g2_nand2_1 _33168_ (.Y(_07446_),
    .A(net5694),
    .B(\u_inv.d_next[147] ));
 sg13g2_a21oi_1 _33169_ (.A1(net5786),
    .A2(_07445_),
    .Y(_07447_),
    .B1(net4982));
 sg13g2_a22oi_1 _33170_ (.Y(_07448_),
    .B1(_07446_),
    .B2(_07447_),
    .A2(_07443_),
    .A1(_07442_));
 sg13g2_xnor2_1 _33171_ (.Y(_07449_),
    .A(net4814),
    .B(_07448_));
 sg13g2_nand2_1 _33172_ (.Y(_07450_),
    .A(_07440_),
    .B(_07449_));
 sg13g2_xnor2_1 _33173_ (.Y(_07451_),
    .A(_04831_),
    .B(_07294_));
 sg13g2_o21ai_1 _33174_ (.B1(net5073),
    .Y(_07452_),
    .A1(net5786),
    .A2(\u_inv.d_next[144] ));
 sg13g2_a21o_1 _33175_ (.A2(_07451_),
    .A1(net5787),
    .B1(_07452_),
    .X(_07453_));
 sg13g2_nor2b_1 _33176_ (.A(_04831_),
    .B_N(_07284_),
    .Y(_07454_));
 sg13g2_xor2_1 _33177_ (.B(_07284_),
    .A(_04831_),
    .X(_07455_));
 sg13g2_o21ai_1 _33178_ (.B1(_07453_),
    .Y(_07456_),
    .A1(net5073),
    .A2(_07455_));
 sg13g2_nand2_1 _33179_ (.Y(_07457_),
    .A(net4761),
    .B(_07456_));
 sg13g2_nand2_1 _33180_ (.Y(_07458_),
    .A(_04828_),
    .B(_04830_));
 sg13g2_a21oi_1 _33181_ (.A1(_04831_),
    .A2(_07294_),
    .Y(_07459_),
    .B1(_07458_));
 sg13g2_or4_1 _33182_ (.A(net5693),
    .B(_06335_),
    .C(_07393_),
    .D(_07459_),
    .X(_07460_));
 sg13g2_a21oi_1 _33183_ (.A1(net5694),
    .A2(net5876),
    .Y(_07461_),
    .B1(net4982));
 sg13g2_nor2_1 _33184_ (.A(_04925_),
    .B(_07454_),
    .Y(_07462_));
 sg13g2_o21ai_1 _33185_ (.B1(net4983),
    .Y(_07463_),
    .A1(_04828_),
    .A2(_07462_));
 sg13g2_a21oi_1 _33186_ (.A1(_04828_),
    .A2(_07462_),
    .Y(_07464_),
    .B1(_07463_));
 sg13g2_a21oi_2 _33187_ (.B1(_07464_),
    .Y(_07465_),
    .A2(_07461_),
    .A1(_07460_));
 sg13g2_inv_1 _33188_ (.Y(_07466_),
    .A(_07465_));
 sg13g2_o21ai_1 _33189_ (.B1(net4761),
    .Y(_07467_),
    .A1(_07456_),
    .A2(_07465_));
 sg13g2_a21oi_1 _33190_ (.A1(net4761),
    .A2(_07448_),
    .Y(_07468_),
    .B1(_07439_));
 sg13g2_o21ai_1 _33191_ (.B1(_07468_),
    .Y(_07469_),
    .A1(_07450_),
    .A2(_07467_));
 sg13g2_nand4_1 _33192_ (.B(_07412_),
    .C(_07432_),
    .A(_07403_),
    .Y(_07470_),
    .D(_07469_));
 sg13g2_o21ai_1 _33193_ (.B1(net4762),
    .Y(_07471_),
    .A1(_07421_),
    .A2(_07429_));
 sg13g2_nand3b_1 _33194_ (.B(_07412_),
    .C(_07403_),
    .Y(_07472_),
    .A_N(_07471_));
 sg13g2_a21oi_1 _33195_ (.A1(net4761),
    .A2(_07411_),
    .Y(_07473_),
    .B1(_07401_));
 sg13g2_and3_1 _33196_ (.X(_07474_),
    .A(_07470_),
    .B(_07472_),
    .C(_07473_));
 sg13g2_nand3_1 _33197_ (.B(_07472_),
    .C(_07473_),
    .A(_07470_),
    .Y(_07475_));
 sg13g2_o21ai_1 _33198_ (.B1(_04911_),
    .Y(_07476_),
    .A1(_04905_),
    .A2(_07282_));
 sg13g2_and2_1 _33199_ (.A(_04838_),
    .B(_07476_),
    .X(_07477_));
 sg13g2_a21oi_1 _33200_ (.A1(_04838_),
    .A2(_07476_),
    .Y(_07478_),
    .B1(_04853_));
 sg13g2_nand2b_1 _33201_ (.Y(_07479_),
    .B(_04860_),
    .A_N(_07478_));
 sg13g2_o21ai_1 _33202_ (.B1(_04842_),
    .Y(_07480_),
    .A1(_04861_),
    .A2(_07478_));
 sg13g2_a21oi_1 _33203_ (.A1(_04857_),
    .A2(_07480_),
    .Y(_07481_),
    .B1(_04848_));
 sg13g2_a21o_1 _33204_ (.A2(_07480_),
    .A1(_04857_),
    .B1(_04848_),
    .X(_07482_));
 sg13g2_nand3_1 _33205_ (.B(_04857_),
    .C(_07480_),
    .A(_04848_),
    .Y(_07483_));
 sg13g2_a21oi_1 _33206_ (.A1(_07482_),
    .A2(_07483_),
    .Y(_07484_),
    .B1(net5072));
 sg13g2_a21o_2 _33207_ (.A2(_07293_),
    .A1(_06295_),
    .B1(_06324_),
    .X(_07485_));
 sg13g2_a21oi_2 _33208_ (.B1(_06326_),
    .Y(_07486_),
    .A2(_07485_),
    .A1(_06296_));
 sg13g2_nor2_1 _33209_ (.A(_06293_),
    .B(_07486_),
    .Y(_07487_));
 sg13g2_or3_1 _33210_ (.A(_04848_),
    .B(_06320_),
    .C(_07487_),
    .X(_07488_));
 sg13g2_o21ai_1 _33211_ (.B1(_04848_),
    .Y(_07489_),
    .A1(_06320_),
    .A2(_07487_));
 sg13g2_nand3_1 _33212_ (.B(_07488_),
    .C(_07489_),
    .A(net5788),
    .Y(_07490_));
 sg13g2_a21oi_1 _33213_ (.A1(net5695),
    .A2(\u_inv.d_next[142] ),
    .Y(_07491_),
    .B1(net4982));
 sg13g2_a21o_2 _33214_ (.A2(_07491_),
    .A1(_07490_),
    .B1(_07484_),
    .X(_07492_));
 sg13g2_nand2b_1 _33215_ (.Y(_07493_),
    .B(net4766),
    .A_N(_07492_));
 sg13g2_inv_1 _33216_ (.Y(_07494_),
    .A(_07493_));
 sg13g2_nand2_1 _33217_ (.Y(_07495_),
    .A(net4816),
    .B(_07492_));
 sg13g2_xnor2_1 _33218_ (.Y(_07496_),
    .A(net4816),
    .B(_07492_));
 sg13g2_o21ai_1 _33219_ (.B1(_04845_),
    .Y(_07497_),
    .A1(_04862_),
    .A2(_07481_));
 sg13g2_or3_1 _33220_ (.A(_04845_),
    .B(_04862_),
    .C(_07481_),
    .X(_07498_));
 sg13g2_nand3_1 _33221_ (.B(_07497_),
    .C(_07498_),
    .A(net4984),
    .Y(_07499_));
 sg13g2_nand2_1 _33222_ (.Y(_07500_),
    .A(_04847_),
    .B(_07489_));
 sg13g2_xnor2_1 _33223_ (.Y(_07501_),
    .A(_04846_),
    .B(_07500_));
 sg13g2_o21ai_1 _33224_ (.B1(net5072),
    .Y(_07502_),
    .A1(net5788),
    .A2(_14206_));
 sg13g2_a21o_1 _33225_ (.A2(_07501_),
    .A1(net5788),
    .B1(_07502_),
    .X(_07503_));
 sg13g2_and3_2 _33226_ (.X(_07504_),
    .A(net4766),
    .B(_07499_),
    .C(_07503_));
 sg13g2_a21oi_1 _33227_ (.A1(_07499_),
    .A2(_07503_),
    .Y(_07505_),
    .B1(net4766));
 sg13g2_nor2_1 _33228_ (.A(_07504_),
    .B(_07505_),
    .Y(_07506_));
 sg13g2_or3_1 _33229_ (.A(_07496_),
    .B(_07504_),
    .C(_07505_),
    .X(_07507_));
 sg13g2_o21ai_1 _33230_ (.B1(_04841_),
    .Y(_07508_),
    .A1(_04861_),
    .A2(_07478_));
 sg13g2_a21o_1 _33231_ (.A2(_07508_),
    .A1(_04856_),
    .B1(_04839_),
    .X(_07509_));
 sg13g2_nand3_1 _33232_ (.B(_04856_),
    .C(_07508_),
    .A(_04839_),
    .Y(_07510_));
 sg13g2_nand3_1 _33233_ (.B(_07509_),
    .C(_07510_),
    .A(net4984),
    .Y(_07511_));
 sg13g2_o21ai_1 _33234_ (.B1(_04840_),
    .Y(_07512_),
    .A1(_04841_),
    .A2(_07486_));
 sg13g2_xnor2_1 _33235_ (.Y(_07513_),
    .A(_04839_),
    .B(_07512_));
 sg13g2_a21oi_1 _33236_ (.A1(net5788),
    .A2(_07513_),
    .Y(_07514_),
    .B1(net4985));
 sg13g2_o21ai_1 _33237_ (.B1(_07514_),
    .Y(_07515_),
    .A1(net5788),
    .A2(_14207_));
 sg13g2_nand2_1 _33238_ (.Y(_07516_),
    .A(_07511_),
    .B(_07515_));
 sg13g2_nand3_1 _33239_ (.B(_07511_),
    .C(_07515_),
    .A(net4766),
    .Y(_07517_));
 sg13g2_a21o_1 _33240_ (.A2(_07515_),
    .A1(_07511_),
    .B1(net4766),
    .X(_07518_));
 sg13g2_and2_1 _33241_ (.A(_07517_),
    .B(_07518_),
    .X(_07519_));
 sg13g2_xnor2_1 _33242_ (.Y(_07520_),
    .A(_04841_),
    .B(_07479_));
 sg13g2_a21oi_1 _33243_ (.A1(_04841_),
    .A2(_07486_),
    .Y(_07521_),
    .B1(net5695));
 sg13g2_o21ai_1 _33244_ (.B1(_07521_),
    .Y(_07522_),
    .A1(_04841_),
    .A2(_07486_));
 sg13g2_a21oi_1 _33245_ (.A1(net5695),
    .A2(\u_inv.d_next[140] ),
    .Y(_07523_),
    .B1(net4984));
 sg13g2_a22oi_1 _33246_ (.Y(_07524_),
    .B1(_07522_),
    .B2(_07523_),
    .A2(_07520_),
    .A1(net4985));
 sg13g2_nand2_1 _33247_ (.Y(_07525_),
    .A(net4766),
    .B(_07524_));
 sg13g2_xnor2_1 _33248_ (.Y(_07526_),
    .A(net4816),
    .B(_07524_));
 sg13g2_nand3_1 _33249_ (.B(_07518_),
    .C(_07526_),
    .A(_07517_),
    .Y(_07527_));
 sg13g2_nor4_1 _33250_ (.A(_07496_),
    .B(_07504_),
    .C(_07505_),
    .D(_07527_),
    .Y(_07528_));
 sg13g2_o21ai_1 _33251_ (.B1(_04858_),
    .Y(_07529_),
    .A1(_04852_),
    .A2(_07477_));
 sg13g2_and2_1 _33252_ (.A(_04850_),
    .B(_07529_),
    .X(_07530_));
 sg13g2_o21ai_1 _33253_ (.B1(net4984),
    .Y(_07531_),
    .A1(_04850_),
    .A2(_07529_));
 sg13g2_a21oi_1 _33254_ (.A1(_04852_),
    .A2(_07485_),
    .Y(_07532_),
    .B1(_04851_));
 sg13g2_xnor2_1 _33255_ (.Y(_07533_),
    .A(_04850_),
    .B(_07532_));
 sg13g2_a21oi_1 _33256_ (.A1(net5789),
    .A2(_07533_),
    .Y(_07534_),
    .B1(net4984));
 sg13g2_o21ai_1 _33257_ (.B1(_07534_),
    .Y(_07535_),
    .A1(net5789),
    .A2(_14208_));
 sg13g2_o21ai_1 _33258_ (.B1(_07535_),
    .Y(_07536_),
    .A1(_07530_),
    .A2(_07531_));
 sg13g2_xnor2_1 _33259_ (.Y(_07537_),
    .A(net4767),
    .B(_07536_));
 sg13g2_xor2_1 _33260_ (.B(_07477_),
    .A(_04852_),
    .X(_07538_));
 sg13g2_xnor2_1 _33261_ (.Y(_07539_),
    .A(_04852_),
    .B(_07485_));
 sg13g2_a21oi_1 _33262_ (.A1(net5695),
    .A2(\u_inv.d_next[138] ),
    .Y(_07540_),
    .B1(net4984));
 sg13g2_o21ai_1 _33263_ (.B1(_07540_),
    .Y(_07541_),
    .A1(net5695),
    .A2(_07539_));
 sg13g2_o21ai_1 _33264_ (.B1(_07541_),
    .Y(_07542_),
    .A1(net5072),
    .A2(_07538_));
 sg13g2_nor2_1 _33265_ (.A(net4816),
    .B(_07542_),
    .Y(_07543_));
 sg13g2_xnor2_1 _33266_ (.Y(_07544_),
    .A(net4767),
    .B(_07542_));
 sg13g2_inv_1 _33267_ (.Y(_07545_),
    .A(_07544_));
 sg13g2_nand2_1 _33268_ (.Y(_07546_),
    .A(_07537_),
    .B(_07544_));
 sg13g2_nand2_1 _33269_ (.Y(_07547_),
    .A(_04909_),
    .B(_07293_));
 sg13g2_xnor2_1 _33270_ (.Y(_07548_),
    .A(_04909_),
    .B(_07293_));
 sg13g2_o21ai_1 _33271_ (.B1(net5072),
    .Y(_07549_),
    .A1(net5788),
    .A2(\u_inv.d_next[136] ));
 sg13g2_a21o_1 _33272_ (.A2(_07548_),
    .A1(net5788),
    .B1(_07549_),
    .X(_07550_));
 sg13g2_xnor2_1 _33273_ (.Y(_07551_),
    .A(_04910_),
    .B(_07283_));
 sg13g2_o21ai_1 _33274_ (.B1(_07550_),
    .Y(_07552_),
    .A1(net5072),
    .A2(_07551_));
 sg13g2_and2_1 _33275_ (.A(net4766),
    .B(_07552_),
    .X(_07553_));
 sg13g2_xnor2_1 _33276_ (.Y(_07554_),
    .A(net4816),
    .B(_07552_));
 sg13g2_xnor2_1 _33277_ (.Y(_07555_),
    .A(net4766),
    .B(_07552_));
 sg13g2_a21o_1 _33278_ (.A2(_07283_),
    .A1(_04910_),
    .B1(_04835_),
    .X(_07556_));
 sg13g2_o21ai_1 _33279_ (.B1(net4984),
    .Y(_07557_),
    .A1(_04907_),
    .A2(_07556_));
 sg13g2_a21oi_1 _33280_ (.A1(_04907_),
    .A2(_07556_),
    .Y(_07558_),
    .B1(_07557_));
 sg13g2_nand3_1 _33281_ (.B(_04908_),
    .C(_07547_),
    .A(_04906_),
    .Y(_07559_));
 sg13g2_a21o_1 _33282_ (.A2(_07547_),
    .A1(_04908_),
    .B1(_04906_),
    .X(_07560_));
 sg13g2_nand3_1 _33283_ (.B(_07559_),
    .C(_07560_),
    .A(net5788),
    .Y(_07561_));
 sg13g2_a21oi_1 _33284_ (.A1(net5695),
    .A2(\u_inv.d_next[137] ),
    .Y(_07562_),
    .B1(net4984));
 sg13g2_a21oi_2 _33285_ (.B1(_07558_),
    .Y(_07563_),
    .A2(_07562_),
    .A1(_07561_));
 sg13g2_inv_1 _33286_ (.Y(_07564_),
    .A(_07563_));
 sg13g2_nand2_1 _33287_ (.Y(_07565_),
    .A(net4816),
    .B(_07564_));
 sg13g2_xnor2_1 _33288_ (.Y(_07566_),
    .A(net4818),
    .B(_07563_));
 sg13g2_nand4_1 _33289_ (.B(_07544_),
    .C(_07554_),
    .A(_07537_),
    .Y(_07567_),
    .D(_07566_));
 sg13g2_a21o_1 _33290_ (.A2(_05690_),
    .A1(_05569_),
    .B1(_05697_),
    .X(_07568_));
 sg13g2_nand2_1 _33291_ (.Y(_07569_),
    .A(_04892_),
    .B(_07568_));
 sg13g2_a21oi_1 _33292_ (.A1(_04892_),
    .A2(_07568_),
    .Y(_07570_),
    .B1(_04886_));
 sg13g2_nor2_1 _33293_ (.A(_04895_),
    .B(_07570_),
    .Y(_07571_));
 sg13g2_o21ai_1 _33294_ (.B1(_04880_),
    .Y(_07572_),
    .A1(_04895_),
    .A2(_07570_));
 sg13g2_a21oi_1 _33295_ (.A1(_04899_),
    .A2(_07572_),
    .Y(_07573_),
    .B1(_04872_));
 sg13g2_o21ai_1 _33296_ (.B1(_04869_),
    .Y(_07574_),
    .A1(_04901_),
    .A2(_07573_));
 sg13g2_or3_1 _33297_ (.A(_04869_),
    .B(_04901_),
    .C(_07573_),
    .X(_07575_));
 sg13g2_nand3_1 _33298_ (.B(_07574_),
    .C(_07575_),
    .A(net4986),
    .Y(_07576_));
 sg13g2_a21oi_1 _33299_ (.A1(_06275_),
    .A2(_06277_),
    .Y(_07577_),
    .B1(_05696_));
 sg13g2_nand2_1 _33300_ (.Y(_07578_),
    .A(_05693_),
    .B(_07577_));
 sg13g2_nand3_1 _33301_ (.B(_06300_),
    .C(_07577_),
    .A(_05693_),
    .Y(_07579_));
 sg13g2_a21o_1 _33302_ (.A2(_07579_),
    .A1(_06311_),
    .B1(_04879_),
    .X(_07580_));
 sg13g2_nand2b_1 _33303_ (.Y(_07581_),
    .B(_04876_),
    .A_N(_07580_));
 sg13g2_a21o_1 _33304_ (.A2(_07581_),
    .A1(_06313_),
    .B1(_04873_),
    .X(_07582_));
 sg13g2_nand3_1 _33305_ (.B(_04871_),
    .C(_07582_),
    .A(_04870_),
    .Y(_07583_));
 sg13g2_a21o_1 _33306_ (.A2(_07582_),
    .A1(_04871_),
    .B1(_04870_),
    .X(_07584_));
 sg13g2_nand3_1 _33307_ (.B(_07583_),
    .C(_07584_),
    .A(net5789),
    .Y(_07585_));
 sg13g2_a21oi_1 _33308_ (.A1(net5695),
    .A2(\u_inv.d_next[135] ),
    .Y(_07586_),
    .B1(net4987));
 sg13g2_nand2_1 _33309_ (.Y(_07587_),
    .A(_07585_),
    .B(_07586_));
 sg13g2_and3_2 _33310_ (.X(_07588_),
    .A(net4771),
    .B(_07576_),
    .C(_07587_));
 sg13g2_a21oi_1 _33311_ (.A1(_07576_),
    .A2(_07587_),
    .Y(_07589_),
    .B1(net4770));
 sg13g2_or2_1 _33312_ (.X(_07590_),
    .B(_07589_),
    .A(_07588_));
 sg13g2_nand3_1 _33313_ (.B(_04899_),
    .C(_07572_),
    .A(_04872_),
    .Y(_07591_));
 sg13g2_nand2b_1 _33314_ (.Y(_07592_),
    .B(_07591_),
    .A_N(_07573_));
 sg13g2_nand3_1 _33315_ (.B(_06313_),
    .C(_07581_),
    .A(_04873_),
    .Y(_07593_));
 sg13g2_and2_1 _33316_ (.A(net5789),
    .B(_07582_),
    .X(_07594_));
 sg13g2_nand2_1 _33317_ (.Y(_07595_),
    .A(net5695),
    .B(\u_inv.d_next[134] ));
 sg13g2_a21oi_1 _33318_ (.A1(_07593_),
    .A2(_07594_),
    .Y(_07596_),
    .B1(net4985));
 sg13g2_a22oi_1 _33319_ (.Y(_07597_),
    .B1(_07595_),
    .B2(_07596_),
    .A2(_07592_),
    .A1(net4987));
 sg13g2_and2_1 _33320_ (.A(net4770),
    .B(_07597_),
    .X(_07598_));
 sg13g2_nand2b_1 _33321_ (.Y(_07599_),
    .B(net4819),
    .A_N(_07597_));
 sg13g2_xnor2_1 _33322_ (.Y(_07600_),
    .A(net4770),
    .B(_07597_));
 sg13g2_nor3_1 _33323_ (.A(_07588_),
    .B(_07589_),
    .C(_07600_),
    .Y(_07601_));
 sg13g2_o21ai_1 _33324_ (.B1(_04879_),
    .Y(_07602_),
    .A1(_04895_),
    .A2(_07570_));
 sg13g2_a21o_1 _33325_ (.A2(_07602_),
    .A1(_04897_),
    .B1(_04875_),
    .X(_07603_));
 sg13g2_nand3_1 _33326_ (.B(_04897_),
    .C(_07602_),
    .A(_04875_),
    .Y(_07604_));
 sg13g2_nand3_1 _33327_ (.B(_07603_),
    .C(_07604_),
    .A(net4985),
    .Y(_07605_));
 sg13g2_nand2_1 _33328_ (.Y(_07606_),
    .A(_04877_),
    .B(_07580_));
 sg13g2_xnor2_1 _33329_ (.Y(_07607_),
    .A(_04875_),
    .B(_07606_));
 sg13g2_a21oi_1 _33330_ (.A1(net5789),
    .A2(_07607_),
    .Y(_07608_),
    .B1(net4985));
 sg13g2_o21ai_1 _33331_ (.B1(_07608_),
    .Y(_07609_),
    .A1(net5789),
    .A2(_14211_));
 sg13g2_and2_1 _33332_ (.A(_07605_),
    .B(_07609_),
    .X(_07610_));
 sg13g2_inv_1 _33333_ (.Y(_07611_),
    .A(_07610_));
 sg13g2_nand3_1 _33334_ (.B(_07605_),
    .C(_07609_),
    .A(net4770),
    .Y(_07612_));
 sg13g2_a21o_1 _33335_ (.A2(_07609_),
    .A1(_07605_),
    .B1(net4770),
    .X(_07613_));
 sg13g2_and2_1 _33336_ (.A(_07612_),
    .B(_07613_),
    .X(_07614_));
 sg13g2_xnor2_1 _33337_ (.Y(_07615_),
    .A(_04878_),
    .B(_07571_));
 sg13g2_nand3_1 _33338_ (.B(_06311_),
    .C(_07579_),
    .A(_04879_),
    .Y(_07616_));
 sg13g2_nand3_1 _33339_ (.B(_07580_),
    .C(_07616_),
    .A(net5789),
    .Y(_07617_));
 sg13g2_a21oi_1 _33340_ (.A1(net5696),
    .A2(\u_inv.d_next[132] ),
    .Y(_07618_),
    .B1(net4985));
 sg13g2_a22oi_1 _33341_ (.Y(_07619_),
    .B1(_07617_),
    .B2(_07618_),
    .A2(_07615_),
    .A1(net4985));
 sg13g2_nand2_1 _33342_ (.Y(_07620_),
    .A(net4770),
    .B(_07619_));
 sg13g2_xnor2_1 _33343_ (.Y(_07621_),
    .A(net4819),
    .B(_07619_));
 sg13g2_nand3_1 _33344_ (.B(_07613_),
    .C(_07621_),
    .A(_07612_),
    .Y(_07622_));
 sg13g2_nor4_1 _33345_ (.A(_07588_),
    .B(_07589_),
    .C(_07600_),
    .D(_07622_),
    .Y(_07623_));
 sg13g2_xnor2_1 _33346_ (.Y(_07624_),
    .A(_04884_),
    .B(_07569_));
 sg13g2_a21o_1 _33347_ (.A2(_07578_),
    .A1(_06308_),
    .B1(_04884_),
    .X(_07625_));
 sg13g2_nand3_1 _33348_ (.B(_06308_),
    .C(_07578_),
    .A(_04884_),
    .Y(_07626_));
 sg13g2_and2_1 _33349_ (.A(_07625_),
    .B(_07626_),
    .X(_07627_));
 sg13g2_nand2_1 _33350_ (.Y(_07628_),
    .A(net5700),
    .B(\u_inv.d_next[130] ));
 sg13g2_a21oi_1 _33351_ (.A1(net5800),
    .A2(_07627_),
    .Y(_07629_),
    .B1(net4994));
 sg13g2_a22oi_1 _33352_ (.Y(_07630_),
    .B1(_07628_),
    .B2(_07629_),
    .A2(_07624_),
    .A1(net4994));
 sg13g2_and2_1 _33353_ (.A(net4770),
    .B(_07630_),
    .X(_07631_));
 sg13g2_nand2b_1 _33354_ (.Y(_07632_),
    .B(net4819),
    .A_N(_07630_));
 sg13g2_nand2b_1 _33355_ (.Y(_07633_),
    .B(_07632_),
    .A_N(_07631_));
 sg13g2_a21oi_1 _33356_ (.A1(_04884_),
    .A2(_07569_),
    .Y(_07634_),
    .B1(_04893_));
 sg13g2_and2_1 _33357_ (.A(net5619),
    .B(_07634_),
    .X(_07635_));
 sg13g2_o21ai_1 _33358_ (.B1(net4994),
    .Y(_07636_),
    .A1(net5619),
    .A2(_07634_));
 sg13g2_nand3_1 _33359_ (.B(_04883_),
    .C(_07625_),
    .A(net5619),
    .Y(_07637_));
 sg13g2_a21o_1 _33360_ (.A2(_07625_),
    .A1(_04883_),
    .B1(net5619),
    .X(_07638_));
 sg13g2_nand3_1 _33361_ (.B(_07637_),
    .C(_07638_),
    .A(net5800),
    .Y(_07639_));
 sg13g2_a21oi_1 _33362_ (.A1(net5700),
    .A2(\u_inv.d_next[131] ),
    .Y(_07640_),
    .B1(net4994));
 sg13g2_nand2_1 _33363_ (.Y(_07641_),
    .A(_07639_),
    .B(_07640_));
 sg13g2_o21ai_1 _33364_ (.B1(_07641_),
    .Y(_07642_),
    .A1(_07635_),
    .A2(_07636_));
 sg13g2_nor2_1 _33365_ (.A(net4819),
    .B(_07642_),
    .Y(_07643_));
 sg13g2_xnor2_1 _33366_ (.Y(_07644_),
    .A(net4770),
    .B(_07642_));
 sg13g2_nand2b_1 _33367_ (.Y(_07645_),
    .B(_07644_),
    .A_N(_07633_));
 sg13g2_nand3b_1 _33368_ (.B(_05692_),
    .C(_05694_),
    .Y(_07646_),
    .A_N(_07577_));
 sg13g2_nor2_1 _33369_ (.A(net5700),
    .B(_06306_),
    .Y(_07647_));
 sg13g2_nand3_1 _33370_ (.B(_07646_),
    .C(_07647_),
    .A(_07578_),
    .Y(_07648_));
 sg13g2_nand2_1 _33371_ (.Y(_07649_),
    .A(net5700),
    .B(\u_inv.d_next[129] ));
 sg13g2_a21oi_1 _33372_ (.A1(_07648_),
    .A2(_07649_),
    .Y(_07650_),
    .B1(net4994));
 sg13g2_o21ai_1 _33373_ (.B1(_04889_),
    .Y(_07651_),
    .A1(_05691_),
    .A2(_05695_));
 sg13g2_xnor2_1 _33374_ (.Y(_07652_),
    .A(_05693_),
    .B(_07651_));
 sg13g2_a21oi_2 _33375_ (.B1(_07650_),
    .Y(_07653_),
    .A2(_07652_),
    .A1(net4994));
 sg13g2_nor2_1 _33376_ (.A(net4819),
    .B(_07653_),
    .Y(_07654_));
 sg13g2_xnor2_1 _33377_ (.Y(_07655_),
    .A(_05695_),
    .B(_06278_));
 sg13g2_o21ai_1 _33378_ (.B1(net5084),
    .Y(_07656_),
    .A1(net5800),
    .A2(\u_inv.d_next[128] ));
 sg13g2_a21o_1 _33379_ (.A2(_07655_),
    .A1(net5800),
    .B1(_07656_),
    .X(_07657_));
 sg13g2_xnor2_1 _33380_ (.Y(_07658_),
    .A(_05691_),
    .B(_05695_));
 sg13g2_o21ai_1 _33381_ (.B1(_07657_),
    .Y(_07659_),
    .A1(net5084),
    .A2(_07658_));
 sg13g2_and2_1 _33382_ (.A(net4772),
    .B(_07659_),
    .X(_07660_));
 sg13g2_nor2_1 _33383_ (.A(_07654_),
    .B(_07660_),
    .Y(_07661_));
 sg13g2_nor2_1 _33384_ (.A(_07631_),
    .B(_07643_),
    .Y(_07662_));
 sg13g2_o21ai_1 _33385_ (.B1(_07662_),
    .Y(_07663_),
    .A1(_07645_),
    .A2(_07661_));
 sg13g2_and2_1 _33386_ (.A(_07612_),
    .B(_07620_),
    .X(_07664_));
 sg13g2_nand2_1 _33387_ (.Y(_07665_),
    .A(_07612_),
    .B(_07620_));
 sg13g2_or2_1 _33388_ (.X(_07666_),
    .B(_07598_),
    .A(_07588_));
 sg13g2_a221oi_1 _33389_ (.B2(_07601_),
    .C1(_07666_),
    .B1(_07665_),
    .A1(_07623_),
    .Y(_07667_),
    .A2(_07663_));
 sg13g2_nor4_1 _33390_ (.A(_07507_),
    .B(_07527_),
    .C(_07567_),
    .D(_07667_),
    .Y(_07668_));
 sg13g2_a21oi_1 _33391_ (.A1(net4767),
    .A2(_07563_),
    .Y(_07669_),
    .B1(_07553_));
 sg13g2_a21o_1 _33392_ (.A2(_07542_),
    .A1(_07536_),
    .B1(net4818),
    .X(_07670_));
 sg13g2_o21ai_1 _33393_ (.B1(_07670_),
    .Y(_07671_),
    .A1(_07546_),
    .A2(_07669_));
 sg13g2_and2_1 _33394_ (.A(_07528_),
    .B(_07671_),
    .X(_07672_));
 sg13g2_and2_1 _33395_ (.A(_07517_),
    .B(_07525_),
    .X(_07673_));
 sg13g2_o21ai_1 _33396_ (.B1(_07493_),
    .Y(_07674_),
    .A1(_07507_),
    .A2(_07673_));
 sg13g2_nor4_2 _33397_ (.A(_07504_),
    .B(_07668_),
    .C(_07672_),
    .Y(_07675_),
    .D(_07674_));
 sg13g2_xnor2_1 _33398_ (.Y(_07676_),
    .A(net4762),
    .B(_07456_));
 sg13g2_xnor2_1 _33399_ (.Y(_07677_),
    .A(net4762),
    .B(_07465_));
 sg13g2_nor3_1 _33400_ (.A(_07450_),
    .B(_07676_),
    .C(_07677_),
    .Y(_07678_));
 sg13g2_inv_1 _33401_ (.Y(_07679_),
    .A(_07678_));
 sg13g2_nand4_1 _33402_ (.B(_07412_),
    .C(_07432_),
    .A(_07403_),
    .Y(_07680_),
    .D(_07678_));
 sg13g2_o21ai_1 _33403_ (.B1(_07474_),
    .Y(_07681_),
    .A1(_07675_),
    .A2(_07680_));
 sg13g2_a21oi_2 _33404_ (.B1(_07380_),
    .Y(_07682_),
    .A2(_07681_),
    .A1(_07385_));
 sg13g2_a21o_2 _33405_ (.A2(_07681_),
    .A1(_07385_),
    .B1(_07380_),
    .X(_07683_));
 sg13g2_a21oi_2 _33406_ (.B1(_05700_),
    .Y(_07684_),
    .A2(_05690_),
    .A1(_05569_));
 sg13g2_nand2b_2 _33407_ (.Y(_07685_),
    .B(_04943_),
    .A_N(_07684_));
 sg13g2_o21ai_1 _33408_ (.B1(_04784_),
    .Y(_07686_),
    .A1(_04944_),
    .A2(_07684_));
 sg13g2_o21ai_1 _33409_ (.B1(_04785_),
    .Y(_07687_),
    .A1(_04944_),
    .A2(_07684_));
 sg13g2_a21oi_2 _33410_ (.B1(_04976_),
    .Y(_07688_),
    .A2(_07685_),
    .A1(_04787_));
 sg13g2_o21ai_1 _33411_ (.B1(_04993_),
    .Y(_07689_),
    .A1(_04732_),
    .A2(_07688_));
 sg13g2_a21oi_1 _33412_ (.A1(_04711_),
    .A2(_07689_),
    .Y(_07690_),
    .B1(_04999_));
 sg13g2_a21o_1 _33413_ (.A2(_07689_),
    .A1(_04711_),
    .B1(_04999_),
    .X(_07691_));
 sg13g2_o21ai_1 _33414_ (.B1(_05002_),
    .Y(_07692_),
    .A1(_04695_),
    .A2(_07690_));
 sg13g2_xor2_1 _33415_ (.B(_07692_),
    .A(_04689_),
    .X(_07693_));
 sg13g2_and2_1 _33416_ (.A(_06305_),
    .B(_06356_),
    .X(_07694_));
 sg13g2_nor3_1 _33417_ (.A(_04779_),
    .B(_04783_),
    .C(_07694_),
    .Y(_07695_));
 sg13g2_a21oi_1 _33418_ (.A1(_06305_),
    .A2(_06356_),
    .Y(_07696_),
    .B1(_05928_));
 sg13g2_a21o_2 _33419_ (.A2(_06356_),
    .A1(_06305_),
    .B1(_05928_),
    .X(_07697_));
 sg13g2_o21ai_1 _33420_ (.B1(_05975_),
    .Y(_07698_),
    .A1(_05913_),
    .A2(_07697_));
 sg13g2_a21oi_2 _33421_ (.B1(_05938_),
    .Y(_07699_),
    .A2(_07698_),
    .A1(_05925_));
 sg13g2_nor2_1 _33422_ (.A(_05917_),
    .B(_07699_),
    .Y(_07700_));
 sg13g2_nor2_1 _33423_ (.A(_05939_),
    .B(_07700_),
    .Y(_07701_));
 sg13g2_nor3_1 _33424_ (.A(_05917_),
    .B(_05918_),
    .C(_07699_),
    .Y(_07702_));
 sg13g2_nor2_1 _33425_ (.A(_05942_),
    .B(_07702_),
    .Y(_07703_));
 sg13g2_o21ai_1 _33426_ (.B1(_05914_),
    .Y(_07704_),
    .A1(_05942_),
    .A2(_07702_));
 sg13g2_nand3_1 _33427_ (.B(_05944_),
    .C(_07704_),
    .A(_04689_),
    .Y(_07705_));
 sg13g2_a21oi_1 _33428_ (.A1(_05944_),
    .A2(_07704_),
    .Y(_07706_),
    .B1(_04689_));
 sg13g2_nor2_1 _33429_ (.A(net5677),
    .B(_07706_),
    .Y(_07707_));
 sg13g2_a21oi_1 _33430_ (.A1(_07705_),
    .A2(_07707_),
    .Y(_07708_),
    .B1(net4959));
 sg13g2_o21ai_1 _33431_ (.B1(_07708_),
    .Y(_07709_),
    .A1(net5761),
    .A2(_14191_));
 sg13g2_o21ai_1 _33432_ (.B1(_07709_),
    .Y(_07710_),
    .A1(net5050),
    .A2(_07693_));
 sg13g2_nand2b_1 _33433_ (.Y(_07711_),
    .B(net4750),
    .A_N(_07710_));
 sg13g2_xnor2_1 _33434_ (.Y(_07712_),
    .A(net4805),
    .B(_07710_));
 sg13g2_a21oi_1 _33435_ (.A1(\u_inv.d_next[190] ),
    .A2(\u_inv.d_reg[190] ),
    .Y(_07713_),
    .B1(_07706_));
 sg13g2_xor2_1 _33436_ (.B(_07713_),
    .A(_04687_),
    .X(_07714_));
 sg13g2_nand2_1 _33437_ (.Y(_07715_),
    .A(net5677),
    .B(\u_inv.d_next[191] ));
 sg13g2_a21oi_1 _33438_ (.A1(net5761),
    .A2(_07714_),
    .Y(_07716_),
    .B1(net4960));
 sg13g2_a21oi_1 _33439_ (.A1(_04689_),
    .A2(_07692_),
    .Y(_07717_),
    .B1(_05003_));
 sg13g2_or2_1 _33440_ (.X(_07718_),
    .B(_07717_),
    .A(_04687_));
 sg13g2_a21oi_1 _33441_ (.A1(_04687_),
    .A2(_07717_),
    .Y(_07719_),
    .B1(net5050));
 sg13g2_a22oi_1 _33442_ (.Y(_07720_),
    .B1(_07718_),
    .B2(_07719_),
    .A2(_07716_),
    .A1(_07715_));
 sg13g2_nand2_1 _33443_ (.Y(_07721_),
    .A(net4750),
    .B(_07720_));
 sg13g2_xnor2_1 _33444_ (.Y(_07722_),
    .A(net4750),
    .B(_07720_));
 sg13g2_xnor2_1 _33445_ (.Y(_07723_),
    .A(_04694_),
    .B(_07690_));
 sg13g2_xnor2_1 _33446_ (.Y(_07724_),
    .A(_04694_),
    .B(_07703_));
 sg13g2_a21oi_1 _33447_ (.A1(net5677),
    .A2(\u_inv.d_next[188] ),
    .Y(_07725_),
    .B1(net4960));
 sg13g2_o21ai_1 _33448_ (.B1(_07725_),
    .Y(_07726_),
    .A1(net5677),
    .A2(_07724_));
 sg13g2_o21ai_1 _33449_ (.B1(_07726_),
    .Y(_07727_),
    .A1(net5050),
    .A2(_07723_));
 sg13g2_nand2b_1 _33450_ (.Y(_07728_),
    .B(net4750),
    .A_N(_07727_));
 sg13g2_xnor2_1 _33451_ (.Y(_07729_),
    .A(net4750),
    .B(_07727_));
 sg13g2_o21ai_1 _33452_ (.B1(_04693_),
    .Y(_07730_),
    .A1(_04694_),
    .A2(_07703_));
 sg13g2_xnor2_1 _33453_ (.Y(_07731_),
    .A(_04691_),
    .B(_07730_));
 sg13g2_nand2_1 _33454_ (.Y(_07732_),
    .A(net5677),
    .B(\u_inv.d_next[189] ));
 sg13g2_a21oi_1 _33455_ (.A1(net5761),
    .A2(_07731_),
    .Y(_07733_),
    .B1(net4960));
 sg13g2_a21o_1 _33456_ (.A2(_07691_),
    .A1(_04694_),
    .B1(_05001_),
    .X(_07734_));
 sg13g2_nand2b_1 _33457_ (.Y(_07735_),
    .B(_04691_),
    .A_N(_07734_));
 sg13g2_a21oi_1 _33458_ (.A1(_04692_),
    .A2(_07734_),
    .Y(_07736_),
    .B1(net5050));
 sg13g2_a22oi_1 _33459_ (.Y(_07737_),
    .B1(_07735_),
    .B2(_07736_),
    .A2(_07733_),
    .A1(_07732_));
 sg13g2_nand2_1 _33460_ (.Y(_07738_),
    .A(net4750),
    .B(_07737_));
 sg13g2_xnor2_1 _33461_ (.Y(_07739_),
    .A(net4806),
    .B(_07737_));
 sg13g2_nand2_1 _33462_ (.Y(_07740_),
    .A(_07729_),
    .B(_07739_));
 sg13g2_inv_1 _33463_ (.Y(_07741_),
    .A(_07740_));
 sg13g2_nor3_1 _33464_ (.A(_07712_),
    .B(_07722_),
    .C(_07740_),
    .Y(_07742_));
 sg13g2_a21oi_1 _33465_ (.A1(_04710_),
    .A2(_07689_),
    .Y(_07743_),
    .B1(_04996_));
 sg13g2_xnor2_1 _33466_ (.Y(_07744_),
    .A(_04701_),
    .B(_07743_));
 sg13g2_o21ai_1 _33467_ (.B1(_04701_),
    .Y(_07745_),
    .A1(_05939_),
    .A2(_07700_));
 sg13g2_xnor2_1 _33468_ (.Y(_07746_),
    .A(_04701_),
    .B(_07701_));
 sg13g2_nand2_1 _33469_ (.Y(_07747_),
    .A(net5677),
    .B(\u_inv.d_next[186] ));
 sg13g2_a21oi_1 _33470_ (.A1(net5761),
    .A2(_07746_),
    .Y(_07748_),
    .B1(net4960));
 sg13g2_a22oi_1 _33471_ (.Y(_07749_),
    .B1(_07747_),
    .B2(_07748_),
    .A2(_07744_),
    .A1(net4960));
 sg13g2_nand2_1 _33472_ (.Y(_07750_),
    .A(net4751),
    .B(_07749_));
 sg13g2_inv_1 _33473_ (.Y(_07751_),
    .A(_07750_));
 sg13g2_xnor2_1 _33474_ (.Y(_07752_),
    .A(net4806),
    .B(_07749_));
 sg13g2_nand3_1 _33475_ (.B(_04700_),
    .C(_07745_),
    .A(_04699_),
    .Y(_07753_));
 sg13g2_a21o_1 _33476_ (.A2(_07745_),
    .A1(_04700_),
    .B1(_04699_),
    .X(_07754_));
 sg13g2_nand3_1 _33477_ (.B(_07753_),
    .C(_07754_),
    .A(net5761),
    .Y(_07755_));
 sg13g2_a21oi_1 _33478_ (.A1(net5679),
    .A2(\u_inv.d_next[187] ),
    .Y(_07756_),
    .B1(net4960));
 sg13g2_o21ai_1 _33479_ (.B1(_04997_),
    .Y(_07757_),
    .A1(_04701_),
    .A2(_07743_));
 sg13g2_nand2b_1 _33480_ (.Y(_07758_),
    .B(_04699_),
    .A_N(_07757_));
 sg13g2_a21oi_1 _33481_ (.A1(_04698_),
    .A2(_07757_),
    .Y(_07759_),
    .B1(net5050));
 sg13g2_a22oi_1 _33482_ (.Y(_07760_),
    .B1(_07758_),
    .B2(_07759_),
    .A2(_07756_),
    .A1(_07755_));
 sg13g2_xnor2_1 _33483_ (.Y(_07761_),
    .A(net4806),
    .B(_07760_));
 sg13g2_o21ai_1 _33484_ (.B1(_04707_),
    .Y(_07762_),
    .A1(_04709_),
    .A2(_07699_));
 sg13g2_a21oi_1 _33485_ (.A1(_04705_),
    .A2(_07762_),
    .Y(_07763_),
    .B1(net5677));
 sg13g2_o21ai_1 _33486_ (.B1(_07763_),
    .Y(_07764_),
    .A1(_04705_),
    .A2(_07762_));
 sg13g2_a21oi_1 _33487_ (.A1(net5677),
    .A2(\u_inv.d_next[185] ),
    .Y(_07765_),
    .B1(net4960));
 sg13g2_a21oi_1 _33488_ (.A1(_04709_),
    .A2(_07689_),
    .Y(_07766_),
    .B1(_04995_));
 sg13g2_nand2b_1 _33489_ (.Y(_07767_),
    .B(_04705_),
    .A_N(_07766_));
 sg13g2_a21oi_1 _33490_ (.A1(_04706_),
    .A2(_07766_),
    .Y(_07768_),
    .B1(net5050));
 sg13g2_a22oi_1 _33491_ (.Y(_07769_),
    .B1(_07767_),
    .B2(_07768_),
    .A2(_07765_),
    .A1(_07764_));
 sg13g2_nand2_1 _33492_ (.Y(_07770_),
    .A(net4751),
    .B(_07769_));
 sg13g2_xnor2_1 _33493_ (.Y(_07771_),
    .A(net4806),
    .B(_07769_));
 sg13g2_inv_1 _33494_ (.Y(_07772_),
    .A(_07771_));
 sg13g2_xnor2_1 _33495_ (.Y(_07773_),
    .A(_04709_),
    .B(_07689_));
 sg13g2_xnor2_1 _33496_ (.Y(_07774_),
    .A(_04709_),
    .B(_07699_));
 sg13g2_o21ai_1 _33497_ (.B1(net5051),
    .Y(_07775_),
    .A1(net5761),
    .A2(\u_inv.d_next[184] ));
 sg13g2_a21o_1 _33498_ (.A2(_07774_),
    .A1(net5761),
    .B1(_07775_),
    .X(_07776_));
 sg13g2_o21ai_1 _33499_ (.B1(_07776_),
    .Y(_07777_),
    .A1(net5051),
    .A2(_07773_));
 sg13g2_nand2_1 _33500_ (.Y(_07778_),
    .A(net4750),
    .B(_07777_));
 sg13g2_xnor2_1 _33501_ (.Y(_07779_),
    .A(net4806),
    .B(_07777_));
 sg13g2_xnor2_1 _33502_ (.Y(_07780_),
    .A(net4750),
    .B(_07777_));
 sg13g2_nand4_1 _33503_ (.B(_07761_),
    .C(_07771_),
    .A(_07752_),
    .Y(_07781_),
    .D(_07779_));
 sg13g2_nor4_1 _33504_ (.A(_07712_),
    .B(_07722_),
    .C(_07740_),
    .D(_07781_),
    .Y(_07782_));
 sg13g2_a21oi_1 _33505_ (.A1(_05924_),
    .A2(_07698_),
    .Y(_07783_),
    .B1(_05931_));
 sg13g2_nand3_1 _33506_ (.B(_05924_),
    .C(_07698_),
    .A(_05923_),
    .Y(_07784_));
 sg13g2_nand2_1 _33507_ (.Y(_07785_),
    .A(_05933_),
    .B(_07784_));
 sg13g2_and2_1 _33508_ (.A(_05921_),
    .B(_07785_),
    .X(_07786_));
 sg13g2_o21ai_1 _33509_ (.B1(_04721_),
    .Y(_07787_),
    .A1(_05936_),
    .A2(_07786_));
 sg13g2_nand3_1 _33510_ (.B(_04720_),
    .C(_07787_),
    .A(_04719_),
    .Y(_07788_));
 sg13g2_a21o_1 _33511_ (.A2(_07787_),
    .A1(_04720_),
    .B1(_04719_),
    .X(_07789_));
 sg13g2_nand3_1 _33512_ (.B(_07788_),
    .C(_07789_),
    .A(net5772),
    .Y(_07790_));
 sg13g2_nand2_1 _33513_ (.Y(_07791_),
    .A(net5685),
    .B(\u_inv.d_next[183] ));
 sg13g2_nand3_1 _33514_ (.B(_07790_),
    .C(_07791_),
    .A(net5060),
    .Y(_07792_));
 sg13g2_o21ai_1 _33515_ (.B1(_04980_),
    .Y(_07793_),
    .A1(_04731_),
    .A2(_07688_));
 sg13g2_nand3b_1 _33516_ (.B(_04730_),
    .C(_04726_),
    .Y(_07794_),
    .A_N(_07688_));
 sg13g2_nand2_1 _33517_ (.Y(_07795_),
    .A(_04983_),
    .B(_07794_));
 sg13g2_a21o_1 _33518_ (.A2(_07794_),
    .A1(_04983_),
    .B1(_04717_),
    .X(_07796_));
 sg13g2_a21o_1 _33519_ (.A2(_07796_),
    .A1(_04988_),
    .B1(_04721_),
    .X(_07797_));
 sg13g2_nand3_1 _33520_ (.B(_04990_),
    .C(_07797_),
    .A(_04719_),
    .Y(_07798_));
 sg13g2_a21o_1 _33521_ (.A2(_07797_),
    .A1(_04990_),
    .B1(_04719_),
    .X(_07799_));
 sg13g2_nand3_1 _33522_ (.B(_07798_),
    .C(_07799_),
    .A(net4969),
    .Y(_07800_));
 sg13g2_nand2_1 _33523_ (.Y(_07801_),
    .A(_07792_),
    .B(_07800_));
 sg13g2_and3_2 _33524_ (.X(_07802_),
    .A(net4755),
    .B(_07792_),
    .C(_07800_));
 sg13g2_a21oi_1 _33525_ (.A1(_07792_),
    .A2(_07800_),
    .Y(_07803_),
    .B1(net4755));
 sg13g2_nor2_1 _33526_ (.A(_07802_),
    .B(_07803_),
    .Y(_07804_));
 sg13g2_nand3_1 _33527_ (.B(_04988_),
    .C(_07796_),
    .A(_04721_),
    .Y(_07805_));
 sg13g2_a21oi_1 _33528_ (.A1(_07797_),
    .A2(_07805_),
    .Y(_07806_),
    .B1(net5060));
 sg13g2_or3_1 _33529_ (.A(_04721_),
    .B(_05936_),
    .C(_07786_),
    .X(_07807_));
 sg13g2_nand3_1 _33530_ (.B(_07787_),
    .C(_07807_),
    .A(net5772),
    .Y(_07808_));
 sg13g2_a21oi_1 _33531_ (.A1(net5685),
    .A2(\u_inv.d_next[182] ),
    .Y(_07809_),
    .B1(net4969));
 sg13g2_a21o_2 _33532_ (.A2(_07809_),
    .A1(_07808_),
    .B1(_07806_),
    .X(_07810_));
 sg13g2_nand2b_1 _33533_ (.Y(_07811_),
    .B(net4755),
    .A_N(_07810_));
 sg13g2_xnor2_1 _33534_ (.Y(_07812_),
    .A(net4755),
    .B(_07810_));
 sg13g2_xnor2_1 _33535_ (.Y(_07813_),
    .A(net4810),
    .B(_07810_));
 sg13g2_nor3_1 _33536_ (.A(_07802_),
    .B(_07803_),
    .C(_07813_),
    .Y(_07814_));
 sg13g2_a21oi_1 _33537_ (.A1(_04715_),
    .A2(_07785_),
    .Y(_07815_),
    .B1(_04714_));
 sg13g2_xnor2_1 _33538_ (.Y(_07816_),
    .A(_04713_),
    .B(_07815_));
 sg13g2_a21oi_1 _33539_ (.A1(net5685),
    .A2(\u_inv.d_next[181] ),
    .Y(_07817_),
    .B1(net4969));
 sg13g2_o21ai_1 _33540_ (.B1(_07817_),
    .Y(_07818_),
    .A1(net5685),
    .A2(_07816_));
 sg13g2_a21o_1 _33541_ (.A2(_07794_),
    .A1(_04983_),
    .B1(_04715_),
    .X(_07819_));
 sg13g2_nand3_1 _33542_ (.B(_04987_),
    .C(_07819_),
    .A(_04713_),
    .Y(_07820_));
 sg13g2_a21o_1 _33543_ (.A2(_07819_),
    .A1(_04987_),
    .B1(_04713_),
    .X(_07821_));
 sg13g2_nand3_1 _33544_ (.B(_07820_),
    .C(_07821_),
    .A(net4969),
    .Y(_07822_));
 sg13g2_nand2_1 _33545_ (.Y(_07823_),
    .A(_07818_),
    .B(_07822_));
 sg13g2_nand3_1 _33546_ (.B(_07818_),
    .C(_07822_),
    .A(net4755),
    .Y(_07824_));
 sg13g2_a21o_1 _33547_ (.A2(_07822_),
    .A1(_07818_),
    .B1(net4755),
    .X(_07825_));
 sg13g2_nand2_1 _33548_ (.Y(_07826_),
    .A(net4755),
    .B(_07823_));
 sg13g2_nand3_1 _33549_ (.B(_07818_),
    .C(_07822_),
    .A(net4810),
    .Y(_07827_));
 sg13g2_nand2_1 _33550_ (.Y(_07828_),
    .A(_07826_),
    .B(_07827_));
 sg13g2_xnor2_1 _33551_ (.Y(_07829_),
    .A(_04715_),
    .B(_07795_));
 sg13g2_xnor2_1 _33552_ (.Y(_07830_),
    .A(_04715_),
    .B(_07785_));
 sg13g2_o21ai_1 _33553_ (.B1(net5061),
    .Y(_07831_),
    .A1(net5772),
    .A2(\u_inv.d_next[180] ));
 sg13g2_a21oi_1 _33554_ (.A1(net5772),
    .A2(_07830_),
    .Y(_07832_),
    .B1(_07831_));
 sg13g2_a21oi_2 _33555_ (.B1(_07832_),
    .Y(_07833_),
    .A2(_07829_),
    .A1(net4969));
 sg13g2_nor2_1 _33556_ (.A(net4810),
    .B(_07833_),
    .Y(_07834_));
 sg13g2_xnor2_1 _33557_ (.Y(_07835_),
    .A(net4755),
    .B(_07833_));
 sg13g2_xnor2_1 _33558_ (.Y(_07836_),
    .A(net4810),
    .B(_07833_));
 sg13g2_nand3_1 _33559_ (.B(_07825_),
    .C(_07835_),
    .A(_07824_),
    .Y(_07837_));
 sg13g2_nor4_1 _33560_ (.A(_07802_),
    .B(_07803_),
    .C(_07813_),
    .D(_07837_),
    .Y(_07838_));
 sg13g2_o21ai_1 _33561_ (.B1(_04724_),
    .Y(_07839_),
    .A1(_04725_),
    .A2(_07783_));
 sg13g2_xnor2_1 _33562_ (.Y(_07840_),
    .A(_04723_),
    .B(_07839_));
 sg13g2_nand2_1 _33563_ (.Y(_07841_),
    .A(net5685),
    .B(\u_inv.d_next[179] ));
 sg13g2_a21oi_1 _33564_ (.A1(net5772),
    .A2(_07840_),
    .Y(_07842_),
    .B1(net4969));
 sg13g2_a21oi_1 _33565_ (.A1(_04725_),
    .A2(_07793_),
    .Y(_07843_),
    .B1(_04982_));
 sg13g2_or2_1 _33566_ (.X(_07844_),
    .B(_07843_),
    .A(_04723_));
 sg13g2_a21oi_1 _33567_ (.A1(_04723_),
    .A2(_07843_),
    .Y(_07845_),
    .B1(net5061));
 sg13g2_a22oi_1 _33568_ (.Y(_07846_),
    .B1(_07844_),
    .B2(_07845_),
    .A2(_07842_),
    .A1(_07841_));
 sg13g2_xnor2_1 _33569_ (.Y(_07847_),
    .A(net4810),
    .B(_07846_));
 sg13g2_xnor2_1 _33570_ (.Y(_07848_),
    .A(_04725_),
    .B(_07793_));
 sg13g2_xor2_1 _33571_ (.B(_07783_),
    .A(_04725_),
    .X(_07849_));
 sg13g2_nand2_1 _33572_ (.Y(_07850_),
    .A(net5685),
    .B(\u_inv.d_next[178] ));
 sg13g2_a21oi_1 _33573_ (.A1(net5772),
    .A2(_07849_),
    .Y(_07851_),
    .B1(net4973));
 sg13g2_a22oi_1 _33574_ (.Y(_07852_),
    .B1(_07850_),
    .B2(_07851_),
    .A2(_07848_),
    .A1(net4969));
 sg13g2_and2_1 _33575_ (.A(net4756),
    .B(_07852_),
    .X(_07853_));
 sg13g2_xnor2_1 _33576_ (.Y(_07854_),
    .A(net4810),
    .B(_07852_));
 sg13g2_nand2_1 _33577_ (.Y(_07855_),
    .A(_07847_),
    .B(_07854_));
 sg13g2_a21oi_1 _33578_ (.A1(_04729_),
    .A2(_07698_),
    .Y(_07856_),
    .B1(_04728_));
 sg13g2_xnor2_1 _33579_ (.Y(_07857_),
    .A(_04727_),
    .B(_07856_));
 sg13g2_o21ai_1 _33580_ (.B1(net5061),
    .Y(_07858_),
    .A1(net5772),
    .A2(_14196_));
 sg13g2_a21oi_1 _33581_ (.A1(net5772),
    .A2(_07857_),
    .Y(_07859_),
    .B1(_07858_));
 sg13g2_o21ai_1 _33582_ (.B1(_04978_),
    .Y(_07860_),
    .A1(_04729_),
    .A2(_07688_));
 sg13g2_o21ai_1 _33583_ (.B1(net4969),
    .Y(_07861_),
    .A1(_04727_),
    .A2(_07860_));
 sg13g2_a21oi_1 _33584_ (.A1(_04727_),
    .A2(_07860_),
    .Y(_07862_),
    .B1(_07861_));
 sg13g2_nor2_2 _33585_ (.A(_07859_),
    .B(_07862_),
    .Y(_07863_));
 sg13g2_inv_1 _33586_ (.Y(_07864_),
    .A(_07863_));
 sg13g2_xnor2_1 _33587_ (.Y(_07865_),
    .A(net4810),
    .B(_07863_));
 sg13g2_xnor2_1 _33588_ (.Y(_07866_),
    .A(_04729_),
    .B(_07688_));
 sg13g2_xor2_1 _33589_ (.B(_07698_),
    .A(_04729_),
    .X(_07867_));
 sg13g2_mux2_1 _33590_ (.A0(\u_inv.d_next[176] ),
    .A1(_07867_),
    .S(net5773),
    .X(_07868_));
 sg13g2_nand2_1 _33591_ (.Y(_07869_),
    .A(net5060),
    .B(_07868_));
 sg13g2_o21ai_1 _33592_ (.B1(_07869_),
    .Y(_07870_),
    .A1(net5061),
    .A2(_07866_));
 sg13g2_nand2_1 _33593_ (.Y(_07871_),
    .A(net4756),
    .B(_07870_));
 sg13g2_xnor2_1 _33594_ (.Y(_07872_),
    .A(net4756),
    .B(_07870_));
 sg13g2_inv_2 _33595_ (.Y(_07873_),
    .A(_07872_));
 sg13g2_and4_1 _33596_ (.A(_07847_),
    .B(_07854_),
    .C(_07865_),
    .D(_07873_),
    .X(_07874_));
 sg13g2_and2_1 _33597_ (.A(_07838_),
    .B(_07874_),
    .X(_07875_));
 sg13g2_and2_1 _33598_ (.A(_07782_),
    .B(_07875_),
    .X(_07876_));
 sg13g2_a21oi_2 _33599_ (.B1(_04961_),
    .Y(_07877_),
    .A2(_07685_),
    .A1(_04786_));
 sg13g2_o21ai_1 _33600_ (.B1(_04972_),
    .Y(_07878_),
    .A1(_04756_),
    .A2(_07877_));
 sg13g2_a21o_1 _33601_ (.A2(_07878_),
    .A1(_04745_),
    .B1(_04964_),
    .X(_07879_));
 sg13g2_xor2_1 _33602_ (.B(_07879_),
    .A(_04738_),
    .X(_07880_));
 sg13g2_nand2b_2 _33603_ (.Y(_07881_),
    .B(_07697_),
    .A_N(_05952_));
 sg13g2_a21oi_2 _33604_ (.B1(_05960_),
    .Y(_07882_),
    .A2(_07696_),
    .A1(_05912_));
 sg13g2_nor2b_1 _33605_ (.A(_07882_),
    .B_N(_04754_),
    .Y(_07883_));
 sg13g2_nand2_1 _33606_ (.Y(_07884_),
    .A(_04753_),
    .B(_07883_));
 sg13g2_nor3_1 _33607_ (.A(_05908_),
    .B(_05909_),
    .C(_07882_),
    .Y(_07885_));
 sg13g2_nand2b_1 _33608_ (.Y(_07886_),
    .B(_05967_),
    .A_N(_07885_));
 sg13g2_o21ai_1 _33609_ (.B1(_05906_),
    .Y(_07887_),
    .A1(_05968_),
    .A2(_07885_));
 sg13g2_nand3_1 _33610_ (.B(_05972_),
    .C(_07887_),
    .A(_04738_),
    .Y(_07888_));
 sg13g2_a21o_1 _33611_ (.A2(_07887_),
    .A1(_05972_),
    .B1(_04738_),
    .X(_07889_));
 sg13g2_nand3_1 _33612_ (.B(_07888_),
    .C(_07889_),
    .A(net5773),
    .Y(_07890_));
 sg13g2_a21oi_1 _33613_ (.A1(net5684),
    .A2(\u_inv.d_next[174] ),
    .Y(_07891_),
    .B1(net4967));
 sg13g2_nand2_1 _33614_ (.Y(_07892_),
    .A(_07890_),
    .B(_07891_));
 sg13g2_o21ai_1 _33615_ (.B1(_07892_),
    .Y(_07893_),
    .A1(net5060),
    .A2(_07880_));
 sg13g2_nand2b_1 _33616_ (.Y(_07894_),
    .B(net4757),
    .A_N(_07893_));
 sg13g2_xnor2_1 _33617_ (.Y(_07895_),
    .A(net4808),
    .B(_07893_));
 sg13g2_nand2_1 _33618_ (.Y(_07896_),
    .A(_04737_),
    .B(_07889_));
 sg13g2_xnor2_1 _33619_ (.Y(_07897_),
    .A(_04736_),
    .B(_07896_));
 sg13g2_a21o_1 _33620_ (.A2(\u_inv.d_next[175] ),
    .A1(net5684),
    .B1(net4968),
    .X(_07898_));
 sg13g2_a21oi_1 _33621_ (.A1(net5773),
    .A2(_07897_),
    .Y(_07899_),
    .B1(_07898_));
 sg13g2_a21oi_1 _33622_ (.A1(_04738_),
    .A2(_07879_),
    .Y(_07900_),
    .B1(_04965_));
 sg13g2_or2_1 _33623_ (.X(_07901_),
    .B(_07900_),
    .A(_04736_));
 sg13g2_a21oi_1 _33624_ (.A1(_04736_),
    .A2(_07900_),
    .Y(_07902_),
    .B1(net5060));
 sg13g2_a21o_2 _33625_ (.A2(_07902_),
    .A1(_07901_),
    .B1(_07899_),
    .X(_07903_));
 sg13g2_xnor2_1 _33626_ (.Y(_07904_),
    .A(net4808),
    .B(_07903_));
 sg13g2_nor2_1 _33627_ (.A(_07895_),
    .B(_07904_),
    .Y(_07905_));
 sg13g2_xnor2_1 _33628_ (.Y(_07906_),
    .A(_04744_),
    .B(_07878_));
 sg13g2_xnor2_1 _33629_ (.Y(_07907_),
    .A(_04744_),
    .B(_07886_));
 sg13g2_a21oi_1 _33630_ (.A1(net5684),
    .A2(\u_inv.d_next[172] ),
    .Y(_07908_),
    .B1(net4968));
 sg13g2_o21ai_1 _33631_ (.B1(_07908_),
    .Y(_07909_),
    .A1(net5684),
    .A2(_07907_));
 sg13g2_o21ai_1 _33632_ (.B1(_07909_),
    .Y(_07910_),
    .A1(net5060),
    .A2(_07906_));
 sg13g2_nor2_1 _33633_ (.A(net4809),
    .B(_07910_),
    .Y(_07911_));
 sg13g2_xnor2_1 _33634_ (.Y(_07912_),
    .A(net4757),
    .B(_07910_));
 sg13g2_inv_1 _33635_ (.Y(_07913_),
    .A(_07912_));
 sg13g2_a21oi_1 _33636_ (.A1(_04744_),
    .A2(_07886_),
    .Y(_07914_),
    .B1(_04742_));
 sg13g2_xnor2_1 _33637_ (.Y(_07915_),
    .A(_04740_),
    .B(_07914_));
 sg13g2_nand2_1 _33638_ (.Y(_07916_),
    .A(net5684),
    .B(\u_inv.d_next[173] ));
 sg13g2_a21oi_1 _33639_ (.A1(net5773),
    .A2(_07915_),
    .Y(_07917_),
    .B1(net4967));
 sg13g2_a21oi_1 _33640_ (.A1(_04743_),
    .A2(_07878_),
    .Y(_07918_),
    .B1(_04962_));
 sg13g2_o21ai_1 _33641_ (.B1(net4968),
    .Y(_07919_),
    .A1(_04741_),
    .A2(_07918_));
 sg13g2_a21oi_1 _33642_ (.A1(_04741_),
    .A2(_07918_),
    .Y(_07920_),
    .B1(_07919_));
 sg13g2_a21oi_2 _33643_ (.B1(_07920_),
    .Y(_07921_),
    .A2(_07917_),
    .A1(_07916_));
 sg13g2_xnor2_1 _33644_ (.Y(_07922_),
    .A(net4809),
    .B(_07921_));
 sg13g2_o21ai_1 _33645_ (.B1(_04968_),
    .Y(_07923_),
    .A1(_04755_),
    .A2(_07877_));
 sg13g2_xnor2_1 _33646_ (.Y(_07924_),
    .A(_04751_),
    .B(_07923_));
 sg13g2_nand3_1 _33647_ (.B(_05964_),
    .C(_07884_),
    .A(_04751_),
    .Y(_07925_));
 sg13g2_a21o_1 _33648_ (.A2(_07884_),
    .A1(_05964_),
    .B1(_04751_),
    .X(_07926_));
 sg13g2_nand3_1 _33649_ (.B(_07925_),
    .C(_07926_),
    .A(net5773),
    .Y(_07927_));
 sg13g2_a21oi_1 _33650_ (.A1(net5684),
    .A2(\u_inv.d_next[170] ),
    .Y(_07928_),
    .B1(net4967));
 sg13g2_a22oi_1 _33651_ (.Y(_07929_),
    .B1(_07927_),
    .B2(_07928_),
    .A2(_07924_),
    .A1(net4967));
 sg13g2_xnor2_1 _33652_ (.Y(_07930_),
    .A(net4808),
    .B(_07929_));
 sg13g2_inv_1 _33653_ (.Y(_07931_),
    .A(_07930_));
 sg13g2_nand3_1 _33654_ (.B(_04750_),
    .C(_07926_),
    .A(_04749_),
    .Y(_07932_));
 sg13g2_a21o_1 _33655_ (.A2(_07926_),
    .A1(_04750_),
    .B1(_04749_),
    .X(_07933_));
 sg13g2_nand3_1 _33656_ (.B(_07932_),
    .C(_07933_),
    .A(net5773),
    .Y(_07934_));
 sg13g2_a21oi_1 _33657_ (.A1(net5684),
    .A2(\u_inv.d_next[171] ),
    .Y(_07935_),
    .B1(net4967));
 sg13g2_a21oi_1 _33658_ (.A1(_04751_),
    .A2(_07923_),
    .Y(_07936_),
    .B1(_04969_));
 sg13g2_o21ai_1 _33659_ (.B1(net4967),
    .Y(_07937_),
    .A1(_04749_),
    .A2(_07936_));
 sg13g2_a21oi_1 _33660_ (.A1(_04749_),
    .A2(_07936_),
    .Y(_07938_),
    .B1(_07937_));
 sg13g2_a21oi_2 _33661_ (.B1(_07938_),
    .Y(_07939_),
    .A2(_07935_),
    .A1(_07934_));
 sg13g2_xnor2_1 _33662_ (.Y(_07940_),
    .A(net4808),
    .B(_07939_));
 sg13g2_nand2_1 _33663_ (.Y(_07941_),
    .A(_07930_),
    .B(_07940_));
 sg13g2_a21o_1 _33664_ (.A2(\u_inv.d_reg[168] ),
    .A1(\u_inv.d_next[168] ),
    .B1(_07883_),
    .X(_07942_));
 sg13g2_xor2_1 _33665_ (.B(_07942_),
    .A(_04753_),
    .X(_07943_));
 sg13g2_nand2_1 _33666_ (.Y(_07944_),
    .A(net5684),
    .B(\u_inv.d_next[169] ));
 sg13g2_a21oi_1 _33667_ (.A1(net5773),
    .A2(_07943_),
    .Y(_07945_),
    .B1(net4967));
 sg13g2_o21ai_1 _33668_ (.B1(_04966_),
    .Y(_07946_),
    .A1(_04754_),
    .A2(_07877_));
 sg13g2_o21ai_1 _33669_ (.B1(net4967),
    .Y(_07947_),
    .A1(_04753_),
    .A2(_07946_));
 sg13g2_a21oi_1 _33670_ (.A1(_04753_),
    .A2(_07946_),
    .Y(_07948_),
    .B1(_07947_));
 sg13g2_a21oi_2 _33671_ (.B1(_07948_),
    .Y(_07949_),
    .A2(_07945_),
    .A1(_07944_));
 sg13g2_inv_1 _33672_ (.Y(_07950_),
    .A(_07949_));
 sg13g2_xnor2_1 _33673_ (.Y(_07951_),
    .A(net4808),
    .B(_07949_));
 sg13g2_xnor2_1 _33674_ (.Y(_07952_),
    .A(_04754_),
    .B(_07877_));
 sg13g2_xor2_1 _33675_ (.B(_07882_),
    .A(_04754_),
    .X(_07953_));
 sg13g2_o21ai_1 _33676_ (.B1(net5060),
    .Y(_07954_),
    .A1(net5774),
    .A2(\u_inv.d_next[168] ));
 sg13g2_a21o_1 _33677_ (.A2(_07953_),
    .A1(net5774),
    .B1(_07954_),
    .X(_07955_));
 sg13g2_o21ai_1 _33678_ (.B1(_07955_),
    .Y(_07956_),
    .A1(net5060),
    .A2(_07952_));
 sg13g2_nand2_1 _33679_ (.Y(_07957_),
    .A(net4757),
    .B(_07956_));
 sg13g2_xnor2_1 _33680_ (.Y(_07958_),
    .A(net4808),
    .B(_07956_));
 sg13g2_and4_1 _33681_ (.A(_07930_),
    .B(_07940_),
    .C(_07951_),
    .D(_07958_),
    .X(_07959_));
 sg13g2_and4_1 _33682_ (.A(_07905_),
    .B(_07912_),
    .C(_07922_),
    .D(_07959_),
    .X(_07960_));
 sg13g2_nand2_1 _33683_ (.Y(_07961_),
    .A(_04952_),
    .B(_07687_));
 sg13g2_a21oi_1 _33684_ (.A1(_04952_),
    .A2(_07687_),
    .Y(_07962_),
    .B1(_04763_));
 sg13g2_nand2b_1 _33685_ (.Y(_07963_),
    .B(_04956_),
    .A_N(_07962_));
 sg13g2_a21oi_1 _33686_ (.A1(_04768_),
    .A2(_07963_),
    .Y(_07964_),
    .B1(_04959_));
 sg13g2_a21oi_1 _33687_ (.A1(_04765_),
    .A2(_07964_),
    .Y(_07965_),
    .B1(net5062));
 sg13g2_o21ai_1 _33688_ (.B1(_07965_),
    .Y(_07966_),
    .A1(_04765_),
    .A2(_07964_));
 sg13g2_nand3_1 _33689_ (.B(_04761_),
    .C(_07881_),
    .A(_04758_),
    .Y(_07967_));
 sg13g2_a21o_1 _33690_ (.A2(_07967_),
    .A1(_05956_),
    .B1(_04768_),
    .X(_07968_));
 sg13g2_nand2_1 _33691_ (.Y(_07969_),
    .A(_04766_),
    .B(_07968_));
 sg13g2_xnor2_1 _33692_ (.Y(_07970_),
    .A(_04764_),
    .B(_07969_));
 sg13g2_a21oi_1 _33693_ (.A1(net5686),
    .A2(\u_inv.d_next[167] ),
    .Y(_07971_),
    .B1(net4970));
 sg13g2_o21ai_1 _33694_ (.B1(_07971_),
    .Y(_07972_),
    .A1(net5686),
    .A2(_07970_));
 sg13g2_nand2_1 _33695_ (.Y(_07973_),
    .A(_07966_),
    .B(_07972_));
 sg13g2_xnor2_1 _33696_ (.Y(_07974_),
    .A(net4759),
    .B(_07973_));
 sg13g2_xnor2_1 _33697_ (.Y(_07975_),
    .A(_04767_),
    .B(_07963_));
 sg13g2_nand3_1 _33698_ (.B(_05956_),
    .C(_07967_),
    .A(_04768_),
    .Y(_07976_));
 sg13g2_nand3_1 _33699_ (.B(_07968_),
    .C(_07976_),
    .A(net5774),
    .Y(_07977_));
 sg13g2_a21oi_1 _33700_ (.A1(net5686),
    .A2(\u_inv.d_next[166] ),
    .Y(_07978_),
    .B1(net4970));
 sg13g2_nand2_1 _33701_ (.Y(_07979_),
    .A(_07977_),
    .B(_07978_));
 sg13g2_o21ai_1 _33702_ (.B1(_07979_),
    .Y(_07980_),
    .A1(net5062),
    .A2(_07975_));
 sg13g2_xnor2_1 _33703_ (.Y(_07981_),
    .A(net4758),
    .B(_07980_));
 sg13g2_nand2_2 _33704_ (.Y(_07982_),
    .A(_07974_),
    .B(_07981_));
 sg13g2_xnor2_1 _33705_ (.Y(_07983_),
    .A(_04761_),
    .B(_07881_));
 sg13g2_o21ai_1 _33706_ (.B1(net5062),
    .Y(_07984_),
    .A1(net5774),
    .A2(\u_inv.d_next[164] ));
 sg13g2_a21o_1 _33707_ (.A2(_07983_),
    .A1(net5774),
    .B1(_07984_),
    .X(_07985_));
 sg13g2_a21oi_1 _33708_ (.A1(_04952_),
    .A2(_07687_),
    .Y(_07986_),
    .B1(_04761_));
 sg13g2_o21ai_1 _33709_ (.B1(net4970),
    .Y(_07987_),
    .A1(_04762_),
    .A2(_07961_));
 sg13g2_o21ai_1 _33710_ (.B1(_07985_),
    .Y(_07988_),
    .A1(_07986_),
    .A2(_07987_));
 sg13g2_and2_1 _33711_ (.A(net4758),
    .B(_07988_),
    .X(_07989_));
 sg13g2_xnor2_1 _33712_ (.Y(_07990_),
    .A(net4811),
    .B(_07988_));
 sg13g2_o21ai_1 _33713_ (.B1(_04758_),
    .Y(_07991_),
    .A1(_04955_),
    .A2(_07986_));
 sg13g2_or3_1 _33714_ (.A(_04758_),
    .B(_04955_),
    .C(_07986_),
    .X(_07992_));
 sg13g2_nand3_1 _33715_ (.B(_07991_),
    .C(_07992_),
    .A(net4970),
    .Y(_07993_));
 sg13g2_a21oi_1 _33716_ (.A1(_04761_),
    .A2(_07881_),
    .Y(_07994_),
    .B1(_04760_));
 sg13g2_xnor2_1 _33717_ (.Y(_07995_),
    .A(_04759_),
    .B(_07994_));
 sg13g2_o21ai_1 _33718_ (.B1(net5062),
    .Y(_07996_),
    .A1(net5686),
    .A2(_07995_));
 sg13g2_a21o_1 _33719_ (.A2(\u_inv.d_next[165] ),
    .A1(net5686),
    .B1(_07996_),
    .X(_07997_));
 sg13g2_nand2_1 _33720_ (.Y(_07998_),
    .A(_07993_),
    .B(_07997_));
 sg13g2_nand3_1 _33721_ (.B(_07993_),
    .C(_07997_),
    .A(net4758),
    .Y(_07999_));
 sg13g2_xnor2_1 _33722_ (.Y(_08000_),
    .A(net4758),
    .B(_07998_));
 sg13g2_nand2_2 _33723_ (.Y(_08001_),
    .A(_07990_),
    .B(_08000_));
 sg13g2_a21o_1 _33724_ (.A2(_07686_),
    .A1(_04946_),
    .B1(_04774_),
    .X(_08002_));
 sg13g2_a21oi_1 _33725_ (.A1(_04948_),
    .A2(_08002_),
    .Y(_08003_),
    .B1(_04772_));
 sg13g2_nand3_1 _33726_ (.B(_04948_),
    .C(_08002_),
    .A(_04772_),
    .Y(_08004_));
 sg13g2_nand2_1 _33727_ (.Y(_08005_),
    .A(net4970),
    .B(_08004_));
 sg13g2_o21ai_1 _33728_ (.B1(_04774_),
    .Y(_08006_),
    .A1(_05950_),
    .A2(_07695_));
 sg13g2_inv_1 _33729_ (.Y(_08007_),
    .A(_08006_));
 sg13g2_nand3_1 _33730_ (.B(_04773_),
    .C(_08006_),
    .A(_04772_),
    .Y(_08008_));
 sg13g2_a21o_1 _33731_ (.A2(_08006_),
    .A1(_04773_),
    .B1(_04772_),
    .X(_08009_));
 sg13g2_nand3_1 _33732_ (.B(_08008_),
    .C(_08009_),
    .A(net5774),
    .Y(_08010_));
 sg13g2_nand2_1 _33733_ (.Y(_08011_),
    .A(net5686),
    .B(\u_inv.d_next[163] ));
 sg13g2_nand3_1 _33734_ (.B(_08010_),
    .C(_08011_),
    .A(net5062),
    .Y(_08012_));
 sg13g2_o21ai_1 _33735_ (.B1(_08012_),
    .Y(_08013_),
    .A1(_08003_),
    .A2(_08005_));
 sg13g2_xnor2_1 _33736_ (.Y(_08014_),
    .A(net4758),
    .B(_08013_));
 sg13g2_nand3_1 _33737_ (.B(_04946_),
    .C(_07686_),
    .A(_04774_),
    .Y(_08015_));
 sg13g2_a21oi_1 _33738_ (.A1(_08002_),
    .A2(_08015_),
    .Y(_08016_),
    .B1(net5062));
 sg13g2_nor3_1 _33739_ (.A(_04774_),
    .B(_05950_),
    .C(_07695_),
    .Y(_08017_));
 sg13g2_nor2_1 _33740_ (.A(_08007_),
    .B(_08017_),
    .Y(_08018_));
 sg13g2_a21o_1 _33741_ (.A2(\u_inv.d_next[162] ),
    .A1(net5686),
    .B1(net4970),
    .X(_08019_));
 sg13g2_a21oi_1 _33742_ (.A1(net5774),
    .A2(_08018_),
    .Y(_08020_),
    .B1(_08019_));
 sg13g2_or2_1 _33743_ (.X(_08021_),
    .B(_08020_),
    .A(_08016_));
 sg13g2_nor2_1 _33744_ (.A(net4811),
    .B(_08021_),
    .Y(_08022_));
 sg13g2_xnor2_1 _33745_ (.Y(_08023_),
    .A(net4758),
    .B(_08021_));
 sg13g2_o21ai_1 _33746_ (.B1(_04779_),
    .Y(_08024_),
    .A1(_04783_),
    .A2(_07694_));
 sg13g2_nor2b_1 _33747_ (.A(_08024_),
    .B_N(_04781_),
    .Y(_08025_));
 sg13g2_o21ai_1 _33748_ (.B1(net5774),
    .Y(_08026_),
    .A1(_04779_),
    .A2(_04781_));
 sg13g2_or3_1 _33749_ (.A(_07695_),
    .B(_08025_),
    .C(_08026_),
    .X(_08027_));
 sg13g2_nand2_1 _33750_ (.Y(_08028_),
    .A(net5686),
    .B(\u_inv.d_next[161] ));
 sg13g2_a21oi_1 _33751_ (.A1(_08027_),
    .A2(_08028_),
    .Y(_08029_),
    .B1(net4970));
 sg13g2_a21oi_1 _33752_ (.A1(_04783_),
    .A2(_07685_),
    .Y(_08030_),
    .B1(_04945_));
 sg13g2_xnor2_1 _33753_ (.Y(_08031_),
    .A(_04779_),
    .B(_08030_));
 sg13g2_a21oi_2 _33754_ (.B1(_08029_),
    .Y(_08032_),
    .A2(_08031_),
    .A1(net4970));
 sg13g2_nor2_1 _33755_ (.A(net4811),
    .B(_08032_),
    .Y(_08033_));
 sg13g2_xnor2_1 _33756_ (.Y(_08034_),
    .A(net4758),
    .B(_08032_));
 sg13g2_xnor2_1 _33757_ (.Y(_08035_),
    .A(_04783_),
    .B(_07685_));
 sg13g2_xnor2_1 _33758_ (.Y(_08036_),
    .A(_04782_),
    .B(_07694_));
 sg13g2_nand2_1 _33759_ (.Y(_08037_),
    .A(net5687),
    .B(\u_inv.d_next[160] ));
 sg13g2_a21oi_1 _33760_ (.A1(net5776),
    .A2(_08036_),
    .Y(_08038_),
    .B1(net4972));
 sg13g2_a22oi_1 _33761_ (.Y(_08039_),
    .B1(_08037_),
    .B2(_08038_),
    .A2(_08035_),
    .A1(net4972));
 sg13g2_nand2_1 _33762_ (.Y(_08040_),
    .A(net4758),
    .B(_08039_));
 sg13g2_xnor2_1 _33763_ (.Y(_08041_),
    .A(net4811),
    .B(_08039_));
 sg13g2_nand4_1 _33764_ (.B(_08023_),
    .C(_08034_),
    .A(_08014_),
    .Y(_08042_),
    .D(_08041_));
 sg13g2_nor3_2 _33765_ (.A(_07982_),
    .B(_08001_),
    .C(_08042_),
    .Y(_08043_));
 sg13g2_inv_1 _33766_ (.Y(_08044_),
    .A(_08043_));
 sg13g2_and3_1 _33767_ (.X(_08045_),
    .A(_07876_),
    .B(_07960_),
    .C(_08043_));
 sg13g2_o21ai_1 _33768_ (.B1(net4756),
    .Y(_08046_),
    .A1(_07863_),
    .A2(_07870_));
 sg13g2_a21oi_1 _33769_ (.A1(net4756),
    .A2(_07846_),
    .Y(_08047_),
    .B1(_07853_));
 sg13g2_o21ai_1 _33770_ (.B1(_08047_),
    .Y(_08048_),
    .A1(_07855_),
    .A2(_08046_));
 sg13g2_inv_1 _33771_ (.Y(_08049_),
    .A(_08048_));
 sg13g2_nand2b_1 _33772_ (.Y(_08050_),
    .B(_07811_),
    .A_N(_07802_));
 sg13g2_o21ai_1 _33773_ (.B1(_07824_),
    .Y(_08051_),
    .A1(net4810),
    .A2(_07833_));
 sg13g2_a221oi_1 _33774_ (.B2(_07814_),
    .C1(_08050_),
    .B1(_08051_),
    .A1(_07838_),
    .Y(_08052_),
    .A2(_08048_));
 sg13g2_nand2b_1 _33775_ (.Y(_08053_),
    .B(_07782_),
    .A_N(_08052_));
 sg13g2_nand2_1 _33776_ (.Y(_08054_),
    .A(_07770_),
    .B(_07778_));
 sg13g2_inv_1 _33777_ (.Y(_08055_),
    .A(_08054_));
 sg13g2_nand3_1 _33778_ (.B(_07761_),
    .C(_08054_),
    .A(_07752_),
    .Y(_08056_));
 sg13g2_o21ai_1 _33779_ (.B1(net4751),
    .Y(_08057_),
    .A1(_07749_),
    .A2(_07760_));
 sg13g2_nand2_2 _33780_ (.Y(_08058_),
    .A(_08056_),
    .B(_08057_));
 sg13g2_and2_1 _33781_ (.A(_07728_),
    .B(_07738_),
    .X(_08059_));
 sg13g2_nor3_1 _33782_ (.A(_07712_),
    .B(_07722_),
    .C(_08059_),
    .Y(_08060_));
 sg13g2_a21oi_1 _33783_ (.A1(_07742_),
    .A2(_08058_),
    .Y(_08061_),
    .B1(_08060_));
 sg13g2_nand4_1 _33784_ (.B(_07721_),
    .C(_08053_),
    .A(_07711_),
    .Y(_08062_),
    .D(_08061_));
 sg13g2_nor2b_1 _33785_ (.A(_07989_),
    .B_N(_07999_),
    .Y(_08063_));
 sg13g2_nor2b_1 _33786_ (.A(_08033_),
    .B_N(_08040_),
    .Y(_08064_));
 sg13g2_nand3b_1 _33787_ (.B(_08023_),
    .C(_08014_),
    .Y(_08065_),
    .A_N(_08064_));
 sg13g2_a21o_1 _33788_ (.A2(_08021_),
    .A1(_08013_),
    .B1(net4811),
    .X(_08066_));
 sg13g2_nand2_1 _33789_ (.Y(_08067_),
    .A(_08065_),
    .B(_08066_));
 sg13g2_a21oi_1 _33790_ (.A1(_08065_),
    .A2(_08066_),
    .Y(_08068_),
    .B1(_08001_));
 sg13g2_nor2b_1 _33791_ (.A(_08068_),
    .B_N(_08063_),
    .Y(_08069_));
 sg13g2_a21o_1 _33792_ (.A2(_07980_),
    .A1(_07973_),
    .B1(net4811),
    .X(_08070_));
 sg13g2_o21ai_1 _33793_ (.B1(_08070_),
    .Y(_08071_),
    .A1(_07982_),
    .A2(_08069_));
 sg13g2_nand2_1 _33794_ (.Y(_08072_),
    .A(_07960_),
    .B(_08071_));
 sg13g2_o21ai_1 _33795_ (.B1(net4757),
    .Y(_08073_),
    .A1(_07949_),
    .A2(_07956_));
 sg13g2_o21ai_1 _33796_ (.B1(net4757),
    .Y(_08074_),
    .A1(_07929_),
    .A2(_07939_));
 sg13g2_o21ai_1 _33797_ (.B1(_08074_),
    .Y(_08075_),
    .A1(_07941_),
    .A2(_08073_));
 sg13g2_inv_1 _33798_ (.Y(_08076_),
    .A(_08075_));
 sg13g2_nand4_1 _33799_ (.B(_07912_),
    .C(_07922_),
    .A(_07905_),
    .Y(_08077_),
    .D(_08075_));
 sg13g2_a21o_1 _33800_ (.A2(_07921_),
    .A1(net4757),
    .B1(_07911_),
    .X(_08078_));
 sg13g2_a21oi_1 _33801_ (.A1(_07893_),
    .A2(_07903_),
    .Y(_08079_),
    .B1(net4809));
 sg13g2_a21oi_1 _33802_ (.A1(_07905_),
    .A2(_08078_),
    .Y(_08080_),
    .B1(_08079_));
 sg13g2_nand3_1 _33803_ (.B(_08077_),
    .C(_08080_),
    .A(_08072_),
    .Y(_08081_));
 sg13g2_a21o_1 _33804_ (.A2(_08081_),
    .A1(_07876_),
    .B1(_08062_),
    .X(_08082_));
 sg13g2_nor3_2 _33805_ (.A(_07982_),
    .B(_08001_),
    .C(_08042_),
    .Y(_08083_));
 sg13g2_nand2_1 _33806_ (.Y(_08084_),
    .A(_07960_),
    .B(_08083_));
 sg13g2_and3_1 _33807_ (.X(_08085_),
    .A(_07876_),
    .B(_07960_),
    .C(_08083_));
 sg13g2_inv_1 _33808_ (.Y(_08086_),
    .A(_08085_));
 sg13g2_a221oi_1 _33809_ (.B2(_07876_),
    .C1(_08062_),
    .B1(_08081_),
    .A1(_07683_),
    .Y(_08087_),
    .A2(_08045_));
 sg13g2_o21ai_1 _33810_ (.B1(_05405_),
    .Y(_08088_),
    .A1(_05314_),
    .A2(_05347_));
 sg13g2_a21o_2 _33811_ (.A2(_05346_),
    .A1(_05315_),
    .B1(_05406_),
    .X(_08089_));
 sg13g2_and2_1 _33812_ (.A(_05684_),
    .B(_08089_),
    .X(_08090_));
 sg13g2_a21oi_2 _33813_ (.B1(_05688_),
    .Y(_08091_),
    .A2(_05567_),
    .A1(_05348_));
 sg13g2_a21o_2 _33814_ (.A2(_05567_),
    .A1(_05348_),
    .B1(_05688_),
    .X(_08092_));
 sg13g2_a21oi_1 _33815_ (.A1(_05512_),
    .A2(_08092_),
    .Y(_08093_),
    .B1(_05654_));
 sg13g2_a21o_2 _33816_ (.A2(_08092_),
    .A1(_05512_),
    .B1(_05654_),
    .X(_08094_));
 sg13g2_a21oi_2 _33817_ (.B1(_05597_),
    .Y(_08095_),
    .A2(_08094_),
    .A1(_05459_));
 sg13g2_nor3_1 _33818_ (.A(_05428_),
    .B(_05436_),
    .C(_08095_),
    .Y(_08096_));
 sg13g2_nor2_1 _33819_ (.A(_05576_),
    .B(_08096_),
    .Y(_08097_));
 sg13g2_o21ai_1 _33820_ (.B1(_05413_),
    .Y(_08098_),
    .A1(_05576_),
    .A2(_08096_));
 sg13g2_nand3_1 _33821_ (.B(_05581_),
    .C(_08098_),
    .A(_05419_),
    .Y(_08099_));
 sg13g2_a21o_1 _33822_ (.A2(_08098_),
    .A1(_05581_),
    .B1(_05419_),
    .X(_08100_));
 sg13g2_a21oi_1 _33823_ (.A1(_08099_),
    .A2(_08100_),
    .Y(_08101_),
    .B1(net5081));
 sg13g2_a21oi_1 _33824_ (.A1(_06115_),
    .A2(_06272_),
    .Y(_08102_),
    .B1(_05508_));
 sg13g2_a21oi_2 _33825_ (.B1(_05997_),
    .Y(_08103_),
    .A2(_06272_),
    .A1(_06115_));
 sg13g2_a21oi_2 _33826_ (.B1(_06031_),
    .Y(_08104_),
    .A2(_08103_),
    .A1(_05995_));
 sg13g2_a21oi_2 _33827_ (.B1(_06046_),
    .Y(_08105_),
    .A2(_06272_),
    .A1(_06115_));
 sg13g2_nor2_1 _33828_ (.A(_06044_),
    .B(_08105_),
    .Y(_08106_));
 sg13g2_o21ai_1 _33829_ (.B1(_05986_),
    .Y(_08107_),
    .A1(_06044_),
    .A2(_08105_));
 sg13g2_a21oi_1 _33830_ (.A1(_06008_),
    .A2(_08107_),
    .Y(_08108_),
    .B1(_05435_));
 sg13g2_and2_1 _33831_ (.A(_05432_),
    .B(_08108_),
    .X(_08109_));
 sg13g2_nor2_1 _33832_ (.A(_06011_),
    .B(_08109_),
    .Y(_08110_));
 sg13g2_a21oi_2 _33833_ (.B1(_06013_),
    .Y(_08111_),
    .A2(_08109_),
    .A1(_05979_));
 sg13g2_o21ai_1 _33834_ (.B1(_06017_),
    .Y(_08112_),
    .A1(_05977_),
    .A2(_08111_));
 sg13g2_xnor2_1 _33835_ (.Y(_08113_),
    .A(_05420_),
    .B(_08112_));
 sg13g2_nand2_1 _33836_ (.Y(_08114_),
    .A(net5705),
    .B(\u_inv.d_next[126] ));
 sg13g2_a21oi_1 _33837_ (.A1(net5800),
    .A2(_08113_),
    .Y(_08115_),
    .B1(net4994));
 sg13g2_a21oi_1 _33838_ (.A1(_08114_),
    .A2(_08115_),
    .Y(_08116_),
    .B1(_08101_));
 sg13g2_and2_1 _33839_ (.A(net4771),
    .B(_08116_),
    .X(_08117_));
 sg13g2_xnor2_1 _33840_ (.Y(_08118_),
    .A(net4771),
    .B(_08116_));
 sg13g2_inv_1 _33841_ (.Y(_08119_),
    .A(_08118_));
 sg13g2_a21oi_1 _33842_ (.A1(_05578_),
    .A2(_08100_),
    .Y(_08120_),
    .B1(_05416_));
 sg13g2_nand3_1 _33843_ (.B(_05578_),
    .C(_08100_),
    .A(_05416_),
    .Y(_08121_));
 sg13g2_nor2_1 _33844_ (.A(net5081),
    .B(_08120_),
    .Y(_08122_));
 sg13g2_a21oi_1 _33845_ (.A1(_05419_),
    .A2(_08112_),
    .Y(_08123_),
    .B1(_05418_));
 sg13g2_xor2_1 _33846_ (.B(_08123_),
    .A(_05416_),
    .X(_08124_));
 sg13g2_nand2_1 _33847_ (.Y(_08125_),
    .A(net5700),
    .B(\u_inv.d_next[127] ));
 sg13g2_a21oi_1 _33848_ (.A1(net5800),
    .A2(_08124_),
    .Y(_08126_),
    .B1(net4994));
 sg13g2_a22oi_1 _33849_ (.Y(_08127_),
    .B1(_08125_),
    .B2(_08126_),
    .A2(_08122_),
    .A1(_08121_));
 sg13g2_xnor2_1 _33850_ (.Y(_08128_),
    .A(net4819),
    .B(_08127_));
 sg13g2_xnor2_1 _33851_ (.Y(_08129_),
    .A(net4771),
    .B(_08127_));
 sg13g2_o21ai_1 _33852_ (.B1(_05579_),
    .Y(_08130_),
    .A1(_05410_),
    .A2(_08097_));
 sg13g2_nand2b_1 _33853_ (.Y(_08131_),
    .B(_05408_),
    .A_N(_08130_));
 sg13g2_a21oi_1 _33854_ (.A1(_05407_),
    .A2(_08130_),
    .Y(_08132_),
    .B1(net5084));
 sg13g2_o21ai_1 _33855_ (.B1(_05409_),
    .Y(_08133_),
    .A1(_05411_),
    .A2(_08111_));
 sg13g2_xnor2_1 _33856_ (.Y(_08134_),
    .A(_05408_),
    .B(_08133_));
 sg13g2_nand2_1 _33857_ (.Y(_08135_),
    .A(net5705),
    .B(\u_inv.d_next[125] ));
 sg13g2_a21oi_1 _33858_ (.A1(net5800),
    .A2(_08134_),
    .Y(_08136_),
    .B1(net4999));
 sg13g2_a22oi_1 _33859_ (.Y(_08137_),
    .B1(_08135_),
    .B2(_08136_),
    .A2(_08132_),
    .A1(_08131_));
 sg13g2_xnor2_1 _33860_ (.Y(_08138_),
    .A(net4820),
    .B(_08137_));
 sg13g2_xnor2_1 _33861_ (.Y(_08139_),
    .A(_05410_),
    .B(_08097_));
 sg13g2_xnor2_1 _33862_ (.Y(_08140_),
    .A(_05410_),
    .B(_08111_));
 sg13g2_nand2_1 _33863_ (.Y(_08141_),
    .A(net5701),
    .B(\u_inv.d_next[124] ));
 sg13g2_a21oi_1 _33864_ (.A1(net5800),
    .A2(_08140_),
    .Y(_08142_),
    .B1(net4993));
 sg13g2_a22oi_1 _33865_ (.Y(_08143_),
    .B1(_08141_),
    .B2(_08142_),
    .A2(_08139_),
    .A1(net4993));
 sg13g2_and2_1 _33866_ (.A(net4771),
    .B(_08143_),
    .X(_08144_));
 sg13g2_xnor2_1 _33867_ (.Y(_08145_),
    .A(net4820),
    .B(_08143_));
 sg13g2_and2_1 _33868_ (.A(_08138_),
    .B(_08145_),
    .X(_08146_));
 sg13g2_nand2_1 _33869_ (.Y(_08147_),
    .A(_08138_),
    .B(_08145_));
 sg13g2_o21ai_1 _33870_ (.B1(_05574_),
    .Y(_08148_),
    .A1(_05436_),
    .A2(_08095_));
 sg13g2_xor2_1 _33871_ (.B(_08148_),
    .A(_05427_),
    .X(_08149_));
 sg13g2_xnor2_1 _33872_ (.Y(_08150_),
    .A(_05427_),
    .B(_08110_));
 sg13g2_a21oi_1 _33873_ (.A1(net5700),
    .A2(\u_inv.d_next[122] ),
    .Y(_08151_),
    .B1(net4993));
 sg13g2_o21ai_1 _33874_ (.B1(_08151_),
    .Y(_08152_),
    .A1(net5700),
    .A2(_08150_));
 sg13g2_o21ai_1 _33875_ (.B1(_08152_),
    .Y(_08153_),
    .A1(net5081),
    .A2(_08149_));
 sg13g2_nand2b_1 _33876_ (.Y(_08154_),
    .B(net4775),
    .A_N(_08153_));
 sg13g2_xnor2_1 _33877_ (.Y(_08155_),
    .A(net4822),
    .B(_08153_));
 sg13g2_inv_1 _33878_ (.Y(_08156_),
    .A(_08155_));
 sg13g2_a21oi_1 _33879_ (.A1(_05427_),
    .A2(_08148_),
    .Y(_08157_),
    .B1(_05571_));
 sg13g2_nand2b_1 _33880_ (.Y(_08158_),
    .B(_05425_),
    .A_N(_08157_));
 sg13g2_a21oi_1 _33881_ (.A1(_05424_),
    .A2(_08157_),
    .Y(_08159_),
    .B1(net5081));
 sg13g2_o21ai_1 _33882_ (.B1(_05426_),
    .Y(_08160_),
    .A1(_05427_),
    .A2(_08110_));
 sg13g2_xnor2_1 _33883_ (.Y(_08161_),
    .A(_05424_),
    .B(_08160_));
 sg13g2_nand2_1 _33884_ (.Y(_08162_),
    .A(net5700),
    .B(\u_inv.d_next[123] ));
 sg13g2_a21oi_1 _33885_ (.A1(net5804),
    .A2(_08161_),
    .Y(_08163_),
    .B1(net4993));
 sg13g2_a22oi_1 _33886_ (.Y(_08164_),
    .B1(_08162_),
    .B2(_08163_),
    .A2(_08159_),
    .A1(_08158_));
 sg13g2_nand2_1 _33887_ (.Y(_08165_),
    .A(net4775),
    .B(_08164_));
 sg13g2_xnor2_1 _33888_ (.Y(_08166_),
    .A(net4822),
    .B(_08164_));
 sg13g2_o21ai_1 _33889_ (.B1(_05572_),
    .Y(_08167_),
    .A1(_05434_),
    .A2(_08095_));
 sg13g2_o21ai_1 _33890_ (.B1(net4993),
    .Y(_08168_),
    .A1(_05432_),
    .A2(_08167_));
 sg13g2_a21oi_1 _33891_ (.A1(_05432_),
    .A2(_08167_),
    .Y(_08169_),
    .B1(_08168_));
 sg13g2_nand2_1 _33892_ (.Y(_08170_),
    .A(_05431_),
    .B(_05433_));
 sg13g2_o21ai_1 _33893_ (.B1(net5804),
    .Y(_08171_),
    .A1(_05431_),
    .A2(_05433_));
 sg13g2_nor2_1 _33894_ (.A(_08109_),
    .B(_08171_),
    .Y(_08172_));
 sg13g2_o21ai_1 _33895_ (.B1(_08172_),
    .Y(_08173_),
    .A1(_08108_),
    .A2(_08170_));
 sg13g2_a21oi_1 _33896_ (.A1(net5702),
    .A2(\u_inv.d_next[121] ),
    .Y(_08174_),
    .B1(net4993));
 sg13g2_a21o_2 _33897_ (.A2(_08174_),
    .A1(_08173_),
    .B1(_08169_),
    .X(_08175_));
 sg13g2_xnor2_1 _33898_ (.Y(_08176_),
    .A(net4775),
    .B(_08175_));
 sg13g2_nand3_1 _33899_ (.B(_06008_),
    .C(_08107_),
    .A(_05435_),
    .Y(_08177_));
 sg13g2_nor2_1 _33900_ (.A(net5702),
    .B(_08108_),
    .Y(_08178_));
 sg13g2_xnor2_1 _33901_ (.Y(_08179_),
    .A(_05434_),
    .B(_08095_));
 sg13g2_a221oi_1 _33902_ (.B2(_08178_),
    .C1(net4993),
    .B1(_08177_),
    .A1(net5702),
    .Y(_08180_),
    .A2(\u_inv.d_next[120] ));
 sg13g2_a21oi_2 _33903_ (.B1(_08180_),
    .Y(_08181_),
    .A2(_08179_),
    .A1(net4993));
 sg13g2_nand2_1 _33904_ (.Y(_08182_),
    .A(net4775),
    .B(_08181_));
 sg13g2_xnor2_1 _33905_ (.Y(_08183_),
    .A(net4775),
    .B(_08181_));
 sg13g2_inv_1 _33906_ (.Y(_08184_),
    .A(_08183_));
 sg13g2_nand4_1 _33907_ (.B(_08166_),
    .C(_08176_),
    .A(_08156_),
    .Y(_08185_),
    .D(_08184_));
 sg13g2_nor4_2 _33908_ (.A(_08118_),
    .B(_08129_),
    .C(_08147_),
    .Y(_08186_),
    .D(_08185_));
 sg13g2_nor3_1 _33909_ (.A(_05451_),
    .B(_05458_),
    .C(_08093_),
    .Y(_08187_));
 sg13g2_or2_1 _33910_ (.X(_08188_),
    .B(_08187_),
    .A(_05590_));
 sg13g2_o21ai_1 _33911_ (.B1(_05441_),
    .Y(_08189_),
    .A1(_05590_),
    .A2(_08187_));
 sg13g2_a21o_1 _33912_ (.A2(_08189_),
    .A1(_05593_),
    .B1(_05443_),
    .X(_08190_));
 sg13g2_a21o_1 _33913_ (.A2(_08190_),
    .A1(_05594_),
    .B1(_05446_),
    .X(_08191_));
 sg13g2_nand3_1 _33914_ (.B(_05594_),
    .C(_08190_),
    .A(_05446_),
    .Y(_08192_));
 sg13g2_nand3_1 _33915_ (.B(_08191_),
    .C(_08192_),
    .A(net4997),
    .Y(_08193_));
 sg13g2_or3_1 _33916_ (.A(_05454_),
    .B(_05457_),
    .C(_08106_),
    .X(_08194_));
 sg13g2_o21ai_1 _33917_ (.B1(_05984_),
    .Y(_08195_),
    .A1(_06044_),
    .A2(_08105_));
 sg13g2_nand2_1 _33918_ (.Y(_08196_),
    .A(_06002_),
    .B(_08195_));
 sg13g2_a21oi_1 _33919_ (.A1(_06002_),
    .A2(_08195_),
    .Y(_08197_),
    .B1(_05440_));
 sg13g2_and2_1 _33920_ (.A(_05439_),
    .B(_08197_),
    .X(_08198_));
 sg13g2_inv_1 _33921_ (.Y(_08199_),
    .A(_08198_));
 sg13g2_o21ai_1 _33922_ (.B1(_05443_),
    .Y(_08200_),
    .A1(_06005_),
    .A2(_08198_));
 sg13g2_nand3_1 _33923_ (.B(_05446_),
    .C(_08200_),
    .A(_05442_),
    .Y(_08201_));
 sg13g2_a21o_1 _33924_ (.A2(_08200_),
    .A1(_05442_),
    .B1(_05446_),
    .X(_08202_));
 sg13g2_nand3_1 _33925_ (.B(_08201_),
    .C(_08202_),
    .A(net5802),
    .Y(_08203_));
 sg13g2_nand2_1 _33926_ (.Y(_08204_),
    .A(net5702),
    .B(\u_inv.d_next[119] ));
 sg13g2_nand3_1 _33927_ (.B(_08203_),
    .C(_08204_),
    .A(net5082),
    .Y(_08205_));
 sg13g2_nand3_1 _33928_ (.B(_08193_),
    .C(_08205_),
    .A(net4773),
    .Y(_08206_));
 sg13g2_a21o_1 _33929_ (.A2(_08205_),
    .A1(_08193_),
    .B1(net4773),
    .X(_08207_));
 sg13g2_and2_1 _33930_ (.A(_08206_),
    .B(_08207_),
    .X(_08208_));
 sg13g2_nand3_1 _33931_ (.B(_05593_),
    .C(_08189_),
    .A(_05443_),
    .Y(_08209_));
 sg13g2_a21oi_1 _33932_ (.A1(_08190_),
    .A2(_08209_),
    .Y(_08210_),
    .B1(net5082));
 sg13g2_or3_1 _33933_ (.A(_05443_),
    .B(_06005_),
    .C(_08198_),
    .X(_08211_));
 sg13g2_nand3_1 _33934_ (.B(_08200_),
    .C(_08211_),
    .A(net5802),
    .Y(_08212_));
 sg13g2_a21oi_1 _33935_ (.A1(net5702),
    .A2(\u_inv.d_next[118] ),
    .Y(_08213_),
    .B1(net4997));
 sg13g2_a21o_2 _33936_ (.A2(_08213_),
    .A1(_08212_),
    .B1(_08210_),
    .X(_08214_));
 sg13g2_nand2b_1 _33937_ (.Y(_08215_),
    .B(net4773),
    .A_N(_08214_));
 sg13g2_xnor2_1 _33938_ (.Y(_08216_),
    .A(net4773),
    .B(_08214_));
 sg13g2_inv_1 _33939_ (.Y(_08217_),
    .A(_08216_));
 sg13g2_nand2_1 _33940_ (.Y(_08218_),
    .A(_08208_),
    .B(_08216_));
 sg13g2_a21o_1 _33941_ (.A2(_08188_),
    .A1(_05440_),
    .B1(_05591_),
    .X(_08219_));
 sg13g2_o21ai_1 _33942_ (.B1(net5002),
    .Y(_08220_),
    .A1(_05439_),
    .A2(_08219_));
 sg13g2_a21oi_1 _33943_ (.A1(_05439_),
    .A2(_08219_),
    .Y(_08221_),
    .B1(_08220_));
 sg13g2_a21oi_1 _33944_ (.A1(\u_inv.d_next[116] ),
    .A2(\u_inv.d_reg[116] ),
    .Y(_08222_),
    .B1(_08197_));
 sg13g2_nand2_1 _33945_ (.Y(_08223_),
    .A(_05438_),
    .B(_08222_));
 sg13g2_nand4_1 _33946_ (.B(_06004_),
    .C(_08199_),
    .A(net5810),
    .Y(_08224_),
    .D(_08223_));
 sg13g2_a21oi_1 _33947_ (.A1(net5708),
    .A2(\u_inv.d_next[117] ),
    .Y(_08225_),
    .B1(net5002));
 sg13g2_a21oi_2 _33948_ (.B1(_08221_),
    .Y(_08226_),
    .A2(_08225_),
    .A1(_08224_));
 sg13g2_xnor2_1 _33949_ (.Y(_08227_),
    .A(net4822),
    .B(_08226_));
 sg13g2_xnor2_1 _33950_ (.Y(_08228_),
    .A(net4773),
    .B(_08226_));
 sg13g2_xor2_1 _33951_ (.B(_08196_),
    .A(_05440_),
    .X(_08229_));
 sg13g2_o21ai_1 _33952_ (.B1(net5089),
    .Y(_08230_),
    .A1(net5802),
    .A2(\u_inv.d_next[116] ));
 sg13g2_a21o_1 _33953_ (.A2(_08229_),
    .A1(net5803),
    .B1(_08230_),
    .X(_08231_));
 sg13g2_xnor2_1 _33954_ (.Y(_08232_),
    .A(_05440_),
    .B(_08188_));
 sg13g2_o21ai_1 _33955_ (.B1(_08231_),
    .Y(_08233_),
    .A1(net5082),
    .A2(_08232_));
 sg13g2_and2_1 _33956_ (.A(net4773),
    .B(_08233_),
    .X(_08234_));
 sg13g2_xnor2_1 _33957_ (.Y(_08235_),
    .A(net4773),
    .B(_08233_));
 sg13g2_o21ai_1 _33958_ (.B1(_05585_),
    .Y(_08236_),
    .A1(_05458_),
    .A2(_08093_));
 sg13g2_a21oi_1 _33959_ (.A1(_05450_),
    .A2(_08236_),
    .Y(_08237_),
    .B1(_05587_));
 sg13g2_or2_1 _33960_ (.X(_08238_),
    .B(_08237_),
    .A(_05449_));
 sg13g2_a21oi_1 _33961_ (.A1(_05449_),
    .A2(_08237_),
    .Y(_08239_),
    .B1(net5082));
 sg13g2_a21oi_1 _33962_ (.A1(_06000_),
    .A2(_08194_),
    .Y(_08240_),
    .B1(_05450_));
 sg13g2_a21oi_1 _33963_ (.A1(\u_inv.d_next[114] ),
    .A2(\u_inv.d_reg[114] ),
    .Y(_08241_),
    .B1(_08240_));
 sg13g2_o21ai_1 _33964_ (.B1(net5803),
    .Y(_08242_),
    .A1(_05449_),
    .A2(_08241_));
 sg13g2_a21o_1 _33965_ (.A2(_08241_),
    .A1(_05449_),
    .B1(_08242_),
    .X(_08243_));
 sg13g2_a21oi_1 _33966_ (.A1(net5704),
    .A2(\u_inv.d_next[115] ),
    .Y(_08244_),
    .B1(net4997));
 sg13g2_a22oi_1 _33967_ (.Y(_08245_),
    .B1(_08243_),
    .B2(_08244_),
    .A2(_08239_),
    .A1(_08238_));
 sg13g2_xnor2_1 _33968_ (.Y(_08246_),
    .A(net4821),
    .B(_08245_));
 sg13g2_xor2_1 _33969_ (.B(_08236_),
    .A(_05450_),
    .X(_08247_));
 sg13g2_and3_1 _33970_ (.X(_08248_),
    .A(_05450_),
    .B(_06000_),
    .C(_08194_));
 sg13g2_nor3_1 _33971_ (.A(net5704),
    .B(_08240_),
    .C(_08248_),
    .Y(_08249_));
 sg13g2_a21oi_1 _33972_ (.A1(net5702),
    .A2(\u_inv.d_next[114] ),
    .Y(_08250_),
    .B1(net4997));
 sg13g2_nand2b_1 _33973_ (.Y(_08251_),
    .B(_08250_),
    .A_N(_08249_));
 sg13g2_o21ai_1 _33974_ (.B1(_08251_),
    .Y(_08252_),
    .A1(net5084),
    .A2(_08247_));
 sg13g2_nor2_1 _33975_ (.A(net4822),
    .B(_08252_),
    .Y(_08253_));
 sg13g2_xnor2_1 _33976_ (.Y(_08254_),
    .A(net4774),
    .B(_08252_));
 sg13g2_a21oi_1 _33977_ (.A1(_05457_),
    .A2(_08094_),
    .Y(_08255_),
    .B1(_05584_));
 sg13g2_o21ai_1 _33978_ (.B1(net4997),
    .Y(_08256_),
    .A1(_05454_),
    .A2(_08255_));
 sg13g2_a21oi_1 _33979_ (.A1(_05454_),
    .A2(_08255_),
    .Y(_08257_),
    .B1(_08256_));
 sg13g2_nor2_1 _33980_ (.A(_05455_),
    .B(_05456_),
    .Y(_08258_));
 sg13g2_o21ai_1 _33981_ (.B1(_08258_),
    .Y(_08259_),
    .A1(_05457_),
    .A2(_08106_));
 sg13g2_a21oi_1 _33982_ (.A1(_05455_),
    .A2(_05456_),
    .Y(_08260_),
    .B1(net5702));
 sg13g2_nand3_1 _33983_ (.B(_08259_),
    .C(_08260_),
    .A(_08194_),
    .Y(_08261_));
 sg13g2_a21oi_1 _33984_ (.A1(net5704),
    .A2(\u_inv.d_next[113] ),
    .Y(_08262_),
    .B1(net4998));
 sg13g2_a21oi_2 _33985_ (.B1(_08257_),
    .Y(_08263_),
    .A2(_08262_),
    .A1(_08261_));
 sg13g2_nor2_1 _33986_ (.A(net4774),
    .B(_08263_),
    .Y(_08264_));
 sg13g2_xnor2_1 _33987_ (.Y(_08265_),
    .A(net4822),
    .B(_08263_));
 sg13g2_xnor2_1 _33988_ (.Y(_08266_),
    .A(_05457_),
    .B(_08106_));
 sg13g2_o21ai_1 _33989_ (.B1(net5083),
    .Y(_08267_),
    .A1(net5803),
    .A2(\u_inv.d_next[112] ));
 sg13g2_a21o_1 _33990_ (.A2(_08266_),
    .A1(net5803),
    .B1(_08267_),
    .X(_08268_));
 sg13g2_xnor2_1 _33991_ (.Y(_08269_),
    .A(_05457_),
    .B(_08094_));
 sg13g2_o21ai_1 _33992_ (.B1(_08268_),
    .Y(_08270_),
    .A1(net5083),
    .A2(_08269_));
 sg13g2_nand2_1 _33993_ (.Y(_08271_),
    .A(net4776),
    .B(_08270_));
 sg13g2_xnor2_1 _33994_ (.Y(_08272_),
    .A(net4822),
    .B(_08270_));
 sg13g2_nand4_1 _33995_ (.B(_08254_),
    .C(_08265_),
    .A(_08246_),
    .Y(_08273_),
    .D(_08272_));
 sg13g2_nor4_2 _33996_ (.A(_08218_),
    .B(_08228_),
    .C(_08235_),
    .Y(_08274_),
    .D(_08273_));
 sg13g2_and2_1 _33997_ (.A(_08186_),
    .B(_08274_),
    .X(_08275_));
 sg13g2_o21ai_1 _33998_ (.B1(_05639_),
    .Y(_08276_),
    .A1(_05511_),
    .A2(_08091_));
 sg13g2_a21oi_2 _33999_ (.B1(_05646_),
    .Y(_08277_),
    .A2(_08276_),
    .A1(_05484_));
 sg13g2_o21ai_1 _34000_ (.B1(_05649_),
    .Y(_08278_),
    .A1(_05471_),
    .A2(_08277_));
 sg13g2_nand2_1 _34001_ (.Y(_08279_),
    .A(_05465_),
    .B(_08278_));
 sg13g2_xor2_1 _34002_ (.B(_08278_),
    .A(_05465_),
    .X(_08280_));
 sg13g2_nor2_1 _34003_ (.A(_05482_),
    .B(_08104_),
    .Y(_08281_));
 sg13g2_nand2_1 _34004_ (.Y(_08282_),
    .A(_05480_),
    .B(_08281_));
 sg13g2_nor3_1 _34005_ (.A(_05991_),
    .B(_05992_),
    .C(_08104_),
    .Y(_08283_));
 sg13g2_o21ai_1 _34006_ (.B1(_05470_),
    .Y(_08284_),
    .A1(_06037_),
    .A2(_08283_));
 sg13g2_o21ai_1 _34007_ (.B1(_05989_),
    .Y(_08285_),
    .A1(_06037_),
    .A2(_08283_));
 sg13g2_and3_1 _34008_ (.X(_08286_),
    .A(_05465_),
    .B(_06041_),
    .C(_08285_));
 sg13g2_a21oi_1 _34009_ (.A1(_06041_),
    .A2(_08285_),
    .Y(_08287_),
    .B1(_05465_));
 sg13g2_nor3_1 _34010_ (.A(net5709),
    .B(_08286_),
    .C(_08287_),
    .Y(_08288_));
 sg13g2_a21oi_1 _34011_ (.A1(net5702),
    .A2(\u_inv.d_next[110] ),
    .Y(_08289_),
    .B1(net4997));
 sg13g2_nand2b_1 _34012_ (.Y(_08290_),
    .B(_08289_),
    .A_N(_08288_));
 sg13g2_o21ai_1 _34013_ (.B1(_08290_),
    .Y(_08291_),
    .A1(net5082),
    .A2(_08280_));
 sg13g2_nand2b_1 _34014_ (.Y(_08292_),
    .B(net4781),
    .A_N(_08291_));
 sg13g2_xnor2_1 _34015_ (.Y(_08293_),
    .A(net4824),
    .B(_08291_));
 sg13g2_inv_1 _34016_ (.Y(_08294_),
    .A(_08293_));
 sg13g2_and2_1 _34017_ (.A(_05650_),
    .B(_08279_),
    .X(_08295_));
 sg13g2_nand2b_1 _34018_ (.Y(_08296_),
    .B(_05462_),
    .A_N(_08295_));
 sg13g2_a21oi_1 _34019_ (.A1(_05463_),
    .A2(_08295_),
    .Y(_08297_),
    .B1(net5082));
 sg13g2_nor2_1 _34020_ (.A(_05464_),
    .B(_08287_),
    .Y(_08298_));
 sg13g2_a21oi_1 _34021_ (.A1(_05463_),
    .A2(_08298_),
    .Y(_08299_),
    .B1(net5709));
 sg13g2_o21ai_1 _34022_ (.B1(_08299_),
    .Y(_08300_),
    .A1(_05463_),
    .A2(_08298_));
 sg13g2_a21oi_1 _34023_ (.A1(net5709),
    .A2(\u_inv.d_next[111] ),
    .Y(_08301_),
    .B1(net4997));
 sg13g2_a22oi_1 _34024_ (.Y(_08302_),
    .B1(_08300_),
    .B2(_08301_),
    .A2(_08297_),
    .A1(_08296_));
 sg13g2_xnor2_1 _34025_ (.Y(_08303_),
    .A(net4781),
    .B(_08302_));
 sg13g2_nor2_1 _34026_ (.A(_08293_),
    .B(_08303_),
    .Y(_08304_));
 sg13g2_nor2_1 _34027_ (.A(_05470_),
    .B(_08277_),
    .Y(_08305_));
 sg13g2_or2_1 _34028_ (.X(_08306_),
    .B(_08305_),
    .A(_05648_));
 sg13g2_or2_1 _34029_ (.X(_08307_),
    .B(_08306_),
    .A(_05469_));
 sg13g2_a21oi_1 _34030_ (.A1(_05469_),
    .A2(_08306_),
    .Y(_08308_),
    .B1(net5082));
 sg13g2_a21oi_1 _34031_ (.A1(\u_inv.d_next[108] ),
    .A2(\u_inv.d_reg[108] ),
    .Y(_08309_),
    .B1(_05469_));
 sg13g2_nand3b_1 _34032_ (.B(_08285_),
    .C(net5812),
    .Y(_08310_),
    .A_N(_06040_));
 sg13g2_a21oi_1 _34033_ (.A1(_08284_),
    .A2(_08309_),
    .Y(_08311_),
    .B1(_08310_));
 sg13g2_a21oi_1 _34034_ (.A1(net5716),
    .A2(\u_inv.d_next[109] ),
    .Y(_08312_),
    .B1(_08311_));
 sg13g2_a22oi_1 _34035_ (.Y(_08313_),
    .B1(_08312_),
    .B2(net5082),
    .A2(_08308_),
    .A1(_08307_));
 sg13g2_xnor2_1 _34036_ (.Y(_08314_),
    .A(net4824),
    .B(_08313_));
 sg13g2_xor2_1 _34037_ (.B(_08277_),
    .A(_05470_),
    .X(_08315_));
 sg13g2_nor3_1 _34038_ (.A(_05470_),
    .B(_06037_),
    .C(_08283_),
    .Y(_08316_));
 sg13g2_nand2_1 _34039_ (.Y(_08317_),
    .A(net5812),
    .B(_08284_));
 sg13g2_a21oi_1 _34040_ (.A1(net5709),
    .A2(\u_inv.d_next[108] ),
    .Y(_08318_),
    .B1(net4997));
 sg13g2_o21ai_1 _34041_ (.B1(_08318_),
    .Y(_08319_),
    .A1(_08316_),
    .A2(_08317_));
 sg13g2_o21ai_1 _34042_ (.B1(_08319_),
    .Y(_08320_),
    .A1(net5091),
    .A2(_08315_));
 sg13g2_nor2_1 _34043_ (.A(net4824),
    .B(_08320_),
    .Y(_08321_));
 sg13g2_xnor2_1 _34044_ (.Y(_08322_),
    .A(net4781),
    .B(_08320_));
 sg13g2_nand2_1 _34045_ (.Y(_08323_),
    .A(_08314_),
    .B(_08322_));
 sg13g2_a21oi_1 _34046_ (.A1(_05483_),
    .A2(_08276_),
    .Y(_08324_),
    .B1(_05643_));
 sg13g2_o21ai_1 _34047_ (.B1(_05644_),
    .Y(_08325_),
    .A1(_05477_),
    .A2(_08324_));
 sg13g2_or2_1 _34048_ (.X(_08326_),
    .B(_08325_),
    .A(_05475_));
 sg13g2_a21oi_1 _34049_ (.A1(_05475_),
    .A2(_08325_),
    .Y(_08327_),
    .B1(net5091));
 sg13g2_a21o_1 _34050_ (.A2(_08282_),
    .A1(_06034_),
    .B1(_05478_),
    .X(_08328_));
 sg13g2_nand3_1 _34051_ (.B(_05476_),
    .C(_08328_),
    .A(_05474_),
    .Y(_08329_));
 sg13g2_a21o_1 _34052_ (.A2(_08328_),
    .A1(_05476_),
    .B1(_05474_),
    .X(_08330_));
 sg13g2_nand3_1 _34053_ (.B(_08329_),
    .C(_08330_),
    .A(net5812),
    .Y(_08331_));
 sg13g2_a21oi_1 _34054_ (.A1(net5709),
    .A2(\u_inv.d_next[107] ),
    .Y(_08332_),
    .B1(net5005));
 sg13g2_a22oi_1 _34055_ (.Y(_08333_),
    .B1(_08331_),
    .B2(_08332_),
    .A2(_08327_),
    .A1(_08326_));
 sg13g2_xnor2_1 _34056_ (.Y(_08334_),
    .A(net4823),
    .B(_08333_));
 sg13g2_xnor2_1 _34057_ (.Y(_08335_),
    .A(_05477_),
    .B(_08324_));
 sg13g2_nand3_1 _34058_ (.B(_06034_),
    .C(_08282_),
    .A(_05478_),
    .Y(_08336_));
 sg13g2_and2_1 _34059_ (.A(net5812),
    .B(_08328_),
    .X(_08337_));
 sg13g2_nand2_1 _34060_ (.Y(_08338_),
    .A(net5709),
    .B(\u_inv.d_next[106] ));
 sg13g2_a21oi_1 _34061_ (.A1(_08336_),
    .A2(_08337_),
    .Y(_08339_),
    .B1(net5005));
 sg13g2_a22oi_1 _34062_ (.Y(_08340_),
    .B1(_08338_),
    .B2(_08339_),
    .A2(_08335_),
    .A1(net5005));
 sg13g2_nand2_1 _34063_ (.Y(_08341_),
    .A(net4779),
    .B(_08340_));
 sg13g2_inv_1 _34064_ (.Y(_08342_),
    .A(_08341_));
 sg13g2_xnor2_1 _34065_ (.Y(_08343_),
    .A(net4823),
    .B(_08340_));
 sg13g2_nand2_1 _34066_ (.Y(_08344_),
    .A(_08334_),
    .B(_08343_));
 sg13g2_xnor2_1 _34067_ (.Y(_08345_),
    .A(_05482_),
    .B(_08104_));
 sg13g2_o21ai_1 _34068_ (.B1(net5091),
    .Y(_08346_),
    .A1(net5812),
    .A2(\u_inv.d_next[104] ));
 sg13g2_a21o_1 _34069_ (.A2(_08345_),
    .A1(net5812),
    .B1(_08346_),
    .X(_08347_));
 sg13g2_xnor2_1 _34070_ (.Y(_08348_),
    .A(_05482_),
    .B(_08276_));
 sg13g2_o21ai_1 _34071_ (.B1(_08347_),
    .Y(_08349_),
    .A1(net5091),
    .A2(_08348_));
 sg13g2_and2_1 _34072_ (.A(net4779),
    .B(_08349_),
    .X(_08350_));
 sg13g2_xnor2_1 _34073_ (.Y(_08351_),
    .A(net4779),
    .B(_08349_));
 sg13g2_nor3_1 _34074_ (.A(_05480_),
    .B(_05481_),
    .C(_08281_),
    .Y(_08352_));
 sg13g2_nand3_1 _34075_ (.B(_06032_),
    .C(_08282_),
    .A(net5812),
    .Y(_08353_));
 sg13g2_nand2_1 _34076_ (.Y(_08354_),
    .A(net5709),
    .B(\u_inv.d_next[105] ));
 sg13g2_o21ai_1 _34077_ (.B1(_08354_),
    .Y(_08355_),
    .A1(_08352_),
    .A2(_08353_));
 sg13g2_a21oi_1 _34078_ (.A1(_05482_),
    .A2(_08276_),
    .Y(_08356_),
    .B1(_05641_));
 sg13g2_or2_1 _34079_ (.X(_08357_),
    .B(_08356_),
    .A(_05480_));
 sg13g2_a21oi_1 _34080_ (.A1(_05480_),
    .A2(_08356_),
    .Y(_08358_),
    .B1(net5091));
 sg13g2_a22oi_1 _34081_ (.Y(_08359_),
    .B1(_08357_),
    .B2(_08358_),
    .A2(_08355_),
    .A1(net5091));
 sg13g2_nor2_1 _34082_ (.A(net4823),
    .B(_08359_),
    .Y(_08360_));
 sg13g2_xnor2_1 _34083_ (.Y(_08361_),
    .A(net4824),
    .B(_08359_));
 sg13g2_or3_1 _34084_ (.A(_08344_),
    .B(_08351_),
    .C(_08361_),
    .X(_08362_));
 sg13g2_inv_1 _34085_ (.Y(_08363_),
    .A(_08362_));
 sg13g2_nor4_1 _34086_ (.A(_08293_),
    .B(_08303_),
    .C(_08323_),
    .D(_08362_),
    .Y(_08364_));
 sg13g2_a21oi_1 _34087_ (.A1(_05510_),
    .A2(_08092_),
    .Y(_08365_),
    .B1(_05631_));
 sg13g2_o21ai_1 _34088_ (.B1(_05637_),
    .Y(_08366_),
    .A1(_05493_),
    .A2(_08365_));
 sg13g2_nand2_1 _34089_ (.Y(_08367_),
    .A(_05489_),
    .B(_08366_));
 sg13g2_xor2_1 _34090_ (.B(_08366_),
    .A(_05489_),
    .X(_08368_));
 sg13g2_nor2_2 _34091_ (.A(_06024_),
    .B(_08103_),
    .Y(_08369_));
 sg13g2_or2_1 _34092_ (.X(_08370_),
    .B(_08369_),
    .A(_05994_));
 sg13g2_and2_1 _34093_ (.A(_06027_),
    .B(_08370_),
    .X(_08371_));
 sg13g2_xnor2_1 _34094_ (.Y(_08372_),
    .A(_05489_),
    .B(_08371_));
 sg13g2_a21oi_1 _34095_ (.A1(net5709),
    .A2(\u_inv.d_next[102] ),
    .Y(_08373_),
    .B1(net5005));
 sg13g2_o21ai_1 _34096_ (.B1(_08373_),
    .Y(_08374_),
    .A1(net5710),
    .A2(_08372_));
 sg13g2_o21ai_1 _34097_ (.B1(_08374_),
    .Y(_08375_),
    .A1(net5092),
    .A2(_08368_));
 sg13g2_nand2b_1 _34098_ (.Y(_08376_),
    .B(net4779),
    .A_N(_08375_));
 sg13g2_inv_1 _34099_ (.Y(_08377_),
    .A(_08376_));
 sg13g2_xnor2_1 _34100_ (.Y(_08378_),
    .A(net4779),
    .B(_08375_));
 sg13g2_and2_1 _34101_ (.A(_05633_),
    .B(_08367_),
    .X(_08379_));
 sg13g2_and2_1 _34102_ (.A(_05487_),
    .B(_08379_),
    .X(_08380_));
 sg13g2_o21ai_1 _34103_ (.B1(net5005),
    .Y(_08381_),
    .A1(_05487_),
    .A2(_08379_));
 sg13g2_o21ai_1 _34104_ (.B1(_05488_),
    .Y(_08382_),
    .A1(_05489_),
    .A2(_08371_));
 sg13g2_xnor2_1 _34105_ (.Y(_08383_),
    .A(_05487_),
    .B(_08382_));
 sg13g2_a21oi_1 _34106_ (.A1(net5813),
    .A2(_08383_),
    .Y(_08384_),
    .B1(net5005));
 sg13g2_o21ai_1 _34107_ (.B1(_08384_),
    .Y(_08385_),
    .A1(net5813),
    .A2(_14218_));
 sg13g2_o21ai_1 _34108_ (.B1(_08385_),
    .Y(_08386_),
    .A1(_08380_),
    .A2(_08381_));
 sg13g2_xnor2_1 _34109_ (.Y(_08387_),
    .A(net4779),
    .B(_08386_));
 sg13g2_nand2_1 _34110_ (.Y(_08388_),
    .A(_08378_),
    .B(_08387_));
 sg13g2_a21o_1 _34111_ (.A2(_08092_),
    .A1(_05509_),
    .B1(_05628_),
    .X(_08389_));
 sg13g2_xor2_1 _34112_ (.B(_08389_),
    .A(_05500_),
    .X(_08390_));
 sg13g2_nand2_1 _34113_ (.Y(_08391_),
    .A(_05505_),
    .B(_08102_));
 sg13g2_a21oi_1 _34114_ (.A1(_06021_),
    .A2(_08391_),
    .Y(_08392_),
    .B1(_05500_));
 sg13g2_nand3_1 _34115_ (.B(_06021_),
    .C(_08391_),
    .A(_05500_),
    .Y(_08393_));
 sg13g2_nand2_1 _34116_ (.Y(_08394_),
    .A(net5817),
    .B(_08393_));
 sg13g2_a21oi_1 _34117_ (.A1(net5714),
    .A2(\u_inv.d_next[98] ),
    .Y(_08395_),
    .B1(net5005));
 sg13g2_o21ai_1 _34118_ (.B1(_08395_),
    .Y(_08396_),
    .A1(_08392_),
    .A2(_08394_));
 sg13g2_o21ai_1 _34119_ (.B1(_08396_),
    .Y(_08397_),
    .A1(net5092),
    .A2(_08390_));
 sg13g2_nand2b_1 _34120_ (.Y(_08398_),
    .B(net4784),
    .A_N(_08397_));
 sg13g2_inv_1 _34121_ (.Y(_08399_),
    .A(_08398_));
 sg13g2_nand2_1 _34122_ (.Y(_08400_),
    .A(net4827),
    .B(_08397_));
 sg13g2_xnor2_1 _34123_ (.Y(_08401_),
    .A(net4827),
    .B(_08397_));
 sg13g2_a21oi_1 _34124_ (.A1(_05500_),
    .A2(_08389_),
    .Y(_08402_),
    .B1(_05629_));
 sg13g2_or2_1 _34125_ (.X(_08403_),
    .B(_08402_),
    .A(_05497_));
 sg13g2_a21oi_1 _34126_ (.A1(_05497_),
    .A2(_08402_),
    .Y(_08404_),
    .B1(net5092));
 sg13g2_a21oi_1 _34127_ (.A1(\u_inv.d_next[98] ),
    .A2(net5870),
    .Y(_08405_),
    .B1(_08392_));
 sg13g2_xnor2_1 _34128_ (.Y(_08406_),
    .A(_05498_),
    .B(_08405_));
 sg13g2_a21o_1 _34129_ (.A2(\u_inv.d_next[99] ),
    .A1(net5710),
    .B1(net5005),
    .X(_08407_));
 sg13g2_a21oi_1 _34130_ (.A1(net5813),
    .A2(_08406_),
    .Y(_08408_),
    .B1(_08407_));
 sg13g2_a21o_2 _34131_ (.A2(_08404_),
    .A1(_08403_),
    .B1(_08408_),
    .X(_08409_));
 sg13g2_xnor2_1 _34132_ (.Y(_08410_),
    .A(net4784),
    .B(_08409_));
 sg13g2_nor2b_1 _34133_ (.A(_08401_),
    .B_N(_08410_),
    .Y(_08411_));
 sg13g2_or3_1 _34134_ (.A(_05505_),
    .B(_05506_),
    .C(_08102_),
    .X(_08412_));
 sg13g2_a21oi_1 _34135_ (.A1(_05505_),
    .A2(_05506_),
    .Y(_08413_),
    .B1(net5710));
 sg13g2_nand3_1 _34136_ (.B(_08412_),
    .C(_08413_),
    .A(_08391_),
    .Y(_08414_));
 sg13g2_a21oi_1 _34137_ (.A1(net5710),
    .A2(\u_inv.d_next[97] ),
    .Y(_08415_),
    .B1(net5006));
 sg13g2_nand2_1 _34138_ (.Y(_08416_),
    .A(_05508_),
    .B(_08092_));
 sg13g2_nand3_1 _34139_ (.B(_05627_),
    .C(_08416_),
    .A(_05504_),
    .Y(_08417_));
 sg13g2_a21oi_1 _34140_ (.A1(_05627_),
    .A2(_08416_),
    .Y(_08418_),
    .B1(_05504_));
 sg13g2_nor2_1 _34141_ (.A(net5092),
    .B(_08418_),
    .Y(_08419_));
 sg13g2_a22oi_1 _34142_ (.Y(_08420_),
    .B1(_08417_),
    .B2(_08419_),
    .A2(_08415_),
    .A1(_08414_));
 sg13g2_inv_1 _34143_ (.Y(_08421_),
    .A(_08420_));
 sg13g2_xnor2_1 _34144_ (.Y(_08422_),
    .A(net4823),
    .B(_08420_));
 sg13g2_nand3_1 _34145_ (.B(_06115_),
    .C(_06272_),
    .A(_05508_),
    .Y(_08423_));
 sg13g2_nand2b_1 _34146_ (.Y(_08424_),
    .B(_08423_),
    .A_N(_08102_));
 sg13g2_o21ai_1 _34147_ (.B1(net5092),
    .Y(_08425_),
    .A1(net5813),
    .A2(\u_inv.d_next[96] ));
 sg13g2_a21o_1 _34148_ (.A2(_08424_),
    .A1(net5813),
    .B1(_08425_),
    .X(_08426_));
 sg13g2_xnor2_1 _34149_ (.Y(_08427_),
    .A(_05507_),
    .B(_08091_));
 sg13g2_o21ai_1 _34150_ (.B1(_08426_),
    .Y(_08428_),
    .A1(net5091),
    .A2(_08427_));
 sg13g2_and2_1 _34151_ (.A(net4780),
    .B(_08428_),
    .X(_08429_));
 sg13g2_xnor2_1 _34152_ (.Y(_08430_),
    .A(net4823),
    .B(_08428_));
 sg13g2_and3_1 _34153_ (.X(_08431_),
    .A(_08411_),
    .B(_08422_),
    .C(_08430_));
 sg13g2_inv_1 _34154_ (.Y(_08432_),
    .A(_08431_));
 sg13g2_nor2b_1 _34155_ (.A(_08369_),
    .B_N(_05492_),
    .Y(_08433_));
 sg13g2_xor2_1 _34156_ (.B(_08369_),
    .A(_05492_),
    .X(_08434_));
 sg13g2_o21ai_1 _34157_ (.B1(net5091),
    .Y(_08435_),
    .A1(net5813),
    .A2(\u_inv.d_next[100] ));
 sg13g2_a21o_1 _34158_ (.A2(_08434_),
    .A1(net5813),
    .B1(_08435_),
    .X(_08436_));
 sg13g2_xnor2_1 _34159_ (.Y(_08437_),
    .A(_05492_),
    .B(_08365_));
 sg13g2_o21ai_1 _34160_ (.B1(_08436_),
    .Y(_08438_),
    .A1(net5092),
    .A2(_08437_));
 sg13g2_nand2_1 _34161_ (.Y(_08439_),
    .A(net4780),
    .B(_08438_));
 sg13g2_xnor2_1 _34162_ (.Y(_08440_),
    .A(net4824),
    .B(_08438_));
 sg13g2_o21ai_1 _34163_ (.B1(_05635_),
    .Y(_08441_),
    .A1(_05492_),
    .A2(_08365_));
 sg13g2_o21ai_1 _34164_ (.B1(net5010),
    .Y(_08442_),
    .A1(_05491_),
    .A2(_08441_));
 sg13g2_a21oi_1 _34165_ (.A1(_05491_),
    .A2(_08441_),
    .Y(_08443_),
    .B1(_08442_));
 sg13g2_a21oi_1 _34166_ (.A1(\u_inv.d_next[100] ),
    .A2(\u_inv.d_reg[100] ),
    .Y(_08444_),
    .B1(_08433_));
 sg13g2_xnor2_1 _34167_ (.Y(_08445_),
    .A(_05491_),
    .B(_08444_));
 sg13g2_nand2_1 _34168_ (.Y(_08446_),
    .A(net5710),
    .B(\u_inv.d_next[101] ));
 sg13g2_a21oi_1 _34169_ (.A1(net5812),
    .A2(_08445_),
    .Y(_08447_),
    .B1(net5006));
 sg13g2_a21oi_2 _34170_ (.B1(_08443_),
    .Y(_08448_),
    .A2(_08447_),
    .A1(_08446_));
 sg13g2_nor2_1 _34171_ (.A(net4779),
    .B(_08448_),
    .Y(_08449_));
 sg13g2_xnor2_1 _34172_ (.Y(_08450_),
    .A(net4823),
    .B(_08448_));
 sg13g2_and2_1 _34173_ (.A(_08440_),
    .B(_08450_),
    .X(_08451_));
 sg13g2_and4_1 _34174_ (.A(_08378_),
    .B(_08387_),
    .C(_08431_),
    .D(_08451_),
    .X(_08452_));
 sg13g2_inv_1 _34175_ (.Y(_08453_),
    .A(_08452_));
 sg13g2_nand2_1 _34176_ (.Y(_08454_),
    .A(_08364_),
    .B(_08452_));
 sg13g2_nand4_1 _34177_ (.B(_08274_),
    .C(_08364_),
    .A(_08186_),
    .Y(_08455_),
    .D(_08452_));
 sg13g2_a21o_2 _34178_ (.A2(_08089_),
    .A1(_05684_),
    .B1(_05565_),
    .X(_08456_));
 sg13g2_a21oi_2 _34179_ (.B1(_05536_),
    .Y(_08457_),
    .A2(_08456_),
    .A1(_05614_));
 sg13g2_nor2_1 _34180_ (.A(_05616_),
    .B(_08457_),
    .Y(_08458_));
 sg13g2_a21oi_2 _34181_ (.B1(_05620_),
    .Y(_08459_),
    .A2(_08457_),
    .A1(_05530_));
 sg13g2_o21ai_1 _34182_ (.B1(_05625_),
    .Y(_08460_),
    .A1(_05523_),
    .A2(_08459_));
 sg13g2_a21oi_1 _34183_ (.A1(_05517_),
    .A2(_08460_),
    .Y(_08461_),
    .B1(_05621_));
 sg13g2_or2_1 _34184_ (.X(_08462_),
    .B(_08461_),
    .A(_05515_));
 sg13g2_a21oi_1 _34185_ (.A1(_05515_),
    .A2(_08461_),
    .Y(_08463_),
    .B1(net5094));
 sg13g2_nand2_1 _34186_ (.Y(_08464_),
    .A(_05402_),
    .B(_06268_));
 sg13g2_nand3_1 _34187_ (.B(_05402_),
    .C(_06268_),
    .A(_05400_),
    .Y(_08465_));
 sg13g2_o21ai_1 _34188_ (.B1(_06269_),
    .Y(_08466_),
    .A1(_06265_),
    .A2(_06267_));
 sg13g2_o21ai_1 _34189_ (.B1(_06074_),
    .Y(_08467_),
    .A1(_06062_),
    .A2(_08466_));
 sg13g2_o21ai_1 _34190_ (.B1(_06273_),
    .Y(_08468_),
    .A1(_06265_),
    .A2(_06267_));
 sg13g2_a21oi_1 _34191_ (.A1(_06088_),
    .A2(_08468_),
    .Y(_08469_),
    .B1(_06054_));
 sg13g2_or2_1 _34192_ (.X(_08470_),
    .B(_08469_),
    .A(_06113_));
 sg13g2_a21oi_1 _34193_ (.A1(_06049_),
    .A2(_08470_),
    .Y(_08471_),
    .B1(_06095_));
 sg13g2_nand2b_1 _34194_ (.Y(_08472_),
    .B(_05522_),
    .A_N(_08471_));
 sg13g2_or2_1 _34195_ (.X(_08473_),
    .B(_08471_),
    .A(_06047_));
 sg13g2_a21o_1 _34196_ (.A2(_08473_),
    .A1(_06098_),
    .B1(_05517_),
    .X(_08474_));
 sg13g2_nand2_1 _34197_ (.Y(_08475_),
    .A(_05516_),
    .B(_08474_));
 sg13g2_xnor2_1 _34198_ (.Y(_08476_),
    .A(_05515_),
    .B(_08475_));
 sg13g2_nand2_1 _34199_ (.Y(_08477_),
    .A(net5712),
    .B(\u_inv.d_next[95] ));
 sg13g2_a21oi_1 _34200_ (.A1(net5815),
    .A2(_08476_),
    .Y(_08478_),
    .B1(net5008));
 sg13g2_a22oi_1 _34201_ (.Y(_08479_),
    .B1(_08477_),
    .B2(_08478_),
    .A2(_08463_),
    .A1(_08462_));
 sg13g2_xnor2_1 _34202_ (.Y(_08480_),
    .A(net4782),
    .B(_08479_));
 sg13g2_xor2_1 _34203_ (.B(_08460_),
    .A(_05517_),
    .X(_08481_));
 sg13g2_nand3_1 _34204_ (.B(_06098_),
    .C(_08473_),
    .A(_05517_),
    .Y(_08482_));
 sg13g2_nand3_1 _34205_ (.B(_08474_),
    .C(_08482_),
    .A(net5815),
    .Y(_08483_));
 sg13g2_a21oi_1 _34206_ (.A1(net5712),
    .A2(\u_inv.d_next[94] ),
    .Y(_08484_),
    .B1(net5007));
 sg13g2_nand2_1 _34207_ (.Y(_08485_),
    .A(_08483_),
    .B(_08484_));
 sg13g2_o21ai_1 _34208_ (.B1(_08485_),
    .Y(_08486_),
    .A1(net5094),
    .A2(_08481_));
 sg13g2_nand2b_1 _34209_ (.Y(_08487_),
    .B(net4782),
    .A_N(_08486_));
 sg13g2_xnor2_1 _34210_ (.Y(_08488_),
    .A(net4826),
    .B(_08486_));
 sg13g2_nor2_1 _34211_ (.A(_08480_),
    .B(_08488_),
    .Y(_08489_));
 sg13g2_o21ai_1 _34212_ (.B1(_05623_),
    .Y(_08490_),
    .A1(_05522_),
    .A2(_08459_));
 sg13g2_or2_1 _34213_ (.X(_08491_),
    .B(_08490_),
    .A(_05520_));
 sg13g2_a21oi_1 _34214_ (.A1(_05520_),
    .A2(_08490_),
    .Y(_08492_),
    .B1(net5095));
 sg13g2_nand3_1 _34215_ (.B(_05521_),
    .C(_08472_),
    .A(_05519_),
    .Y(_08493_));
 sg13g2_nand4_1 _34216_ (.B(_06096_),
    .C(_08473_),
    .A(net5815),
    .Y(_08494_),
    .D(_08493_));
 sg13g2_a21oi_1 _34217_ (.A1(net5712),
    .A2(\u_inv.d_next[93] ),
    .Y(_08495_),
    .B1(net5007));
 sg13g2_a22oi_1 _34218_ (.Y(_08496_),
    .B1(_08494_),
    .B2(_08495_),
    .A2(_08492_),
    .A1(_08491_));
 sg13g2_nand2_1 _34219_ (.Y(_08497_),
    .A(net4784),
    .B(_08496_));
 sg13g2_xnor2_1 _34220_ (.Y(_08498_),
    .A(net4827),
    .B(_08496_));
 sg13g2_xor2_1 _34221_ (.B(_08459_),
    .A(_05522_),
    .X(_08499_));
 sg13g2_xor2_1 _34222_ (.B(_08471_),
    .A(_05522_),
    .X(_08500_));
 sg13g2_a21oi_1 _34223_ (.A1(net5715),
    .A2(\u_inv.d_next[92] ),
    .Y(_08501_),
    .B1(net5007));
 sg13g2_o21ai_1 _34224_ (.B1(_08501_),
    .Y(_08502_),
    .A1(net5712),
    .A2(_08500_));
 sg13g2_o21ai_1 _34225_ (.B1(_08502_),
    .Y(_08503_),
    .A1(net5094),
    .A2(_08499_));
 sg13g2_nand2b_1 _34226_ (.Y(_08504_),
    .B(net4784),
    .A_N(_08503_));
 sg13g2_xnor2_1 _34227_ (.Y(_08505_),
    .A(net4828),
    .B(_08503_));
 sg13g2_inv_1 _34228_ (.Y(_08506_),
    .A(_08505_));
 sg13g2_nand2_1 _34229_ (.Y(_08507_),
    .A(_08498_),
    .B(_08506_));
 sg13g2_nand3b_1 _34230_ (.B(_05533_),
    .C(_08470_),
    .Y(_08508_),
    .A_N(_05531_));
 sg13g2_a21o_1 _34231_ (.A2(_08508_),
    .A1(_06092_),
    .B1(_05529_),
    .X(_08509_));
 sg13g2_and2_1 _34232_ (.A(_05528_),
    .B(_08509_),
    .X(_08510_));
 sg13g2_xnor2_1 _34233_ (.Y(_08511_),
    .A(_05526_),
    .B(_08510_));
 sg13g2_a21oi_1 _34234_ (.A1(net5714),
    .A2(\u_inv.d_next[91] ),
    .Y(_08512_),
    .B1(net5009));
 sg13g2_o21ai_1 _34235_ (.B1(_08512_),
    .Y(_08513_),
    .A1(net5714),
    .A2(_08511_));
 sg13g2_o21ai_1 _34236_ (.B1(_05529_),
    .Y(_08514_),
    .A1(_05616_),
    .A2(_08457_));
 sg13g2_nand2b_1 _34237_ (.Y(_08515_),
    .B(_08514_),
    .A_N(_05617_));
 sg13g2_and2_1 _34238_ (.A(_05527_),
    .B(_08515_),
    .X(_08516_));
 sg13g2_o21ai_1 _34239_ (.B1(net5009),
    .Y(_08517_),
    .A1(_05527_),
    .A2(_08515_));
 sg13g2_o21ai_1 _34240_ (.B1(_08513_),
    .Y(_08518_),
    .A1(_08516_),
    .A2(_08517_));
 sg13g2_xnor2_1 _34241_ (.Y(_08519_),
    .A(net4785),
    .B(_08518_));
 sg13g2_xnor2_1 _34242_ (.Y(_08520_),
    .A(_05529_),
    .B(_08458_));
 sg13g2_and3_1 _34243_ (.X(_08521_),
    .A(_05529_),
    .B(_06092_),
    .C(_08508_));
 sg13g2_nand2_1 _34244_ (.Y(_08522_),
    .A(net5817),
    .B(_08509_));
 sg13g2_a21oi_1 _34245_ (.A1(net5714),
    .A2(\u_inv.d_next[90] ),
    .Y(_08523_),
    .B1(net5009));
 sg13g2_o21ai_1 _34246_ (.B1(_08523_),
    .Y(_08524_),
    .A1(_08521_),
    .A2(_08522_));
 sg13g2_o21ai_1 _34247_ (.B1(_08524_),
    .Y(_08525_),
    .A1(net5095),
    .A2(_08520_));
 sg13g2_nor2_1 _34248_ (.A(net4827),
    .B(_08525_),
    .Y(_08526_));
 sg13g2_xnor2_1 _34249_ (.Y(_08527_),
    .A(net4784),
    .B(_08525_));
 sg13g2_a21oi_1 _34250_ (.A1(_05614_),
    .A2(_08456_),
    .Y(_08528_),
    .B1(_05533_));
 sg13g2_a21oi_1 _34251_ (.A1(\u_inv.d_next[88] ),
    .A2(_14721_),
    .Y(_08529_),
    .B1(_08528_));
 sg13g2_and2_1 _34252_ (.A(_05531_),
    .B(_08529_),
    .X(_08530_));
 sg13g2_o21ai_1 _34253_ (.B1(net5009),
    .Y(_08531_),
    .A1(_05531_),
    .A2(_08529_));
 sg13g2_nand2_1 _34254_ (.Y(_08532_),
    .A(_05531_),
    .B(_05532_));
 sg13g2_a21oi_1 _34255_ (.A1(_05533_),
    .A2(_08470_),
    .Y(_08533_),
    .B1(_08532_));
 sg13g2_nand3b_1 _34256_ (.B(_08508_),
    .C(net5817),
    .Y(_08534_),
    .A_N(_06091_));
 sg13g2_a21oi_1 _34257_ (.A1(net5714),
    .A2(\u_inv.d_next[89] ),
    .Y(_08535_),
    .B1(net5010));
 sg13g2_o21ai_1 _34258_ (.B1(_08535_),
    .Y(_08536_),
    .A1(_08533_),
    .A2(_08534_));
 sg13g2_o21ai_1 _34259_ (.B1(_08536_),
    .Y(_08537_),
    .A1(_08530_),
    .A2(_08531_));
 sg13g2_nor2_1 _34260_ (.A(net4827),
    .B(_08537_),
    .Y(_08538_));
 sg13g2_xnor2_1 _34261_ (.Y(_08539_),
    .A(net4784),
    .B(_08537_));
 sg13g2_nand3_1 _34262_ (.B(_05614_),
    .C(_08456_),
    .A(_05533_),
    .Y(_08540_));
 sg13g2_nand2b_1 _34263_ (.Y(_08541_),
    .B(_08540_),
    .A_N(_08528_));
 sg13g2_xnor2_1 _34264_ (.Y(_08542_),
    .A(_05533_),
    .B(_08470_));
 sg13g2_o21ai_1 _34265_ (.B1(net5095),
    .Y(_08543_),
    .A1(net5815),
    .A2(\u_inv.d_next[88] ));
 sg13g2_a21o_1 _34266_ (.A2(_08542_),
    .A1(net5816),
    .B1(_08543_),
    .X(_08544_));
 sg13g2_o21ai_1 _34267_ (.B1(_08544_),
    .Y(_08545_),
    .A1(net5094),
    .A2(_08541_));
 sg13g2_nand2_1 _34268_ (.Y(_08546_),
    .A(net4785),
    .B(_08545_));
 sg13g2_xnor2_1 _34269_ (.Y(_08547_),
    .A(net4827),
    .B(_08545_));
 sg13g2_and4_1 _34270_ (.A(_08519_),
    .B(_08527_),
    .C(_08539_),
    .D(_08547_),
    .X(_08548_));
 sg13g2_nand4_1 _34271_ (.B(_08527_),
    .C(_08539_),
    .A(_08519_),
    .Y(_08549_),
    .D(_08547_));
 sg13g2_nor4_1 _34272_ (.A(_08480_),
    .B(_08488_),
    .C(_08507_),
    .D(_08549_),
    .Y(_08550_));
 sg13g2_nor2_1 _34273_ (.A(_05561_),
    .B(_08090_),
    .Y(_08551_));
 sg13g2_a21oi_1 _34274_ (.A1(_05684_),
    .A2(_08089_),
    .Y(_08552_),
    .B1(_05563_));
 sg13g2_a21oi_1 _34275_ (.A1(_05684_),
    .A2(_08089_),
    .Y(_08553_),
    .B1(_05564_));
 sg13g2_nand2b_1 _34276_ (.Y(_08554_),
    .B(_05604_),
    .A_N(_08553_));
 sg13g2_o21ai_1 _34277_ (.B1(_05549_),
    .Y(_08555_),
    .A1(_05605_),
    .A2(_08553_));
 sg13g2_and3_1 _34278_ (.X(_08556_),
    .A(_05543_),
    .B(_05611_),
    .C(_08555_));
 sg13g2_a21oi_1 _34279_ (.A1(_05611_),
    .A2(_08555_),
    .Y(_08557_),
    .B1(_05543_));
 sg13g2_or2_1 _34280_ (.X(_08558_),
    .B(_08557_),
    .A(_08556_));
 sg13g2_a21oi_1 _34281_ (.A1(_06088_),
    .A2(_08468_),
    .Y(_08559_),
    .B1(_05562_));
 sg13g2_a221oi_1 _34282_ (.B2(_08468_),
    .C1(_05562_),
    .B1(_06088_),
    .A1(_05557_),
    .Y(_08560_),
    .A2(_05558_));
 sg13g2_nand2_1 _34283_ (.Y(_08561_),
    .A(net5616),
    .B(_08559_));
 sg13g2_a21oi_2 _34284_ (.B1(_06108_),
    .Y(_08562_),
    .A2(_08560_),
    .A1(_06053_));
 sg13g2_nor2_1 _34285_ (.A(_06051_),
    .B(_08562_),
    .Y(_08563_));
 sg13g2_nor3_1 _34286_ (.A(_05543_),
    .B(_06110_),
    .C(_08563_),
    .Y(_08564_));
 sg13g2_o21ai_1 _34287_ (.B1(_05543_),
    .Y(_08565_),
    .A1(_06110_),
    .A2(_08563_));
 sg13g2_nor2b_1 _34288_ (.A(_08564_),
    .B_N(_08565_),
    .Y(_08566_));
 sg13g2_nand2_1 _34289_ (.Y(_08567_),
    .A(net5712),
    .B(\u_inv.d_next[86] ));
 sg13g2_a21oi_1 _34290_ (.A1(net5816),
    .A2(_08566_),
    .Y(_08568_),
    .B1(net5008));
 sg13g2_a22oi_1 _34291_ (.Y(_08569_),
    .B1(_08567_),
    .B2(_08568_),
    .A2(_08558_),
    .A1(net5008));
 sg13g2_and2_1 _34292_ (.A(net4782),
    .B(_08569_),
    .X(_08570_));
 sg13g2_nand2b_1 _34293_ (.Y(_08571_),
    .B(net4828),
    .A_N(_08569_));
 sg13g2_nand2b_1 _34294_ (.Y(_08572_),
    .B(_08571_),
    .A_N(_08570_));
 sg13g2_nor2b_1 _34295_ (.A(_05542_),
    .B_N(_08565_),
    .Y(_08573_));
 sg13g2_xnor2_1 _34296_ (.Y(_08574_),
    .A(_05541_),
    .B(_08573_));
 sg13g2_nand2_1 _34297_ (.Y(_08575_),
    .A(net5713),
    .B(\u_inv.d_next[87] ));
 sg13g2_a21oi_1 _34298_ (.A1(net5816),
    .A2(_08574_),
    .Y(_08576_),
    .B1(net5008));
 sg13g2_o21ai_1 _34299_ (.B1(_05541_),
    .Y(_08577_),
    .A1(_05606_),
    .A2(_08557_));
 sg13g2_nor3_1 _34300_ (.A(_05541_),
    .B(_05606_),
    .C(_08557_),
    .Y(_08578_));
 sg13g2_nor2_1 _34301_ (.A(net5094),
    .B(_08578_),
    .Y(_08579_));
 sg13g2_a22oi_1 _34302_ (.Y(_08580_),
    .B1(_08577_),
    .B2(_08579_),
    .A2(_08576_),
    .A1(_08575_));
 sg13g2_xnor2_1 _34303_ (.Y(_08581_),
    .A(net4782),
    .B(_08580_));
 sg13g2_nor2_1 _34304_ (.A(_08572_),
    .B(_08581_),
    .Y(_08582_));
 sg13g2_or2_1 _34305_ (.X(_08583_),
    .B(_08581_),
    .A(_08572_));
 sg13g2_nor2_1 _34306_ (.A(_05548_),
    .B(_08562_),
    .Y(_08584_));
 sg13g2_a21oi_1 _34307_ (.A1(\u_inv.d_next[84] ),
    .A2(\u_inv.d_reg[84] ),
    .Y(_08585_),
    .B1(_08584_));
 sg13g2_xnor2_1 _34308_ (.Y(_08586_),
    .A(_05546_),
    .B(_08585_));
 sg13g2_nand2_1 _34309_ (.Y(_08587_),
    .A(net5816),
    .B(_08586_));
 sg13g2_a21oi_1 _34310_ (.A1(net5713),
    .A2(\u_inv.d_next[85] ),
    .Y(_08588_),
    .B1(net5008));
 sg13g2_a21o_1 _34311_ (.A2(_08554_),
    .A1(_05548_),
    .B1(_05609_),
    .X(_08589_));
 sg13g2_o21ai_1 _34312_ (.B1(net5009),
    .Y(_08590_),
    .A1(_05546_),
    .A2(_08589_));
 sg13g2_a21oi_1 _34313_ (.A1(_05546_),
    .A2(_08589_),
    .Y(_08591_),
    .B1(_08590_));
 sg13g2_a21oi_2 _34314_ (.B1(_08591_),
    .Y(_08592_),
    .A2(_08588_),
    .A1(_08587_));
 sg13g2_inv_1 _34315_ (.Y(_08593_),
    .A(_08592_));
 sg13g2_xnor2_1 _34316_ (.Y(_08594_),
    .A(net4828),
    .B(_08592_));
 sg13g2_xnor2_1 _34317_ (.Y(_08595_),
    .A(_05548_),
    .B(_08554_));
 sg13g2_a21oi_1 _34318_ (.A1(_05548_),
    .A2(_08562_),
    .Y(_08596_),
    .B1(net5713));
 sg13g2_nand2b_1 _34319_ (.Y(_08597_),
    .B(_08596_),
    .A_N(_08584_));
 sg13g2_a21oi_1 _34320_ (.A1(net5713),
    .A2(\u_inv.d_next[84] ),
    .Y(_08598_),
    .B1(net5008));
 sg13g2_a22oi_1 _34321_ (.Y(_08599_),
    .B1(_08597_),
    .B2(_08598_),
    .A2(_08595_),
    .A1(net5008));
 sg13g2_nand2_1 _34322_ (.Y(_08600_),
    .A(net4783),
    .B(_08599_));
 sg13g2_xnor2_1 _34323_ (.Y(_08601_),
    .A(net4826),
    .B(_08599_));
 sg13g2_nand2_1 _34324_ (.Y(_08602_),
    .A(_08594_),
    .B(_08601_));
 sg13g2_xnor2_1 _34325_ (.Y(_08603_),
    .A(_05562_),
    .B(_08090_));
 sg13g2_nand3_1 _34326_ (.B(_06088_),
    .C(_08468_),
    .A(_05562_),
    .Y(_08604_));
 sg13g2_nand2b_1 _34327_ (.Y(_08605_),
    .B(_08604_),
    .A_N(_08559_));
 sg13g2_o21ai_1 _34328_ (.B1(net5094),
    .Y(_08606_),
    .A1(net5815),
    .A2(\u_inv.d_next[80] ));
 sg13g2_a21oi_1 _34329_ (.A1(net5815),
    .A2(_08605_),
    .Y(_08607_),
    .B1(_08606_));
 sg13g2_a21o_1 _34330_ (.A2(_08603_),
    .A1(net5007),
    .B1(_08607_),
    .X(_08608_));
 sg13g2_and2_1 _34331_ (.A(net4782),
    .B(_08608_),
    .X(_08609_));
 sg13g2_xnor2_1 _34332_ (.Y(_08610_),
    .A(net4782),
    .B(_08608_));
 sg13g2_nor2_1 _34333_ (.A(_05601_),
    .B(_08552_),
    .Y(_08611_));
 sg13g2_o21ai_1 _34334_ (.B1(_05554_),
    .Y(_08612_),
    .A1(_05601_),
    .A2(_08552_));
 sg13g2_xnor2_1 _34335_ (.Y(_08613_),
    .A(_05554_),
    .B(_08611_));
 sg13g2_nand3_1 _34336_ (.B(_06105_),
    .C(_08561_),
    .A(_05554_),
    .Y(_08614_));
 sg13g2_a21o_1 _34337_ (.A2(_08561_),
    .A1(_06105_),
    .B1(_05554_),
    .X(_08615_));
 sg13g2_nand3_1 _34338_ (.B(_08614_),
    .C(_08615_),
    .A(net5815),
    .Y(_08616_));
 sg13g2_a21oi_1 _34339_ (.A1(net5712),
    .A2(\u_inv.d_next[82] ),
    .Y(_08617_),
    .B1(net5007));
 sg13g2_nand2_1 _34340_ (.Y(_08618_),
    .A(_08616_),
    .B(_08617_));
 sg13g2_o21ai_1 _34341_ (.B1(_08618_),
    .Y(_08619_),
    .A1(net5094),
    .A2(_08613_));
 sg13g2_nor2_1 _34342_ (.A(net4826),
    .B(_08619_),
    .Y(_08620_));
 sg13g2_xnor2_1 _34343_ (.Y(_08621_),
    .A(net4826),
    .B(_08619_));
 sg13g2_nand3_1 _34344_ (.B(_05553_),
    .C(_08615_),
    .A(_05551_),
    .Y(_08622_));
 sg13g2_a21o_1 _34345_ (.A2(_08615_),
    .A1(_05553_),
    .B1(_05551_),
    .X(_08623_));
 sg13g2_nand3_1 _34346_ (.B(_08622_),
    .C(_08623_),
    .A(net5816),
    .Y(_08624_));
 sg13g2_nand2_1 _34347_ (.Y(_08625_),
    .A(net5712),
    .B(\u_inv.d_next[83] ));
 sg13g2_nand3_1 _34348_ (.B(_08624_),
    .C(_08625_),
    .A(net5094),
    .Y(_08626_));
 sg13g2_nand3_1 _34349_ (.B(_05602_),
    .C(_08612_),
    .A(_05551_),
    .Y(_08627_));
 sg13g2_a21oi_1 _34350_ (.A1(_05602_),
    .A2(_08612_),
    .Y(_08628_),
    .B1(_05551_));
 sg13g2_nand2_1 _34351_ (.Y(_08629_),
    .A(net5007),
    .B(_08627_));
 sg13g2_o21ai_1 _34352_ (.B1(_08626_),
    .Y(_08630_),
    .A1(_08628_),
    .A2(_08629_));
 sg13g2_xnor2_1 _34353_ (.Y(_08631_),
    .A(net4782),
    .B(_08630_));
 sg13g2_nand2b_1 _34354_ (.Y(_08632_),
    .B(_08631_),
    .A_N(_08621_));
 sg13g2_o21ai_1 _34355_ (.B1(net5616),
    .Y(_08633_),
    .A1(_05599_),
    .A2(_08551_));
 sg13g2_or3_1 _34356_ (.A(net5616),
    .B(_05599_),
    .C(_08551_),
    .X(_08634_));
 sg13g2_and3_1 _34357_ (.X(_08635_),
    .A(net5007),
    .B(_08633_),
    .C(_08634_));
 sg13g2_or3_1 _34358_ (.A(net5616),
    .B(_05560_),
    .C(_08559_),
    .X(_08636_));
 sg13g2_nand4_1 _34359_ (.B(_06103_),
    .C(_08561_),
    .A(net5815),
    .Y(_08637_),
    .D(_08636_));
 sg13g2_a21oi_1 _34360_ (.A1(net5712),
    .A2(\u_inv.d_next[81] ),
    .Y(_08638_),
    .B1(net5007));
 sg13g2_a21oi_1 _34361_ (.A1(_08637_),
    .A2(_08638_),
    .Y(_08639_),
    .B1(_08635_));
 sg13g2_a21o_1 _34362_ (.A2(_08638_),
    .A1(_08637_),
    .B1(_08635_),
    .X(_08640_));
 sg13g2_xnor2_1 _34363_ (.Y(_08641_),
    .A(net4826),
    .B(_08639_));
 sg13g2_nand2b_1 _34364_ (.Y(_08642_),
    .B(_08641_),
    .A_N(_08632_));
 sg13g2_or2_1 _34365_ (.X(_08643_),
    .B(_08642_),
    .A(_08610_));
 sg13g2_nor4_1 _34366_ (.A(_08583_),
    .B(_08602_),
    .C(_08610_),
    .D(_08642_),
    .Y(_08644_));
 sg13g2_inv_1 _34367_ (.Y(_08645_),
    .A(_08644_));
 sg13g2_and2_1 _34368_ (.A(_08550_),
    .B(_08644_),
    .X(_08646_));
 sg13g2_and2_1 _34369_ (.A(_05668_),
    .B(_08088_),
    .X(_08647_));
 sg13g2_a21o_2 _34370_ (.A2(_08088_),
    .A1(_05668_),
    .B1(_05374_),
    .X(_08648_));
 sg13g2_a21oi_1 _34371_ (.A1(_05677_),
    .A2(_08648_),
    .Y(_08649_),
    .B1(_05366_));
 sg13g2_a21oi_1 _34372_ (.A1(net5877),
    .A2(_14735_),
    .Y(_08650_),
    .B1(_08649_));
 sg13g2_a21o_1 _34373_ (.A2(_08648_),
    .A1(_05677_),
    .B1(_05368_),
    .X(_08651_));
 sg13g2_a21o_1 _34374_ (.A2(_08651_),
    .A1(_05680_),
    .B1(_05360_),
    .X(_08652_));
 sg13g2_nand2_1 _34375_ (.Y(_08653_),
    .A(_05671_),
    .B(_08652_));
 sg13g2_a21oi_1 _34376_ (.A1(_05671_),
    .A2(_08652_),
    .Y(_08654_),
    .B1(_05353_));
 sg13g2_xnor2_1 _34377_ (.Y(_08655_),
    .A(_05353_),
    .B(_08653_));
 sg13g2_nand2_1 _34378_ (.Y(_08656_),
    .A(_06058_),
    .B(_08467_));
 sg13g2_nand4_1 _34379_ (.B(_05366_),
    .C(_06058_),
    .A(_05365_),
    .Y(_08657_),
    .D(_08467_));
 sg13g2_nand2b_2 _34380_ (.Y(_08658_),
    .B(_08657_),
    .A_N(_06087_));
 sg13g2_nand3_1 _34381_ (.B(_05358_),
    .C(_08658_),
    .A(_05355_),
    .Y(_08659_));
 sg13g2_nand3_1 _34382_ (.B(_06078_),
    .C(_08659_),
    .A(_05352_),
    .Y(_08660_));
 sg13g2_a21o_1 _34383_ (.A2(_08659_),
    .A1(_06078_),
    .B1(_05352_),
    .X(_08661_));
 sg13g2_nand3_1 _34384_ (.B(_08660_),
    .C(_08661_),
    .A(net5814),
    .Y(_08662_));
 sg13g2_a21oi_1 _34385_ (.A1(net5711),
    .A2(\u_inv.d_next[78] ),
    .Y(_08663_),
    .B1(net5006));
 sg13g2_nand2_1 _34386_ (.Y(_08664_),
    .A(_08662_),
    .B(_08663_));
 sg13g2_o21ai_1 _34387_ (.B1(_08664_),
    .Y(_08665_),
    .A1(net5093),
    .A2(_08655_));
 sg13g2_nor2_1 _34388_ (.A(net4825),
    .B(_08665_),
    .Y(_08666_));
 sg13g2_nand2_1 _34389_ (.Y(_08667_),
    .A(net4825),
    .B(_08665_));
 sg13g2_xnor2_1 _34390_ (.Y(_08668_),
    .A(net4825),
    .B(_08665_));
 sg13g2_o21ai_1 _34391_ (.B1(_05350_),
    .Y(_08669_),
    .A1(_05672_),
    .A2(_08654_));
 sg13g2_or3_1 _34392_ (.A(_05350_),
    .B(_05672_),
    .C(_08654_),
    .X(_08670_));
 sg13g2_nand3_1 _34393_ (.B(_08669_),
    .C(_08670_),
    .A(net5006),
    .Y(_08671_));
 sg13g2_a21o_1 _34394_ (.A2(_08661_),
    .A1(_05351_),
    .B1(_05349_),
    .X(_08672_));
 sg13g2_nand3_1 _34395_ (.B(_05351_),
    .C(_08661_),
    .A(_05349_),
    .Y(_08673_));
 sg13g2_nand3_1 _34396_ (.B(_08672_),
    .C(_08673_),
    .A(net5814),
    .Y(_08674_));
 sg13g2_nand2_1 _34397_ (.Y(_08675_),
    .A(net5711),
    .B(\u_inv.d_next[79] ));
 sg13g2_nand3_1 _34398_ (.B(_08674_),
    .C(_08675_),
    .A(net5093),
    .Y(_08676_));
 sg13g2_and3_1 _34399_ (.X(_08677_),
    .A(net4778),
    .B(_08671_),
    .C(_08676_));
 sg13g2_a21oi_1 _34400_ (.A1(_08671_),
    .A2(_08676_),
    .Y(_08678_),
    .B1(net4778));
 sg13g2_nor2_1 _34401_ (.A(_08677_),
    .B(_08678_),
    .Y(_08679_));
 sg13g2_nor3_1 _34402_ (.A(_08668_),
    .B(_08677_),
    .C(_08678_),
    .Y(_08680_));
 sg13g2_a21oi_1 _34403_ (.A1(_05680_),
    .A2(_08651_),
    .Y(_08681_),
    .B1(_05358_));
 sg13g2_o21ai_1 _34404_ (.B1(_05355_),
    .Y(_08682_),
    .A1(_05670_),
    .A2(_08681_));
 sg13g2_nor3_1 _34405_ (.A(_05355_),
    .B(_05670_),
    .C(_08681_),
    .Y(_08683_));
 sg13g2_nand2_1 _34406_ (.Y(_08684_),
    .A(net5006),
    .B(_08682_));
 sg13g2_a21oi_1 _34407_ (.A1(_05358_),
    .A2(_08658_),
    .Y(_08685_),
    .B1(_05357_));
 sg13g2_xnor2_1 _34408_ (.Y(_08686_),
    .A(_05356_),
    .B(_08685_));
 sg13g2_a21oi_1 _34409_ (.A1(net5711),
    .A2(\u_inv.d_next[77] ),
    .Y(_08687_),
    .B1(net5006));
 sg13g2_o21ai_1 _34410_ (.B1(_08687_),
    .Y(_08688_),
    .A1(net5711),
    .A2(_08686_));
 sg13g2_o21ai_1 _34411_ (.B1(_08688_),
    .Y(_08689_),
    .A1(_08683_),
    .A2(_08684_));
 sg13g2_nor2_1 _34412_ (.A(net4825),
    .B(_08689_),
    .Y(_08690_));
 sg13g2_xnor2_1 _34413_ (.Y(_08691_),
    .A(net4778),
    .B(_08689_));
 sg13g2_xnor2_1 _34414_ (.Y(_08692_),
    .A(_05358_),
    .B(_08658_));
 sg13g2_o21ai_1 _34415_ (.B1(net5093),
    .Y(_08693_),
    .A1(net5814),
    .A2(\u_inv.d_next[76] ));
 sg13g2_a21oi_1 _34416_ (.A1(net5814),
    .A2(_08692_),
    .Y(_08694_),
    .B1(_08693_));
 sg13g2_and3_1 _34417_ (.X(_08695_),
    .A(_05358_),
    .B(_05680_),
    .C(_08651_));
 sg13g2_nor2_1 _34418_ (.A(_08681_),
    .B(_08695_),
    .Y(_08696_));
 sg13g2_a21o_2 _34419_ (.A2(_08696_),
    .A1(net5006),
    .B1(_08694_),
    .X(_08697_));
 sg13g2_nand2_1 _34420_ (.Y(_08698_),
    .A(net4778),
    .B(_08697_));
 sg13g2_xnor2_1 _34421_ (.Y(_08699_),
    .A(net4825),
    .B(_08697_));
 sg13g2_nand3_1 _34422_ (.B(_05677_),
    .C(_08648_),
    .A(_05366_),
    .Y(_08700_));
 sg13g2_nand2b_1 _34423_ (.Y(_08701_),
    .B(_08700_),
    .A_N(_08649_));
 sg13g2_nand3_1 _34424_ (.B(_06084_),
    .C(_08656_),
    .A(_05367_),
    .Y(_08702_));
 sg13g2_a21o_1 _34425_ (.A2(_08656_),
    .A1(_06084_),
    .B1(_05367_),
    .X(_08703_));
 sg13g2_nand3_1 _34426_ (.B(_08702_),
    .C(_08703_),
    .A(net5802),
    .Y(_08704_));
 sg13g2_a21oi_1 _34427_ (.A1(net5711),
    .A2(net5877),
    .Y(_08705_),
    .B1(net4996));
 sg13g2_a22oi_1 _34428_ (.Y(_08706_),
    .B1(_08704_),
    .B2(_08705_),
    .A2(_08701_),
    .A1(net4996));
 sg13g2_and2_1 _34429_ (.A(net4777),
    .B(_08706_),
    .X(_08707_));
 sg13g2_xnor2_1 _34430_ (.Y(_08708_),
    .A(net4777),
    .B(_08706_));
 sg13g2_o21ai_1 _34431_ (.B1(_08703_),
    .Y(_08709_),
    .A1(_14224_),
    .A2(_14735_));
 sg13g2_xnor2_1 _34432_ (.Y(_08710_),
    .A(_05364_),
    .B(_08709_));
 sg13g2_nand2_1 _34433_ (.Y(_08711_),
    .A(net5814),
    .B(_08710_));
 sg13g2_a21oi_1 _34434_ (.A1(net5711),
    .A2(\u_inv.d_next[75] ),
    .Y(_08712_),
    .B1(net4998));
 sg13g2_xnor2_1 _34435_ (.Y(_08713_),
    .A(_05365_),
    .B(_08650_));
 sg13g2_a22oi_1 _34436_ (.Y(_08714_),
    .B1(_08713_),
    .B2(net4998),
    .A2(_08712_),
    .A1(_08711_));
 sg13g2_xnor2_1 _34437_ (.Y(_08715_),
    .A(net4825),
    .B(_08714_));
 sg13g2_nand2b_1 _34438_ (.Y(_08716_),
    .B(_08715_),
    .A_N(_08708_));
 sg13g2_xnor2_1 _34439_ (.Y(_08717_),
    .A(_05372_),
    .B(_08467_));
 sg13g2_o21ai_1 _34440_ (.B1(net5083),
    .Y(_08718_),
    .A1(net5802),
    .A2(net5878));
 sg13g2_a21o_1 _34441_ (.A2(_08717_),
    .A1(net5802),
    .B1(_08718_),
    .X(_08719_));
 sg13g2_xnor2_1 _34442_ (.Y(_08720_),
    .A(_05372_),
    .B(_08647_));
 sg13g2_o21ai_1 _34443_ (.B1(_08719_),
    .Y(_08721_),
    .A1(net5083),
    .A2(_08720_));
 sg13g2_nand2_1 _34444_ (.Y(_08722_),
    .A(net4777),
    .B(_08721_));
 sg13g2_xnor2_1 _34445_ (.Y(_08723_),
    .A(net4777),
    .B(_08721_));
 sg13g2_a21oi_1 _34446_ (.A1(\u_inv.d_next[72] ),
    .A2(_14737_),
    .Y(_08724_),
    .B1(_05370_));
 sg13g2_o21ai_1 _34447_ (.B1(_08724_),
    .Y(_08725_),
    .A1(_05372_),
    .A2(_08647_));
 sg13g2_nand3b_1 _34448_ (.B(_08648_),
    .C(_08725_),
    .Y(_08726_),
    .A_N(_05676_));
 sg13g2_a21oi_1 _34449_ (.A1(_05372_),
    .A2(_08467_),
    .Y(_08727_),
    .B1(_05371_));
 sg13g2_xnor2_1 _34450_ (.Y(_08728_),
    .A(_05370_),
    .B(_08727_));
 sg13g2_or2_1 _34451_ (.X(_08729_),
    .B(_08728_),
    .A(net5703));
 sg13g2_a21oi_1 _34452_ (.A1(net5703),
    .A2(\u_inv.d_next[73] ),
    .Y(_08730_),
    .B1(net4998));
 sg13g2_a22oi_1 _34453_ (.Y(_08731_),
    .B1(_08729_),
    .B2(_08730_),
    .A2(_08726_),
    .A1(net4996));
 sg13g2_inv_1 _34454_ (.Y(_08732_),
    .A(_08731_));
 sg13g2_xnor2_1 _34455_ (.Y(_08733_),
    .A(net4777),
    .B(_08731_));
 sg13g2_nor3_1 _34456_ (.A(_08716_),
    .B(_08723_),
    .C(_08733_),
    .Y(_08734_));
 sg13g2_inv_1 _34457_ (.Y(_08735_),
    .A(_08734_));
 sg13g2_nand4_1 _34458_ (.B(_08691_),
    .C(_08699_),
    .A(_08680_),
    .Y(_08736_),
    .D(_08734_));
 sg13g2_o21ai_1 _34459_ (.B1(_05404_),
    .Y(_08737_),
    .A1(_05314_),
    .A2(_05347_));
 sg13g2_and2_1 _34460_ (.A(_05656_),
    .B(_08737_),
    .X(_08738_));
 sg13g2_a21oi_1 _34461_ (.A1(_05656_),
    .A2(_08737_),
    .Y(_08739_),
    .B1(_05397_));
 sg13g2_or2_1 _34462_ (.X(_08740_),
    .B(_08739_),
    .A(_05659_));
 sg13g2_o21ai_1 _34463_ (.B1(_05389_),
    .Y(_08741_),
    .A1(_05659_),
    .A2(_08739_));
 sg13g2_nand2_1 _34464_ (.Y(_08742_),
    .A(_05663_),
    .B(_08741_));
 sg13g2_a21oi_1 _34465_ (.A1(_05663_),
    .A2(_08741_),
    .Y(_08743_),
    .B1(_05380_));
 sg13g2_xnor2_1 _34466_ (.Y(_08744_),
    .A(_05380_),
    .B(_08742_));
 sg13g2_nand2b_2 _34467_ (.Y(_08745_),
    .B(_08466_),
    .A_N(_06069_));
 sg13g2_a221oi_1 _34468_ (.B2(_08745_),
    .C1(_05383_),
    .B1(_06060_),
    .A1(_05382_),
    .Y(_08746_),
    .A2(_05386_));
 sg13g2_xor2_1 _34469_ (.B(_08746_),
    .A(_05380_),
    .X(_08747_));
 sg13g2_a21oi_1 _34470_ (.A1(net5703),
    .A2(net5879),
    .Y(_08748_),
    .B1(net4996));
 sg13g2_o21ai_1 _34471_ (.B1(_08748_),
    .Y(_08749_),
    .A1(net5703),
    .A2(_08747_));
 sg13g2_o21ai_1 _34472_ (.B1(_08749_),
    .Y(_08750_),
    .A1(net5083),
    .A2(_08744_));
 sg13g2_nand2b_1 _34473_ (.Y(_08751_),
    .B(net4776),
    .A_N(_08750_));
 sg13g2_xnor2_1 _34474_ (.Y(_08752_),
    .A(net4821),
    .B(_08750_));
 sg13g2_inv_1 _34475_ (.Y(_08753_),
    .A(_08752_));
 sg13g2_o21ai_1 _34476_ (.B1(_05377_),
    .Y(_08754_),
    .A1(_05665_),
    .A2(_08743_));
 sg13g2_nor3_1 _34477_ (.A(_05377_),
    .B(_05665_),
    .C(_08743_),
    .Y(_08755_));
 sg13g2_nand2_1 _34478_ (.Y(_08756_),
    .A(net4996),
    .B(_08754_));
 sg13g2_o21ai_1 _34479_ (.B1(_05378_),
    .Y(_08757_),
    .A1(_05379_),
    .A2(_08746_));
 sg13g2_xnor2_1 _34480_ (.Y(_08758_),
    .A(_05377_),
    .B(_08757_));
 sg13g2_a21oi_1 _34481_ (.A1(net5703),
    .A2(\u_inv.d_next[71] ),
    .Y(_08759_),
    .B1(net4996));
 sg13g2_o21ai_1 _34482_ (.B1(_08759_),
    .Y(_08760_),
    .A1(net5703),
    .A2(_08758_));
 sg13g2_o21ai_1 _34483_ (.B1(_08760_),
    .Y(_08761_),
    .A1(_08755_),
    .A2(_08756_));
 sg13g2_xnor2_1 _34484_ (.Y(_08762_),
    .A(net4776),
    .B(_08761_));
 sg13g2_and2_1 _34485_ (.A(_08753_),
    .B(_08762_),
    .X(_08763_));
 sg13g2_nand2_1 _34486_ (.Y(_08764_),
    .A(_05388_),
    .B(_08740_));
 sg13g2_a21oi_1 _34487_ (.A1(_05661_),
    .A2(_08764_),
    .Y(_08765_),
    .B1(_05385_));
 sg13g2_nand3_1 _34488_ (.B(_05661_),
    .C(_08764_),
    .A(_05385_),
    .Y(_08766_));
 sg13g2_nand2_1 _34489_ (.Y(_08767_),
    .A(net4996),
    .B(_08766_));
 sg13g2_a21oi_1 _34490_ (.A1(_05387_),
    .A2(_08745_),
    .Y(_08768_),
    .B1(_05386_));
 sg13g2_xnor2_1 _34491_ (.Y(_08769_),
    .A(_05385_),
    .B(_08768_));
 sg13g2_a21oi_1 _34492_ (.A1(net5703),
    .A2(\u_inv.d_next[69] ),
    .Y(_08770_),
    .B1(net4996));
 sg13g2_o21ai_1 _34493_ (.B1(_08770_),
    .Y(_08771_),
    .A1(net5703),
    .A2(_08769_));
 sg13g2_o21ai_1 _34494_ (.B1(_08771_),
    .Y(_08772_),
    .A1(_08765_),
    .A2(_08767_));
 sg13g2_nand2_1 _34495_ (.Y(_08773_),
    .A(net4821),
    .B(_08772_));
 sg13g2_xnor2_1 _34496_ (.Y(_08774_),
    .A(net4776),
    .B(_08772_));
 sg13g2_xnor2_1 _34497_ (.Y(_08775_),
    .A(_05387_),
    .B(_08745_));
 sg13g2_o21ai_1 _34498_ (.B1(net5083),
    .Y(_08776_),
    .A1(net5802),
    .A2(\u_inv.d_next[68] ));
 sg13g2_a21o_1 _34499_ (.A2(_08775_),
    .A1(net5802),
    .B1(_08776_),
    .X(_08777_));
 sg13g2_xnor2_1 _34500_ (.Y(_08778_),
    .A(_05388_),
    .B(_08740_));
 sg13g2_o21ai_1 _34501_ (.B1(_08777_),
    .Y(_08779_),
    .A1(net5083),
    .A2(_08778_));
 sg13g2_and2_1 _34502_ (.A(net4776),
    .B(_08779_),
    .X(_08780_));
 sg13g2_inv_1 _34503_ (.Y(_08781_),
    .A(_08780_));
 sg13g2_xnor2_1 _34504_ (.Y(_08782_),
    .A(net4821),
    .B(_08779_));
 sg13g2_and4_1 _34505_ (.A(_08753_),
    .B(_08762_),
    .C(_08774_),
    .D(_08782_),
    .X(_08783_));
 sg13g2_xnor2_1 _34506_ (.Y(_08784_),
    .A(_05396_),
    .B(_08738_));
 sg13g2_a21o_1 _34507_ (.A2(_08465_),
    .A1(_06066_),
    .B1(_05396_),
    .X(_08785_));
 sg13g2_nand3_1 _34508_ (.B(_06066_),
    .C(_08465_),
    .A(_05396_),
    .Y(_08786_));
 sg13g2_nand3_1 _34509_ (.B(_08785_),
    .C(_08786_),
    .A(net5801),
    .Y(_08787_));
 sg13g2_a21oi_1 _34510_ (.A1(net5701),
    .A2(net5880),
    .Y(_08788_),
    .B1(net4995));
 sg13g2_nand2_1 _34511_ (.Y(_08789_),
    .A(_08787_),
    .B(_08788_));
 sg13g2_o21ai_1 _34512_ (.B1(_08789_),
    .Y(_08790_),
    .A1(net5081),
    .A2(_08784_));
 sg13g2_nor2_1 _34513_ (.A(net4821),
    .B(_08790_),
    .Y(_08791_));
 sg13g2_xnor2_1 _34514_ (.Y(_08792_),
    .A(net4776),
    .B(_08790_));
 sg13g2_o21ai_1 _34515_ (.B1(_05658_),
    .Y(_08793_),
    .A1(_05395_),
    .A2(_08738_));
 sg13g2_o21ai_1 _34516_ (.B1(net4995),
    .Y(_08794_),
    .A1(_05394_),
    .A2(_08793_));
 sg13g2_a21oi_1 _34517_ (.A1(_05394_),
    .A2(_08793_),
    .Y(_08795_),
    .B1(_08794_));
 sg13g2_o21ai_1 _34518_ (.B1(_08785_),
    .Y(_08796_),
    .A1(_14225_),
    .A2(_14743_));
 sg13g2_xnor2_1 _34519_ (.Y(_08797_),
    .A(_05393_),
    .B(_08796_));
 sg13g2_nand2_1 _34520_ (.Y(_08798_),
    .A(net5701),
    .B(\u_inv.d_next[67] ));
 sg13g2_a21oi_1 _34521_ (.A1(net5801),
    .A2(_08797_),
    .Y(_08799_),
    .B1(net4995));
 sg13g2_a21o_1 _34522_ (.A2(_08799_),
    .A1(_08798_),
    .B1(_08795_),
    .X(_08800_));
 sg13g2_xnor2_1 _34523_ (.Y(_08801_),
    .A(net4776),
    .B(_08800_));
 sg13g2_nand2_1 _34524_ (.Y(_08802_),
    .A(_08792_),
    .B(_08801_));
 sg13g2_nor2_1 _34525_ (.A(_05400_),
    .B(_05401_),
    .Y(_08803_));
 sg13g2_nand3b_1 _34526_ (.B(_08465_),
    .C(net5801),
    .Y(_08804_),
    .A_N(_06064_));
 sg13g2_a21oi_1 _34527_ (.A1(_08464_),
    .A2(_08803_),
    .Y(_08805_),
    .B1(_08804_));
 sg13g2_nand2_1 _34528_ (.Y(_08806_),
    .A(net5701),
    .B(\u_inv.d_next[65] ));
 sg13g2_nor2_1 _34529_ (.A(net4995),
    .B(_08805_),
    .Y(_08807_));
 sg13g2_a21oi_1 _34530_ (.A1(_05348_),
    .A2(_05403_),
    .Y(_08808_),
    .B1(_05655_));
 sg13g2_xnor2_1 _34531_ (.Y(_08809_),
    .A(_05400_),
    .B(_08808_));
 sg13g2_a22oi_1 _34532_ (.Y(_08810_),
    .B1(_08809_),
    .B2(net4995),
    .A2(_08807_),
    .A1(_08806_));
 sg13g2_inv_1 _34533_ (.Y(_08811_),
    .A(_08810_));
 sg13g2_xnor2_1 _34534_ (.Y(_08812_),
    .A(_05402_),
    .B(_06268_));
 sg13g2_o21ai_1 _34535_ (.B1(net5081),
    .Y(_08813_),
    .A1(net5801),
    .A2(\u_inv.d_next[64] ));
 sg13g2_a21o_1 _34536_ (.A2(_08812_),
    .A1(net5801),
    .B1(_08813_),
    .X(_08814_));
 sg13g2_xnor2_1 _34537_ (.Y(_08815_),
    .A(_05348_),
    .B(_05403_));
 sg13g2_o21ai_1 _34538_ (.B1(_08814_),
    .Y(_08816_),
    .A1(net5081),
    .A2(_08815_));
 sg13g2_nand2_1 _34539_ (.Y(_08817_),
    .A(net4772),
    .B(_08816_));
 sg13g2_o21ai_1 _34540_ (.B1(net4772),
    .Y(_08818_),
    .A1(_08810_),
    .A2(_08816_));
 sg13g2_a21o_1 _34541_ (.A2(_08800_),
    .A1(_08790_),
    .B1(net4821),
    .X(_08819_));
 sg13g2_o21ai_1 _34542_ (.B1(_08819_),
    .Y(_08820_),
    .A1(_08802_),
    .A2(_08818_));
 sg13g2_o21ai_1 _34543_ (.B1(_08751_),
    .Y(_08821_),
    .A1(net4821),
    .A2(_08761_));
 sg13g2_o21ai_1 _34544_ (.B1(_08781_),
    .Y(_08822_),
    .A1(net4821),
    .A2(_08772_));
 sg13g2_a221oi_1 _34545_ (.B2(_08763_),
    .C1(_08821_),
    .B1(_08822_),
    .A1(_08783_),
    .Y(_08823_),
    .A2(_08820_));
 sg13g2_nor2_2 _34546_ (.A(_08736_),
    .B(_08823_),
    .Y(_08824_));
 sg13g2_nor2b_1 _34547_ (.A(_08690_),
    .B_N(_08698_),
    .Y(_08825_));
 sg13g2_nand2b_1 _34548_ (.Y(_08826_),
    .B(_08680_),
    .A_N(_08825_));
 sg13g2_nor2_1 _34549_ (.A(_08666_),
    .B(_08677_),
    .Y(_08827_));
 sg13g2_o21ai_1 _34550_ (.B1(net4777),
    .Y(_08828_),
    .A1(_08721_),
    .A2(_08731_));
 sg13g2_a21oi_1 _34551_ (.A1(net4777),
    .A2(_08714_),
    .Y(_08829_),
    .B1(_08707_));
 sg13g2_o21ai_1 _34552_ (.B1(_08829_),
    .Y(_08830_),
    .A1(_08716_),
    .A2(_08828_));
 sg13g2_nand4_1 _34553_ (.B(_08691_),
    .C(_08699_),
    .A(_08680_),
    .Y(_08831_),
    .D(_08830_));
 sg13g2_nand3_1 _34554_ (.B(_08827_),
    .C(_08831_),
    .A(_08826_),
    .Y(_08832_));
 sg13g2_nor2_2 _34555_ (.A(_08824_),
    .B(_08832_),
    .Y(_08833_));
 sg13g2_o21ai_1 _34556_ (.B1(_08646_),
    .Y(_08834_),
    .A1(_08824_),
    .A2(_08832_));
 sg13g2_a21oi_1 _34557_ (.A1(net4782),
    .A2(_08639_),
    .Y(_08835_),
    .B1(_08609_));
 sg13g2_a21o_1 _34558_ (.A2(_08630_),
    .A1(_08619_),
    .B1(net4826),
    .X(_08836_));
 sg13g2_o21ai_1 _34559_ (.B1(_08836_),
    .Y(_08837_),
    .A1(_08632_),
    .A2(_08835_));
 sg13g2_nand4_1 _34560_ (.B(_08594_),
    .C(_08601_),
    .A(_08582_),
    .Y(_08838_),
    .D(_08837_));
 sg13g2_o21ai_1 _34561_ (.B1(net4783),
    .Y(_08839_),
    .A1(_08592_),
    .A2(_08599_));
 sg13g2_a21oi_1 _34562_ (.A1(net4783),
    .A2(_08580_),
    .Y(_08840_),
    .B1(_08570_));
 sg13g2_o21ai_1 _34563_ (.B1(_08840_),
    .Y(_08841_),
    .A1(_08583_),
    .A2(_08839_));
 sg13g2_nand2b_2 _34564_ (.Y(_08842_),
    .B(_08838_),
    .A_N(_08841_));
 sg13g2_nand2_1 _34565_ (.Y(_08843_),
    .A(_08550_),
    .B(_08842_));
 sg13g2_nor2b_1 _34566_ (.A(_08538_),
    .B_N(_08546_),
    .Y(_08844_));
 sg13g2_nand3b_1 _34567_ (.B(_08527_),
    .C(_08519_),
    .Y(_08845_),
    .A_N(_08844_));
 sg13g2_a21oi_1 _34568_ (.A1(_08518_),
    .A2(_08525_),
    .Y(_08846_),
    .B1(net4828));
 sg13g2_nor2b_2 _34569_ (.A(_08846_),
    .B_N(_08845_),
    .Y(_08847_));
 sg13g2_nor4_1 _34570_ (.A(_08480_),
    .B(_08488_),
    .C(_08507_),
    .D(_08847_),
    .Y(_08848_));
 sg13g2_nand2_1 _34571_ (.Y(_08849_),
    .A(_08497_),
    .B(_08504_));
 sg13g2_a221oi_1 _34572_ (.B2(_08849_),
    .C1(_08848_),
    .B1(_08489_),
    .A1(net4783),
    .Y(_08850_),
    .A2(_08479_));
 sg13g2_and4_1 _34573_ (.A(_08487_),
    .B(_08834_),
    .C(_08843_),
    .D(_08850_),
    .X(_08851_));
 sg13g2_o21ai_1 _34574_ (.B1(_05327_),
    .Y(_08852_),
    .A1(_05259_),
    .A2(_05263_));
 sg13g2_a221oi_1 _34575_ (.B2(_05262_),
    .C1(net5617),
    .B1(_05261_),
    .A1(_05230_),
    .Y(_08853_),
    .A2(_05258_));
 sg13g2_nor2_1 _34576_ (.A(_05328_),
    .B(_08853_),
    .Y(_08854_));
 sg13g2_o21ai_1 _34577_ (.B1(_05311_),
    .Y(_08855_),
    .A1(_05328_),
    .A2(_08853_));
 sg13g2_a21oi_1 _34578_ (.A1(_05326_),
    .A2(_08855_),
    .Y(_08856_),
    .B1(_05283_));
 sg13g2_a21o_1 _34579_ (.A2(_08855_),
    .A1(_05326_),
    .B1(_05283_),
    .X(_08857_));
 sg13g2_o21ai_1 _34580_ (.B1(_05288_),
    .Y(_08858_),
    .A1(_05336_),
    .A2(_08856_));
 sg13g2_a21oi_1 _34581_ (.A1(_05337_),
    .A2(_08857_),
    .Y(_08859_),
    .B1(_05290_));
 sg13g2_o21ai_1 _34582_ (.B1(_05278_),
    .Y(_08860_),
    .A1(_05340_),
    .A2(_08859_));
 sg13g2_nand2_1 _34583_ (.Y(_08861_),
    .A(_05331_),
    .B(_08860_));
 sg13g2_a21oi_1 _34584_ (.A1(_05331_),
    .A2(_08860_),
    .Y(_08862_),
    .B1(_05270_));
 sg13g2_xnor2_1 _34585_ (.Y(_08863_),
    .A(_05270_),
    .B(_08861_));
 sg13g2_o21ai_1 _34586_ (.B1(_06151_),
    .Y(_08864_),
    .A1(_06261_),
    .A2(_06264_));
 sg13g2_nand2_1 _34587_ (.Y(_08865_),
    .A(_06129_),
    .B(_08864_));
 sg13g2_o21ai_1 _34588_ (.B1(_06136_),
    .Y(_08866_),
    .A1(_06123_),
    .A2(_08864_));
 sg13g2_nand2_1 _34589_ (.Y(_08867_),
    .A(_06119_),
    .B(_08866_));
 sg13g2_nand3_1 _34590_ (.B(_06119_),
    .C(_08866_),
    .A(_06118_),
    .Y(_08868_));
 sg13g2_a21oi_1 _34591_ (.A1(_06142_),
    .A2(_08868_),
    .Y(_08869_),
    .B1(_05277_));
 sg13g2_nor2b_1 _34592_ (.A(_05274_),
    .B_N(_08869_),
    .Y(_08870_));
 sg13g2_nor3_1 _34593_ (.A(_05270_),
    .B(_06147_),
    .C(_08870_),
    .Y(_08871_));
 sg13g2_o21ai_1 _34594_ (.B1(_05270_),
    .Y(_08872_),
    .A1(_06147_),
    .A2(_08870_));
 sg13g2_nand2_1 _34595_ (.Y(_08873_),
    .A(net5801),
    .B(_08872_));
 sg13g2_a21oi_1 _34596_ (.A1(net5701),
    .A2(\u_inv.d_next[62] ),
    .Y(_08874_),
    .B1(net4995));
 sg13g2_o21ai_1 _34597_ (.B1(_08874_),
    .Y(_08875_),
    .A1(_08871_),
    .A2(_08873_));
 sg13g2_o21ai_1 _34598_ (.B1(_08875_),
    .Y(_08876_),
    .A1(net5071),
    .A2(_08863_));
 sg13g2_nand2b_1 _34599_ (.Y(_08877_),
    .B(net4769),
    .A_N(_08876_));
 sg13g2_xnor2_1 _34600_ (.Y(_08878_),
    .A(net4820),
    .B(_08876_));
 sg13g2_o21ai_1 _34601_ (.B1(_05267_),
    .Y(_08879_),
    .A1(_05333_),
    .A2(_08862_));
 sg13g2_or3_1 _34602_ (.A(_05267_),
    .B(_05333_),
    .C(_08862_),
    .X(_08880_));
 sg13g2_nand3_1 _34603_ (.B(_08879_),
    .C(_08880_),
    .A(net4995),
    .Y(_08881_));
 sg13g2_nand3_1 _34604_ (.B(_05269_),
    .C(_08872_),
    .A(_05268_),
    .Y(_08882_));
 sg13g2_a21o_1 _34605_ (.A2(_08872_),
    .A1(_05269_),
    .B1(_05268_),
    .X(_08883_));
 sg13g2_nand3_1 _34606_ (.B(_08882_),
    .C(_08883_),
    .A(net5801),
    .Y(_08884_));
 sg13g2_nand2_1 _34607_ (.Y(_08885_),
    .A(net5701),
    .B(\u_inv.d_next[63] ));
 sg13g2_nand3_1 _34608_ (.B(_08884_),
    .C(_08885_),
    .A(net5081),
    .Y(_08886_));
 sg13g2_and3_2 _34609_ (.X(_08887_),
    .A(net4769),
    .B(_08881_),
    .C(_08886_));
 sg13g2_nand3_1 _34610_ (.B(_08881_),
    .C(_08886_),
    .A(net4769),
    .Y(_08888_));
 sg13g2_a21oi_1 _34611_ (.A1(_08881_),
    .A2(_08886_),
    .Y(_08889_),
    .B1(net4769));
 sg13g2_nor2_1 _34612_ (.A(_08887_),
    .B(_08889_),
    .Y(_08890_));
 sg13g2_nor3_1 _34613_ (.A(_08878_),
    .B(_08887_),
    .C(_08889_),
    .Y(_08891_));
 sg13g2_or3_1 _34614_ (.A(_08878_),
    .B(_08887_),
    .C(_08889_),
    .X(_08892_));
 sg13g2_a221oi_1 _34615_ (.B2(_08858_),
    .C1(_05284_),
    .B1(_05339_),
    .A1(_05275_),
    .Y(_08893_),
    .A2(_05276_));
 sg13g2_o21ai_1 _34616_ (.B1(_05277_),
    .Y(_08894_),
    .A1(_05340_),
    .A2(_08859_));
 sg13g2_a21o_1 _34617_ (.A2(_08894_),
    .A1(_05329_),
    .B1(_05274_),
    .X(_08895_));
 sg13g2_nand3_1 _34618_ (.B(_05329_),
    .C(_08894_),
    .A(_05274_),
    .Y(_08896_));
 sg13g2_nand3_1 _34619_ (.B(_08895_),
    .C(_08896_),
    .A(net4986),
    .Y(_08897_));
 sg13g2_nand3b_1 _34620_ (.B(_05274_),
    .C(_05275_),
    .Y(_08898_),
    .A_N(_08869_));
 sg13g2_o21ai_1 _34621_ (.B1(net5801),
    .Y(_08899_),
    .A1(_05274_),
    .A2(_05275_));
 sg13g2_nor2_1 _34622_ (.A(_08870_),
    .B(_08899_),
    .Y(_08900_));
 sg13g2_a22oi_1 _34623_ (.Y(_08901_),
    .B1(_08898_),
    .B2(_08900_),
    .A2(\u_inv.d_next[61] ),
    .A1(net5701));
 sg13g2_nand2_1 _34624_ (.Y(_08902_),
    .A(net5071),
    .B(_08901_));
 sg13g2_nand3_1 _34625_ (.B(_08897_),
    .C(_08902_),
    .A(net4769),
    .Y(_08903_));
 sg13g2_a21oi_1 _34626_ (.A1(_08897_),
    .A2(_08902_),
    .Y(_08904_),
    .B1(net4769));
 sg13g2_a21o_1 _34627_ (.A2(_08902_),
    .A1(_08897_),
    .B1(net4769),
    .X(_08905_));
 sg13g2_and2_1 _34628_ (.A(_08903_),
    .B(_08905_),
    .X(_08906_));
 sg13g2_nand3_1 _34629_ (.B(_06142_),
    .C(_08868_),
    .A(_05277_),
    .Y(_08907_));
 sg13g2_nand2_1 _34630_ (.Y(_08908_),
    .A(net5696),
    .B(\u_inv.d_next[60] ));
 sg13g2_nand2_1 _34631_ (.Y(_08909_),
    .A(net5790),
    .B(_08907_));
 sg13g2_o21ai_1 _34632_ (.B1(_08908_),
    .Y(_08910_),
    .A1(_08869_),
    .A2(_08909_));
 sg13g2_nor3_1 _34633_ (.A(_05277_),
    .B(_05340_),
    .C(_08859_),
    .Y(_08911_));
 sg13g2_nor3_1 _34634_ (.A(net5071),
    .B(_08893_),
    .C(_08911_),
    .Y(_08912_));
 sg13g2_a21o_1 _34635_ (.A2(_08910_),
    .A1(net5071),
    .B1(_08912_),
    .X(_08913_));
 sg13g2_nand2_1 _34636_ (.Y(_08914_),
    .A(net4769),
    .B(_08913_));
 sg13g2_xnor2_1 _34637_ (.Y(_08915_),
    .A(net4820),
    .B(_08913_));
 sg13g2_nand3_1 _34638_ (.B(_08905_),
    .C(_08915_),
    .A(_08903_),
    .Y(_08916_));
 sg13g2_nor4_1 _34639_ (.A(_08878_),
    .B(_08887_),
    .C(_08889_),
    .D(_08916_),
    .Y(_08917_));
 sg13g2_nand3b_1 _34640_ (.B(_05337_),
    .C(_08857_),
    .Y(_08918_),
    .A_N(_05288_));
 sg13g2_nand2_1 _34641_ (.Y(_08919_),
    .A(_08858_),
    .B(_08918_));
 sg13g2_nand2b_1 _34642_ (.Y(_08920_),
    .B(_08867_),
    .A_N(_06138_));
 sg13g2_a21o_1 _34643_ (.A2(_08867_),
    .A1(_06139_),
    .B1(_05288_),
    .X(_08921_));
 sg13g2_nand3_1 _34644_ (.B(_06139_),
    .C(_08867_),
    .A(_05288_),
    .Y(_08922_));
 sg13g2_nand3_1 _34645_ (.B(_08921_),
    .C(_08922_),
    .A(net5790),
    .Y(_08923_));
 sg13g2_a21oi_1 _34646_ (.A1(net5696),
    .A2(\u_inv.d_next[58] ),
    .Y(_08924_),
    .B1(net4986));
 sg13g2_a22oi_1 _34647_ (.Y(_08925_),
    .B1(_08923_),
    .B2(_08924_),
    .A2(_08919_),
    .A1(net4986));
 sg13g2_and2_1 _34648_ (.A(net4764),
    .B(_08925_),
    .X(_08926_));
 sg13g2_xnor2_1 _34649_ (.Y(_08927_),
    .A(net4764),
    .B(_08925_));
 sg13g2_a21oi_1 _34650_ (.A1(_05338_),
    .A2(_08858_),
    .Y(_08928_),
    .B1(_05286_));
 sg13g2_nand3_1 _34651_ (.B(_05338_),
    .C(_08858_),
    .A(_05286_),
    .Y(_08929_));
 sg13g2_nor2_1 _34652_ (.A(net5071),
    .B(_08928_),
    .Y(_08930_));
 sg13g2_nand2_1 _34653_ (.Y(_08931_),
    .A(_05287_),
    .B(_08921_));
 sg13g2_xnor2_1 _34654_ (.Y(_08932_),
    .A(_05286_),
    .B(_08931_));
 sg13g2_nand2_1 _34655_ (.Y(_08933_),
    .A(net5790),
    .B(_08932_));
 sg13g2_a21oi_1 _34656_ (.A1(net5696),
    .A2(\u_inv.d_next[59] ),
    .Y(_08934_),
    .B1(net4986));
 sg13g2_a22oi_1 _34657_ (.Y(_08935_),
    .B1(_08933_),
    .B2(_08934_),
    .A2(_08930_),
    .A1(_08929_));
 sg13g2_xnor2_1 _34658_ (.Y(_08936_),
    .A(net4817),
    .B(_08935_));
 sg13g2_nand2b_1 _34659_ (.Y(_08937_),
    .B(_08936_),
    .A_N(_08927_));
 sg13g2_o21ai_1 _34660_ (.B1(net5071),
    .Y(_08938_),
    .A1(net5790),
    .A2(\u_inv.d_next[57] ));
 sg13g2_nand2_1 _34661_ (.Y(_08939_),
    .A(_05280_),
    .B(_05281_));
 sg13g2_a21oi_1 _34662_ (.A1(_05282_),
    .A2(_08866_),
    .Y(_08940_),
    .B1(_08939_));
 sg13g2_o21ai_1 _34663_ (.B1(net5790),
    .Y(_08941_),
    .A1(_08920_),
    .A2(_08940_));
 sg13g2_nand2b_1 _34664_ (.Y(_08942_),
    .B(_08941_),
    .A_N(_08938_));
 sg13g2_a21oi_1 _34665_ (.A1(_05326_),
    .A2(_08855_),
    .Y(_08943_),
    .B1(_05282_));
 sg13g2_nor2_1 _34666_ (.A(_05334_),
    .B(_08943_),
    .Y(_08944_));
 sg13g2_xor2_1 _34667_ (.B(_08944_),
    .A(_05280_),
    .X(_08945_));
 sg13g2_o21ai_1 _34668_ (.B1(_08942_),
    .Y(_08946_),
    .A1(net5072),
    .A2(_08945_));
 sg13g2_inv_1 _34669_ (.Y(_08947_),
    .A(_08946_));
 sg13g2_xor2_1 _34670_ (.B(_08866_),
    .A(_05282_),
    .X(_08948_));
 sg13g2_mux2_1 _34671_ (.A0(\u_inv.d_next[56] ),
    .A1(_08948_),
    .S(net5790),
    .X(_08949_));
 sg13g2_nand2_1 _34672_ (.Y(_08950_),
    .A(net5071),
    .B(_08949_));
 sg13g2_nand3_1 _34673_ (.B(_05326_),
    .C(_08855_),
    .A(_05282_),
    .Y(_08951_));
 sg13g2_nand2b_1 _34674_ (.Y(_08952_),
    .B(_08951_),
    .A_N(_08943_));
 sg13g2_o21ai_1 _34675_ (.B1(_08950_),
    .Y(_08953_),
    .A1(net5071),
    .A2(_08952_));
 sg13g2_and2_1 _34676_ (.A(net4764),
    .B(_08953_),
    .X(_08954_));
 sg13g2_o21ai_1 _34677_ (.B1(net4765),
    .Y(_08955_),
    .A1(_08946_),
    .A2(_08953_));
 sg13g2_a21oi_1 _34678_ (.A1(net4765),
    .A2(_08935_),
    .Y(_08956_),
    .B1(_08926_));
 sg13g2_o21ai_1 _34679_ (.B1(_08956_),
    .Y(_08957_),
    .A1(_08937_),
    .A2(_08955_));
 sg13g2_and2_1 _34680_ (.A(_08903_),
    .B(_08914_),
    .X(_08958_));
 sg13g2_nand2_1 _34681_ (.Y(_08959_),
    .A(_08903_),
    .B(_08914_));
 sg13g2_nand2_1 _34682_ (.Y(_08960_),
    .A(_08877_),
    .B(_08888_));
 sg13g2_a221oi_1 _34683_ (.B2(_08891_),
    .C1(_08960_),
    .B1(_08959_),
    .A1(_08917_),
    .Y(_08961_),
    .A2(_08957_));
 sg13g2_xnor2_1 _34684_ (.Y(_08962_),
    .A(net4765),
    .B(_08946_));
 sg13g2_xnor2_1 _34685_ (.Y(_08963_),
    .A(net4765),
    .B(_08953_));
 sg13g2_or3_1 _34686_ (.A(_08937_),
    .B(_08962_),
    .C(_08963_),
    .X(_08964_));
 sg13g2_or3_1 _34687_ (.A(_08892_),
    .B(_08916_),
    .C(_08964_),
    .X(_08965_));
 sg13g2_nor2_1 _34688_ (.A(_05305_),
    .B(_08854_),
    .Y(_08966_));
 sg13g2_o21ai_1 _34689_ (.B1(_05310_),
    .Y(_08967_),
    .A1(_05328_),
    .A2(_08853_));
 sg13g2_a21oi_2 _34690_ (.B1(_05302_),
    .Y(_08968_),
    .A2(_08967_),
    .A1(_05317_));
 sg13g2_a21oi_1 _34691_ (.A1(_05300_),
    .A2(_08968_),
    .Y(_08969_),
    .B1(_05320_));
 sg13g2_o21ai_1 _34692_ (.B1(_05322_),
    .Y(_08970_),
    .A1(_05296_),
    .A2(_08969_));
 sg13g2_and2_1 _34693_ (.A(_05293_),
    .B(_08970_),
    .X(_08971_));
 sg13g2_o21ai_1 _34694_ (.B1(net4986),
    .Y(_08972_),
    .A1(_05293_),
    .A2(_08970_));
 sg13g2_nand2b_1 _34695_ (.Y(_08973_),
    .B(_08865_),
    .A_N(_06121_));
 sg13g2_and2_1 _34696_ (.A(_06132_),
    .B(_08973_),
    .X(_08974_));
 sg13g2_o21ai_1 _34697_ (.B1(_05294_),
    .Y(_08975_),
    .A1(_05297_),
    .A2(_08974_));
 sg13g2_xnor2_1 _34698_ (.Y(_08976_),
    .A(_05293_),
    .B(_08975_));
 sg13g2_a21oi_1 _34699_ (.A1(net5696),
    .A2(\u_inv.d_next[55] ),
    .Y(_08977_),
    .B1(net4986));
 sg13g2_o21ai_1 _34700_ (.B1(_08977_),
    .Y(_08978_),
    .A1(net5696),
    .A2(_08976_));
 sg13g2_o21ai_1 _34701_ (.B1(_08978_),
    .Y(_08979_),
    .A1(_08971_),
    .A2(_08972_));
 sg13g2_nor2_1 _34702_ (.A(net4817),
    .B(_08979_),
    .Y(_08980_));
 sg13g2_xnor2_1 _34703_ (.Y(_08981_),
    .A(net4817),
    .B(_08979_));
 sg13g2_xnor2_1 _34704_ (.Y(_08982_),
    .A(_05296_),
    .B(_08969_));
 sg13g2_xnor2_1 _34705_ (.Y(_08983_),
    .A(_05296_),
    .B(_08974_));
 sg13g2_nand2_1 _34706_ (.Y(_08984_),
    .A(net5693),
    .B(\u_inv.d_next[54] ));
 sg13g2_a21oi_1 _34707_ (.A1(net5790),
    .A2(_08983_),
    .Y(_08985_),
    .B1(net4981));
 sg13g2_a22oi_1 _34708_ (.Y(_08986_),
    .B1(_08984_),
    .B2(_08985_),
    .A2(_08982_),
    .A1(net4981));
 sg13g2_and2_1 _34709_ (.A(net4764),
    .B(_08986_),
    .X(_08987_));
 sg13g2_xnor2_1 _34710_ (.Y(_08988_),
    .A(net4764),
    .B(_08986_));
 sg13g2_or2_1 _34711_ (.X(_08989_),
    .B(_08988_),
    .A(_08981_));
 sg13g2_xnor2_1 _34712_ (.Y(_08990_),
    .A(_05302_),
    .B(_08865_));
 sg13g2_o21ai_1 _34713_ (.B1(net5070),
    .Y(_08991_),
    .A1(net5787),
    .A2(\u_inv.d_next[52] ));
 sg13g2_a21oi_1 _34714_ (.A1(net5787),
    .A2(_08990_),
    .Y(_08992_),
    .B1(_08991_));
 sg13g2_nand3_1 _34715_ (.B(_05317_),
    .C(_08967_),
    .A(_05302_),
    .Y(_08993_));
 sg13g2_nor2_1 _34716_ (.A(net5070),
    .B(_08968_),
    .Y(_08994_));
 sg13g2_a21o_2 _34717_ (.A2(_08994_),
    .A1(_08993_),
    .B1(_08992_),
    .X(_08995_));
 sg13g2_and2_1 _34718_ (.A(net4764),
    .B(_08995_),
    .X(_08996_));
 sg13g2_xnor2_1 _34719_ (.Y(_08997_),
    .A(net4764),
    .B(_08995_));
 sg13g2_o21ai_1 _34720_ (.B1(_05299_),
    .Y(_08998_),
    .A1(_05318_),
    .A2(_08968_));
 sg13g2_or3_1 _34721_ (.A(_05299_),
    .B(_05318_),
    .C(_08968_),
    .X(_08999_));
 sg13g2_nand3_1 _34722_ (.B(_08998_),
    .C(_08999_),
    .A(net4981),
    .Y(_09000_));
 sg13g2_a21oi_1 _34723_ (.A1(_05302_),
    .A2(_08865_),
    .Y(_09001_),
    .B1(_05301_));
 sg13g2_xnor2_1 _34724_ (.Y(_09002_),
    .A(_05300_),
    .B(_09001_));
 sg13g2_nor2_1 _34725_ (.A(net5787),
    .B(_14230_),
    .Y(_09003_));
 sg13g2_o21ai_1 _34726_ (.B1(net5070),
    .Y(_09004_),
    .A1(net5693),
    .A2(_09002_));
 sg13g2_o21ai_1 _34727_ (.B1(_09000_),
    .Y(_09005_),
    .A1(_09003_),
    .A2(_09004_));
 sg13g2_nor2_1 _34728_ (.A(net4817),
    .B(_09005_),
    .Y(_09006_));
 sg13g2_nand2_1 _34729_ (.Y(_09007_),
    .A(net4817),
    .B(_09005_));
 sg13g2_xnor2_1 _34730_ (.Y(_09008_),
    .A(net4764),
    .B(_09005_));
 sg13g2_nor2b_1 _34731_ (.A(_08997_),
    .B_N(_09008_),
    .Y(_09009_));
 sg13g2_xnor2_1 _34732_ (.Y(_09010_),
    .A(_05305_),
    .B(_08854_));
 sg13g2_o21ai_1 _34733_ (.B1(_05263_),
    .Y(_09011_),
    .A1(_06261_),
    .A2(_06264_));
 sg13g2_nand2b_1 _34734_ (.Y(_09012_),
    .B(net5617),
    .A_N(_09011_));
 sg13g2_and2_1 _34735_ (.A(_06125_),
    .B(_09012_),
    .X(_09013_));
 sg13g2_xnor2_1 _34736_ (.Y(_09014_),
    .A(_05305_),
    .B(_09013_));
 sg13g2_nand2_1 _34737_ (.Y(_09015_),
    .A(net5693),
    .B(\u_inv.d_next[50] ));
 sg13g2_a21oi_1 _34738_ (.A1(net5787),
    .A2(_09014_),
    .Y(_09016_),
    .B1(net4981));
 sg13g2_a22oi_1 _34739_ (.Y(_09017_),
    .B1(_09015_),
    .B2(_09016_),
    .A2(_09010_),
    .A1(net4983));
 sg13g2_and2_1 _34740_ (.A(net4763),
    .B(_09017_),
    .X(_09018_));
 sg13g2_xnor2_1 _34741_ (.Y(_09019_),
    .A(net4815),
    .B(_09017_));
 sg13g2_xnor2_1 _34742_ (.Y(_09020_),
    .A(net4763),
    .B(_09017_));
 sg13g2_o21ai_1 _34743_ (.B1(_05309_),
    .Y(_09021_),
    .A1(_05316_),
    .A2(_08966_));
 sg13g2_or3_1 _34744_ (.A(_05309_),
    .B(_05316_),
    .C(_08966_),
    .X(_09022_));
 sg13g2_nand3_1 _34745_ (.B(_09021_),
    .C(_09022_),
    .A(net4983),
    .Y(_09023_));
 sg13g2_o21ai_1 _34746_ (.B1(_05304_),
    .Y(_09024_),
    .A1(_05306_),
    .A2(_09013_));
 sg13g2_xnor2_1 _34747_ (.Y(_09025_),
    .A(_05309_),
    .B(_09024_));
 sg13g2_nor2b_1 _34748_ (.A(net5787),
    .B_N(\u_inv.d_next[51] ),
    .Y(_09026_));
 sg13g2_o21ai_1 _34749_ (.B1(net5070),
    .Y(_09027_),
    .A1(net5693),
    .A2(_09025_));
 sg13g2_o21ai_1 _34750_ (.B1(_09023_),
    .Y(_09028_),
    .A1(_09026_),
    .A2(_09027_));
 sg13g2_nor2_1 _34751_ (.A(net4815),
    .B(_09028_),
    .Y(_09029_));
 sg13g2_xnor2_1 _34752_ (.Y(_09030_),
    .A(net4815),
    .B(_09028_));
 sg13g2_nand3b_1 _34753_ (.B(_09011_),
    .C(_05261_),
    .Y(_09031_),
    .A_N(net5617));
 sg13g2_a21oi_1 _34754_ (.A1(_05260_),
    .A2(net5617),
    .Y(_09032_),
    .B1(net5693));
 sg13g2_nand3_1 _34755_ (.B(_09031_),
    .C(_09032_),
    .A(_09012_),
    .Y(_09033_));
 sg13g2_a21oi_1 _34756_ (.A1(net5693),
    .A2(\u_inv.d_next[49] ),
    .Y(_09034_),
    .B1(net4981));
 sg13g2_o21ai_1 _34757_ (.B1(net4981),
    .Y(_09035_),
    .A1(net5617),
    .A2(_08852_));
 sg13g2_a21oi_1 _34758_ (.A1(net5617),
    .A2(_08852_),
    .Y(_09036_),
    .B1(_09035_));
 sg13g2_a21oi_2 _34759_ (.B1(_09036_),
    .Y(_09037_),
    .A2(_09034_),
    .A1(_09033_));
 sg13g2_nor3_1 _34760_ (.A(_05263_),
    .B(_06261_),
    .C(_06264_),
    .Y(_09038_));
 sg13g2_nand3b_1 _34761_ (.B(net5787),
    .C(_09011_),
    .Y(_09039_),
    .A_N(_09038_));
 sg13g2_xnor2_1 _34762_ (.Y(_09040_),
    .A(_05259_),
    .B(_05263_));
 sg13g2_a21oi_1 _34763_ (.A1(net5693),
    .A2(\u_inv.d_next[48] ),
    .Y(_09041_),
    .B1(net4981));
 sg13g2_a22oi_1 _34764_ (.Y(_09042_),
    .B1(_09041_),
    .B2(_09039_),
    .A2(_09040_),
    .A1(net4981));
 sg13g2_nand2_1 _34765_ (.Y(_09043_),
    .A(net4763),
    .B(_09042_));
 sg13g2_o21ai_1 _34766_ (.B1(net4763),
    .Y(_09044_),
    .A1(_09037_),
    .A2(_09042_));
 sg13g2_nor3_1 _34767_ (.A(_09020_),
    .B(_09030_),
    .C(_09044_),
    .Y(_09045_));
 sg13g2_or2_1 _34768_ (.X(_09046_),
    .B(_09029_),
    .A(_09018_));
 sg13g2_nor2_1 _34769_ (.A(_09045_),
    .B(_09046_),
    .Y(_09047_));
 sg13g2_o21ai_1 _34770_ (.B1(_09009_),
    .Y(_09048_),
    .A1(_09045_),
    .A2(_09046_));
 sg13g2_nor2_1 _34771_ (.A(_08996_),
    .B(_09006_),
    .Y(_09049_));
 sg13g2_or2_1 _34772_ (.X(_09050_),
    .B(_09006_),
    .A(_08996_));
 sg13g2_a21oi_1 _34773_ (.A1(_09048_),
    .A2(_09049_),
    .Y(_09051_),
    .B1(_08989_));
 sg13g2_nor3_2 _34774_ (.A(_08980_),
    .B(_08987_),
    .C(_09051_),
    .Y(_09052_));
 sg13g2_o21ai_1 _34775_ (.B1(_08961_),
    .Y(_09053_),
    .A1(_08965_),
    .A2(_09052_));
 sg13g2_a221oi_1 _34776_ (.B2(_05221_),
    .C1(_05220_),
    .B1(_05231_),
    .A1(_05172_),
    .Y(_09054_),
    .A2(_05226_));
 sg13g2_inv_1 _34777_ (.Y(_09055_),
    .A(_09054_));
 sg13g2_o21ai_1 _34778_ (.B1(_05237_),
    .Y(_09056_),
    .A1(_05219_),
    .A2(_09054_));
 sg13g2_a21o_1 _34779_ (.A2(_09056_),
    .A1(_05215_),
    .B1(_05241_),
    .X(_09057_));
 sg13g2_xnor2_1 _34780_ (.Y(_09058_),
    .A(_05208_),
    .B(_09057_));
 sg13g2_a21oi_1 _34781_ (.A1(_06206_),
    .A2(net1070),
    .Y(_09059_),
    .B1(_05225_));
 sg13g2_and2_1 _34782_ (.A(net5618),
    .B(_09059_),
    .X(_09060_));
 sg13g2_nand2_1 _34783_ (.Y(_09061_),
    .A(net5618),
    .B(_09059_));
 sg13g2_a21oi_2 _34784_ (.B1(_06167_),
    .Y(_09062_),
    .A2(_09060_),
    .A1(_06249_));
 sg13g2_nor2_1 _34785_ (.A(_06159_),
    .B(_09062_),
    .Y(_09063_));
 sg13g2_nor2_1 _34786_ (.A(_06169_),
    .B(_09063_),
    .Y(_09064_));
 sg13g2_xor2_1 _34787_ (.B(_09064_),
    .A(_05208_),
    .X(_09065_));
 sg13g2_nand2_1 _34788_ (.Y(_09066_),
    .A(net5675),
    .B(\u_inv.d_next[38] ));
 sg13g2_a21oi_1 _34789_ (.A1(net5758),
    .A2(_09065_),
    .Y(_09067_),
    .B1(net4957));
 sg13g2_a22oi_1 _34790_ (.Y(_09068_),
    .B1(_09066_),
    .B2(_09067_),
    .A2(_09058_),
    .A1(net4957));
 sg13g2_nand2_1 _34791_ (.Y(_09069_),
    .A(net4748),
    .B(_09068_));
 sg13g2_xnor2_1 _34792_ (.Y(_09070_),
    .A(net4803),
    .B(_09068_));
 sg13g2_a21oi_1 _34793_ (.A1(_05208_),
    .A2(_09057_),
    .Y(_09071_),
    .B1(_05242_));
 sg13g2_o21ai_1 _34794_ (.B1(net4957),
    .Y(_09072_),
    .A1(_05205_),
    .A2(_09071_));
 sg13g2_a21oi_1 _34795_ (.A1(_05205_),
    .A2(_09071_),
    .Y(_09073_),
    .B1(_09072_));
 sg13g2_o21ai_1 _34796_ (.B1(_05206_),
    .Y(_09074_),
    .A1(_05208_),
    .A2(_09064_));
 sg13g2_xnor2_1 _34797_ (.Y(_09075_),
    .A(_05205_),
    .B(_09074_));
 sg13g2_nand2_1 _34798_ (.Y(_09076_),
    .A(net5675),
    .B(\u_inv.d_next[39] ));
 sg13g2_a21oi_1 _34799_ (.A1(net5758),
    .A2(_09075_),
    .Y(_09077_),
    .B1(net4958));
 sg13g2_a21oi_2 _34800_ (.B1(_09073_),
    .Y(_09078_),
    .A2(_09077_),
    .A1(_09076_));
 sg13g2_xnor2_1 _34801_ (.Y(_09079_),
    .A(net4803),
    .B(_09078_));
 sg13g2_nand2_1 _34802_ (.Y(_09080_),
    .A(_09070_),
    .B(_09079_));
 sg13g2_xnor2_1 _34803_ (.Y(_09081_),
    .A(_05214_),
    .B(_09062_));
 sg13g2_o21ai_1 _34804_ (.B1(net5048),
    .Y(_09082_),
    .A1(net5758),
    .A2(\u_inv.d_next[36] ));
 sg13g2_a21o_1 _34805_ (.A2(_09081_),
    .A1(net5759),
    .B1(_09082_),
    .X(_09083_));
 sg13g2_xnor2_1 _34806_ (.Y(_09084_),
    .A(_05214_),
    .B(_09056_));
 sg13g2_o21ai_1 _34807_ (.B1(_09083_),
    .Y(_09085_),
    .A1(net5048),
    .A2(_09084_));
 sg13g2_nand2_1 _34808_ (.Y(_09086_),
    .A(net4748),
    .B(_09085_));
 sg13g2_o21ai_1 _34809_ (.B1(_05212_),
    .Y(_09087_),
    .A1(_05214_),
    .A2(_09062_));
 sg13g2_nand2_1 _34810_ (.Y(_09088_),
    .A(_05211_),
    .B(_09087_));
 sg13g2_nor2_1 _34811_ (.A(_05211_),
    .B(_09087_),
    .Y(_09089_));
 sg13g2_nor2_1 _34812_ (.A(net5675),
    .B(_09089_),
    .Y(_09090_));
 sg13g2_a221oi_1 _34813_ (.B2(_09090_),
    .C1(net4958),
    .B1(_09088_),
    .A1(net5675),
    .Y(_09091_),
    .A2(\u_inv.d_next[37] ));
 sg13g2_a21o_1 _34814_ (.A2(_09056_),
    .A1(_05214_),
    .B1(_05239_),
    .X(_09092_));
 sg13g2_o21ai_1 _34815_ (.B1(net4957),
    .Y(_09093_),
    .A1(_05211_),
    .A2(_09092_));
 sg13g2_a21oi_1 _34816_ (.A1(_05211_),
    .A2(_09092_),
    .Y(_09094_),
    .B1(_09093_));
 sg13g2_nor2_2 _34817_ (.A(_09091_),
    .B(_09094_),
    .Y(_09095_));
 sg13g2_o21ai_1 _34818_ (.B1(net4748),
    .Y(_09096_),
    .A1(_09085_),
    .A2(_09095_));
 sg13g2_xnor2_1 _34819_ (.Y(_09097_),
    .A(net4748),
    .B(_09085_));
 sg13g2_inv_1 _34820_ (.Y(_09098_),
    .A(_09097_));
 sg13g2_nand2b_1 _34821_ (.Y(_09099_),
    .B(net4804),
    .A_N(_09095_));
 sg13g2_xnor2_1 _34822_ (.Y(_09100_),
    .A(net4804),
    .B(_09095_));
 sg13g2_nor2b_1 _34823_ (.A(_09097_),
    .B_N(_09100_),
    .Y(_09101_));
 sg13g2_a21oi_1 _34824_ (.A1(_05217_),
    .A2(_09055_),
    .Y(_09102_),
    .B1(_05234_));
 sg13g2_a21oi_1 _34825_ (.A1(_05218_),
    .A2(_09102_),
    .Y(_09103_),
    .B1(net5048));
 sg13g2_o21ai_1 _34826_ (.B1(_09103_),
    .Y(_09104_),
    .A1(_05218_),
    .A2(_09102_));
 sg13g2_a21o_1 _34827_ (.A2(_09061_),
    .A1(_06164_),
    .B1(_05217_),
    .X(_09105_));
 sg13g2_o21ai_1 _34828_ (.B1(_09105_),
    .Y(_09106_),
    .A1(_14235_),
    .A2(_14775_));
 sg13g2_xor2_1 _34829_ (.B(_09106_),
    .A(_05218_),
    .X(_09107_));
 sg13g2_a21oi_1 _34830_ (.A1(net5675),
    .A2(\u_inv.d_next[35] ),
    .Y(_09108_),
    .B1(net4957));
 sg13g2_o21ai_1 _34831_ (.B1(_09108_),
    .Y(_09109_),
    .A1(net5675),
    .A2(_09107_));
 sg13g2_nand2_2 _34832_ (.Y(_09110_),
    .A(_09104_),
    .B(_09109_));
 sg13g2_xnor2_1 _34833_ (.Y(_09111_),
    .A(net4803),
    .B(_09110_));
 sg13g2_xnor2_1 _34834_ (.Y(_09112_),
    .A(_05217_),
    .B(_09054_));
 sg13g2_and3_1 _34835_ (.X(_09113_),
    .A(_05217_),
    .B(_06164_),
    .C(_09061_));
 sg13g2_nand2_1 _34836_ (.Y(_09114_),
    .A(net5758),
    .B(_09105_));
 sg13g2_a21oi_1 _34837_ (.A1(net5675),
    .A2(\u_inv.d_next[34] ),
    .Y(_09115_),
    .B1(net4957));
 sg13g2_o21ai_1 _34838_ (.B1(_09115_),
    .Y(_09116_),
    .A1(_09113_),
    .A2(_09114_));
 sg13g2_o21ai_1 _34839_ (.B1(_09116_),
    .Y(_09117_),
    .A1(net5048),
    .A2(_09112_));
 sg13g2_xnor2_1 _34840_ (.Y(_09118_),
    .A(net4803),
    .B(_09117_));
 sg13g2_or2_1 _34841_ (.X(_09119_),
    .B(_09118_),
    .A(_09111_));
 sg13g2_inv_1 _34842_ (.Y(_09120_),
    .A(_09119_));
 sg13g2_nor3_1 _34843_ (.A(net5618),
    .B(_05223_),
    .C(_09059_),
    .Y(_09121_));
 sg13g2_or3_1 _34844_ (.A(_06162_),
    .B(_09060_),
    .C(_09121_),
    .X(_09122_));
 sg13g2_o21ai_1 _34845_ (.B1(net5048),
    .Y(_09123_),
    .A1(net5758),
    .A2(\u_inv.d_next[33] ));
 sg13g2_a21oi_1 _34846_ (.A1(net5758),
    .A2(_09122_),
    .Y(_09124_),
    .B1(_09123_));
 sg13g2_a21oi_1 _34847_ (.A1(_05172_),
    .A2(_05225_),
    .Y(_09125_),
    .B1(_05231_));
 sg13g2_xor2_1 _34848_ (.B(_09125_),
    .A(net5618),
    .X(_09126_));
 sg13g2_a21oi_2 _34849_ (.B1(_09124_),
    .Y(_09127_),
    .A2(_09126_),
    .A1(net4957));
 sg13g2_xnor2_1 _34850_ (.Y(_09128_),
    .A(_05224_),
    .B(_06248_));
 sg13g2_o21ai_1 _34851_ (.B1(net5048),
    .Y(_09129_),
    .A1(net5758),
    .A2(\u_inv.d_next[32] ));
 sg13g2_a21oi_1 _34852_ (.A1(net5758),
    .A2(_09128_),
    .Y(_09130_),
    .B1(_09129_));
 sg13g2_xnor2_1 _34853_ (.Y(_09131_),
    .A(_05172_),
    .B(_05224_));
 sg13g2_a21oi_2 _34854_ (.B1(_09130_),
    .Y(_09132_),
    .A2(_09131_),
    .A1(net4957));
 sg13g2_a21o_1 _34855_ (.A2(_09132_),
    .A1(net4803),
    .B1(_09127_),
    .X(_09133_));
 sg13g2_nor3_1 _34856_ (.A(_09111_),
    .B(_09118_),
    .C(_09133_),
    .Y(_09134_));
 sg13g2_a21oi_1 _34857_ (.A1(_09110_),
    .A2(_09117_),
    .Y(_09135_),
    .B1(net4803));
 sg13g2_nor2_1 _34858_ (.A(_09134_),
    .B(_09135_),
    .Y(_09136_));
 sg13g2_inv_1 _34859_ (.Y(_09137_),
    .A(_09136_));
 sg13g2_o21ai_1 _34860_ (.B1(_09101_),
    .Y(_09138_),
    .A1(_09134_),
    .A2(_09135_));
 sg13g2_a21oi_1 _34861_ (.A1(_09096_),
    .A2(_09138_),
    .Y(_09139_),
    .B1(_09080_));
 sg13g2_o21ai_1 _34862_ (.B1(net4748),
    .Y(_09140_),
    .A1(_09068_),
    .A2(_09078_));
 sg13g2_nand2b_2 _34863_ (.Y(_09141_),
    .B(_09140_),
    .A_N(_09139_));
 sg13g2_a21oi_2 _34864_ (.B1(_05244_),
    .Y(_09142_),
    .A2(_05227_),
    .A1(_05172_));
 sg13g2_o21ai_1 _34865_ (.B1(_05253_),
    .Y(_09143_),
    .A1(_05192_),
    .A2(_09142_));
 sg13g2_a21oi_2 _34866_ (.B1(_05255_),
    .Y(_09144_),
    .A2(_09143_),
    .A1(_05200_));
 sg13g2_inv_1 _34867_ (.Y(_09145_),
    .A(_09144_));
 sg13g2_o21ai_1 _34868_ (.B1(_05247_),
    .Y(_09146_),
    .A1(_05185_),
    .A2(_09144_));
 sg13g2_xnor2_1 _34869_ (.Y(_09147_),
    .A(_05177_),
    .B(_09146_));
 sg13g2_nor2_1 _34870_ (.A(_06156_),
    .B(_06251_),
    .Y(_09148_));
 sg13g2_a21oi_1 _34871_ (.A1(_06157_),
    .A2(_09148_),
    .Y(_09149_),
    .B1(_06259_));
 sg13g2_a21o_1 _34872_ (.A2(_09148_),
    .A1(_06157_),
    .B1(_06259_),
    .X(_09150_));
 sg13g2_a21oi_1 _34873_ (.A1(_06154_),
    .A2(_09150_),
    .Y(_09151_),
    .B1(_06252_));
 sg13g2_xor2_1 _34874_ (.B(_09151_),
    .A(_05177_),
    .X(_09152_));
 sg13g2_nand2_1 _34875_ (.Y(_09153_),
    .A(net5678),
    .B(\u_inv.d_next[46] ));
 sg13g2_a21oi_1 _34876_ (.A1(net5760),
    .A2(_09152_),
    .Y(_09154_),
    .B1(net4959));
 sg13g2_a22oi_1 _34877_ (.Y(_09155_),
    .B1(_09153_),
    .B2(_09154_),
    .A2(_09147_),
    .A1(net4959));
 sg13g2_and2_1 _34878_ (.A(net4749),
    .B(_09155_),
    .X(_09156_));
 sg13g2_xnor2_1 _34879_ (.Y(_09157_),
    .A(net4749),
    .B(_09155_));
 sg13g2_a21oi_1 _34880_ (.A1(_05177_),
    .A2(_09146_),
    .Y(_09158_),
    .B1(_05248_));
 sg13g2_or2_1 _34881_ (.X(_09159_),
    .B(_09158_),
    .A(_05175_));
 sg13g2_a21oi_1 _34882_ (.A1(_05175_),
    .A2(_09158_),
    .Y(_09160_),
    .B1(net5049));
 sg13g2_o21ai_1 _34883_ (.B1(_05176_),
    .Y(_09161_),
    .A1(_05177_),
    .A2(_09151_));
 sg13g2_xnor2_1 _34884_ (.Y(_09162_),
    .A(_05175_),
    .B(_09161_));
 sg13g2_nand2_1 _34885_ (.Y(_09163_),
    .A(net5678),
    .B(\u_inv.d_next[47] ));
 sg13g2_a21oi_1 _34886_ (.A1(net5760),
    .A2(_09162_),
    .Y(_09164_),
    .B1(net4959));
 sg13g2_a22oi_1 _34887_ (.Y(_09165_),
    .B1(_09163_),
    .B2(_09164_),
    .A2(_09160_),
    .A1(_09159_));
 sg13g2_xnor2_1 _34888_ (.Y(_09166_),
    .A(net4805),
    .B(_09165_));
 sg13g2_nand2b_1 _34889_ (.Y(_09167_),
    .B(_09166_),
    .A_N(_09157_));
 sg13g2_xnor2_1 _34890_ (.Y(_09168_),
    .A(_05184_),
    .B(_09149_));
 sg13g2_o21ai_1 _34891_ (.B1(net5049),
    .Y(_09169_),
    .A1(net5760),
    .A2(\u_inv.d_next[44] ));
 sg13g2_a21o_1 _34892_ (.A2(_09168_),
    .A1(net5760),
    .B1(_09169_),
    .X(_09170_));
 sg13g2_xor2_1 _34893_ (.B(_09144_),
    .A(_05184_),
    .X(_09171_));
 sg13g2_o21ai_1 _34894_ (.B1(_09170_),
    .Y(_09172_),
    .A1(net5049),
    .A2(_09171_));
 sg13g2_and2_1 _34895_ (.A(net4749),
    .B(_09172_),
    .X(_09173_));
 sg13g2_inv_1 _34896_ (.Y(_09174_),
    .A(_09173_));
 sg13g2_xnor2_1 _34897_ (.Y(_09175_),
    .A(net4805),
    .B(_09172_));
 sg13g2_inv_1 _34898_ (.Y(_09176_),
    .A(_09175_));
 sg13g2_a21o_1 _34899_ (.A2(_09145_),
    .A1(_05184_),
    .B1(_05246_),
    .X(_09177_));
 sg13g2_nand2b_1 _34900_ (.Y(_09178_),
    .B(_05182_),
    .A_N(_09177_));
 sg13g2_a21oi_1 _34901_ (.A1(_05181_),
    .A2(_09177_),
    .Y(_09179_),
    .B1(net5050));
 sg13g2_o21ai_1 _34902_ (.B1(_05183_),
    .Y(_09180_),
    .A1(_05184_),
    .A2(_09149_));
 sg13g2_xnor2_1 _34903_ (.Y(_09181_),
    .A(_05182_),
    .B(_09180_));
 sg13g2_nand2_1 _34904_ (.Y(_09182_),
    .A(net5678),
    .B(\u_inv.d_next[45] ));
 sg13g2_a21oi_1 _34905_ (.A1(net5760),
    .A2(_09181_),
    .Y(_09183_),
    .B1(net4959));
 sg13g2_a22oi_1 _34906_ (.Y(_09184_),
    .B1(_09182_),
    .B2(_09183_),
    .A2(_09179_),
    .A1(_09178_));
 sg13g2_nand2_1 _34907_ (.Y(_09185_),
    .A(net4749),
    .B(_09184_));
 sg13g2_nor2_1 _34908_ (.A(net4752),
    .B(_09184_),
    .Y(_09186_));
 sg13g2_xnor2_1 _34909_ (.Y(_09187_),
    .A(net4805),
    .B(_09184_));
 sg13g2_and2_1 _34910_ (.A(_09175_),
    .B(_09187_),
    .X(_09188_));
 sg13g2_nand2_1 _34911_ (.Y(_09189_),
    .A(_05199_),
    .B(_09143_));
 sg13g2_xor2_1 _34912_ (.B(_09143_),
    .A(_05199_),
    .X(_09190_));
 sg13g2_o21ai_1 _34913_ (.B1(_06256_),
    .Y(_09191_),
    .A1(_06156_),
    .A2(_06251_));
 sg13g2_xor2_1 _34914_ (.B(_09191_),
    .A(_05199_),
    .X(_09192_));
 sg13g2_a21oi_1 _34915_ (.A1(net5678),
    .A2(\u_inv.d_next[42] ),
    .Y(_09193_),
    .B1(net4959));
 sg13g2_o21ai_1 _34916_ (.B1(_09193_),
    .Y(_09194_),
    .A1(net5678),
    .A2(_09192_));
 sg13g2_o21ai_1 _34917_ (.B1(_09194_),
    .Y(_09195_),
    .A1(net5049),
    .A2(_09190_));
 sg13g2_xnor2_1 _34918_ (.Y(_09196_),
    .A(net4749),
    .B(_09195_));
 sg13g2_nand2_1 _34919_ (.Y(_09197_),
    .A(_05254_),
    .B(_09189_));
 sg13g2_and2_1 _34920_ (.A(_05195_),
    .B(_09197_),
    .X(_09198_));
 sg13g2_o21ai_1 _34921_ (.B1(net4959),
    .Y(_09199_),
    .A1(_05195_),
    .A2(_09197_));
 sg13g2_a21o_1 _34922_ (.A2(_09191_),
    .A1(_05198_),
    .B1(_05196_),
    .X(_09200_));
 sg13g2_xnor2_1 _34923_ (.Y(_09201_),
    .A(_05195_),
    .B(_09200_));
 sg13g2_a21oi_1 _34924_ (.A1(net5678),
    .A2(\u_inv.d_next[43] ),
    .Y(_09202_),
    .B1(net4959));
 sg13g2_o21ai_1 _34925_ (.B1(_09202_),
    .Y(_09203_),
    .A1(net5678),
    .A2(_09201_));
 sg13g2_o21ai_1 _34926_ (.B1(_09203_),
    .Y(_09204_),
    .A1(_09198_),
    .A2(_09199_));
 sg13g2_xnor2_1 _34927_ (.Y(_09205_),
    .A(net4749),
    .B(_09204_));
 sg13g2_nand2_1 _34928_ (.Y(_09206_),
    .A(_09196_),
    .B(_09205_));
 sg13g2_nor2_1 _34929_ (.A(_05190_),
    .B(_09142_),
    .Y(_09207_));
 sg13g2_nor2_1 _34930_ (.A(_05252_),
    .B(_09207_),
    .Y(_09208_));
 sg13g2_a21oi_1 _34931_ (.A1(_05187_),
    .A2(_09208_),
    .Y(_09209_),
    .B1(net5049));
 sg13g2_o21ai_1 _34932_ (.B1(_09209_),
    .Y(_09210_),
    .A1(_05187_),
    .A2(_09208_));
 sg13g2_o21ai_1 _34933_ (.B1(_05189_),
    .Y(_09211_),
    .A1(_05191_),
    .A2(_06251_));
 sg13g2_xnor2_1 _34934_ (.Y(_09212_),
    .A(_05188_),
    .B(_09211_));
 sg13g2_nor2b_1 _34935_ (.A(net5760),
    .B_N(\u_inv.d_next[41] ),
    .Y(_09213_));
 sg13g2_o21ai_1 _34936_ (.B1(net5049),
    .Y(_09214_),
    .A1(net5678),
    .A2(_09212_));
 sg13g2_o21ai_1 _34937_ (.B1(_09210_),
    .Y(_09215_),
    .A1(_09213_),
    .A2(_09214_));
 sg13g2_nor2_1 _34938_ (.A(net4805),
    .B(_09215_),
    .Y(_09216_));
 sg13g2_nand2_1 _34939_ (.Y(_09217_),
    .A(net4805),
    .B(_09215_));
 sg13g2_nor2b_1 _34940_ (.A(_09216_),
    .B_N(_09217_),
    .Y(_09218_));
 sg13g2_xnor2_1 _34941_ (.Y(_09219_),
    .A(_05191_),
    .B(_06251_));
 sg13g2_o21ai_1 _34942_ (.B1(net5049),
    .Y(_09220_),
    .A1(net5760),
    .A2(\u_inv.d_next[40] ));
 sg13g2_a21o_1 _34943_ (.A2(_09219_),
    .A1(net5760),
    .B1(_09220_),
    .X(_09221_));
 sg13g2_xnor2_1 _34944_ (.Y(_09222_),
    .A(_05190_),
    .B(_09142_));
 sg13g2_o21ai_1 _34945_ (.B1(_09221_),
    .Y(_09223_),
    .A1(net5049),
    .A2(_09222_));
 sg13g2_and2_1 _34946_ (.A(net4749),
    .B(_09223_),
    .X(_09224_));
 sg13g2_xnor2_1 _34947_ (.Y(_09225_),
    .A(net4749),
    .B(_09223_));
 sg13g2_inv_1 _34948_ (.Y(_09226_),
    .A(_09225_));
 sg13g2_and4_1 _34949_ (.A(_09196_),
    .B(_09205_),
    .C(_09218_),
    .D(_09226_),
    .X(_09227_));
 sg13g2_nand3b_1 _34950_ (.B(_09188_),
    .C(_09227_),
    .Y(_09228_),
    .A_N(_09167_));
 sg13g2_inv_1 _34951_ (.Y(_09229_),
    .A(_09228_));
 sg13g2_nor2_1 _34952_ (.A(_09216_),
    .B(_09224_),
    .Y(_09230_));
 sg13g2_a21o_1 _34953_ (.A2(_09204_),
    .A1(_09195_),
    .B1(net4805),
    .X(_09231_));
 sg13g2_o21ai_1 _34954_ (.B1(_09231_),
    .Y(_09232_),
    .A1(_09206_),
    .A2(_09230_));
 sg13g2_inv_1 _34955_ (.Y(_09233_),
    .A(_09232_));
 sg13g2_a221oi_1 _34956_ (.B2(_09232_),
    .C1(_09173_),
    .B1(_09188_),
    .A1(net4752),
    .Y(_09234_),
    .A2(_09184_));
 sg13g2_a21oi_1 _34957_ (.A1(net4752),
    .A2(_09165_),
    .Y(_09235_),
    .B1(_09156_));
 sg13g2_o21ai_1 _34958_ (.B1(_09235_),
    .Y(_09236_),
    .A1(_09167_),
    .A2(_09234_));
 sg13g2_a21o_2 _34959_ (.A2(_09229_),
    .A1(_09141_),
    .B1(_09236_),
    .X(_09237_));
 sg13g2_nand2b_1 _34960_ (.Y(_09238_),
    .B(net4815),
    .A_N(_09037_));
 sg13g2_xnor2_1 _34961_ (.Y(_09239_),
    .A(net4763),
    .B(_09037_));
 sg13g2_xnor2_1 _34962_ (.Y(_09240_),
    .A(net4763),
    .B(_09042_));
 sg13g2_nor4_1 _34963_ (.A(_09020_),
    .B(_09030_),
    .C(_09239_),
    .D(_09240_),
    .Y(_09241_));
 sg13g2_nand3b_1 _34964_ (.B(_09009_),
    .C(_09241_),
    .Y(_09242_),
    .A_N(_08989_));
 sg13g2_inv_1 _34965_ (.Y(_09243_),
    .A(_09242_));
 sg13g2_nor4_2 _34966_ (.A(_08892_),
    .B(_08916_),
    .C(_08964_),
    .Y(_09244_),
    .D(_09242_));
 sg13g2_a21o_2 _34967_ (.A2(_09244_),
    .A1(_09237_),
    .B1(_09053_),
    .X(_09245_));
 sg13g2_a21o_1 _34968_ (.A2(_05167_),
    .A1(_05079_),
    .B1(_05045_),
    .X(_09246_));
 sg13g2_nor2_1 _34969_ (.A(_05013_),
    .B(_09246_),
    .Y(_09247_));
 sg13g2_nor2_1 _34970_ (.A(_05015_),
    .B(_09247_),
    .Y(_09248_));
 sg13g2_o21ai_1 _34971_ (.B1(_05029_),
    .Y(_09249_),
    .A1(_05015_),
    .A2(_09247_));
 sg13g2_nand2b_1 _34972_ (.Y(_09250_),
    .B(_09249_),
    .A_N(_05040_));
 sg13g2_o21ai_1 _34973_ (.B1(_05042_),
    .Y(_09251_),
    .A1(_05030_),
    .A2(_09249_));
 sg13g2_a21o_1 _34974_ (.A2(_09251_),
    .A1(_05026_),
    .B1(_05036_),
    .X(_09252_));
 sg13g2_xnor2_1 _34975_ (.Y(_09253_),
    .A(_05020_),
    .B(_09252_));
 sg13g2_o21ai_1 _34976_ (.B1(_05163_),
    .Y(_09254_),
    .A1(_06229_),
    .A2(_06241_));
 sg13g2_or2_1 _34977_ (.X(_09255_),
    .B(_09254_),
    .A(_05161_));
 sg13g2_o21ai_1 _34978_ (.B1(_06244_),
    .Y(_09256_),
    .A1(_06229_),
    .A2(_06241_));
 sg13g2_nand2_2 _34979_ (.Y(_09257_),
    .A(_06188_),
    .B(_09256_));
 sg13g2_o21ai_1 _34980_ (.B1(_06195_),
    .Y(_09258_),
    .A1(_06181_),
    .A2(_09256_));
 sg13g2_and2_1 _34981_ (.A(_05045_),
    .B(_09258_),
    .X(_09259_));
 sg13g2_nand2_1 _34982_ (.Y(_09260_),
    .A(_05013_),
    .B(_09259_));
 sg13g2_a21oi_1 _34983_ (.A1(_06178_),
    .A2(_09258_),
    .Y(_09261_),
    .B1(_06203_));
 sg13g2_nor3_1 _34984_ (.A(_05023_),
    .B(_05025_),
    .C(_09261_),
    .Y(_09262_));
 sg13g2_nor2_1 _34985_ (.A(_06197_),
    .B(_09262_),
    .Y(_09263_));
 sg13g2_xor2_1 _34986_ (.B(_09263_),
    .A(_05020_),
    .X(_09264_));
 sg13g2_nand2_1 _34987_ (.Y(_09265_),
    .A(net5670),
    .B(\u_inv.d_next[30] ));
 sg13g2_a21oi_1 _34988_ (.A1(net5746),
    .A2(_09264_),
    .Y(_09266_),
    .B1(net4947));
 sg13g2_a22oi_1 _34989_ (.Y(_09267_),
    .B1(_09265_),
    .B2(_09266_),
    .A2(_09253_),
    .A1(net4947));
 sg13g2_nand2_1 _34990_ (.Y(_09268_),
    .A(net4744),
    .B(_09267_));
 sg13g2_inv_1 _34991_ (.Y(_09269_),
    .A(_09268_));
 sg13g2_xnor2_1 _34992_ (.Y(_09270_),
    .A(net4801),
    .B(_09267_));
 sg13g2_a21oi_1 _34993_ (.A1(_05020_),
    .A2(_09252_),
    .Y(_09271_),
    .B1(_05038_));
 sg13g2_o21ai_1 _34994_ (.B1(net4947),
    .Y(_09272_),
    .A1(_05018_),
    .A2(_09271_));
 sg13g2_a21oi_1 _34995_ (.A1(_05018_),
    .A2(_09271_),
    .Y(_09273_),
    .B1(_09272_));
 sg13g2_o21ai_1 _34996_ (.B1(_05019_),
    .Y(_09274_),
    .A1(_05020_),
    .A2(_09263_));
 sg13g2_xnor2_1 _34997_ (.Y(_09275_),
    .A(_05018_),
    .B(_09274_));
 sg13g2_nand2_1 _34998_ (.Y(_09276_),
    .A(net5670),
    .B(\u_inv.d_next[31] ));
 sg13g2_a21oi_1 _34999_ (.A1(net5746),
    .A2(_09275_),
    .Y(_09277_),
    .B1(net4947));
 sg13g2_a21oi_1 _35000_ (.A1(_09276_),
    .A2(_09277_),
    .Y(_09278_),
    .B1(_09273_));
 sg13g2_xnor2_1 _35001_ (.Y(_09279_),
    .A(net4801),
    .B(_09278_));
 sg13g2_and2_1 _35002_ (.A(_09270_),
    .B(_09279_),
    .X(_09280_));
 sg13g2_xnor2_1 _35003_ (.Y(_09281_),
    .A(_05025_),
    .B(_09261_));
 sg13g2_o21ai_1 _35004_ (.B1(net5039),
    .Y(_09282_),
    .A1(net5746),
    .A2(\u_inv.d_next[28] ));
 sg13g2_a21o_1 _35005_ (.A2(_09281_),
    .A1(net5746),
    .B1(_09282_),
    .X(_09283_));
 sg13g2_xnor2_1 _35006_ (.Y(_09284_),
    .A(_05025_),
    .B(_09251_));
 sg13g2_o21ai_1 _35007_ (.B1(_09283_),
    .Y(_09285_),
    .A1(net5039),
    .A2(_09284_));
 sg13g2_nand2_1 _35008_ (.Y(_09286_),
    .A(net4744),
    .B(_09285_));
 sg13g2_a21oi_1 _35009_ (.A1(_05025_),
    .A2(_09251_),
    .Y(_09287_),
    .B1(_05035_));
 sg13g2_o21ai_1 _35010_ (.B1(net4949),
    .Y(_09288_),
    .A1(_05023_),
    .A2(_09287_));
 sg13g2_a21oi_1 _35011_ (.A1(_05023_),
    .A2(_09287_),
    .Y(_09289_),
    .B1(_09288_));
 sg13g2_o21ai_1 _35012_ (.B1(_05024_),
    .Y(_09290_),
    .A1(_05025_),
    .A2(_09261_));
 sg13g2_xnor2_1 _35013_ (.Y(_09291_),
    .A(_05023_),
    .B(_09290_));
 sg13g2_nand2_1 _35014_ (.Y(_09292_),
    .A(net5670),
    .B(\u_inv.d_next[29] ));
 sg13g2_a21oi_1 _35015_ (.A1(net5746),
    .A2(_09291_),
    .Y(_09293_),
    .B1(net4947));
 sg13g2_a21oi_2 _35016_ (.B1(_09289_),
    .Y(_09294_),
    .A2(_09293_),
    .A1(_09292_));
 sg13g2_o21ai_1 _35017_ (.B1(net4744),
    .Y(_09295_),
    .A1(_09285_),
    .A2(_09294_));
 sg13g2_xnor2_1 _35018_ (.Y(_09296_),
    .A(net4746),
    .B(_09285_));
 sg13g2_nor2_1 _35019_ (.A(net4746),
    .B(_09294_),
    .Y(_09297_));
 sg13g2_xnor2_1 _35020_ (.Y(_09298_),
    .A(net4801),
    .B(_09294_));
 sg13g2_nor2b_1 _35021_ (.A(_09296_),
    .B_N(_09298_),
    .Y(_09299_));
 sg13g2_nand2b_1 _35022_ (.Y(_09300_),
    .B(_09298_),
    .A_N(_09296_));
 sg13g2_a21o_1 _35023_ (.A2(_09260_),
    .A1(_06200_),
    .B1(_05029_),
    .X(_09301_));
 sg13g2_nand2_1 _35024_ (.Y(_09302_),
    .A(_05028_),
    .B(_09301_));
 sg13g2_xnor2_1 _35025_ (.Y(_09303_),
    .A(_05031_),
    .B(_09302_));
 sg13g2_nand2_1 _35026_ (.Y(_09304_),
    .A(net5746),
    .B(_09303_));
 sg13g2_a21oi_1 _35027_ (.A1(net5670),
    .A2(\u_inv.d_next[27] ),
    .Y(_09305_),
    .B1(net4947));
 sg13g2_or2_1 _35028_ (.X(_09306_),
    .B(_09250_),
    .A(_05032_));
 sg13g2_a21oi_1 _35029_ (.A1(_05032_),
    .A2(_09250_),
    .Y(_09307_),
    .B1(net5039));
 sg13g2_a22oi_1 _35030_ (.Y(_09308_),
    .B1(_09306_),
    .B2(_09307_),
    .A2(_09305_),
    .A1(_09304_));
 sg13g2_xnor2_1 _35031_ (.Y(_09309_),
    .A(net4801),
    .B(_09308_));
 sg13g2_xor2_1 _35032_ (.B(_09248_),
    .A(_05029_),
    .X(_09310_));
 sg13g2_nand3_1 _35033_ (.B(_06200_),
    .C(_09260_),
    .A(_05029_),
    .Y(_09311_));
 sg13g2_nand3_1 _35034_ (.B(_09301_),
    .C(_09311_),
    .A(net5746),
    .Y(_09312_));
 sg13g2_a21oi_1 _35035_ (.A1(net5670),
    .A2(\u_inv.d_next[26] ),
    .Y(_09313_),
    .B1(net4947));
 sg13g2_a22oi_1 _35036_ (.Y(_09314_),
    .B1(_09312_),
    .B2(_09313_),
    .A2(_09310_),
    .A1(net4947));
 sg13g2_nand2_1 _35037_ (.Y(_09315_),
    .A(net4744),
    .B(_09314_));
 sg13g2_xnor2_1 _35038_ (.Y(_09316_),
    .A(net4801),
    .B(_09314_));
 sg13g2_xnor2_1 _35039_ (.Y(_09317_),
    .A(net4744),
    .B(_09314_));
 sg13g2_nand2_1 _35040_ (.Y(_09318_),
    .A(_09309_),
    .B(_09316_));
 sg13g2_nand3_1 _35041_ (.B(_05079_),
    .C(_05167_),
    .A(_05045_),
    .Y(_09319_));
 sg13g2_and2_1 _35042_ (.A(net4946),
    .B(_09319_),
    .X(_09320_));
 sg13g2_xnor2_1 _35043_ (.Y(_09321_),
    .A(_05045_),
    .B(_09258_));
 sg13g2_nor2_1 _35044_ (.A(net5744),
    .B(\u_inv.d_next[24] ),
    .Y(_09322_));
 sg13g2_a21oi_1 _35045_ (.A1(net5744),
    .A2(_09321_),
    .Y(_09323_),
    .B1(_09322_));
 sg13g2_a22oi_1 _35046_ (.Y(_09324_),
    .B1(_09323_),
    .B2(net5038),
    .A2(_09320_),
    .A1(_09246_));
 sg13g2_nor2_1 _35047_ (.A(net4799),
    .B(_09324_),
    .Y(_09325_));
 sg13g2_a21oi_1 _35048_ (.A1(\u_inv.d_next[24] ),
    .A2(\u_inv.d_reg[24] ),
    .Y(_09326_),
    .B1(_09259_));
 sg13g2_xnor2_1 _35049_ (.Y(_09327_),
    .A(_05013_),
    .B(_09326_));
 sg13g2_nand2_1 _35050_ (.Y(_09328_),
    .A(net5668),
    .B(\u_inv.d_next[25] ));
 sg13g2_a21oi_1 _35051_ (.A1(net5744),
    .A2(_09327_),
    .Y(_09329_),
    .B1(net4946));
 sg13g2_nand2_1 _35052_ (.Y(_09330_),
    .A(_05014_),
    .B(_09246_));
 sg13g2_o21ai_1 _35053_ (.B1(net4946),
    .Y(_09331_),
    .A1(_05013_),
    .A2(_09330_));
 sg13g2_a21oi_1 _35054_ (.A1(_05013_),
    .A2(_09330_),
    .Y(_09332_),
    .B1(_09331_));
 sg13g2_a21oi_1 _35055_ (.A1(_09328_),
    .A2(_09329_),
    .Y(_09333_),
    .B1(_09332_));
 sg13g2_inv_1 _35056_ (.Y(_09334_),
    .A(_09333_));
 sg13g2_a21oi_1 _35057_ (.A1(_09324_),
    .A2(_09334_),
    .Y(_09335_),
    .B1(net4801));
 sg13g2_nand3_1 _35058_ (.B(_09316_),
    .C(_09335_),
    .A(_09309_),
    .Y(_09336_));
 sg13g2_o21ai_1 _35059_ (.B1(net4744),
    .Y(_09337_),
    .A1(_09308_),
    .A2(_09314_));
 sg13g2_and2_1 _35060_ (.A(_09336_),
    .B(_09337_),
    .X(_09338_));
 sg13g2_o21ai_1 _35061_ (.B1(_09295_),
    .Y(_09339_),
    .A1(_09300_),
    .A2(_09338_));
 sg13g2_a221oi_1 _35062_ (.B2(_09339_),
    .C1(_09269_),
    .B1(_09280_),
    .A1(net4744),
    .Y(_09340_),
    .A2(_09278_));
 sg13g2_xnor2_1 _35063_ (.Y(_09341_),
    .A(net4799),
    .B(_09324_));
 sg13g2_nand2_1 _35064_ (.Y(_09342_),
    .A(net4801),
    .B(_09334_));
 sg13g2_xnor2_1 _35065_ (.Y(_09343_),
    .A(net4744),
    .B(_09333_));
 sg13g2_nor3_1 _35066_ (.A(_09318_),
    .B(_09341_),
    .C(_09343_),
    .Y(_09344_));
 sg13g2_nand3_1 _35067_ (.B(_09299_),
    .C(_09344_),
    .A(_09280_),
    .Y(_09345_));
 sg13g2_nor2_1 _35068_ (.A(_06214_),
    .B(_06219_),
    .Y(_09346_));
 sg13g2_o21ai_1 _35069_ (.B1(_05120_),
    .Y(_09347_),
    .A1(_06214_),
    .A2(_06219_));
 sg13g2_nand2_1 _35070_ (.Y(_09348_),
    .A(_05119_),
    .B(_09347_));
 sg13g2_xnor2_1 _35071_ (.Y(_09349_),
    .A(_06215_),
    .B(_09348_));
 sg13g2_nand2_1 _35072_ (.Y(_09350_),
    .A(net5733),
    .B(_09349_));
 sg13g2_a21oi_1 _35073_ (.A1(net5657),
    .A2(\u_inv.d_next[7] ),
    .Y(_09351_),
    .B1(net4930));
 sg13g2_nor2_1 _35074_ (.A(_05120_),
    .B(_05144_),
    .Y(_09352_));
 sg13g2_nor2_1 _35075_ (.A(_05117_),
    .B(_09352_),
    .Y(_09353_));
 sg13g2_xnor2_1 _35076_ (.Y(_09354_),
    .A(_06216_),
    .B(_09353_));
 sg13g2_a22oi_1 _35077_ (.Y(_09355_),
    .B1(_09354_),
    .B2(net4930),
    .A2(_09351_),
    .A1(_09350_));
 sg13g2_xnor2_1 _35078_ (.Y(_09356_),
    .A(net4793),
    .B(_09355_));
 sg13g2_xnor2_1 _35079_ (.Y(_09357_),
    .A(_05120_),
    .B(_09346_));
 sg13g2_xnor2_1 _35080_ (.Y(_09358_),
    .A(_05120_),
    .B(_05144_));
 sg13g2_nand2_1 _35081_ (.Y(_09359_),
    .A(net5657),
    .B(\u_inv.d_next[6] ));
 sg13g2_a21oi_1 _35082_ (.A1(net5733),
    .A2(_09357_),
    .Y(_09360_),
    .B1(net4930));
 sg13g2_a22oi_1 _35083_ (.Y(_09361_),
    .B1(_09359_),
    .B2(_09360_),
    .A2(_09358_),
    .A1(net4930));
 sg13g2_nand2_1 _35084_ (.Y(_09362_),
    .A(net4793),
    .B(_09361_));
 sg13g2_xnor2_1 _35085_ (.Y(_09363_),
    .A(net4741),
    .B(_09361_));
 sg13g2_nor2b_1 _35086_ (.A(_09356_),
    .B_N(_09363_),
    .Y(_09364_));
 sg13g2_nand3_1 _35087_ (.B(_05142_),
    .C(_06212_),
    .A(_05136_),
    .Y(_09365_));
 sg13g2_o21ai_1 _35088_ (.B1(net5733),
    .Y(_09366_),
    .A1(_05136_),
    .A2(_05142_));
 sg13g2_nor2_1 _35089_ (.A(_06214_),
    .B(_09366_),
    .Y(_09367_));
 sg13g2_xnor2_1 _35090_ (.Y(_09368_),
    .A(_05139_),
    .B(_05142_));
 sg13g2_a221oi_1 _35091_ (.B2(_09367_),
    .C1(net4924),
    .B1(_09365_),
    .A1(net5657),
    .Y(_09369_),
    .A2(\u_inv.d_next[5] ));
 sg13g2_a21o_2 _35092_ (.A2(_09368_),
    .A1(net4924),
    .B1(_09369_),
    .X(_09370_));
 sg13g2_xnor2_1 _35093_ (.Y(_09371_),
    .A(_05135_),
    .B(_05138_));
 sg13g2_nor2_1 _35094_ (.A(_05137_),
    .B(_06211_),
    .Y(_09372_));
 sg13g2_nand2_1 _35095_ (.Y(_09373_),
    .A(net5721),
    .B(_06212_));
 sg13g2_a21oi_1 _35096_ (.A1(net5654),
    .A2(\u_inv.d_next[4] ),
    .Y(_09374_),
    .B1(net4924));
 sg13g2_o21ai_1 _35097_ (.B1(_09374_),
    .Y(_09375_),
    .A1(_09372_),
    .A2(_09373_));
 sg13g2_o21ai_1 _35098_ (.B1(_09375_),
    .Y(_09376_),
    .A1(net5020),
    .A2(_09371_));
 sg13g2_inv_1 _35099_ (.Y(_09377_),
    .A(_09376_));
 sg13g2_a21oi_1 _35100_ (.A1(net4791),
    .A2(_09376_),
    .Y(_09378_),
    .B1(_09370_));
 sg13g2_xnor2_1 _35101_ (.Y(_09379_),
    .A(net4791),
    .B(_09377_));
 sg13g2_xnor2_1 _35102_ (.Y(_09380_),
    .A(_05125_),
    .B(_05134_));
 sg13g2_xnor2_1 _35103_ (.Y(_09381_),
    .A(_05125_),
    .B(_06210_));
 sg13g2_a21oi_1 _35104_ (.A1(net5721),
    .A2(_09381_),
    .Y(_09382_),
    .B1(net4924));
 sg13g2_o21ai_1 _35105_ (.B1(_09382_),
    .Y(_09383_),
    .A1(net5721),
    .A2(\u_inv.d_next[3] ));
 sg13g2_o21ai_1 _35106_ (.B1(_09383_),
    .Y(_09384_),
    .A1(net5020),
    .A2(_09380_));
 sg13g2_a221oi_1 _35107_ (.B2(_06440_),
    .C1(_09384_),
    .B1(_06438_),
    .A1(_05834_),
    .Y(_09385_),
    .A2(_05835_));
 sg13g2_nand2_1 _35108_ (.Y(_09386_),
    .A(net4737),
    .B(_09384_));
 sg13g2_nand3_1 _35109_ (.B(net5349),
    .C(_06461_),
    .A(_06448_),
    .Y(_09387_));
 sg13g2_inv_1 _35110_ (.Y(_09388_),
    .A(_09387_));
 sg13g2_a221oi_1 _35111_ (.B2(_06462_),
    .C1(_06441_),
    .B1(_06452_),
    .A1(_05834_),
    .Y(_09389_),
    .A2(_05835_));
 sg13g2_or2_1 _35112_ (.X(_09390_),
    .B(_09389_),
    .A(_09388_));
 sg13g2_or3_1 _35113_ (.A(_09385_),
    .B(_09388_),
    .C(_09389_),
    .X(_09391_));
 sg13g2_nand2_1 _35114_ (.Y(_09392_),
    .A(_09386_),
    .B(_09391_));
 sg13g2_a21oi_1 _35115_ (.A1(_09386_),
    .A2(_09391_),
    .Y(_09393_),
    .B1(_09379_));
 sg13g2_nand2_1 _35116_ (.Y(_09394_),
    .A(net4737),
    .B(_09370_));
 sg13g2_nand2b_1 _35117_ (.Y(_09395_),
    .B(net4791),
    .A_N(_09370_));
 sg13g2_nand2_1 _35118_ (.Y(_09396_),
    .A(_09394_),
    .B(_09395_));
 sg13g2_a221oi_1 _35119_ (.B2(_09395_),
    .C1(_09379_),
    .B1(_09394_),
    .A1(_09386_),
    .Y(_09397_),
    .A2(_09391_));
 sg13g2_or2_1 _35120_ (.X(_09398_),
    .B(_09397_),
    .A(_09378_));
 sg13g2_o21ai_1 _35121_ (.B1(_09364_),
    .Y(_09399_),
    .A1(_09378_),
    .A2(_09397_));
 sg13g2_o21ai_1 _35122_ (.B1(net4793),
    .Y(_09400_),
    .A1(_09355_),
    .A2(_09361_));
 sg13g2_and2_1 _35123_ (.A(_05151_),
    .B(_06223_),
    .X(_09401_));
 sg13g2_and2_1 _35124_ (.A(_05149_),
    .B(_09401_),
    .X(_09402_));
 sg13g2_or2_1 _35125_ (.X(_09403_),
    .B(_09402_),
    .A(_06232_));
 sg13g2_a21o_1 _35126_ (.A2(_09403_),
    .A1(_05107_),
    .B1(_05106_),
    .X(_09404_));
 sg13g2_a21oi_1 _35127_ (.A1(_05104_),
    .A2(_09404_),
    .Y(_09405_),
    .B1(net5657));
 sg13g2_o21ai_1 _35128_ (.B1(_09405_),
    .Y(_09406_),
    .A1(_05104_),
    .A2(_09404_));
 sg13g2_a21oi_1 _35129_ (.A1(net5657),
    .A2(\u_inv.d_next[11] ),
    .Y(_09407_),
    .B1(net4931));
 sg13g2_nor2_1 _35130_ (.A(_05107_),
    .B(_05153_),
    .Y(_09408_));
 sg13g2_a21oi_1 _35131_ (.A1(\u_inv.d_next[10] ),
    .A2(_14799_),
    .Y(_09409_),
    .B1(_09408_));
 sg13g2_o21ai_1 _35132_ (.B1(net4931),
    .Y(_09410_),
    .A1(_05103_),
    .A2(_09409_));
 sg13g2_a21oi_1 _35133_ (.A1(_05103_),
    .A2(_09409_),
    .Y(_09411_),
    .B1(_09410_));
 sg13g2_a21o_2 _35134_ (.A2(_09407_),
    .A1(_09406_),
    .B1(_09411_),
    .X(_09412_));
 sg13g2_xnor2_1 _35135_ (.Y(_09413_),
    .A(net4793),
    .B(_09412_));
 sg13g2_xnor2_1 _35136_ (.Y(_09414_),
    .A(_05107_),
    .B(_05153_));
 sg13g2_a21oi_1 _35137_ (.A1(_05107_),
    .A2(_09403_),
    .Y(_09415_),
    .B1(net5657));
 sg13g2_o21ai_1 _35138_ (.B1(_09415_),
    .Y(_09416_),
    .A1(_05107_),
    .A2(_09403_));
 sg13g2_a21oi_1 _35139_ (.A1(net5658),
    .A2(\u_inv.d_next[10] ),
    .Y(_09417_),
    .B1(net4931));
 sg13g2_a22oi_1 _35140_ (.Y(_09418_),
    .B1(_09416_),
    .B2(_09417_),
    .A2(_09414_),
    .A1(net4931));
 sg13g2_nand2_1 _35141_ (.Y(_09419_),
    .A(net4741),
    .B(_09418_));
 sg13g2_xnor2_1 _35142_ (.Y(_09420_),
    .A(net4741),
    .B(_09418_));
 sg13g2_nor2_1 _35143_ (.A(_09413_),
    .B(_09420_),
    .Y(_09421_));
 sg13g2_nor3_1 _35144_ (.A(_05122_),
    .B(_05145_),
    .C(_05151_),
    .Y(_09422_));
 sg13g2_xor2_1 _35145_ (.B(_05151_),
    .A(_05147_),
    .X(_09423_));
 sg13g2_nor2_1 _35146_ (.A(net5657),
    .B(_09401_),
    .Y(_09424_));
 sg13g2_o21ai_1 _35147_ (.B1(_09424_),
    .Y(_09425_),
    .A1(_05151_),
    .A2(_06223_));
 sg13g2_a21oi_1 _35148_ (.A1(net5657),
    .A2(\u_inv.d_next[8] ),
    .Y(_09426_),
    .B1(net4930));
 sg13g2_a22oi_1 _35149_ (.Y(_09427_),
    .B1(_09425_),
    .B2(_09426_),
    .A2(_09423_),
    .A1(net4930));
 sg13g2_nand2_1 _35150_ (.Y(_09428_),
    .A(net4793),
    .B(_09427_));
 sg13g2_xnor2_1 _35151_ (.Y(_09429_),
    .A(net4793),
    .B(_09427_));
 sg13g2_nand2_1 _35152_ (.Y(_09430_),
    .A(_05148_),
    .B(_05150_));
 sg13g2_o21ai_1 _35153_ (.B1(net5733),
    .Y(_09431_),
    .A1(_05148_),
    .A2(_05150_));
 sg13g2_nor2_1 _35154_ (.A(_09402_),
    .B(_09431_),
    .Y(_09432_));
 sg13g2_o21ai_1 _35155_ (.B1(_09432_),
    .Y(_09433_),
    .A1(_09401_),
    .A2(_09430_));
 sg13g2_a21oi_1 _35156_ (.A1(net5658),
    .A2(\u_inv.d_next[9] ),
    .Y(_09434_),
    .B1(net4930));
 sg13g2_nor2_1 _35157_ (.A(_05112_),
    .B(_09422_),
    .Y(_09435_));
 sg13g2_o21ai_1 _35158_ (.B1(net4930),
    .Y(_09436_),
    .A1(_05148_),
    .A2(_09435_));
 sg13g2_a21oi_1 _35159_ (.A1(_05148_),
    .A2(_09435_),
    .Y(_09437_),
    .B1(_09436_));
 sg13g2_a21oi_2 _35160_ (.B1(_09437_),
    .Y(_09438_),
    .A2(_09434_),
    .A1(_09433_));
 sg13g2_nand2_1 _35161_ (.Y(_09439_),
    .A(net4794),
    .B(_09438_));
 sg13g2_nor2_1 _35162_ (.A(net4793),
    .B(_09438_),
    .Y(_09440_));
 sg13g2_xnor2_1 _35163_ (.Y(_09441_),
    .A(net4793),
    .B(_09438_));
 sg13g2_or4_1 _35164_ (.A(_09413_),
    .B(_09420_),
    .C(_09429_),
    .D(_09441_),
    .X(_09442_));
 sg13g2_a21oi_2 _35165_ (.B1(_09442_),
    .Y(_09443_),
    .A2(_09400_),
    .A1(_09399_));
 sg13g2_a21o_1 _35166_ (.A2(_05154_),
    .A1(_05108_),
    .B1(_05099_),
    .X(_09444_));
 sg13g2_a21o_1 _35167_ (.A2(_09444_),
    .A1(_05095_),
    .B1(_05090_),
    .X(_09445_));
 sg13g2_o21ai_1 _35168_ (.B1(_05086_),
    .Y(_09446_),
    .A1(_05091_),
    .A2(_09445_));
 sg13g2_and2_1 _35169_ (.A(_05080_),
    .B(_09446_),
    .X(_09447_));
 sg13g2_o21ai_1 _35170_ (.B1(net4933),
    .Y(_09448_),
    .A1(_05082_),
    .A2(_09447_));
 sg13g2_a21oi_1 _35171_ (.A1(_05082_),
    .A2(_09447_),
    .Y(_09449_),
    .B1(_09448_));
 sg13g2_a21oi_2 _35172_ (.B1(_06234_),
    .Y(_09450_),
    .A2(_09402_),
    .A1(_06226_));
 sg13g2_o21ai_1 _35173_ (.B1(_06237_),
    .Y(_09451_),
    .A1(_06224_),
    .A2(_09450_));
 sg13g2_nand2_1 _35174_ (.Y(_09452_),
    .A(_05085_),
    .B(_09451_));
 sg13g2_nand3_1 _35175_ (.B(_05083_),
    .C(_09452_),
    .A(_05082_),
    .Y(_09453_));
 sg13g2_a21oi_1 _35176_ (.A1(_05083_),
    .A2(_09452_),
    .Y(_09454_),
    .B1(_05082_));
 sg13g2_nor2_1 _35177_ (.A(net5661),
    .B(_09454_),
    .Y(_09455_));
 sg13g2_a221oi_1 _35178_ (.B2(_09455_),
    .C1(net4933),
    .B1(_09453_),
    .A1(net5661),
    .Y(_09456_),
    .A2(\u_inv.d_next[15] ));
 sg13g2_or2_1 _35179_ (.X(_09457_),
    .B(_09456_),
    .A(_09449_));
 sg13g2_xnor2_1 _35180_ (.Y(_09458_),
    .A(net4740),
    .B(_09457_));
 sg13g2_or3_1 _35181_ (.A(_05086_),
    .B(_05091_),
    .C(_09445_),
    .X(_09459_));
 sg13g2_nand2_1 _35182_ (.Y(_09460_),
    .A(_09446_),
    .B(_09459_));
 sg13g2_xnor2_1 _35183_ (.Y(_09461_),
    .A(_05086_),
    .B(_09451_));
 sg13g2_nand2_1 _35184_ (.Y(_09462_),
    .A(net5661),
    .B(\u_inv.d_next[14] ));
 sg13g2_a21oi_1 _35185_ (.A1(net5731),
    .A2(_09461_),
    .Y(_09463_),
    .B1(net4933));
 sg13g2_a22oi_1 _35186_ (.Y(_09464_),
    .B1(_09462_),
    .B2(_09463_),
    .A2(_09460_),
    .A1(net4933));
 sg13g2_nand2_1 _35187_ (.Y(_09465_),
    .A(net4740),
    .B(_09464_));
 sg13g2_xnor2_1 _35188_ (.Y(_09466_),
    .A(net4795),
    .B(_09464_));
 sg13g2_and2_1 _35189_ (.A(_09458_),
    .B(_09466_),
    .X(_09467_));
 sg13g2_or2_1 _35190_ (.X(_09468_),
    .B(_09444_),
    .A(_05094_));
 sg13g2_a21oi_1 _35191_ (.A1(_05094_),
    .A2(_09444_),
    .Y(_09469_),
    .B1(net5030));
 sg13g2_xnor2_1 _35192_ (.Y(_09470_),
    .A(_05094_),
    .B(_09450_));
 sg13g2_nor2_1 _35193_ (.A(net5733),
    .B(\u_inv.d_next[12] ),
    .Y(_09471_));
 sg13g2_a21oi_1 _35194_ (.A1(net5731),
    .A2(_09470_),
    .Y(_09472_),
    .B1(_09471_));
 sg13g2_a22oi_1 _35195_ (.Y(_09473_),
    .B1(_09472_),
    .B2(net5030),
    .A2(_09469_),
    .A1(_09468_));
 sg13g2_or2_1 _35196_ (.X(_09474_),
    .B(_09473_),
    .A(net4794));
 sg13g2_xnor2_1 _35197_ (.Y(_09475_),
    .A(net4741),
    .B(_09473_));
 sg13g2_and2_1 _35198_ (.A(_05088_),
    .B(_05089_),
    .X(_09476_));
 sg13g2_o21ai_1 _35199_ (.B1(_05092_),
    .Y(_09477_),
    .A1(_05094_),
    .A2(_09450_));
 sg13g2_or2_1 _35200_ (.X(_09478_),
    .B(_09477_),
    .A(_05088_));
 sg13g2_a21oi_1 _35201_ (.A1(_05088_),
    .A2(_09477_),
    .Y(_09479_),
    .B1(net5661));
 sg13g2_a221oi_1 _35202_ (.B2(_09479_),
    .C1(net4933),
    .B1(_09478_),
    .A1(net5661),
    .Y(_09480_),
    .A2(\u_inv.d_next[13] ));
 sg13g2_a221oi_1 _35203_ (.B2(_09476_),
    .C1(_09480_),
    .B1(_09469_),
    .A1(net4933),
    .Y(_09481_),
    .A2(_09445_));
 sg13g2_nand2_1 _35204_ (.Y(_09482_),
    .A(net4740),
    .B(_09481_));
 sg13g2_nand2b_1 _35205_ (.Y(_09483_),
    .B(net4795),
    .A_N(_09481_));
 sg13g2_and2_1 _35206_ (.A(_09482_),
    .B(_09483_),
    .X(_09484_));
 sg13g2_and2_1 _35207_ (.A(_09475_),
    .B(_09484_),
    .X(_09485_));
 sg13g2_and2_1 _35208_ (.A(_09467_),
    .B(_09485_),
    .X(_09486_));
 sg13g2_and2_1 _35209_ (.A(_09474_),
    .B(_09482_),
    .X(_09487_));
 sg13g2_inv_1 _35210_ (.Y(_09488_),
    .A(_09487_));
 sg13g2_nand2_1 _35211_ (.Y(_09489_),
    .A(_09428_),
    .B(_09439_));
 sg13g2_o21ai_1 _35212_ (.B1(_09419_),
    .Y(_09490_),
    .A1(net4794),
    .A2(_09412_));
 sg13g2_a21o_2 _35213_ (.A2(_09489_),
    .A1(_09421_),
    .B1(_09490_),
    .X(_09491_));
 sg13g2_a21o_1 _35214_ (.A2(_09491_),
    .A1(_09485_),
    .B1(_09488_),
    .X(_09492_));
 sg13g2_o21ai_1 _35215_ (.B1(_09465_),
    .Y(_09493_),
    .A1(net4795),
    .A2(_09457_));
 sg13g2_a221oi_1 _35216_ (.B2(_09467_),
    .C1(_09493_),
    .B1(_09492_),
    .A1(_09443_),
    .Y(_09494_),
    .A2(_09486_));
 sg13g2_nand2_1 _35217_ (.Y(_09495_),
    .A(_06184_),
    .B(_09255_));
 sg13g2_a21oi_1 _35218_ (.A1(_06184_),
    .A2(_09255_),
    .Y(_09496_),
    .B1(_05062_));
 sg13g2_xor2_1 _35219_ (.B(_09495_),
    .A(_05062_),
    .X(_09497_));
 sg13g2_o21ai_1 _35220_ (.B1(net5029),
    .Y(_09498_),
    .A1(net5731),
    .A2(\u_inv.d_next[18] ));
 sg13g2_a21oi_1 _35221_ (.A1(net5731),
    .A2(_09497_),
    .Y(_09499_),
    .B1(_09498_));
 sg13g2_a21oi_1 _35222_ (.A1(_05157_),
    .A2(_05159_),
    .Y(_09500_),
    .B1(_05165_));
 sg13g2_or2_1 _35223_ (.X(_09501_),
    .B(_09500_),
    .A(_05067_));
 sg13g2_nand2_1 _35224_ (.Y(_09502_),
    .A(_05062_),
    .B(_09501_));
 sg13g2_xor2_1 _35225_ (.B(_09501_),
    .A(_05062_),
    .X(_09503_));
 sg13g2_a21oi_2 _35226_ (.B1(_09499_),
    .Y(_09504_),
    .A2(_09503_),
    .A1(net4933));
 sg13g2_nor2_1 _35227_ (.A(net4795),
    .B(_09504_),
    .Y(_09505_));
 sg13g2_xnor2_1 _35228_ (.Y(_09506_),
    .A(net4795),
    .B(_09504_));
 sg13g2_nand2_1 _35229_ (.Y(_09507_),
    .A(_05068_),
    .B(_09502_));
 sg13g2_o21ai_1 _35230_ (.B1(net4933),
    .Y(_09508_),
    .A1(_05061_),
    .A2(_09507_));
 sg13g2_a21oi_1 _35231_ (.A1(_05061_),
    .A2(_09507_),
    .Y(_09509_),
    .B1(_09508_));
 sg13g2_a21oi_1 _35232_ (.A1(\u_inv.d_next[18] ),
    .A2(\u_inv.d_reg[18] ),
    .Y(_09510_),
    .B1(_09496_));
 sg13g2_xnor2_1 _35233_ (.Y(_09511_),
    .A(_05061_),
    .B(_09510_));
 sg13g2_nand2_1 _35234_ (.Y(_09512_),
    .A(net5731),
    .B(_09511_));
 sg13g2_a21oi_1 _35235_ (.A1(net5661),
    .A2(\u_inv.d_next[19] ),
    .Y(_09513_),
    .B1(net4934));
 sg13g2_a21o_1 _35236_ (.A2(_09513_),
    .A1(_09512_),
    .B1(_09509_),
    .X(_09514_));
 sg13g2_xnor2_1 _35237_ (.Y(_09515_),
    .A(net4795),
    .B(_09514_));
 sg13g2_nand3_1 _35238_ (.B(_05162_),
    .C(_09254_),
    .A(_05161_),
    .Y(_09516_));
 sg13g2_nor2_1 _35239_ (.A(net5661),
    .B(_06182_),
    .Y(_09517_));
 sg13g2_nand3_1 _35240_ (.B(_09516_),
    .C(_09517_),
    .A(_09255_),
    .Y(_09518_));
 sg13g2_a21oi_1 _35241_ (.A1(net5661),
    .A2(\u_inv.d_next[17] ),
    .Y(_09519_),
    .B1(net4934));
 sg13g2_nor2_1 _35242_ (.A(_05160_),
    .B(_05163_),
    .Y(_09520_));
 sg13g2_nor2_1 _35243_ (.A(_05065_),
    .B(_09520_),
    .Y(_09521_));
 sg13g2_o21ai_1 _35244_ (.B1(net4934),
    .Y(_09522_),
    .A1(_05161_),
    .A2(_09521_));
 sg13g2_a21oi_1 _35245_ (.A1(_05161_),
    .A2(_09521_),
    .Y(_09523_),
    .B1(_09522_));
 sg13g2_a21oi_2 _35246_ (.B1(_09523_),
    .Y(_09524_),
    .A2(_09519_),
    .A1(_09518_));
 sg13g2_nor2_1 _35247_ (.A(net4740),
    .B(_09524_),
    .Y(_09525_));
 sg13g2_xnor2_1 _35248_ (.Y(_09526_),
    .A(net4795),
    .B(_09524_));
 sg13g2_xnor2_1 _35249_ (.Y(_09527_),
    .A(_05164_),
    .B(_06242_));
 sg13g2_a21oi_1 _35250_ (.A1(net5731),
    .A2(_09527_),
    .Y(_09528_),
    .B1(net4934));
 sg13g2_o21ai_1 _35251_ (.B1(_09528_),
    .Y(_09529_),
    .A1(net5731),
    .A2(\u_inv.d_next[16] ));
 sg13g2_a21o_1 _35252_ (.A2(_05163_),
    .A1(_05160_),
    .B1(net5029),
    .X(_09530_));
 sg13g2_o21ai_1 _35253_ (.B1(_09529_),
    .Y(_09531_),
    .A1(_09520_),
    .A2(_09530_));
 sg13g2_nand2_1 _35254_ (.Y(_09532_),
    .A(net4740),
    .B(_09531_));
 sg13g2_xnor2_1 _35255_ (.Y(_09533_),
    .A(net4796),
    .B(_09531_));
 sg13g2_nand2_1 _35256_ (.Y(_09534_),
    .A(_09526_),
    .B(_09533_));
 sg13g2_nor3_1 _35257_ (.A(_09506_),
    .B(_09515_),
    .C(_09534_),
    .Y(_09535_));
 sg13g2_xnor2_1 _35258_ (.Y(_09536_),
    .A(_05056_),
    .B(_09257_));
 sg13g2_o21ai_1 _35259_ (.B1(net5038),
    .Y(_09537_),
    .A1(net5744),
    .A2(\u_inv.d_next[20] ));
 sg13g2_a21o_1 _35260_ (.A2(_09536_),
    .A1(net5744),
    .B1(_09537_),
    .X(_09538_));
 sg13g2_a21oi_1 _35261_ (.A1(_05063_),
    .A2(_09501_),
    .Y(_09539_),
    .B1(_05069_));
 sg13g2_nor2_1 _35262_ (.A(_05056_),
    .B(_09539_),
    .Y(_09540_));
 sg13g2_a21o_1 _35263_ (.A2(_09539_),
    .A1(_05056_),
    .B1(net5038),
    .X(_09541_));
 sg13g2_o21ai_1 _35264_ (.B1(_09538_),
    .Y(_09542_),
    .A1(_09540_),
    .A2(_09541_));
 sg13g2_nand2_1 _35265_ (.Y(_09543_),
    .A(net4743),
    .B(_09542_));
 sg13g2_xnor2_1 _35266_ (.Y(_09544_),
    .A(net4743),
    .B(_09542_));
 sg13g2_a21oi_1 _35267_ (.A1(_05056_),
    .A2(_09257_),
    .Y(_09545_),
    .B1(_05055_));
 sg13g2_xnor2_1 _35268_ (.Y(_09546_),
    .A(_05054_),
    .B(_09545_));
 sg13g2_o21ai_1 _35269_ (.B1(net5038),
    .Y(_09547_),
    .A1(net5744),
    .A2(_14237_));
 sg13g2_a21oi_1 _35270_ (.A1(net5744),
    .A2(_09546_),
    .Y(_09548_),
    .B1(_09547_));
 sg13g2_nor2_1 _35271_ (.A(_05075_),
    .B(_09540_),
    .Y(_09549_));
 sg13g2_a21oi_1 _35272_ (.A1(_05053_),
    .A2(_09549_),
    .Y(_09550_),
    .B1(net5038));
 sg13g2_o21ai_1 _35273_ (.B1(_09550_),
    .Y(_09551_),
    .A1(_05053_),
    .A2(_09549_));
 sg13g2_nand2b_2 _35274_ (.Y(_09552_),
    .B(_09551_),
    .A_N(_09548_));
 sg13g2_inv_1 _35275_ (.Y(_09553_),
    .A(_09552_));
 sg13g2_nand2_1 _35276_ (.Y(_09554_),
    .A(net4799),
    .B(_09552_));
 sg13g2_xnor2_1 _35277_ (.Y(_09555_),
    .A(net4743),
    .B(_09552_));
 sg13g2_nor2b_1 _35278_ (.A(_09544_),
    .B_N(_09555_),
    .Y(_09556_));
 sg13g2_o21ai_1 _35279_ (.B1(_05076_),
    .Y(_09557_),
    .A1(_05057_),
    .A2(_09539_));
 sg13g2_nand2_1 _35280_ (.Y(_09558_),
    .A(_05051_),
    .B(_09557_));
 sg13g2_xor2_1 _35281_ (.B(_09557_),
    .A(_05051_),
    .X(_09559_));
 sg13g2_a21oi_1 _35282_ (.A1(_06180_),
    .A2(_09257_),
    .Y(_09560_),
    .B1(_06190_));
 sg13g2_and2_1 _35283_ (.A(_05051_),
    .B(_09560_),
    .X(_09561_));
 sg13g2_or2_1 _35284_ (.X(_09562_),
    .B(_09560_),
    .A(_05051_));
 sg13g2_nand2_1 _35285_ (.Y(_09563_),
    .A(net5744),
    .B(_09562_));
 sg13g2_a21oi_1 _35286_ (.A1(net5668),
    .A2(\u_inv.d_next[22] ),
    .Y(_09564_),
    .B1(net4946));
 sg13g2_o21ai_1 _35287_ (.B1(_09564_),
    .Y(_09565_),
    .A1(_09561_),
    .A2(_09563_));
 sg13g2_o21ai_1 _35288_ (.B1(_09565_),
    .Y(_09566_),
    .A1(net5038),
    .A2(_09559_));
 sg13g2_nor2_1 _35289_ (.A(net4799),
    .B(_09566_),
    .Y(_09567_));
 sg13g2_and2_1 _35290_ (.A(net4799),
    .B(_09566_),
    .X(_09568_));
 sg13g2_nor2_1 _35291_ (.A(_09567_),
    .B(_09568_),
    .Y(_09569_));
 sg13g2_nand2_1 _35292_ (.Y(_09570_),
    .A(_05071_),
    .B(_09558_));
 sg13g2_o21ai_1 _35293_ (.B1(net4946),
    .Y(_09571_),
    .A1(_05048_),
    .A2(_09570_));
 sg13g2_a21oi_1 _35294_ (.A1(_05048_),
    .A2(_09570_),
    .Y(_09572_),
    .B1(_09571_));
 sg13g2_nand2_1 _35295_ (.Y(_09573_),
    .A(_05049_),
    .B(_09562_));
 sg13g2_xnor2_1 _35296_ (.Y(_09574_),
    .A(_05047_),
    .B(_09573_));
 sg13g2_nand2_1 _35297_ (.Y(_09575_),
    .A(net5668),
    .B(\u_inv.d_next[23] ));
 sg13g2_a21oi_1 _35298_ (.A1(net5745),
    .A2(_09574_),
    .Y(_09576_),
    .B1(net4946));
 sg13g2_a21o_2 _35299_ (.A2(_09576_),
    .A1(_09575_),
    .B1(_09572_),
    .X(_09577_));
 sg13g2_xnor2_1 _35300_ (.Y(_09578_),
    .A(net4799),
    .B(_09577_));
 sg13g2_nor3_2 _35301_ (.A(_09567_),
    .B(_09568_),
    .C(_09578_),
    .Y(_09579_));
 sg13g2_nand3_1 _35302_ (.B(_09556_),
    .C(_09579_),
    .A(_09535_),
    .Y(_09580_));
 sg13g2_or2_1 _35303_ (.X(_09581_),
    .B(_09580_),
    .A(_09494_));
 sg13g2_o21ai_1 _35304_ (.B1(net4743),
    .Y(_09582_),
    .A1(_09542_),
    .A2(_09553_));
 sg13g2_o21ai_1 _35305_ (.B1(net4740),
    .Y(_09583_),
    .A1(_09524_),
    .A2(_09531_));
 sg13g2_nor3_1 _35306_ (.A(_09506_),
    .B(_09515_),
    .C(_09583_),
    .Y(_09584_));
 sg13g2_a21oi_1 _35307_ (.A1(_09504_),
    .A2(_09514_),
    .Y(_09585_),
    .B1(net4795));
 sg13g2_o21ai_1 _35308_ (.B1(_09556_),
    .Y(_09586_),
    .A1(_09584_),
    .A2(_09585_));
 sg13g2_nand2_1 _35309_ (.Y(_09587_),
    .A(_09582_),
    .B(_09586_));
 sg13g2_a21oi_1 _35310_ (.A1(_09566_),
    .A2(_09577_),
    .Y(_09588_),
    .B1(net4799));
 sg13g2_a21oi_2 _35311_ (.B1(_09588_),
    .Y(_09589_),
    .A2(_09587_),
    .A1(_09579_));
 sg13g2_and2_1 _35312_ (.A(_09340_),
    .B(_09589_),
    .X(_09590_));
 sg13g2_a22oi_1 _35313_ (.Y(_09591_),
    .B1(_09581_),
    .B2(_09590_),
    .A2(_09345_),
    .A1(_09340_));
 sg13g2_xnor2_1 _35314_ (.Y(_09592_),
    .A(net4803),
    .B(_09127_));
 sg13g2_xnor2_1 _35315_ (.Y(_09593_),
    .A(net4748),
    .B(_09132_));
 sg13g2_nor2_1 _35316_ (.A(_09592_),
    .B(_09593_),
    .Y(_09594_));
 sg13g2_nand2_1 _35317_ (.Y(_09595_),
    .A(_09101_),
    .B(_09594_));
 sg13g2_nor3_1 _35318_ (.A(_09080_),
    .B(_09119_),
    .C(_09595_),
    .Y(_09596_));
 sg13g2_inv_1 _35319_ (.Y(_09597_),
    .A(_09596_));
 sg13g2_nor2b_1 _35320_ (.A(_09228_),
    .B_N(_09596_),
    .Y(_09598_));
 sg13g2_inv_1 _35321_ (.Y(_09599_),
    .A(_09598_));
 sg13g2_nand2_1 _35322_ (.Y(_09600_),
    .A(_09244_),
    .B(_09598_));
 sg13g2_a221oi_1 _35323_ (.B2(_09590_),
    .C1(_09600_),
    .B1(_09581_),
    .A1(_09340_),
    .Y(_09601_),
    .A2(_09345_));
 sg13g2_nor2_2 _35324_ (.A(_09245_),
    .B(net1064),
    .Y(_09602_));
 sg13g2_nand2_1 _35325_ (.Y(_09603_),
    .A(net4820),
    .B(_08811_));
 sg13g2_xnor2_1 _35326_ (.Y(_09604_),
    .A(net4820),
    .B(_08810_));
 sg13g2_inv_1 _35327_ (.Y(_09605_),
    .A(_09604_));
 sg13g2_xnor2_1 _35328_ (.Y(_09606_),
    .A(net4772),
    .B(_08816_));
 sg13g2_nor3_1 _35329_ (.A(_08802_),
    .B(_09605_),
    .C(_09606_),
    .Y(_09607_));
 sg13g2_and2_1 _35330_ (.A(_08783_),
    .B(_09607_),
    .X(_09608_));
 sg13g2_nor2b_1 _35331_ (.A(_08736_),
    .B_N(_09608_),
    .Y(_09609_));
 sg13g2_and2_1 _35332_ (.A(_08646_),
    .B(_09609_),
    .X(_09610_));
 sg13g2_o21ai_1 _35333_ (.B1(_09610_),
    .Y(_09611_),
    .A1(_09245_),
    .A2(net1064));
 sg13g2_nand2_1 _35334_ (.Y(_09612_),
    .A(_08851_),
    .B(_09611_));
 sg13g2_a21o_2 _35335_ (.A2(_09611_),
    .A1(_08851_),
    .B1(_08455_),
    .X(_09613_));
 sg13g2_o21ai_1 _35336_ (.B1(net4780),
    .Y(_09614_),
    .A1(_08438_),
    .A2(_08448_));
 sg13g2_a21oi_1 _35337_ (.A1(net4780),
    .A2(_08420_),
    .Y(_09615_),
    .B1(_08429_));
 sg13g2_nor2b_1 _35338_ (.A(_09615_),
    .B_N(_08411_),
    .Y(_09616_));
 sg13g2_a21oi_1 _35339_ (.A1(_08397_),
    .A2(_08409_),
    .Y(_09617_),
    .B1(net4827));
 sg13g2_or2_1 _35340_ (.X(_09618_),
    .B(_09617_),
    .A(_09616_));
 sg13g2_o21ai_1 _35341_ (.B1(_08451_),
    .Y(_09619_),
    .A1(_09616_),
    .A2(_09617_));
 sg13g2_a21oi_1 _35342_ (.A1(_09614_),
    .A2(_09619_),
    .Y(_09620_),
    .B1(_08388_));
 sg13g2_o21ai_1 _35343_ (.B1(_08376_),
    .Y(_09621_),
    .A1(net4823),
    .A2(_08386_));
 sg13g2_or2_1 _35344_ (.X(_09622_),
    .B(_09621_),
    .A(_09620_));
 sg13g2_o21ai_1 _35345_ (.B1(_08364_),
    .Y(_09623_),
    .A1(_09620_),
    .A2(_09621_));
 sg13g2_nor2_1 _35346_ (.A(_08350_),
    .B(_08360_),
    .Y(_09624_));
 sg13g2_o21ai_1 _35347_ (.B1(net4779),
    .Y(_09625_),
    .A1(_08333_),
    .A2(_08340_));
 sg13g2_o21ai_1 _35348_ (.B1(_09625_),
    .Y(_09626_),
    .A1(_08344_),
    .A2(_09624_));
 sg13g2_inv_1 _35349_ (.Y(_09627_),
    .A(_09626_));
 sg13g2_nand4_1 _35350_ (.B(_08314_),
    .C(_08322_),
    .A(_08304_),
    .Y(_09628_),
    .D(_09626_));
 sg13g2_a21o_1 _35351_ (.A2(_08313_),
    .A1(net4781),
    .B1(_08321_),
    .X(_09629_));
 sg13g2_a22oi_1 _35352_ (.Y(_09630_),
    .B1(_08304_),
    .B2(_09629_),
    .A2(_08302_),
    .A1(net4781));
 sg13g2_nand4_1 _35353_ (.B(_09623_),
    .C(_09628_),
    .A(_08292_),
    .Y(_09631_),
    .D(_09630_));
 sg13g2_o21ai_1 _35354_ (.B1(net4774),
    .Y(_09632_),
    .A1(_08263_),
    .A2(_08270_));
 sg13g2_nand3b_1 _35355_ (.B(_08254_),
    .C(_08246_),
    .Y(_09633_),
    .A_N(_09632_));
 sg13g2_nand2b_1 _35356_ (.Y(_09634_),
    .B(_09633_),
    .A_N(_08253_));
 sg13g2_a21oi_1 _35357_ (.A1(net4774),
    .A2(_08245_),
    .Y(_09635_),
    .B1(_09634_));
 sg13g2_or4_1 _35358_ (.A(_08218_),
    .B(_08228_),
    .C(_08235_),
    .D(_09635_),
    .X(_09636_));
 sg13g2_a21o_1 _35359_ (.A2(_08226_),
    .A1(net4773),
    .B1(_08234_),
    .X(_09637_));
 sg13g2_nand2b_1 _35360_ (.Y(_09638_),
    .B(_09637_),
    .A_N(_08218_));
 sg13g2_nand4_1 _35361_ (.B(_08215_),
    .C(_09636_),
    .A(_08206_),
    .Y(_09639_),
    .D(_09638_));
 sg13g2_inv_2 _35362_ (.Y(_09640_),
    .A(_09639_));
 sg13g2_o21ai_1 _35363_ (.B1(_08182_),
    .Y(_09641_),
    .A1(net4822),
    .A2(_08175_));
 sg13g2_nand3_1 _35364_ (.B(_08166_),
    .C(_09641_),
    .A(_08156_),
    .Y(_09642_));
 sg13g2_nand3_1 _35365_ (.B(_08165_),
    .C(_09642_),
    .A(_08154_),
    .Y(_09643_));
 sg13g2_nand4_1 _35366_ (.B(_08128_),
    .C(_08146_),
    .A(_08119_),
    .Y(_09644_),
    .D(_09643_));
 sg13g2_a21oi_1 _35367_ (.A1(net4771),
    .A2(_08127_),
    .Y(_09645_),
    .B1(_08117_));
 sg13g2_a21oi_1 _35368_ (.A1(net4771),
    .A2(_08137_),
    .Y(_09646_),
    .B1(_08144_));
 sg13g2_nand3b_1 _35369_ (.B(_08128_),
    .C(_08119_),
    .Y(_09647_),
    .A_N(_09646_));
 sg13g2_nand3_1 _35370_ (.B(_09645_),
    .C(_09647_),
    .A(_09644_),
    .Y(_09648_));
 sg13g2_a221oi_1 _35371_ (.B2(_08186_),
    .C1(_09648_),
    .B1(_09639_),
    .A1(_08275_),
    .Y(_09649_),
    .A2(_09631_));
 sg13g2_xnor2_1 _35372_ (.Y(_09650_),
    .A(net4820),
    .B(_07653_));
 sg13g2_xnor2_1 _35373_ (.Y(_09651_),
    .A(net4772),
    .B(_07659_));
 sg13g2_nor3_1 _35374_ (.A(_07645_),
    .B(_09650_),
    .C(_09651_),
    .Y(_09652_));
 sg13g2_inv_1 _35375_ (.Y(_09653_),
    .A(_09652_));
 sg13g2_nand2_1 _35376_ (.Y(_09654_),
    .A(_07623_),
    .B(_09652_));
 sg13g2_or4_1 _35377_ (.A(_07507_),
    .B(_07527_),
    .C(_07567_),
    .D(_09654_),
    .X(_09655_));
 sg13g2_or3_1 _35378_ (.A(_07386_),
    .B(_07680_),
    .C(_09655_),
    .X(_09656_));
 sg13g2_a21oi_2 _35379_ (.B1(_09656_),
    .Y(_09657_),
    .A2(_09649_),
    .A1(_09613_));
 sg13g2_a21o_2 _35380_ (.A2(_09649_),
    .A1(_09613_),
    .B1(_09656_),
    .X(_09658_));
 sg13g2_a221oi_1 _35381_ (.B2(_09657_),
    .C1(_08082_),
    .B1(_08085_),
    .A1(_07683_),
    .Y(_09659_),
    .A2(_08045_));
 sg13g2_o21ai_1 _35382_ (.B1(_08087_),
    .Y(_09660_),
    .A1(_08086_),
    .A2(_09658_));
 sg13g2_a21o_2 _35383_ (.A2(_09660_),
    .A1(_07281_),
    .B1(_07271_),
    .X(_09661_));
 sg13g2_xnor2_1 _35384_ (.Y(_09662_),
    .A(_04449_),
    .B(_06437_));
 sg13g2_a21oi_1 _35385_ (.A1(net5720),
    .A2(_09662_),
    .Y(_09663_),
    .B1(_06439_));
 sg13g2_or3_1 _35386_ (.A(_04448_),
    .B(_05704_),
    .C(_05833_),
    .X(_09664_));
 sg13g2_nand3_1 _35387_ (.B(_05834_),
    .C(_09664_),
    .A(net4924),
    .Y(_09665_));
 sg13g2_nand2b_2 _35388_ (.Y(_09666_),
    .B(_09665_),
    .A_N(_09663_));
 sg13g2_inv_1 _35389_ (.Y(_09667_),
    .A(_09666_));
 sg13g2_xnor2_1 _35390_ (.Y(_09668_),
    .A(net4737),
    .B(_09666_));
 sg13g2_and3_2 _35391_ (.X(_09669_),
    .A(net5390),
    .B(_09661_),
    .C(_09668_));
 sg13g2_nand3_1 _35392_ (.B(net5391),
    .C(_09668_),
    .A(_09661_),
    .Y(_09670_));
 sg13g2_o21ai_1 _35393_ (.B1(net4791),
    .Y(_09671_),
    .A1(net5349),
    .A2(_09666_));
 sg13g2_a21oi_2 _35394_ (.B1(net4737),
    .Y(_09672_),
    .A2(_09667_),
    .A1(net5390));
 sg13g2_nor2_2 _35395_ (.A(net4634),
    .B(net4635),
    .Y(_09673_));
 sg13g2_nand2_1 _35396_ (.Y(_09674_),
    .A(net4629),
    .B(net4637));
 sg13g2_nor3_1 _35397_ (.A(_06464_),
    .B(net4634),
    .C(net4635),
    .Y(_09675_));
 sg13g2_o21ai_1 _35398_ (.B1(_06464_),
    .Y(_09676_),
    .A1(net4634),
    .A2(net4635));
 sg13g2_nand2b_2 _35399_ (.Y(_09677_),
    .B(_09676_),
    .A_N(_09675_));
 sg13g2_a21o_1 _35400_ (.A2(_09677_),
    .A1(_19007_),
    .B1(net4451),
    .X(_09678_));
 sg13g2_a21oi_2 _35401_ (.B1(_06466_),
    .Y(_09679_),
    .A2(_09678_),
    .A1(net4691));
 sg13g2_a22oi_1 _35402_ (.Y(_00774_),
    .B1(_09679_),
    .B2(net5590),
    .A2(net4126),
    .A1(_14242_));
 sg13g2_nor2b_1 _35403_ (.A(_09385_),
    .B_N(_09386_),
    .Y(_09680_));
 sg13g2_xnor2_1 _35404_ (.Y(_09681_),
    .A(_09390_),
    .B(_09680_));
 sg13g2_mux2_1 _35405_ (.A0(_09384_),
    .A1(_09681_),
    .S(net5391),
    .X(_09682_));
 sg13g2_inv_1 _35406_ (.Y(_09683_),
    .A(_09682_));
 sg13g2_nor3_1 _35407_ (.A(net4646),
    .B(_06461_),
    .C(net4580),
    .Y(_09684_));
 sg13g2_xnor2_1 _35408_ (.Y(_09685_),
    .A(_09682_),
    .B(_09684_));
 sg13g2_o21ai_1 _35409_ (.B1(net5590),
    .Y(_09686_),
    .A1(net4384),
    .A2(_06463_));
 sg13g2_a21oi_1 _35410_ (.A1(net4384),
    .A2(_09685_),
    .Y(_09687_),
    .B1(_09686_));
 sg13g2_a21o_1 _35411_ (.A2(net4125),
    .A1(net2398),
    .B1(_09687_),
    .X(_00775_));
 sg13g2_xnor2_1 _35412_ (.Y(_09688_),
    .A(_09379_),
    .B(_09392_));
 sg13g2_nand2_1 _35413_ (.Y(_09689_),
    .A(net5390),
    .B(_09688_));
 sg13g2_o21ai_1 _35414_ (.B1(_09689_),
    .Y(_09690_),
    .A1(net5390),
    .A2(_09376_));
 sg13g2_nand3_1 _35415_ (.B(net4636),
    .C(_09690_),
    .A(net4628),
    .Y(_09691_));
 sg13g2_a21o_1 _35416_ (.A2(net4636),
    .A1(net4628),
    .B1(_09690_),
    .X(_09692_));
 sg13g2_nand2_1 _35417_ (.Y(_09693_),
    .A(_09691_),
    .B(_09692_));
 sg13g2_o21ai_1 _35418_ (.B1(_09683_),
    .Y(_09694_),
    .A1(net4634),
    .A2(net4635));
 sg13g2_nor2_1 _35419_ (.A(net4536),
    .B(_09683_),
    .Y(_09695_));
 sg13g2_nand3_1 _35420_ (.B(net4636),
    .C(_09682_),
    .A(net4628),
    .Y(_09696_));
 sg13g2_a21oi_1 _35421_ (.A1(net4689),
    .A2(_09676_),
    .Y(_09697_),
    .B1(_09675_));
 sg13g2_nor2b_1 _35422_ (.A(_09697_),
    .B_N(_09694_),
    .Y(_09698_));
 sg13g2_o21ai_1 _35423_ (.B1(_09693_),
    .Y(_09699_),
    .A1(_09695_),
    .A2(_09698_));
 sg13g2_nor3_1 _35424_ (.A(_09693_),
    .B(_09695_),
    .C(_09698_),
    .Y(_09700_));
 sg13g2_nand3b_1 _35425_ (.B(net4689),
    .C(_09699_),
    .Y(_09701_),
    .A_N(_09700_));
 sg13g2_o21ai_1 _35426_ (.B1(_09701_),
    .Y(_09702_),
    .A1(net4689),
    .A2(_09690_));
 sg13g2_o21ai_1 _35427_ (.B1(net5590),
    .Y(_09703_),
    .A1(net4385),
    .A2(_09682_));
 sg13g2_a21oi_1 _35428_ (.A1(net4385),
    .A2(_09702_),
    .Y(_09704_),
    .B1(_09703_));
 sg13g2_a21o_1 _35429_ (.A2(net4125),
    .A1(net2430),
    .B1(_09704_),
    .X(_00776_));
 sg13g2_a21oi_1 _35430_ (.A1(net4791),
    .A2(_09377_),
    .Y(_09705_),
    .B1(_09393_));
 sg13g2_xnor2_1 _35431_ (.Y(_09706_),
    .A(_09396_),
    .B(_09705_));
 sg13g2_nand2_1 _35432_ (.Y(_09707_),
    .A(net5390),
    .B(_09706_));
 sg13g2_o21ai_1 _35433_ (.B1(_09707_),
    .Y(_09708_),
    .A1(net5390),
    .A2(_09370_));
 sg13g2_nand4_1 _35434_ (.B(_09692_),
    .C(_09694_),
    .A(_09691_),
    .Y(_09709_),
    .D(_09696_));
 sg13g2_and2_1 _35435_ (.A(_09691_),
    .B(_09696_),
    .X(_09710_));
 sg13g2_o21ai_1 _35436_ (.B1(_09710_),
    .Y(_09711_),
    .A1(_09697_),
    .A2(_09709_));
 sg13g2_nor2_1 _35437_ (.A(net4580),
    .B(_09708_),
    .Y(_09712_));
 sg13g2_nand2_1 _35438_ (.Y(_09713_),
    .A(net4536),
    .B(_09708_));
 sg13g2_xnor2_1 _35439_ (.Y(_09714_),
    .A(net4536),
    .B(_09708_));
 sg13g2_inv_1 _35440_ (.Y(_09715_),
    .A(_09714_));
 sg13g2_nand2_1 _35441_ (.Y(_09716_),
    .A(_09711_),
    .B(_09715_));
 sg13g2_nand2b_1 _35442_ (.Y(_09717_),
    .B(_09714_),
    .A_N(_09711_));
 sg13g2_a21o_1 _35443_ (.A2(_09717_),
    .A1(_09716_),
    .B1(net4646),
    .X(_09718_));
 sg13g2_o21ai_1 _35444_ (.B1(_09718_),
    .Y(_09719_),
    .A1(net4689),
    .A2(_09708_));
 sg13g2_o21ai_1 _35445_ (.B1(net5590),
    .Y(_09720_),
    .A1(net4385),
    .A2(_09690_));
 sg13g2_a21oi_1 _35446_ (.A1(net4384),
    .A2(_09719_),
    .Y(_09721_),
    .B1(_09720_));
 sg13g2_a21o_1 _35447_ (.A2(net4125),
    .A1(net2563),
    .B1(_09721_),
    .X(_00777_));
 sg13g2_nand2_1 _35448_ (.Y(_09722_),
    .A(net2781),
    .B(net4135));
 sg13g2_nand2_1 _35449_ (.Y(_09723_),
    .A(_09363_),
    .B(_09398_));
 sg13g2_nor2_1 _35450_ (.A(_09363_),
    .B(_09398_),
    .Y(_09724_));
 sg13g2_nor2_1 _35451_ (.A(net5350),
    .B(_09724_),
    .Y(_09725_));
 sg13g2_a22oi_1 _35452_ (.Y(_09726_),
    .B1(_09723_),
    .B2(_09725_),
    .A2(_09361_),
    .A1(net5350));
 sg13g2_xnor2_1 _35453_ (.Y(_09727_),
    .A(net4536),
    .B(_09726_));
 sg13g2_nand2_1 _35454_ (.Y(_09728_),
    .A(_09713_),
    .B(_09716_));
 sg13g2_xnor2_1 _35455_ (.Y(_09729_),
    .A(_09727_),
    .B(_09728_));
 sg13g2_o21ai_1 _35456_ (.B1(net4390),
    .Y(_09730_),
    .A1(net4694),
    .A2(_09726_));
 sg13g2_a21oi_1 _35457_ (.A1(net4694),
    .A2(_09729_),
    .Y(_09731_),
    .B1(_09730_));
 sg13g2_o21ai_1 _35458_ (.B1(net5590),
    .Y(_09732_),
    .A1(net4385),
    .A2(_09708_));
 sg13g2_o21ai_1 _35459_ (.B1(_09722_),
    .Y(_00778_),
    .A1(_09731_),
    .A2(_09732_));
 sg13g2_nand2_1 _35460_ (.Y(_09733_),
    .A(_09362_),
    .B(_09723_));
 sg13g2_xor2_1 _35461_ (.B(_09733_),
    .A(_09356_),
    .X(_09734_));
 sg13g2_nand2_1 _35462_ (.Y(_09735_),
    .A(net5393),
    .B(_09734_));
 sg13g2_o21ai_1 _35463_ (.B1(_09735_),
    .Y(_09736_),
    .A1(net5393),
    .A2(_09355_));
 sg13g2_nand2_1 _35464_ (.Y(_09737_),
    .A(net4647),
    .B(_09736_));
 sg13g2_nor2_1 _35465_ (.A(net4582),
    .B(_09736_),
    .Y(_09738_));
 sg13g2_nand2_1 _35466_ (.Y(_09739_),
    .A(net4582),
    .B(_09736_));
 sg13g2_xnor2_1 _35467_ (.Y(_09740_),
    .A(net4582),
    .B(_09736_));
 sg13g2_nor2_1 _35468_ (.A(_09712_),
    .B(_09726_),
    .Y(_09741_));
 sg13g2_a21oi_1 _35469_ (.A1(_09711_),
    .A2(_09715_),
    .Y(_09742_),
    .B1(_09741_));
 sg13g2_a21oi_1 _35470_ (.A1(net4539),
    .A2(_09726_),
    .Y(_09743_),
    .B1(_09742_));
 sg13g2_xnor2_1 _35471_ (.Y(_09744_),
    .A(_09740_),
    .B(_09743_));
 sg13g2_o21ai_1 _35472_ (.B1(_09737_),
    .Y(_09745_),
    .A1(net4647),
    .A2(_09744_));
 sg13g2_nand2_1 _35473_ (.Y(_09746_),
    .A(net4390),
    .B(_09745_));
 sg13g2_a21oi_1 _35474_ (.A1(net4354),
    .A2(_09726_),
    .Y(_09747_),
    .B1(net5529));
 sg13g2_a22oi_1 _35475_ (.Y(_09748_),
    .B1(_09746_),
    .B2(_09747_),
    .A2(net4135),
    .A1(net2862));
 sg13g2_inv_1 _35476_ (.Y(_00779_),
    .A(_09748_));
 sg13g2_nand3_1 _35477_ (.B(_09400_),
    .C(_09429_),
    .A(_09399_),
    .Y(_09749_));
 sg13g2_a21o_1 _35478_ (.A2(_09400_),
    .A1(_09399_),
    .B1(_09429_),
    .X(_09750_));
 sg13g2_and3_1 _35479_ (.X(_09751_),
    .A(net5393),
    .B(_09749_),
    .C(_09750_));
 sg13g2_a21oi_2 _35480_ (.B1(_09751_),
    .Y(_09752_),
    .A2(_09427_),
    .A1(net5350));
 sg13g2_xnor2_1 _35481_ (.Y(_09753_),
    .A(net4582),
    .B(_09752_));
 sg13g2_a21oi_1 _35482_ (.A1(_09739_),
    .A2(_09743_),
    .Y(_09754_),
    .B1(_09738_));
 sg13g2_xor2_1 _35483_ (.B(_09754_),
    .A(_09753_),
    .X(_09755_));
 sg13g2_o21ai_1 _35484_ (.B1(net4390),
    .Y(_09756_),
    .A1(net4694),
    .A2(_09752_));
 sg13g2_a21o_1 _35485_ (.A2(_09755_),
    .A1(net4694),
    .B1(_09756_),
    .X(_09757_));
 sg13g2_a21oi_1 _35486_ (.A1(net4354),
    .A2(_09736_),
    .Y(_09758_),
    .B1(net5529));
 sg13g2_a22oi_1 _35487_ (.Y(_09759_),
    .B1(_09757_),
    .B2(_09758_),
    .A2(net4135),
    .A1(net2543));
 sg13g2_inv_1 _35488_ (.Y(_00780_),
    .A(_09759_));
 sg13g2_nand2_1 _35489_ (.Y(_09760_),
    .A(_09428_),
    .B(_09750_));
 sg13g2_xor2_1 _35490_ (.B(_09760_),
    .A(_09441_),
    .X(_09761_));
 sg13g2_nand2_1 _35491_ (.Y(_09762_),
    .A(net5393),
    .B(_09761_));
 sg13g2_o21ai_1 _35492_ (.B1(_09762_),
    .Y(_09763_),
    .A1(net5393),
    .A2(_09438_));
 sg13g2_nand2_1 _35493_ (.Y(_09764_),
    .A(net4647),
    .B(_09763_));
 sg13g2_nor2_1 _35494_ (.A(net4582),
    .B(_09763_),
    .Y(_09765_));
 sg13g2_xnor2_1 _35495_ (.Y(_09766_),
    .A(net4539),
    .B(_09763_));
 sg13g2_nor2_1 _35496_ (.A(_09740_),
    .B(_09753_),
    .Y(_09767_));
 sg13g2_nor4_1 _35497_ (.A(_09714_),
    .B(_09727_),
    .C(_09740_),
    .D(_09753_),
    .Y(_09768_));
 sg13g2_a21oi_1 _35498_ (.A1(_09736_),
    .A2(_09752_),
    .Y(_09769_),
    .B1(net4582));
 sg13g2_a221oi_1 _35499_ (.B2(_09711_),
    .C1(_09769_),
    .B1(_09768_),
    .A1(_09741_),
    .Y(_09770_),
    .A2(_09767_));
 sg13g2_nor2b_1 _35500_ (.A(_09770_),
    .B_N(_09766_),
    .Y(_09771_));
 sg13g2_xnor2_1 _35501_ (.Y(_09772_),
    .A(_09766_),
    .B(_09770_));
 sg13g2_o21ai_1 _35502_ (.B1(_09764_),
    .Y(_09773_),
    .A1(net4647),
    .A2(_09772_));
 sg13g2_nand2_1 _35503_ (.Y(_09774_),
    .A(net4390),
    .B(_09773_));
 sg13g2_a21oi_1 _35504_ (.A1(net4354),
    .A2(_09752_),
    .Y(_09775_),
    .B1(net5529));
 sg13g2_a22oi_1 _35505_ (.Y(_09776_),
    .B1(_09774_),
    .B2(_09775_),
    .A2(net4135),
    .A1(net2426));
 sg13g2_inv_1 _35506_ (.Y(_00781_),
    .A(_09776_));
 sg13g2_nor2b_1 _35507_ (.A(_09489_),
    .B_N(_09750_),
    .Y(_09777_));
 sg13g2_or3_1 _35508_ (.A(_09420_),
    .B(_09440_),
    .C(_09777_),
    .X(_09778_));
 sg13g2_o21ai_1 _35509_ (.B1(_09420_),
    .Y(_09779_),
    .A1(_09440_),
    .A2(_09777_));
 sg13g2_and3_1 _35510_ (.X(_09780_),
    .A(net5393),
    .B(_09778_),
    .C(_09779_));
 sg13g2_a21oi_2 _35511_ (.B1(_09780_),
    .Y(_09781_),
    .A2(_09418_),
    .A1(net5350));
 sg13g2_nand2_1 _35512_ (.Y(_09782_),
    .A(net4647),
    .B(_09781_));
 sg13g2_nand2_1 _35513_ (.Y(_09783_),
    .A(net4582),
    .B(_09781_));
 sg13g2_xnor2_1 _35514_ (.Y(_09784_),
    .A(net4582),
    .B(_09781_));
 sg13g2_nor2_1 _35515_ (.A(_09765_),
    .B(_09771_),
    .Y(_09785_));
 sg13g2_xor2_1 _35516_ (.B(_09785_),
    .A(_09784_),
    .X(_09786_));
 sg13g2_o21ai_1 _35517_ (.B1(_09782_),
    .Y(_09787_),
    .A1(net4647),
    .A2(_09786_));
 sg13g2_nand2_1 _35518_ (.Y(_09788_),
    .A(net4390),
    .B(_09787_));
 sg13g2_a21oi_1 _35519_ (.A1(net4354),
    .A2(_09763_),
    .Y(_09789_),
    .B1(net5529));
 sg13g2_a22oi_1 _35520_ (.Y(_09790_),
    .B1(_09788_),
    .B2(_09789_),
    .A2(net4135),
    .A1(net2604));
 sg13g2_inv_1 _35521_ (.Y(_00782_),
    .A(_09790_));
 sg13g2_nor2_1 _35522_ (.A(net5396),
    .B(_09412_),
    .Y(_09791_));
 sg13g2_nand2_1 _35523_ (.Y(_09792_),
    .A(_09419_),
    .B(_09778_));
 sg13g2_xnor2_1 _35524_ (.Y(_09793_),
    .A(_09413_),
    .B(_09792_));
 sg13g2_a21oi_1 _35525_ (.A1(net5393),
    .A2(_09793_),
    .Y(_09794_),
    .B1(_09791_));
 sg13g2_or3_1 _35526_ (.A(net4634),
    .B(net4635),
    .C(_09794_),
    .X(_09795_));
 sg13g2_o21ai_1 _35527_ (.B1(_09794_),
    .Y(_09796_),
    .A1(net4634),
    .A2(net4635));
 sg13g2_nand2_1 _35528_ (.Y(_09797_),
    .A(_09795_),
    .B(_09796_));
 sg13g2_a21o_1 _35529_ (.A2(_09781_),
    .A1(_09763_),
    .B1(net4583),
    .X(_09798_));
 sg13g2_nand2b_1 _35530_ (.Y(_09799_),
    .B(_09798_),
    .A_N(_09771_));
 sg13g2_nand2_1 _35531_ (.Y(_09800_),
    .A(_09783_),
    .B(_09799_));
 sg13g2_a21oi_1 _35532_ (.A1(_09797_),
    .A2(_09800_),
    .Y(_09801_),
    .B1(net4647));
 sg13g2_o21ai_1 _35533_ (.B1(_09801_),
    .Y(_09802_),
    .A1(_09797_),
    .A2(_09800_));
 sg13g2_or2_1 _35534_ (.X(_09803_),
    .B(_09794_),
    .A(net4694));
 sg13g2_nand3_1 _35535_ (.B(_09802_),
    .C(_09803_),
    .A(net4390),
    .Y(_09804_));
 sg13g2_a21oi_1 _35536_ (.A1(net4354),
    .A2(_09781_),
    .Y(_09805_),
    .B1(net5529));
 sg13g2_a22oi_1 _35537_ (.Y(_09806_),
    .B1(_09804_),
    .B2(_09805_),
    .A2(net4135),
    .A1(net2503));
 sg13g2_inv_1 _35538_ (.Y(_00783_),
    .A(_09806_));
 sg13g2_nor2_1 _35539_ (.A(net5393),
    .B(_09473_),
    .Y(_09807_));
 sg13g2_o21ai_1 _35540_ (.B1(_09475_),
    .Y(_09808_),
    .A1(_09443_),
    .A2(_09491_));
 sg13g2_nor3_1 _35541_ (.A(_09443_),
    .B(_09475_),
    .C(_09491_),
    .Y(_09809_));
 sg13g2_nor2_1 _35542_ (.A(net5350),
    .B(_09809_),
    .Y(_09810_));
 sg13g2_a21o_2 _35543_ (.A2(_09810_),
    .A1(_09808_),
    .B1(_09807_),
    .X(_09811_));
 sg13g2_nor2_1 _35544_ (.A(net4694),
    .B(_09811_),
    .Y(_09812_));
 sg13g2_nand3_1 _35545_ (.B(net4636),
    .C(_09811_),
    .A(net4628),
    .Y(_09813_));
 sg13g2_a21o_1 _35546_ (.A2(net4636),
    .A1(net4628),
    .B1(_09811_),
    .X(_09814_));
 sg13g2_nand2_1 _35547_ (.Y(_09815_),
    .A(_09813_),
    .B(_09814_));
 sg13g2_o21ai_1 _35548_ (.B1(_09795_),
    .Y(_09816_),
    .A1(_09797_),
    .A2(_09800_));
 sg13g2_o21ai_1 _35549_ (.B1(net4694),
    .Y(_09817_),
    .A1(_09815_),
    .A2(_09816_));
 sg13g2_a21oi_1 _35550_ (.A1(_09815_),
    .A2(_09816_),
    .Y(_09818_),
    .B1(_09817_));
 sg13g2_o21ai_1 _35551_ (.B1(net4391),
    .Y(_09819_),
    .A1(_09812_),
    .A2(_09818_));
 sg13g2_a21oi_1 _35552_ (.A1(net4354),
    .A2(_09794_),
    .Y(_09820_),
    .B1(net5529));
 sg13g2_a22oi_1 _35553_ (.Y(_09821_),
    .B1(_09819_),
    .B2(_09820_),
    .A2(net4135),
    .A1(net3093));
 sg13g2_inv_1 _35554_ (.Y(_00784_),
    .A(_09821_));
 sg13g2_nand2_1 _35555_ (.Y(_09822_),
    .A(net5350),
    .B(_09481_));
 sg13g2_nand2_1 _35556_ (.Y(_09823_),
    .A(_09474_),
    .B(_09808_));
 sg13g2_xnor2_1 _35557_ (.Y(_09824_),
    .A(_09484_),
    .B(_09823_));
 sg13g2_o21ai_1 _35558_ (.B1(_09822_),
    .Y(_09825_),
    .A1(net5350),
    .A2(_09824_));
 sg13g2_nand2_1 _35559_ (.Y(_09826_),
    .A(net4583),
    .B(_09825_));
 sg13g2_xnor2_1 _35560_ (.Y(_09827_),
    .A(net4539),
    .B(_09825_));
 sg13g2_nand4_1 _35561_ (.B(_09796_),
    .C(_09813_),
    .A(_09795_),
    .Y(_09828_),
    .D(_09814_));
 sg13g2_and2_1 _35562_ (.A(_09795_),
    .B(_09813_),
    .X(_09829_));
 sg13g2_o21ai_1 _35563_ (.B1(_09829_),
    .Y(_09830_),
    .A1(_09798_),
    .A2(_09828_));
 sg13g2_nor2_1 _35564_ (.A(_09784_),
    .B(_09828_),
    .Y(_09831_));
 sg13g2_nand2_1 _35565_ (.Y(_09832_),
    .A(_09766_),
    .B(_09831_));
 sg13g2_nor2_1 _35566_ (.A(_09770_),
    .B(_09832_),
    .Y(_09833_));
 sg13g2_o21ai_1 _35567_ (.B1(_09827_),
    .Y(_09834_),
    .A1(_09830_),
    .A2(_09833_));
 sg13g2_or3_1 _35568_ (.A(_09827_),
    .B(_09830_),
    .C(_09833_),
    .X(_09835_));
 sg13g2_a21o_1 _35569_ (.A2(_09835_),
    .A1(_09834_),
    .B1(net4647),
    .X(_09836_));
 sg13g2_o21ai_1 _35570_ (.B1(_09836_),
    .Y(_09837_),
    .A1(net4694),
    .A2(_09825_));
 sg13g2_o21ai_1 _35571_ (.B1(net5594),
    .Y(_09838_),
    .A1(net4390),
    .A2(_09811_));
 sg13g2_a21oi_1 _35572_ (.A1(net4390),
    .A2(_09837_),
    .Y(_09839_),
    .B1(_09838_));
 sg13g2_a21o_1 _35573_ (.A2(net4135),
    .A1(net3215),
    .B1(_09839_),
    .X(_00785_));
 sg13g2_nand2_1 _35574_ (.Y(_09840_),
    .A(_09487_),
    .B(_09808_));
 sg13g2_nand3_1 _35575_ (.B(_09483_),
    .C(_09840_),
    .A(_09466_),
    .Y(_09841_));
 sg13g2_a21oi_1 _35576_ (.A1(_09483_),
    .A2(_09840_),
    .Y(_09842_),
    .B1(_09466_));
 sg13g2_nor2_1 _35577_ (.A(net5352),
    .B(_09842_),
    .Y(_09843_));
 sg13g2_a22oi_1 _35578_ (.Y(_09844_),
    .B1(_09841_),
    .B2(_09843_),
    .A2(_09464_),
    .A1(net5352));
 sg13g2_inv_1 _35579_ (.Y(_09845_),
    .A(_09844_));
 sg13g2_nand2_1 _35580_ (.Y(_09846_),
    .A(net4649),
    .B(_09844_));
 sg13g2_xnor2_1 _35581_ (.Y(_09847_),
    .A(net4584),
    .B(_09844_));
 sg13g2_nand2_1 _35582_ (.Y(_09848_),
    .A(_09826_),
    .B(_09834_));
 sg13g2_xor2_1 _35583_ (.B(_09848_),
    .A(_09847_),
    .X(_09849_));
 sg13g2_o21ai_1 _35584_ (.B1(_09846_),
    .Y(_09850_),
    .A1(net4649),
    .A2(_09849_));
 sg13g2_o21ai_1 _35585_ (.B1(net5593),
    .Y(_09851_),
    .A1(net4392),
    .A2(_09825_));
 sg13g2_a21oi_1 _35586_ (.A1(net4392),
    .A2(_09850_),
    .Y(_09852_),
    .B1(_09851_));
 sg13g2_a21o_1 _35587_ (.A2(net4137),
    .A1(net2523),
    .B1(_09852_),
    .X(_00786_));
 sg13g2_and3_1 _35588_ (.X(_09853_),
    .A(_09458_),
    .B(_09465_),
    .C(_09841_));
 sg13g2_a21oi_1 _35589_ (.A1(_09465_),
    .A2(_09841_),
    .Y(_09854_),
    .B1(_09458_));
 sg13g2_o21ai_1 _35590_ (.B1(net5395),
    .Y(_09855_),
    .A1(_09853_),
    .A2(_09854_));
 sg13g2_o21ai_1 _35591_ (.B1(_09855_),
    .Y(_09856_),
    .A1(net5395),
    .A2(_09457_));
 sg13g2_nand2_1 _35592_ (.Y(_09857_),
    .A(net4584),
    .B(_09856_));
 sg13g2_xnor2_1 _35593_ (.Y(_09858_),
    .A(net4538),
    .B(_09856_));
 sg13g2_o21ai_1 _35594_ (.B1(net4584),
    .Y(_09859_),
    .A1(_09825_),
    .A2(_09845_));
 sg13g2_inv_1 _35595_ (.Y(_09860_),
    .A(_09859_));
 sg13g2_a22oi_1 _35596_ (.Y(_09861_),
    .B1(_09859_),
    .B2(_09834_),
    .A2(_09844_),
    .A1(net4538));
 sg13g2_nand2_1 _35597_ (.Y(_09862_),
    .A(_09858_),
    .B(_09861_));
 sg13g2_or2_1 _35598_ (.X(_09863_),
    .B(_09861_),
    .A(_09858_));
 sg13g2_a21o_1 _35599_ (.A2(_09863_),
    .A1(_09862_),
    .B1(net4649),
    .X(_09864_));
 sg13g2_o21ai_1 _35600_ (.B1(_09864_),
    .Y(_09865_),
    .A1(net4692),
    .A2(_09856_));
 sg13g2_nand2_1 _35601_ (.Y(_09866_),
    .A(net4392),
    .B(_09865_));
 sg13g2_a21oi_1 _35602_ (.A1(net4355),
    .A2(_09844_),
    .Y(_09867_),
    .B1(net5530));
 sg13g2_a22oi_1 _35603_ (.Y(_09868_),
    .B1(_09866_),
    .B2(_09867_),
    .A2(net4137),
    .A1(net2508));
 sg13g2_inv_1 _35604_ (.Y(_00787_),
    .A(_09868_));
 sg13g2_nand2_1 _35605_ (.Y(_09869_),
    .A(net5352),
    .B(_09531_));
 sg13g2_nand2b_1 _35606_ (.Y(_09870_),
    .B(_09533_),
    .A_N(_09494_));
 sg13g2_xor2_1 _35607_ (.B(_09533_),
    .A(_09494_),
    .X(_09871_));
 sg13g2_o21ai_1 _35608_ (.B1(_09869_),
    .Y(_09872_),
    .A1(net5352),
    .A2(_09871_));
 sg13g2_nand2_1 _35609_ (.Y(_09873_),
    .A(net4584),
    .B(_09872_));
 sg13g2_xnor2_1 _35610_ (.Y(_09874_),
    .A(net4538),
    .B(_09872_));
 sg13g2_nand3_1 _35611_ (.B(_09862_),
    .C(_09874_),
    .A(_09857_),
    .Y(_09875_));
 sg13g2_a21oi_1 _35612_ (.A1(_09857_),
    .A2(_09862_),
    .Y(_09876_),
    .B1(_09874_));
 sg13g2_nand3b_1 _35613_ (.B(net4692),
    .C(_09875_),
    .Y(_09877_),
    .A_N(_09876_));
 sg13g2_o21ai_1 _35614_ (.B1(_09877_),
    .Y(_09878_),
    .A1(net4692),
    .A2(_09872_));
 sg13g2_o21ai_1 _35615_ (.B1(net5593),
    .Y(_09879_),
    .A1(net4392),
    .A2(_09856_));
 sg13g2_a21oi_1 _35616_ (.A1(net4392),
    .A2(_09878_),
    .Y(_09880_),
    .B1(_09879_));
 sg13g2_a21o_1 _35617_ (.A2(net4137),
    .A1(net2441),
    .B1(_09880_),
    .X(_00788_));
 sg13g2_nor2_1 _35618_ (.A(net5395),
    .B(_09524_),
    .Y(_09881_));
 sg13g2_nand2_1 _35619_ (.Y(_09882_),
    .A(_09532_),
    .B(_09870_));
 sg13g2_xnor2_1 _35620_ (.Y(_09883_),
    .A(_09526_),
    .B(_09882_));
 sg13g2_a21oi_2 _35621_ (.B1(_09881_),
    .Y(_09884_),
    .A2(_09883_),
    .A1(net5395));
 sg13g2_nand2_1 _35622_ (.Y(_09885_),
    .A(net4584),
    .B(_09884_));
 sg13g2_xnor2_1 _35623_ (.Y(_09886_),
    .A(net4538),
    .B(_09884_));
 sg13g2_and2_1 _35624_ (.A(_09858_),
    .B(_09874_),
    .X(_09887_));
 sg13g2_nand2_1 _35625_ (.Y(_09888_),
    .A(_09857_),
    .B(_09873_));
 sg13g2_and4_1 _35626_ (.A(_09827_),
    .B(_09847_),
    .C(_09858_),
    .D(_09874_),
    .X(_09889_));
 sg13g2_a221oi_1 _35627_ (.B2(_09830_),
    .C1(_09888_),
    .B1(_09889_),
    .A1(_09860_),
    .Y(_09890_),
    .A2(_09887_));
 sg13g2_nand3_1 _35628_ (.B(_09831_),
    .C(_09889_),
    .A(_09766_),
    .Y(_09891_));
 sg13g2_o21ai_1 _35629_ (.B1(_09890_),
    .Y(_09892_),
    .A1(_09770_),
    .A2(_09891_));
 sg13g2_nor2_1 _35630_ (.A(_09886_),
    .B(_09892_),
    .Y(_09893_));
 sg13g2_nand2_1 _35631_ (.Y(_09894_),
    .A(_09886_),
    .B(_09892_));
 sg13g2_nor2_1 _35632_ (.A(net4649),
    .B(_09893_),
    .Y(_09895_));
 sg13g2_a22oi_1 _35633_ (.Y(_09896_),
    .B1(_09894_),
    .B2(_09895_),
    .A2(_09884_),
    .A1(net4649));
 sg13g2_o21ai_1 _35634_ (.B1(net5593),
    .Y(_09897_),
    .A1(net4393),
    .A2(_09872_));
 sg13g2_a21oi_1 _35635_ (.A1(net4393),
    .A2(_09896_),
    .Y(_09898_),
    .B1(_09897_));
 sg13g2_a21o_1 _35636_ (.A2(net4138),
    .A1(net2619),
    .B1(_09898_),
    .X(_00789_));
 sg13g2_nor2_1 _35637_ (.A(net5395),
    .B(_09504_),
    .Y(_09899_));
 sg13g2_and2_1 _35638_ (.A(_09583_),
    .B(_09870_),
    .X(_09900_));
 sg13g2_nor2_1 _35639_ (.A(_09525_),
    .B(_09900_),
    .Y(_09901_));
 sg13g2_nor3_1 _35640_ (.A(_09506_),
    .B(_09525_),
    .C(_09900_),
    .Y(_09902_));
 sg13g2_xnor2_1 _35641_ (.Y(_09903_),
    .A(_09506_),
    .B(_09901_));
 sg13g2_a21oi_2 _35642_ (.B1(_09899_),
    .Y(_09904_),
    .A2(_09903_),
    .A1(net5395));
 sg13g2_inv_1 _35643_ (.Y(_09905_),
    .A(_09904_));
 sg13g2_nand2_1 _35644_ (.Y(_09906_),
    .A(net4649),
    .B(_09904_));
 sg13g2_nor2_1 _35645_ (.A(net4584),
    .B(_09905_),
    .Y(_09907_));
 sg13g2_xnor2_1 _35646_ (.Y(_09908_),
    .A(net4584),
    .B(_09904_));
 sg13g2_nand2_1 _35647_ (.Y(_09909_),
    .A(_09885_),
    .B(_09894_));
 sg13g2_xor2_1 _35648_ (.B(_09909_),
    .A(_09908_),
    .X(_09910_));
 sg13g2_o21ai_1 _35649_ (.B1(_09906_),
    .Y(_09911_),
    .A1(net4649),
    .A2(_09910_));
 sg13g2_o21ai_1 _35650_ (.B1(net5593),
    .Y(_09912_),
    .A1(net4393),
    .A2(_09884_));
 sg13g2_a21oi_1 _35651_ (.A1(net4393),
    .A2(_09911_),
    .Y(_09913_),
    .B1(_09912_));
 sg13g2_a21o_1 _35652_ (.A2(net4137),
    .A1(net2934),
    .B1(_09913_),
    .X(_00790_));
 sg13g2_nor2_1 _35653_ (.A(_09505_),
    .B(_09902_),
    .Y(_09914_));
 sg13g2_and2_1 _35654_ (.A(net5352),
    .B(_09514_),
    .X(_09915_));
 sg13g2_xnor2_1 _35655_ (.Y(_09916_),
    .A(_09515_),
    .B(_09914_));
 sg13g2_a21oi_2 _35656_ (.B1(_09915_),
    .Y(_09917_),
    .A2(_09916_),
    .A1(net5395));
 sg13g2_nand3_1 _35657_ (.B(net4636),
    .C(_09917_),
    .A(net4628),
    .Y(_09918_));
 sg13g2_nor2_1 _35658_ (.A(net4586),
    .B(_09917_),
    .Y(_09919_));
 sg13g2_a21o_1 _35659_ (.A2(net4636),
    .A1(net4628),
    .B1(_09917_),
    .X(_09920_));
 sg13g2_and2_1 _35660_ (.A(_09918_),
    .B(_09920_),
    .X(_09921_));
 sg13g2_o21ai_1 _35661_ (.B1(net4584),
    .Y(_09922_),
    .A1(_09884_),
    .A2(_09905_));
 sg13g2_a21o_1 _35662_ (.A2(_09922_),
    .A1(_09894_),
    .B1(_09907_),
    .X(_09923_));
 sg13g2_xor2_1 _35663_ (.B(_09923_),
    .A(_09921_),
    .X(_09924_));
 sg13g2_nand2_1 _35664_ (.Y(_09925_),
    .A(net4692),
    .B(_09924_));
 sg13g2_o21ai_1 _35665_ (.B1(_09925_),
    .Y(_09926_),
    .A1(net4692),
    .A2(_09917_));
 sg13g2_nand2_1 _35666_ (.Y(_09927_),
    .A(net4392),
    .B(_09926_));
 sg13g2_a21oi_1 _35667_ (.A1(net4355),
    .A2(_09904_),
    .Y(_09928_),
    .B1(net5530));
 sg13g2_a22oi_1 _35668_ (.Y(_09929_),
    .B1(_09927_),
    .B2(_09928_),
    .A2(net4137),
    .A1(net2787));
 sg13g2_inv_1 _35669_ (.Y(_00791_),
    .A(_09929_));
 sg13g2_nand2_1 _35670_ (.Y(_09930_),
    .A(net5354),
    .B(_09542_));
 sg13g2_nor2b_1 _35671_ (.A(_09494_),
    .B_N(_09535_),
    .Y(_09931_));
 sg13g2_or3_1 _35672_ (.A(_09584_),
    .B(_09585_),
    .C(_09931_),
    .X(_09932_));
 sg13g2_nand2b_1 _35673_ (.Y(_09933_),
    .B(_09932_),
    .A_N(_09544_));
 sg13g2_xor2_1 _35674_ (.B(_09932_),
    .A(_09544_),
    .X(_09934_));
 sg13g2_o21ai_1 _35675_ (.B1(_09930_),
    .Y(_09935_),
    .A1(net5354),
    .A2(_09934_));
 sg13g2_nand3_1 _35676_ (.B(net4636),
    .C(_09935_),
    .A(net4628),
    .Y(_09936_));
 sg13g2_a21o_1 _35677_ (.A2(net4638),
    .A1(net4630),
    .B1(_09935_),
    .X(_09937_));
 sg13g2_and2_1 _35678_ (.A(_09936_),
    .B(_09937_),
    .X(_09938_));
 sg13g2_o21ai_1 _35679_ (.B1(_09918_),
    .Y(_09939_),
    .A1(_09919_),
    .A2(_09923_));
 sg13g2_xnor2_1 _35680_ (.Y(_09940_),
    .A(_09938_),
    .B(_09939_));
 sg13g2_nand2_1 _35681_ (.Y(_09941_),
    .A(net4697),
    .B(_09940_));
 sg13g2_o21ai_1 _35682_ (.B1(_09941_),
    .Y(_09942_),
    .A1(net4692),
    .A2(_09935_));
 sg13g2_o21ai_1 _35683_ (.B1(net5593),
    .Y(_09943_),
    .A1(net4392),
    .A2(_09917_));
 sg13g2_a21oi_1 _35684_ (.A1(net4392),
    .A2(_09942_),
    .Y(_09944_),
    .B1(_09943_));
 sg13g2_a21o_1 _35685_ (.A2(net4137),
    .A1(net2704),
    .B1(_09944_),
    .X(_00792_));
 sg13g2_nand2_1 _35686_ (.Y(_09945_),
    .A(_09543_),
    .B(_09933_));
 sg13g2_xor2_1 _35687_ (.B(_09945_),
    .A(_09555_),
    .X(_09946_));
 sg13g2_nor2_1 _35688_ (.A(net5354),
    .B(_09946_),
    .Y(_09947_));
 sg13g2_a21oi_2 _35689_ (.B1(_09947_),
    .Y(_09948_),
    .A2(_09552_),
    .A1(net5354));
 sg13g2_nand2_1 _35690_ (.Y(_09949_),
    .A(net4590),
    .B(_09948_));
 sg13g2_xnor2_1 _35691_ (.Y(_09950_),
    .A(net4541),
    .B(_09948_));
 sg13g2_nand4_1 _35692_ (.B(_09920_),
    .C(_09936_),
    .A(_09918_),
    .Y(_09951_),
    .D(_09937_));
 sg13g2_and2_1 _35693_ (.A(_09918_),
    .B(_09936_),
    .X(_09952_));
 sg13g2_o21ai_1 _35694_ (.B1(_09952_),
    .Y(_09953_),
    .A1(_09922_),
    .A2(_09951_));
 sg13g2_and2_1 _35695_ (.A(_09886_),
    .B(_09908_),
    .X(_09954_));
 sg13g2_nand4_1 _35696_ (.B(_09921_),
    .C(_09938_),
    .A(_09892_),
    .Y(_09955_),
    .D(_09954_));
 sg13g2_nor2b_1 _35697_ (.A(_09953_),
    .B_N(_09955_),
    .Y(_09956_));
 sg13g2_nand2b_1 _35698_ (.Y(_09957_),
    .B(_09950_),
    .A_N(_09956_));
 sg13g2_nand2b_1 _35699_ (.Y(_09958_),
    .B(_09956_),
    .A_N(_09950_));
 sg13g2_a21o_1 _35700_ (.A2(_09958_),
    .A1(_09957_),
    .B1(net4653),
    .X(_09959_));
 sg13g2_o21ai_1 _35701_ (.B1(_09959_),
    .Y(_09960_),
    .A1(net4697),
    .A2(_09948_));
 sg13g2_o21ai_1 _35702_ (.B1(net5595),
    .Y(_09961_),
    .A1(net4397),
    .A2(_09935_));
 sg13g2_a21oi_1 _35703_ (.A1(net4397),
    .A2(_09960_),
    .Y(_09962_),
    .B1(_09961_));
 sg13g2_a21o_1 _35704_ (.A2(net4152),
    .A1(net2904),
    .B1(_09962_),
    .X(_00793_));
 sg13g2_nor2_1 _35705_ (.A(net5397),
    .B(_09566_),
    .Y(_09963_));
 sg13g2_nand2_1 _35706_ (.Y(_09964_),
    .A(_09582_),
    .B(_09933_));
 sg13g2_nand3_1 _35707_ (.B(_09569_),
    .C(_09964_),
    .A(_09554_),
    .Y(_09965_));
 sg13g2_a21oi_1 _35708_ (.A1(_09554_),
    .A2(_09964_),
    .Y(_09966_),
    .B1(_09569_));
 sg13g2_nor2_1 _35709_ (.A(net5354),
    .B(_09966_),
    .Y(_09967_));
 sg13g2_a21oi_2 _35710_ (.B1(_09963_),
    .Y(_09968_),
    .A2(_09967_),
    .A1(_09965_));
 sg13g2_nand2_1 _35711_ (.Y(_09969_),
    .A(net4653),
    .B(_09968_));
 sg13g2_nand2_1 _35712_ (.Y(_09970_),
    .A(net4541),
    .B(_09968_));
 sg13g2_xnor2_1 _35713_ (.Y(_09971_),
    .A(net4590),
    .B(_09968_));
 sg13g2_nand2_1 _35714_ (.Y(_09972_),
    .A(_09949_),
    .B(_09957_));
 sg13g2_xor2_1 _35715_ (.B(_09972_),
    .A(_09971_),
    .X(_09973_));
 sg13g2_o21ai_1 _35716_ (.B1(_09969_),
    .Y(_09974_),
    .A1(net4653),
    .A2(_09973_));
 sg13g2_o21ai_1 _35717_ (.B1(net5595),
    .Y(_09975_),
    .A1(net4397),
    .A2(_09948_));
 sg13g2_a21oi_1 _35718_ (.A1(net4397),
    .A2(_09974_),
    .Y(_09976_),
    .B1(_09975_));
 sg13g2_a21o_1 _35719_ (.A2(net4152),
    .A1(net2596),
    .B1(_09976_),
    .X(_00794_));
 sg13g2_nand2_1 _35720_ (.Y(_09977_),
    .A(net4356),
    .B(_09968_));
 sg13g2_nand2b_1 _35721_ (.Y(_09978_),
    .B(_09965_),
    .A_N(_09567_));
 sg13g2_xnor2_1 _35722_ (.Y(_09979_),
    .A(_09578_),
    .B(_09978_));
 sg13g2_nor2_1 _35723_ (.A(net5354),
    .B(_09979_),
    .Y(_09980_));
 sg13g2_a21oi_2 _35724_ (.B1(_09980_),
    .Y(_09981_),
    .A2(_09577_),
    .A1(net5354));
 sg13g2_nand2_1 _35725_ (.Y(_09982_),
    .A(net4590),
    .B(_09981_));
 sg13g2_xnor2_1 _35726_ (.Y(_09983_),
    .A(net4541),
    .B(_09981_));
 sg13g2_o21ai_1 _35727_ (.B1(_09949_),
    .Y(_09984_),
    .A1(net4541),
    .A2(_09968_));
 sg13g2_nand2b_1 _35728_ (.Y(_09985_),
    .B(_09957_),
    .A_N(_09984_));
 sg13g2_a21o_1 _35729_ (.A2(_09985_),
    .A1(_09970_),
    .B1(_09983_),
    .X(_09986_));
 sg13g2_nand3_1 _35730_ (.B(_09983_),
    .C(_09985_),
    .A(_09970_),
    .Y(_09987_));
 sg13g2_and2_1 _35731_ (.A(net4697),
    .B(_09987_),
    .X(_09988_));
 sg13g2_a22oi_1 _35732_ (.Y(_09989_),
    .B1(_09986_),
    .B2(_09988_),
    .A2(_09981_),
    .A1(net4653));
 sg13g2_a21oi_1 _35733_ (.A1(net4397),
    .A2(_09989_),
    .Y(_09990_),
    .B1(net5538));
 sg13g2_a22oi_1 _35734_ (.Y(_09991_),
    .B1(_09977_),
    .B2(_09990_),
    .A2(net4152),
    .A1(net2299));
 sg13g2_inv_1 _35735_ (.Y(_00795_),
    .A(_09991_));
 sg13g2_nand2_1 _35736_ (.Y(_09992_),
    .A(net2308),
    .B(net4152));
 sg13g2_nor2_1 _35737_ (.A(net5397),
    .B(_09324_),
    .Y(_09993_));
 sg13g2_and2_1 _35738_ (.A(_09581_),
    .B(_09589_),
    .X(_09994_));
 sg13g2_nor2_1 _35739_ (.A(_09341_),
    .B(_09994_),
    .Y(_09995_));
 sg13g2_xor2_1 _35740_ (.B(_09994_),
    .A(_09341_),
    .X(_09996_));
 sg13g2_a21oi_2 _35741_ (.B1(_09993_),
    .Y(_09997_),
    .A2(_09996_),
    .A1(net5397));
 sg13g2_xnor2_1 _35742_ (.Y(_09998_),
    .A(net4590),
    .B(_09997_));
 sg13g2_nand2_1 _35743_ (.Y(_09999_),
    .A(_09982_),
    .B(_09987_));
 sg13g2_xor2_1 _35744_ (.B(_09999_),
    .A(_09998_),
    .X(_10000_));
 sg13g2_o21ai_1 _35745_ (.B1(net4397),
    .Y(_10001_),
    .A1(net4697),
    .A2(_09997_));
 sg13g2_a21oi_1 _35746_ (.A1(net4697),
    .A2(_10000_),
    .Y(_10002_),
    .B1(_10001_));
 sg13g2_o21ai_1 _35747_ (.B1(net5595),
    .Y(_10003_),
    .A1(net4397),
    .A2(_09981_));
 sg13g2_o21ai_1 _35748_ (.B1(_09992_),
    .Y(_00796_),
    .A1(_10002_),
    .A2(_10003_));
 sg13g2_o21ai_1 _35749_ (.B1(_09343_),
    .Y(_10004_),
    .A1(_09325_),
    .A2(_09995_));
 sg13g2_nor3_1 _35750_ (.A(_09325_),
    .B(_09343_),
    .C(_09995_),
    .Y(_10005_));
 sg13g2_nor2_1 _35751_ (.A(net5357),
    .B(_10005_),
    .Y(_10006_));
 sg13g2_a22oi_1 _35752_ (.Y(_10007_),
    .B1(_10004_),
    .B2(_10006_),
    .A2(_09334_),
    .A1(net5357));
 sg13g2_nand2_1 _35753_ (.Y(_10008_),
    .A(net4592),
    .B(_10007_));
 sg13g2_xnor2_1 _35754_ (.Y(_10009_),
    .A(net4592),
    .B(_10007_));
 sg13g2_and2_1 _35755_ (.A(_09983_),
    .B(_09998_),
    .X(_10010_));
 sg13g2_and4_1 _35756_ (.A(_09950_),
    .B(_09971_),
    .C(_09983_),
    .D(_09998_),
    .X(_10011_));
 sg13g2_o21ai_1 _35757_ (.B1(_09982_),
    .Y(_10012_),
    .A1(net4541),
    .A2(_09997_));
 sg13g2_a221oi_1 _35758_ (.B2(_09953_),
    .C1(_10012_),
    .B1(_10011_),
    .A1(_09984_),
    .Y(_10013_),
    .A2(_10010_));
 sg13g2_and4_1 _35759_ (.A(_09921_),
    .B(_09938_),
    .C(_09954_),
    .D(_10011_),
    .X(_10014_));
 sg13g2_nand2_1 _35760_ (.Y(_10015_),
    .A(_09892_),
    .B(_10014_));
 sg13g2_and2_1 _35761_ (.A(_10013_),
    .B(_10015_),
    .X(_10016_));
 sg13g2_a21oi_1 _35762_ (.A1(_10009_),
    .A2(_10016_),
    .Y(_10017_),
    .B1(net4654));
 sg13g2_o21ai_1 _35763_ (.B1(_10017_),
    .Y(_10018_),
    .A1(_10009_),
    .A2(_10016_));
 sg13g2_nand2_1 _35764_ (.Y(_10019_),
    .A(net4654),
    .B(_10007_));
 sg13g2_nand3_1 _35765_ (.B(_10018_),
    .C(_10019_),
    .A(net4397),
    .Y(_10020_));
 sg13g2_a21oi_1 _35766_ (.A1(net4356),
    .A2(_09997_),
    .Y(_10021_),
    .B1(net5538));
 sg13g2_a22oi_1 _35767_ (.Y(_10022_),
    .B1(_10020_),
    .B2(_10021_),
    .A2(net4152),
    .A1(net3055));
 sg13g2_inv_1 _35768_ (.Y(_00797_),
    .A(_10022_));
 sg13g2_nand2_1 _35769_ (.Y(_10023_),
    .A(net2473),
    .B(net4152));
 sg13g2_o21ai_1 _35770_ (.B1(_09342_),
    .Y(_10024_),
    .A1(_09335_),
    .A2(_09995_));
 sg13g2_xnor2_1 _35771_ (.Y(_10025_),
    .A(_09317_),
    .B(_10024_));
 sg13g2_nor2_1 _35772_ (.A(net5357),
    .B(_10025_),
    .Y(_10026_));
 sg13g2_a21oi_2 _35773_ (.B1(_10026_),
    .Y(_10027_),
    .A2(_09314_),
    .A1(net5357));
 sg13g2_inv_1 _35774_ (.Y(_10028_),
    .A(_10027_));
 sg13g2_nand2_1 _35775_ (.Y(_10029_),
    .A(net4654),
    .B(_10027_));
 sg13g2_xnor2_1 _35776_ (.Y(_10030_),
    .A(net4543),
    .B(_10027_));
 sg13g2_o21ai_1 _35777_ (.B1(_10008_),
    .Y(_10031_),
    .A1(_10009_),
    .A2(_10016_));
 sg13g2_a21oi_1 _35778_ (.A1(_10030_),
    .A2(_10031_),
    .Y(_10032_),
    .B1(net4654));
 sg13g2_o21ai_1 _35779_ (.B1(_10032_),
    .Y(_10033_),
    .A1(_10030_),
    .A2(_10031_));
 sg13g2_a21oi_1 _35780_ (.A1(_10029_),
    .A2(_10033_),
    .Y(_10034_),
    .B1(net4356));
 sg13g2_o21ai_1 _35781_ (.B1(net5595),
    .Y(_10035_),
    .A1(net4399),
    .A2(_10007_));
 sg13g2_o21ai_1 _35782_ (.B1(_10023_),
    .Y(_00798_),
    .A1(_10034_),
    .A2(_10035_));
 sg13g2_nand2_1 _35783_ (.Y(_10036_),
    .A(net4356),
    .B(_10027_));
 sg13g2_o21ai_1 _35784_ (.B1(_09315_),
    .Y(_10037_),
    .A1(_09317_),
    .A2(_10024_));
 sg13g2_xnor2_1 _35785_ (.Y(_10038_),
    .A(_09309_),
    .B(_10037_));
 sg13g2_nand2_1 _35786_ (.Y(_10039_),
    .A(net5398),
    .B(_10038_));
 sg13g2_o21ai_1 _35787_ (.B1(_10039_),
    .Y(_10040_),
    .A1(net5398),
    .A2(_09308_));
 sg13g2_nand2_1 _35788_ (.Y(_10041_),
    .A(net4654),
    .B(_10040_));
 sg13g2_nand3b_1 _35789_ (.B(net4629),
    .C(net4637),
    .Y(_10042_),
    .A_N(_10040_));
 sg13g2_o21ai_1 _35790_ (.B1(_10040_),
    .Y(_10043_),
    .A1(net4634),
    .A2(net4635));
 sg13g2_and2_1 _35791_ (.A(_10042_),
    .B(_10043_),
    .X(_10044_));
 sg13g2_inv_1 _35792_ (.Y(_10045_),
    .A(_10044_));
 sg13g2_o21ai_1 _35793_ (.B1(net4592),
    .Y(_10046_),
    .A1(_10007_),
    .A2(_10028_));
 sg13g2_o21ai_1 _35794_ (.B1(_10046_),
    .Y(_10047_),
    .A1(_10009_),
    .A2(_10016_));
 sg13g2_o21ai_1 _35795_ (.B1(_10047_),
    .Y(_10048_),
    .A1(net4592),
    .A2(_10028_));
 sg13g2_xnor2_1 _35796_ (.Y(_10049_),
    .A(_10044_),
    .B(_10048_));
 sg13g2_o21ai_1 _35797_ (.B1(_10041_),
    .Y(_10050_),
    .A1(net4654),
    .A2(_10049_));
 sg13g2_a21oi_1 _35798_ (.A1(net4401),
    .A2(_10050_),
    .Y(_10051_),
    .B1(net5539));
 sg13g2_a22oi_1 _35799_ (.Y(_10052_),
    .B1(_10036_),
    .B2(_10051_),
    .A2(net4154),
    .A1(net1612));
 sg13g2_inv_1 _35800_ (.Y(_00799_),
    .A(_10052_));
 sg13g2_nand2_1 _35801_ (.Y(_10053_),
    .A(net5357),
    .B(_09285_));
 sg13g2_nand2b_1 _35802_ (.Y(_10054_),
    .B(_09344_),
    .A_N(_09994_));
 sg13g2_and2_1 _35803_ (.A(_09338_),
    .B(_10054_),
    .X(_10055_));
 sg13g2_or2_1 _35804_ (.X(_10056_),
    .B(_10055_),
    .A(_09296_));
 sg13g2_xnor2_1 _35805_ (.Y(_10057_),
    .A(_09296_),
    .B(_10055_));
 sg13g2_o21ai_1 _35806_ (.B1(_10053_),
    .Y(_10058_),
    .A1(net5357),
    .A2(_10057_));
 sg13g2_nand3_1 _35807_ (.B(net4637),
    .C(_10058_),
    .A(net4629),
    .Y(_10059_));
 sg13g2_a21o_1 _35808_ (.A2(net4637),
    .A1(net4629),
    .B1(_10058_),
    .X(_10060_));
 sg13g2_and2_1 _35809_ (.A(_10059_),
    .B(_10060_),
    .X(_10061_));
 sg13g2_o21ai_1 _35810_ (.B1(_10042_),
    .Y(_10062_),
    .A1(_10045_),
    .A2(_10048_));
 sg13g2_xnor2_1 _35811_ (.Y(_10063_),
    .A(_10061_),
    .B(_10062_));
 sg13g2_a21oi_1 _35812_ (.A1(net4654),
    .A2(_10058_),
    .Y(_10064_),
    .B1(net4357));
 sg13g2_o21ai_1 _35813_ (.B1(_10064_),
    .Y(_10065_),
    .A1(net4654),
    .A2(_10063_));
 sg13g2_a21oi_1 _35814_ (.A1(net4357),
    .A2(_10040_),
    .Y(_10066_),
    .B1(net5539));
 sg13g2_a22oi_1 _35815_ (.Y(_10067_),
    .B1(_10065_),
    .B2(_10066_),
    .A2(net4154),
    .A1(net2840));
 sg13g2_inv_1 _35816_ (.Y(_00800_),
    .A(_10067_));
 sg13g2_nor2_1 _35817_ (.A(net5398),
    .B(_09294_),
    .Y(_10068_));
 sg13g2_nand2_1 _35818_ (.Y(_10069_),
    .A(_09286_),
    .B(_10056_));
 sg13g2_xnor2_1 _35819_ (.Y(_10070_),
    .A(_09298_),
    .B(_10069_));
 sg13g2_a21oi_2 _35820_ (.B1(_10068_),
    .Y(_10071_),
    .A2(_10070_),
    .A1(net5398));
 sg13g2_nand2_1 _35821_ (.Y(_10072_),
    .A(net4592),
    .B(_10071_));
 sg13g2_xnor2_1 _35822_ (.Y(_10073_),
    .A(net4592),
    .B(_10071_));
 sg13g2_nand4_1 _35823_ (.B(_10043_),
    .C(_10059_),
    .A(_10042_),
    .Y(_10074_),
    .D(_10060_));
 sg13g2_and2_1 _35824_ (.A(_10042_),
    .B(_10059_),
    .X(_10075_));
 sg13g2_o21ai_1 _35825_ (.B1(_10075_),
    .Y(_10076_),
    .A1(_10046_),
    .A2(_10074_));
 sg13g2_nor3_1 _35826_ (.A(_10009_),
    .B(_10030_),
    .C(_10074_),
    .Y(_10077_));
 sg13g2_nor2b_1 _35827_ (.A(_10016_),
    .B_N(_10077_),
    .Y(_10078_));
 sg13g2_nor2_1 _35828_ (.A(_10076_),
    .B(_10078_),
    .Y(_10079_));
 sg13g2_nor2_1 _35829_ (.A(_10073_),
    .B(_10079_),
    .Y(_10080_));
 sg13g2_and2_1 _35830_ (.A(_10073_),
    .B(_10079_),
    .X(_10081_));
 sg13g2_o21ai_1 _35831_ (.B1(net4698),
    .Y(_10082_),
    .A1(_10080_),
    .A2(_10081_));
 sg13g2_o21ai_1 _35832_ (.B1(_10082_),
    .Y(_10083_),
    .A1(net4698),
    .A2(_10071_));
 sg13g2_o21ai_1 _35833_ (.B1(net5596),
    .Y(_10084_),
    .A1(net4401),
    .A2(_10058_));
 sg13g2_a21oi_1 _35834_ (.A1(net4401),
    .A2(_10083_),
    .Y(_10085_),
    .B1(_10084_));
 sg13g2_a21o_1 _35835_ (.A2(net4154),
    .A1(net2970),
    .B1(_10085_),
    .X(_00801_));
 sg13g2_a21oi_1 _35836_ (.A1(_09295_),
    .A2(_10056_),
    .Y(_10086_),
    .B1(_09297_));
 sg13g2_o21ai_1 _35837_ (.B1(net5398),
    .Y(_10087_),
    .A1(_09270_),
    .A2(_10086_));
 sg13g2_a21oi_1 _35838_ (.A1(_09270_),
    .A2(_10086_),
    .Y(_10088_),
    .B1(_10087_));
 sg13g2_a21oi_2 _35839_ (.B1(_10088_),
    .Y(_10089_),
    .A2(_09267_),
    .A1(net5357));
 sg13g2_nand2_1 _35840_ (.Y(_10090_),
    .A(net4655),
    .B(_10089_));
 sg13g2_nand2_1 _35841_ (.Y(_10091_),
    .A(net4543),
    .B(_10089_));
 sg13g2_xnor2_1 _35842_ (.Y(_10092_),
    .A(net4543),
    .B(_10089_));
 sg13g2_o21ai_1 _35843_ (.B1(_10072_),
    .Y(_10093_),
    .A1(_10073_),
    .A2(_10079_));
 sg13g2_xnor2_1 _35844_ (.Y(_10094_),
    .A(_10092_),
    .B(_10093_));
 sg13g2_o21ai_1 _35845_ (.B1(_10090_),
    .Y(_10095_),
    .A1(net4655),
    .A2(_10094_));
 sg13g2_o21ai_1 _35846_ (.B1(net5596),
    .Y(_10096_),
    .A1(net4401),
    .A2(_10071_));
 sg13g2_a21oi_1 _35847_ (.A1(net4401),
    .A2(_10095_),
    .Y(_10097_),
    .B1(_10096_));
 sg13g2_a21o_1 _35848_ (.A2(net4154),
    .A1(net1597),
    .B1(_10097_),
    .X(_00802_));
 sg13g2_nand2_1 _35849_ (.Y(_10098_),
    .A(net4362),
    .B(_10089_));
 sg13g2_nor2_1 _35850_ (.A(net5398),
    .B(_09278_),
    .Y(_10099_));
 sg13g2_a21o_1 _35851_ (.A2(_10086_),
    .A1(_09270_),
    .B1(_09269_),
    .X(_10100_));
 sg13g2_xnor2_1 _35852_ (.Y(_10101_),
    .A(_09279_),
    .B(_10100_));
 sg13g2_a21oi_2 _35853_ (.B1(_10099_),
    .Y(_10102_),
    .A2(_10101_),
    .A1(net5398));
 sg13g2_nand2_1 _35854_ (.Y(_10103_),
    .A(net4592),
    .B(_10102_));
 sg13g2_xnor2_1 _35855_ (.Y(_10104_),
    .A(net4592),
    .B(_10102_));
 sg13g2_o21ai_1 _35856_ (.B1(_10072_),
    .Y(_10105_),
    .A1(net4543),
    .A2(_10089_));
 sg13g2_o21ai_1 _35857_ (.B1(_10091_),
    .Y(_10106_),
    .A1(_10080_),
    .A2(_10105_));
 sg13g2_xnor2_1 _35858_ (.Y(_10107_),
    .A(_10104_),
    .B(_10106_));
 sg13g2_nand2_1 _35859_ (.Y(_10108_),
    .A(net4698),
    .B(_10107_));
 sg13g2_o21ai_1 _35860_ (.B1(_10108_),
    .Y(_10109_),
    .A1(net4698),
    .A2(_10102_));
 sg13g2_a21oi_1 _35861_ (.A1(net4401),
    .A2(_10109_),
    .Y(_10110_),
    .B1(net5539));
 sg13g2_a22oi_1 _35862_ (.Y(_10111_),
    .B1(_10098_),
    .B2(_10110_),
    .A2(net4154),
    .A1(net2273));
 sg13g2_inv_1 _35863_ (.Y(_00803_),
    .A(_10111_));
 sg13g2_nand2_1 _35864_ (.Y(_10112_),
    .A(net2055),
    .B(net4154));
 sg13g2_nor2_1 _35865_ (.A(net5401),
    .B(_09132_),
    .Y(_10113_));
 sg13g2_nand2b_1 _35866_ (.Y(_10114_),
    .B(_09591_),
    .A_N(_09593_));
 sg13g2_xnor2_1 _35867_ (.Y(_10115_),
    .A(_09591_),
    .B(_09593_));
 sg13g2_a21oi_2 _35868_ (.B1(_10113_),
    .Y(_10116_),
    .A2(_10115_),
    .A1(net5401));
 sg13g2_nand2_1 _35869_ (.Y(_10117_),
    .A(net4655),
    .B(_10116_));
 sg13g2_xnor2_1 _35870_ (.Y(_10118_),
    .A(net4543),
    .B(_10116_));
 sg13g2_o21ai_1 _35871_ (.B1(_10103_),
    .Y(_10119_),
    .A1(_10104_),
    .A2(_10106_));
 sg13g2_xnor2_1 _35872_ (.Y(_10120_),
    .A(_10118_),
    .B(_10119_));
 sg13g2_o21ai_1 _35873_ (.B1(_10117_),
    .Y(_10121_),
    .A1(net4655),
    .A2(_10120_));
 sg13g2_a21oi_1 _35874_ (.A1(net4401),
    .A2(_10121_),
    .Y(_10122_),
    .B1(net5539));
 sg13g2_o21ai_1 _35875_ (.B1(_10122_),
    .Y(_10123_),
    .A1(net4401),
    .A2(_10102_));
 sg13g2_nand2_1 _35876_ (.Y(_00804_),
    .A(_10112_),
    .B(_10123_));
 sg13g2_nor2_1 _35877_ (.A(net5401),
    .B(_09127_),
    .Y(_10124_));
 sg13g2_o21ai_1 _35878_ (.B1(_10114_),
    .Y(_10125_),
    .A1(net4748),
    .A2(_09132_));
 sg13g2_xnor2_1 _35879_ (.Y(_10126_),
    .A(_09592_),
    .B(_10125_));
 sg13g2_a21oi_2 _35880_ (.B1(_10124_),
    .Y(_10127_),
    .A2(_10126_),
    .A1(net5401));
 sg13g2_nand2_1 _35881_ (.Y(_10128_),
    .A(net4657),
    .B(_10127_));
 sg13g2_nor2_1 _35882_ (.A(_10104_),
    .B(_10118_),
    .Y(_10129_));
 sg13g2_nor4_2 _35883_ (.A(_10073_),
    .B(_10092_),
    .C(_10104_),
    .Y(_10130_),
    .D(_10118_));
 sg13g2_nand2_1 _35884_ (.Y(_10131_),
    .A(_10077_),
    .B(_10130_));
 sg13g2_and3_1 _35885_ (.X(_10132_),
    .A(_10014_),
    .B(_10077_),
    .C(_10130_));
 sg13g2_o21ai_1 _35886_ (.B1(_10103_),
    .Y(_10133_),
    .A1(net4543),
    .A2(_10116_));
 sg13g2_a221oi_1 _35887_ (.B2(_10076_),
    .C1(_10133_),
    .B1(_10130_),
    .A1(_10105_),
    .Y(_10134_),
    .A2(_10129_));
 sg13g2_o21ai_1 _35888_ (.B1(_10134_),
    .Y(_10135_),
    .A1(_10013_),
    .A2(_10131_));
 sg13g2_a21oi_2 _35889_ (.B1(_10135_),
    .Y(_10136_),
    .A2(_10132_),
    .A1(_09892_));
 sg13g2_or2_1 _35890_ (.X(_10137_),
    .B(_10127_),
    .A(net4595));
 sg13g2_xnor2_1 _35891_ (.Y(_10138_),
    .A(net4595),
    .B(_10127_));
 sg13g2_xor2_1 _35892_ (.B(_10138_),
    .A(_10136_),
    .X(_10139_));
 sg13g2_o21ai_1 _35893_ (.B1(_10128_),
    .Y(_10140_),
    .A1(net4657),
    .A2(_10139_));
 sg13g2_nand2_1 _35894_ (.Y(_10141_),
    .A(net4403),
    .B(_10140_));
 sg13g2_a21oi_1 _35895_ (.A1(net4358),
    .A2(_10116_),
    .Y(_10142_),
    .B1(net5547));
 sg13g2_a22oi_1 _35896_ (.Y(_10143_),
    .B1(_10141_),
    .B2(_10142_),
    .A2(net4170),
    .A1(net2130));
 sg13g2_inv_1 _35897_ (.Y(_00805_),
    .A(_10143_));
 sg13g2_nor2_1 _35898_ (.A(net5401),
    .B(_09117_),
    .Y(_10144_));
 sg13g2_nand2_1 _35899_ (.Y(_10145_),
    .A(_09591_),
    .B(_09594_));
 sg13g2_a21o_1 _35900_ (.A2(_10145_),
    .A1(_09133_),
    .B1(_09118_),
    .X(_10146_));
 sg13g2_nand3_1 _35901_ (.B(_09133_),
    .C(_10145_),
    .A(_09118_),
    .Y(_10147_));
 sg13g2_nand3_1 _35902_ (.B(_10146_),
    .C(_10147_),
    .A(net5401),
    .Y(_10148_));
 sg13g2_nor2b_2 _35903_ (.A(_10144_),
    .B_N(_10148_),
    .Y(_10149_));
 sg13g2_nand2_1 _35904_ (.Y(_10150_),
    .A(net4657),
    .B(_10149_));
 sg13g2_o21ai_1 _35905_ (.B1(_10137_),
    .Y(_10151_),
    .A1(_10136_),
    .A2(_10138_));
 sg13g2_nand2_1 _35906_ (.Y(_10152_),
    .A(net4545),
    .B(_10149_));
 sg13g2_xnor2_1 _35907_ (.Y(_10153_),
    .A(net4545),
    .B(_10149_));
 sg13g2_xnor2_1 _35908_ (.Y(_10154_),
    .A(_10151_),
    .B(_10153_));
 sg13g2_o21ai_1 _35909_ (.B1(_10150_),
    .Y(_10155_),
    .A1(net4657),
    .A2(_10154_));
 sg13g2_nand2_1 _35910_ (.Y(_10156_),
    .A(net4403),
    .B(_10155_));
 sg13g2_a21oi_1 _35911_ (.A1(net4358),
    .A2(_10127_),
    .Y(_10157_),
    .B1(net5547));
 sg13g2_a22oi_1 _35912_ (.Y(_10158_),
    .B1(_10156_),
    .B2(_10157_),
    .A2(net4170),
    .A1(net2689));
 sg13g2_inv_1 _35913_ (.Y(_00806_),
    .A(_10158_));
 sg13g2_nand2_1 _35914_ (.Y(_10159_),
    .A(net5359),
    .B(_09110_));
 sg13g2_o21ai_1 _35915_ (.B1(_10146_),
    .Y(_10160_),
    .A1(net4803),
    .A2(_09117_));
 sg13g2_xnor2_1 _35916_ (.Y(_10161_),
    .A(_09111_),
    .B(_10160_));
 sg13g2_o21ai_1 _35917_ (.B1(_10159_),
    .Y(_10162_),
    .A1(net5359),
    .A2(_10161_));
 sg13g2_nand2_1 _35918_ (.Y(_10163_),
    .A(net4657),
    .B(_10162_));
 sg13g2_nand3b_1 _35919_ (.B(net4629),
    .C(net4637),
    .Y(_10164_),
    .A_N(_10162_));
 sg13g2_o21ai_1 _35920_ (.B1(_10162_),
    .Y(_10165_),
    .A1(net4634),
    .A2(net4635));
 sg13g2_nand2_1 _35921_ (.Y(_10166_),
    .A(_10164_),
    .B(_10165_));
 sg13g2_a21o_1 _35922_ (.A2(_10127_),
    .A1(net4545),
    .B1(_10149_),
    .X(_10167_));
 sg13g2_o21ai_1 _35923_ (.B1(_10167_),
    .Y(_10168_),
    .A1(_10136_),
    .A2(_10138_));
 sg13g2_nand2_1 _35924_ (.Y(_10169_),
    .A(_10152_),
    .B(_10168_));
 sg13g2_xor2_1 _35925_ (.B(_10169_),
    .A(_10166_),
    .X(_10170_));
 sg13g2_o21ai_1 _35926_ (.B1(_10163_),
    .Y(_10171_),
    .A1(net4657),
    .A2(_10170_));
 sg13g2_nand2_1 _35927_ (.Y(_10172_),
    .A(net4403),
    .B(_10171_));
 sg13g2_a21oi_1 _35928_ (.A1(net4358),
    .A2(_10149_),
    .Y(_10173_),
    .B1(net5547));
 sg13g2_a22oi_1 _35929_ (.Y(_10174_),
    .B1(_10172_),
    .B2(_10173_),
    .A2(net4170),
    .A1(net2984));
 sg13g2_inv_1 _35930_ (.Y(_00807_),
    .A(_10174_));
 sg13g2_and3_1 _35931_ (.X(_10175_),
    .A(_09120_),
    .B(_09591_),
    .C(_09594_));
 sg13g2_o21ai_1 _35932_ (.B1(_09098_),
    .Y(_10176_),
    .A1(_09137_),
    .A2(_10175_));
 sg13g2_or3_1 _35933_ (.A(_09098_),
    .B(_09137_),
    .C(_10175_),
    .X(_10177_));
 sg13g2_and2_1 _35934_ (.A(_10176_),
    .B(_10177_),
    .X(_10178_));
 sg13g2_mux2_1 _35935_ (.A0(_09085_),
    .A1(_10178_),
    .S(net5401),
    .X(_10179_));
 sg13g2_nand3_1 _35936_ (.B(net4637),
    .C(_10179_),
    .A(net4629),
    .Y(_10180_));
 sg13g2_a21o_1 _35937_ (.A2(net4637),
    .A1(net4629),
    .B1(_10179_),
    .X(_10181_));
 sg13g2_and2_1 _35938_ (.A(_10180_),
    .B(_10181_),
    .X(_10182_));
 sg13g2_o21ai_1 _35939_ (.B1(_10164_),
    .Y(_10183_),
    .A1(_10166_),
    .A2(_10169_));
 sg13g2_xnor2_1 _35940_ (.Y(_10184_),
    .A(_10182_),
    .B(_10183_));
 sg13g2_nand2_1 _35941_ (.Y(_10185_),
    .A(net4700),
    .B(_10184_));
 sg13g2_o21ai_1 _35942_ (.B1(_10185_),
    .Y(_10186_),
    .A1(net4700),
    .A2(_10179_));
 sg13g2_nand2_1 _35943_ (.Y(_10187_),
    .A(net4403),
    .B(_10186_));
 sg13g2_a21oi_1 _35944_ (.A1(net4358),
    .A2(_10162_),
    .Y(_10188_),
    .B1(net5547));
 sg13g2_a22oi_1 _35945_ (.Y(_10189_),
    .B1(_10187_),
    .B2(_10188_),
    .A2(net4170),
    .A1(net2588));
 sg13g2_inv_1 _35946_ (.Y(_00808_),
    .A(_10189_));
 sg13g2_nor2_1 _35947_ (.A(net5401),
    .B(_09095_),
    .Y(_10190_));
 sg13g2_nand2_1 _35948_ (.Y(_10191_),
    .A(_09086_),
    .B(_10176_));
 sg13g2_xnor2_1 _35949_ (.Y(_10192_),
    .A(_09100_),
    .B(_10191_));
 sg13g2_a21oi_2 _35950_ (.B1(_10190_),
    .Y(_10193_),
    .A2(_10192_),
    .A1(net5402));
 sg13g2_nand2_1 _35951_ (.Y(_10194_),
    .A(net4595),
    .B(_10193_));
 sg13g2_xnor2_1 _35952_ (.Y(_10195_),
    .A(net4595),
    .B(_10193_));
 sg13g2_nand4_1 _35953_ (.B(_10165_),
    .C(_10180_),
    .A(_10164_),
    .Y(_10196_),
    .D(_10181_));
 sg13g2_and2_1 _35954_ (.A(_10164_),
    .B(_10180_),
    .X(_10197_));
 sg13g2_o21ai_1 _35955_ (.B1(_10197_),
    .Y(_10198_),
    .A1(_10167_),
    .A2(_10196_));
 sg13g2_nor3_1 _35956_ (.A(_10138_),
    .B(_10153_),
    .C(_10196_),
    .Y(_10199_));
 sg13g2_nor2b_1 _35957_ (.A(_10136_),
    .B_N(_10199_),
    .Y(_10200_));
 sg13g2_nor2_1 _35958_ (.A(_10198_),
    .B(_10200_),
    .Y(_10201_));
 sg13g2_nor2_1 _35959_ (.A(_10195_),
    .B(_10201_),
    .Y(_10202_));
 sg13g2_xnor2_1 _35960_ (.Y(_10203_),
    .A(_10195_),
    .B(_10201_));
 sg13g2_nand2_1 _35961_ (.Y(_10204_),
    .A(net4700),
    .B(_10203_));
 sg13g2_o21ai_1 _35962_ (.B1(_10204_),
    .Y(_10205_),
    .A1(net4700),
    .A2(_10193_));
 sg13g2_o21ai_1 _35963_ (.B1(net5598),
    .Y(_10206_),
    .A1(net4403),
    .A2(_10179_));
 sg13g2_a21oi_1 _35964_ (.A1(net4403),
    .A2(_10205_),
    .Y(_10207_),
    .B1(_10206_));
 sg13g2_a21o_1 _35965_ (.A2(net4171),
    .A1(net2581),
    .B1(_10207_),
    .X(_00809_));
 sg13g2_nand2_1 _35966_ (.Y(_10208_),
    .A(_09096_),
    .B(_10176_));
 sg13g2_nand3_1 _35967_ (.B(_09099_),
    .C(_10208_),
    .A(_09070_),
    .Y(_10209_));
 sg13g2_a21oi_1 _35968_ (.A1(_09099_),
    .A2(_10208_),
    .Y(_10210_),
    .B1(_09070_));
 sg13g2_nor2_1 _35969_ (.A(net5359),
    .B(_10210_),
    .Y(_10211_));
 sg13g2_a22oi_1 _35970_ (.Y(_10212_),
    .B1(_10209_),
    .B2(_10211_),
    .A2(_09068_),
    .A1(net5359));
 sg13g2_nand2_1 _35971_ (.Y(_10213_),
    .A(net4657),
    .B(_10212_));
 sg13g2_nand2_1 _35972_ (.Y(_10214_),
    .A(net4545),
    .B(_10212_));
 sg13g2_xnor2_1 _35973_ (.Y(_10215_),
    .A(net4545),
    .B(_10212_));
 sg13g2_a21oi_1 _35974_ (.A1(net4595),
    .A2(_10193_),
    .Y(_10216_),
    .B1(_10202_));
 sg13g2_xor2_1 _35975_ (.B(_10216_),
    .A(_10215_),
    .X(_10217_));
 sg13g2_o21ai_1 _35976_ (.B1(_10213_),
    .Y(_10218_),
    .A1(net4657),
    .A2(_10217_));
 sg13g2_o21ai_1 _35977_ (.B1(net5598),
    .Y(_10219_),
    .A1(net4404),
    .A2(_10193_));
 sg13g2_a21oi_1 _35978_ (.A1(net4404),
    .A2(_10218_),
    .Y(_10220_),
    .B1(_10219_));
 sg13g2_a21o_1 _35979_ (.A2(net4170),
    .A1(net3217),
    .B1(_10220_),
    .X(_00810_));
 sg13g2_nand2_1 _35980_ (.Y(_10221_),
    .A(net4358),
    .B(_10212_));
 sg13g2_or2_1 _35981_ (.X(_10222_),
    .B(_09078_),
    .A(net5402));
 sg13g2_nand2_1 _35982_ (.Y(_10223_),
    .A(_09069_),
    .B(_10209_));
 sg13g2_xor2_1 _35983_ (.B(_10223_),
    .A(_09079_),
    .X(_10224_));
 sg13g2_o21ai_1 _35984_ (.B1(_10222_),
    .Y(_10225_),
    .A1(net5359),
    .A2(_10224_));
 sg13g2_nand2_1 _35985_ (.Y(_10226_),
    .A(net4660),
    .B(_10225_));
 sg13g2_or2_1 _35986_ (.X(_10227_),
    .B(_10225_),
    .A(net4545));
 sg13g2_xnor2_1 _35987_ (.Y(_10228_),
    .A(net4545),
    .B(_10225_));
 sg13g2_o21ai_1 _35988_ (.B1(_10194_),
    .Y(_10229_),
    .A1(net4545),
    .A2(_10212_));
 sg13g2_o21ai_1 _35989_ (.B1(_10214_),
    .Y(_10230_),
    .A1(_10202_),
    .A2(_10229_));
 sg13g2_xor2_1 _35990_ (.B(_10230_),
    .A(_10228_),
    .X(_10231_));
 sg13g2_o21ai_1 _35991_ (.B1(_10226_),
    .Y(_10232_),
    .A1(net4660),
    .A2(_10231_));
 sg13g2_a21oi_1 _35992_ (.A1(net4403),
    .A2(_10232_),
    .Y(_10233_),
    .B1(net5547));
 sg13g2_a22oi_1 _35993_ (.Y(_10234_),
    .B1(_10221_),
    .B2(_10233_),
    .A2(net4170),
    .A1(net2864));
 sg13g2_inv_1 _35994_ (.Y(_00811_),
    .A(_10234_));
 sg13g2_nand2_1 _35995_ (.Y(_10235_),
    .A(net5361),
    .B(_09223_));
 sg13g2_a221oi_1 _35996_ (.B2(_09590_),
    .C1(_09597_),
    .B1(_09581_),
    .A1(_09340_),
    .Y(_10236_),
    .A2(_09345_));
 sg13g2_nor2_1 _35997_ (.A(_09141_),
    .B(_10236_),
    .Y(_10237_));
 sg13g2_nor2_1 _35998_ (.A(_09225_),
    .B(_10237_),
    .Y(_10238_));
 sg13g2_xnor2_1 _35999_ (.Y(_10239_),
    .A(_09225_),
    .B(_10237_));
 sg13g2_o21ai_1 _36000_ (.B1(_10235_),
    .Y(_10240_),
    .A1(net5361),
    .A2(_10239_));
 sg13g2_nand2_1 _36001_ (.Y(_10241_),
    .A(net4595),
    .B(_10240_));
 sg13g2_xnor2_1 _36002_ (.Y(_10242_),
    .A(net4595),
    .B(_10240_));
 sg13g2_o21ai_1 _36003_ (.B1(_10227_),
    .Y(_10243_),
    .A1(_10228_),
    .A2(_10230_));
 sg13g2_xor2_1 _36004_ (.B(_10243_),
    .A(_10242_),
    .X(_10244_));
 sg13g2_nand2_1 _36005_ (.Y(_10245_),
    .A(net4700),
    .B(_10244_));
 sg13g2_o21ai_1 _36006_ (.B1(_10245_),
    .Y(_10246_),
    .A1(net4700),
    .A2(_10240_));
 sg13g2_nand2_1 _36007_ (.Y(_10247_),
    .A(net4403),
    .B(_10246_));
 sg13g2_a21oi_1 _36008_ (.A1(net4358),
    .A2(_10225_),
    .Y(_10248_),
    .B1(net5547));
 sg13g2_a22oi_1 _36009_ (.Y(_10249_),
    .B1(_10247_),
    .B2(_10248_),
    .A2(net4170),
    .A1(net2268));
 sg13g2_inv_1 _36010_ (.Y(_00812_),
    .A(_10249_));
 sg13g2_nor2_1 _36011_ (.A(_09224_),
    .B(_10238_),
    .Y(_10250_));
 sg13g2_xnor2_1 _36012_ (.Y(_10251_),
    .A(_09218_),
    .B(_10250_));
 sg13g2_nor2_1 _36013_ (.A(net5361),
    .B(_10251_),
    .Y(_10252_));
 sg13g2_a21oi_2 _36014_ (.B1(_10252_),
    .Y(_10253_),
    .A2(_09215_),
    .A1(net5361));
 sg13g2_nand2_1 _36015_ (.Y(_10254_),
    .A(net4597),
    .B(_10253_));
 sg13g2_xnor2_1 _36016_ (.Y(_10255_),
    .A(net4597),
    .B(_10253_));
 sg13g2_nor2_1 _36017_ (.A(_10228_),
    .B(_10242_),
    .Y(_10256_));
 sg13g2_nor4_1 _36018_ (.A(_10195_),
    .B(_10215_),
    .C(_10228_),
    .D(_10242_),
    .Y(_10257_));
 sg13g2_nand2_1 _36019_ (.Y(_10258_),
    .A(_10227_),
    .B(_10241_));
 sg13g2_a221oi_1 _36020_ (.B2(_10198_),
    .C1(_10258_),
    .B1(_10257_),
    .A1(_10229_),
    .Y(_10259_),
    .A2(_10256_));
 sg13g2_nand2_2 _36021_ (.Y(_10260_),
    .A(_10199_),
    .B(_10257_));
 sg13g2_o21ai_1 _36022_ (.B1(_10259_),
    .Y(_10261_),
    .A1(_10136_),
    .A2(_10260_));
 sg13g2_nand2b_1 _36023_ (.Y(_10262_),
    .B(_10261_),
    .A_N(_10255_));
 sg13g2_nand2b_1 _36024_ (.Y(_10263_),
    .B(_10255_),
    .A_N(_10261_));
 sg13g2_a21o_1 _36025_ (.A2(_10263_),
    .A1(_10262_),
    .B1(net4662),
    .X(_10264_));
 sg13g2_o21ai_1 _36026_ (.B1(_10264_),
    .Y(_10265_),
    .A1(net4701),
    .A2(_10253_));
 sg13g2_o21ai_1 _36027_ (.B1(net5597),
    .Y(_10266_),
    .A1(net4405),
    .A2(_10240_));
 sg13g2_a21oi_1 _36028_ (.A1(net4405),
    .A2(_10265_),
    .Y(_10267_),
    .B1(_10266_));
 sg13g2_a21o_1 _36029_ (.A2(net4172),
    .A1(net2261),
    .B1(_10267_),
    .X(_00813_));
 sg13g2_nor2_1 _36030_ (.A(net5405),
    .B(_09195_),
    .Y(_10268_));
 sg13g2_o21ai_1 _36031_ (.B1(_09230_),
    .Y(_10269_),
    .A1(_09225_),
    .A2(_10237_));
 sg13g2_nand3_1 _36032_ (.B(_09217_),
    .C(_10269_),
    .A(_09196_),
    .Y(_10270_));
 sg13g2_a21oi_1 _36033_ (.A1(_09217_),
    .A2(_10269_),
    .Y(_10271_),
    .B1(_09196_));
 sg13g2_nor2_1 _36034_ (.A(net5361),
    .B(_10271_),
    .Y(_10272_));
 sg13g2_a21oi_2 _36035_ (.B1(_10268_),
    .Y(_10273_),
    .A2(_10272_),
    .A1(_10270_));
 sg13g2_inv_1 _36036_ (.Y(_10274_),
    .A(_10273_));
 sg13g2_nand2_1 _36037_ (.Y(_10275_),
    .A(net4662),
    .B(_10273_));
 sg13g2_xnor2_1 _36038_ (.Y(_10276_),
    .A(net4547),
    .B(_10273_));
 sg13g2_nand2_1 _36039_ (.Y(_10277_),
    .A(_10254_),
    .B(_10262_));
 sg13g2_xnor2_1 _36040_ (.Y(_10278_),
    .A(_10276_),
    .B(_10277_));
 sg13g2_o21ai_1 _36041_ (.B1(_10275_),
    .Y(_10279_),
    .A1(net4662),
    .A2(_10278_));
 sg13g2_o21ai_1 _36042_ (.B1(net5597),
    .Y(_10280_),
    .A1(net4405),
    .A2(_10253_));
 sg13g2_a21oi_1 _36043_ (.A1(net4405),
    .A2(_10279_),
    .Y(_10281_),
    .B1(_10280_));
 sg13g2_a21o_1 _36044_ (.A2(net4172),
    .A1(net2885),
    .B1(_10281_),
    .X(_00814_));
 sg13g2_and2_1 _36045_ (.A(net5361),
    .B(_09204_),
    .X(_10282_));
 sg13g2_o21ai_1 _36046_ (.B1(_10270_),
    .Y(_10283_),
    .A1(net4805),
    .A2(_09195_));
 sg13g2_xnor2_1 _36047_ (.Y(_10284_),
    .A(_09205_),
    .B(_10283_));
 sg13g2_a21oi_2 _36048_ (.B1(_10282_),
    .Y(_10285_),
    .A2(_10284_),
    .A1(net5405));
 sg13g2_nand3_1 _36049_ (.B(net4637),
    .C(_10285_),
    .A(net4629),
    .Y(_10286_));
 sg13g2_a21o_1 _36050_ (.A2(net4638),
    .A1(net4630),
    .B1(_10285_),
    .X(_10287_));
 sg13g2_and2_1 _36051_ (.A(_10286_),
    .B(_10287_),
    .X(_10288_));
 sg13g2_o21ai_1 _36052_ (.B1(net4597),
    .Y(_10289_),
    .A1(_10253_),
    .A2(_10274_));
 sg13g2_a22oi_1 _36053_ (.Y(_10290_),
    .B1(_10289_),
    .B2(_10262_),
    .A2(_10273_),
    .A1(net4547));
 sg13g2_nand2_1 _36054_ (.Y(_10291_),
    .A(_10288_),
    .B(_10290_));
 sg13g2_xnor2_1 _36055_ (.Y(_10292_),
    .A(_10288_),
    .B(_10290_));
 sg13g2_nand2_1 _36056_ (.Y(_10293_),
    .A(net4701),
    .B(_10292_));
 sg13g2_o21ai_1 _36057_ (.B1(_10293_),
    .Y(_10294_),
    .A1(net4701),
    .A2(_10285_));
 sg13g2_nand2_1 _36058_ (.Y(_10295_),
    .A(net4405),
    .B(_10294_));
 sg13g2_a21oi_1 _36059_ (.A1(net4360),
    .A2(_10273_),
    .Y(_10296_),
    .B1(net5549));
 sg13g2_a22oi_1 _36060_ (.Y(_10297_),
    .B1(_10295_),
    .B2(_10296_),
    .A2(net4172),
    .A1(net2415));
 sg13g2_inv_1 _36061_ (.Y(_00815_),
    .A(_10297_));
 sg13g2_o21ai_1 _36062_ (.B1(_09227_),
    .Y(_10298_),
    .A1(_09141_),
    .A2(_10236_));
 sg13g2_a21o_1 _36063_ (.A2(_10298_),
    .A1(_09233_),
    .B1(_09176_),
    .X(_10299_));
 sg13g2_nand3_1 _36064_ (.B(_09233_),
    .C(_10298_),
    .A(_09176_),
    .Y(_10300_));
 sg13g2_and2_1 _36065_ (.A(net5405),
    .B(_10300_),
    .X(_10301_));
 sg13g2_a22oi_1 _36066_ (.Y(_10302_),
    .B1(_10299_),
    .B2(_10301_),
    .A2(_09172_),
    .A1(net5361));
 sg13g2_inv_1 _36067_ (.Y(_10303_),
    .A(_10302_));
 sg13g2_nand2_1 _36068_ (.Y(_10304_),
    .A(net4662),
    .B(_10302_));
 sg13g2_nand3_1 _36069_ (.B(net4638),
    .C(_10303_),
    .A(net4630),
    .Y(_10305_));
 sg13g2_o21ai_1 _36070_ (.B1(_10302_),
    .Y(_10306_),
    .A1(_09669_),
    .A2(_09672_));
 sg13g2_and2_1 _36071_ (.A(_10305_),
    .B(_10306_),
    .X(_10307_));
 sg13g2_and2_1 _36072_ (.A(_10286_),
    .B(_10291_),
    .X(_10308_));
 sg13g2_xnor2_1 _36073_ (.Y(_10309_),
    .A(_10307_),
    .B(_10308_));
 sg13g2_o21ai_1 _36074_ (.B1(_10304_),
    .Y(_10310_),
    .A1(net4662),
    .A2(_10309_));
 sg13g2_o21ai_1 _36075_ (.B1(net5597),
    .Y(_10311_),
    .A1(net4405),
    .A2(_10285_));
 sg13g2_a21oi_1 _36076_ (.A1(net4405),
    .A2(_10310_),
    .Y(_10312_),
    .B1(_10311_));
 sg13g2_a21o_1 _36077_ (.A2(net4172),
    .A1(net2343),
    .B1(_10312_),
    .X(_00816_));
 sg13g2_nand2_1 _36078_ (.Y(_10313_),
    .A(net2213),
    .B(net4172));
 sg13g2_nand4_1 _36079_ (.B(_10287_),
    .C(_10305_),
    .A(_10286_),
    .Y(_10314_),
    .D(_10306_));
 sg13g2_and2_1 _36080_ (.A(_10286_),
    .B(_10305_),
    .X(_10315_));
 sg13g2_o21ai_1 _36081_ (.B1(_10315_),
    .Y(_10316_),
    .A1(_10289_),
    .A2(_10314_));
 sg13g2_or3_1 _36082_ (.A(_10255_),
    .B(_10276_),
    .C(_10314_),
    .X(_10317_));
 sg13g2_nor2b_1 _36083_ (.A(_10317_),
    .B_N(_10261_),
    .Y(_10318_));
 sg13g2_nor2_1 _36084_ (.A(_10316_),
    .B(_10318_),
    .Y(_10319_));
 sg13g2_nand2_1 _36085_ (.Y(_10320_),
    .A(_09174_),
    .B(_10299_));
 sg13g2_a21o_1 _36086_ (.A2(_10299_),
    .A1(_09174_),
    .B1(_09186_),
    .X(_10321_));
 sg13g2_o21ai_1 _36087_ (.B1(net5405),
    .Y(_10322_),
    .A1(_09187_),
    .A2(_10320_));
 sg13g2_a21oi_1 _36088_ (.A1(_09187_),
    .A2(_10320_),
    .Y(_10323_),
    .B1(_10322_));
 sg13g2_a21oi_2 _36089_ (.B1(_10323_),
    .Y(_10324_),
    .A2(_09184_),
    .A1(net5362));
 sg13g2_nor2_1 _36090_ (.A(net4547),
    .B(_10324_),
    .Y(_10325_));
 sg13g2_xnor2_1 _36091_ (.Y(_10326_),
    .A(net4597),
    .B(_10324_));
 sg13g2_nor2b_1 _36092_ (.A(_10319_),
    .B_N(_10326_),
    .Y(_10327_));
 sg13g2_xnor2_1 _36093_ (.Y(_10328_),
    .A(_10319_),
    .B(_10326_));
 sg13g2_o21ai_1 _36094_ (.B1(net4407),
    .Y(_10329_),
    .A1(net4701),
    .A2(_10324_));
 sg13g2_a21oi_1 _36095_ (.A1(net4701),
    .A2(_10328_),
    .Y(_10330_),
    .B1(_10329_));
 sg13g2_o21ai_1 _36096_ (.B1(net5597),
    .Y(_10331_),
    .A1(net4407),
    .A2(_10303_));
 sg13g2_o21ai_1 _36097_ (.B1(_10313_),
    .Y(_00817_),
    .A1(_10330_),
    .A2(_10331_));
 sg13g2_a21oi_1 _36098_ (.A1(_09185_),
    .A2(_10321_),
    .Y(_10332_),
    .B1(_09157_));
 sg13g2_and3_1 _36099_ (.X(_10333_),
    .A(_09157_),
    .B(_09185_),
    .C(_10321_));
 sg13g2_nor3_1 _36100_ (.A(net5362),
    .B(_10332_),
    .C(_10333_),
    .Y(_10334_));
 sg13g2_a21oi_2 _36101_ (.B1(_10334_),
    .Y(_10335_),
    .A2(_09155_),
    .A1(net5362));
 sg13g2_nand2_1 _36102_ (.Y(_10336_),
    .A(net4662),
    .B(_10335_));
 sg13g2_nand2_1 _36103_ (.Y(_10337_),
    .A(net4550),
    .B(_10335_));
 sg13g2_xnor2_1 _36104_ (.Y(_10338_),
    .A(net4597),
    .B(_10335_));
 sg13g2_nor2_1 _36105_ (.A(_10325_),
    .B(_10327_),
    .Y(_10339_));
 sg13g2_xnor2_1 _36106_ (.Y(_10340_),
    .A(_10338_),
    .B(_10339_));
 sg13g2_o21ai_1 _36107_ (.B1(_10336_),
    .Y(_10341_),
    .A1(net4665),
    .A2(_10340_));
 sg13g2_nand2_1 _36108_ (.Y(_10342_),
    .A(net4407),
    .B(_10341_));
 sg13g2_a21oi_1 _36109_ (.A1(net4360),
    .A2(_10324_),
    .Y(_10343_),
    .B1(net5549));
 sg13g2_a22oi_1 _36110_ (.Y(_10344_),
    .B1(_10342_),
    .B2(_10343_),
    .A2(net4172),
    .A1(net2407));
 sg13g2_inv_1 _36111_ (.Y(_00818_),
    .A(_10344_));
 sg13g2_o21ai_1 _36112_ (.B1(_09166_),
    .Y(_10345_),
    .A1(_09156_),
    .A2(_10332_));
 sg13g2_nor3_1 _36113_ (.A(_09156_),
    .B(_09166_),
    .C(_10332_),
    .Y(_10346_));
 sg13g2_nor2_1 _36114_ (.A(net5362),
    .B(_10346_),
    .Y(_10347_));
 sg13g2_a22oi_1 _36115_ (.Y(_10348_),
    .B1(_10345_),
    .B2(_10347_),
    .A2(_09165_),
    .A1(net5361));
 sg13g2_nand2_1 _36116_ (.Y(_10349_),
    .A(net4665),
    .B(_10348_));
 sg13g2_nor2_1 _36117_ (.A(net4550),
    .B(_10348_),
    .Y(_10350_));
 sg13g2_xnor2_1 _36118_ (.Y(_10351_),
    .A(net4601),
    .B(_10348_));
 sg13g2_a21oi_1 _36119_ (.A1(_10324_),
    .A2(_10335_),
    .Y(_10352_),
    .B1(net4547));
 sg13g2_o21ai_1 _36120_ (.B1(_10337_),
    .Y(_10353_),
    .A1(_10327_),
    .A2(_10352_));
 sg13g2_inv_1 _36121_ (.Y(_10354_),
    .A(_10353_));
 sg13g2_xnor2_1 _36122_ (.Y(_10355_),
    .A(_10351_),
    .B(_10353_));
 sg13g2_o21ai_1 _36123_ (.B1(_10349_),
    .Y(_10356_),
    .A1(net4665),
    .A2(_10355_));
 sg13g2_nand2_1 _36124_ (.Y(_10357_),
    .A(net4405),
    .B(_10356_));
 sg13g2_a21oi_1 _36125_ (.A1(net4360),
    .A2(_10335_),
    .Y(_10358_),
    .B1(net5549));
 sg13g2_a22oi_1 _36126_ (.Y(_10359_),
    .B1(_10357_),
    .B2(_10358_),
    .A2(net4172),
    .A1(net2104));
 sg13g2_inv_1 _36127_ (.Y(_00819_),
    .A(_10359_));
 sg13g2_nand2_1 _36128_ (.Y(_10360_),
    .A(net5369),
    .B(_09042_));
 sg13g2_a221oi_1 _36129_ (.B2(_09590_),
    .C1(_09599_),
    .B1(_09581_),
    .A1(_09340_),
    .Y(_10361_),
    .A2(_09345_));
 sg13g2_nor2_1 _36130_ (.A(_09237_),
    .B(_10361_),
    .Y(_10362_));
 sg13g2_xnor2_1 _36131_ (.Y(_10363_),
    .A(_09240_),
    .B(_10362_));
 sg13g2_o21ai_1 _36132_ (.B1(_10360_),
    .Y(_10364_),
    .A1(net5369),
    .A2(_10363_));
 sg13g2_xnor2_1 _36133_ (.Y(_10365_),
    .A(net4550),
    .B(_10364_));
 sg13g2_a21oi_1 _36134_ (.A1(_10351_),
    .A2(_10354_),
    .Y(_10366_),
    .B1(_10350_));
 sg13g2_a21oi_1 _36135_ (.A1(_10365_),
    .A2(_10366_),
    .Y(_10367_),
    .B1(net4665));
 sg13g2_o21ai_1 _36136_ (.B1(_10367_),
    .Y(_10368_),
    .A1(_10365_),
    .A2(_10366_));
 sg13g2_o21ai_1 _36137_ (.B1(_10368_),
    .Y(_10369_),
    .A1(net4704),
    .A2(_10364_));
 sg13g2_nand2_1 _36138_ (.Y(_10370_),
    .A(net4410),
    .B(_10369_));
 sg13g2_a21oi_1 _36139_ (.A1(net4360),
    .A2(_10348_),
    .Y(_10371_),
    .B1(net5557));
 sg13g2_a22oi_1 _36140_ (.Y(_10372_),
    .B1(_10370_),
    .B2(_10371_),
    .A2(net4190),
    .A1(net2325));
 sg13g2_inv_1 _36141_ (.Y(_00820_),
    .A(_10372_));
 sg13g2_o21ai_1 _36142_ (.B1(_09043_),
    .Y(_10373_),
    .A1(_09240_),
    .A2(_10362_));
 sg13g2_xnor2_1 _36143_ (.Y(_10374_),
    .A(_09239_),
    .B(_10373_));
 sg13g2_mux2_1 _36144_ (.A0(_09037_),
    .A1(_10374_),
    .S(net5413),
    .X(_10375_));
 sg13g2_xnor2_1 _36145_ (.Y(_10376_),
    .A(net4605),
    .B(_10375_));
 sg13g2_and2_1 _36146_ (.A(_10351_),
    .B(_10365_),
    .X(_10377_));
 sg13g2_and4_1 _36147_ (.A(_10326_),
    .B(_10338_),
    .C(_10351_),
    .D(_10365_),
    .X(_10378_));
 sg13g2_nand2b_1 _36148_ (.Y(_10379_),
    .B(_10378_),
    .A_N(_10317_));
 sg13g2_a21o_1 _36149_ (.A2(_10364_),
    .A1(net4601),
    .B1(_10350_),
    .X(_10380_));
 sg13g2_a221oi_1 _36150_ (.B2(_10316_),
    .C1(_10380_),
    .B1(_10378_),
    .A1(_10352_),
    .Y(_10381_),
    .A2(_10377_));
 sg13g2_o21ai_1 _36151_ (.B1(_10381_),
    .Y(_10382_),
    .A1(_10259_),
    .A2(_10379_));
 sg13g2_or2_1 _36152_ (.X(_10383_),
    .B(_10379_),
    .A(_10260_));
 sg13g2_nor2_1 _36153_ (.A(_10136_),
    .B(_10383_),
    .Y(_10384_));
 sg13g2_nor2_2 _36154_ (.A(_10382_),
    .B(_10384_),
    .Y(_10385_));
 sg13g2_inv_1 _36155_ (.Y(_10386_),
    .A(_10385_));
 sg13g2_nor2_1 _36156_ (.A(_10376_),
    .B(_10385_),
    .Y(_10387_));
 sg13g2_and2_1 _36157_ (.A(_10376_),
    .B(_10385_),
    .X(_10388_));
 sg13g2_o21ai_1 _36158_ (.B1(net4708),
    .Y(_10389_),
    .A1(_10387_),
    .A2(_10388_));
 sg13g2_o21ai_1 _36159_ (.B1(_10389_),
    .Y(_10390_),
    .A1(net4708),
    .A2(_10375_));
 sg13g2_o21ai_1 _36160_ (.B1(net5600),
    .Y(_10391_),
    .A1(net4415),
    .A2(_10364_));
 sg13g2_a21oi_1 _36161_ (.A1(net4418),
    .A2(_10390_),
    .Y(_10392_),
    .B1(_10391_));
 sg13g2_a21o_1 _36162_ (.A2(net4192),
    .A1(net2479),
    .B1(_10392_),
    .X(_00821_));
 sg13g2_o21ai_1 _36163_ (.B1(_09044_),
    .Y(_10393_),
    .A1(_09240_),
    .A2(_10362_));
 sg13g2_and3_1 _36164_ (.X(_10394_),
    .A(_09019_),
    .B(_09238_),
    .C(_10393_));
 sg13g2_a21oi_1 _36165_ (.A1(_09238_),
    .A2(_10393_),
    .Y(_10395_),
    .B1(_09019_));
 sg13g2_nor3_1 _36166_ (.A(net5369),
    .B(_10394_),
    .C(_10395_),
    .Y(_10396_));
 sg13g2_a21o_2 _36167_ (.A2(_09017_),
    .A1(net5369),
    .B1(_10396_),
    .X(_10397_));
 sg13g2_a21oi_1 _36168_ (.A1(net4605),
    .A2(_10375_),
    .Y(_10398_),
    .B1(_10387_));
 sg13g2_xnor2_1 _36169_ (.Y(_10399_),
    .A(net4605),
    .B(_10397_));
 sg13g2_xnor2_1 _36170_ (.Y(_10400_),
    .A(_10398_),
    .B(_10399_));
 sg13g2_nand2_1 _36171_ (.Y(_10401_),
    .A(net4708),
    .B(_10400_));
 sg13g2_o21ai_1 _36172_ (.B1(_10401_),
    .Y(_10402_),
    .A1(net4708),
    .A2(_10397_));
 sg13g2_o21ai_1 _36173_ (.B1(net5603),
    .Y(_10403_),
    .A1(net4418),
    .A2(_10375_));
 sg13g2_a21oi_1 _36174_ (.A1(net4418),
    .A2(_10402_),
    .Y(_10404_),
    .B1(_10403_));
 sg13g2_a21o_1 _36175_ (.A2(net4210),
    .A1(net2881),
    .B1(_10404_),
    .X(_00822_));
 sg13g2_and2_1 _36176_ (.A(net5369),
    .B(_09028_),
    .X(_10405_));
 sg13g2_nor2_1 _36177_ (.A(_09018_),
    .B(_10394_),
    .Y(_10406_));
 sg13g2_xnor2_1 _36178_ (.Y(_10407_),
    .A(_09030_),
    .B(_10406_));
 sg13g2_a21oi_2 _36179_ (.B1(_10405_),
    .Y(_10408_),
    .A2(_10407_),
    .A1(net5413));
 sg13g2_nand3_1 _36180_ (.B(net4641),
    .C(_10408_),
    .A(net4633),
    .Y(_10409_));
 sg13g2_a21o_1 _36181_ (.A2(net4641),
    .A1(net4633),
    .B1(_10408_),
    .X(_10410_));
 sg13g2_nand2_1 _36182_ (.Y(_10411_),
    .A(_10409_),
    .B(_10410_));
 sg13g2_o21ai_1 _36183_ (.B1(net4605),
    .Y(_10412_),
    .A1(_10375_),
    .A2(_10397_));
 sg13g2_o21ai_1 _36184_ (.B1(_10412_),
    .Y(_10413_),
    .A1(_10376_),
    .A2(_10385_));
 sg13g2_o21ai_1 _36185_ (.B1(_10413_),
    .Y(_10414_),
    .A1(net4605),
    .A2(_10397_));
 sg13g2_xnor2_1 _36186_ (.Y(_10415_),
    .A(_10411_),
    .B(_10414_));
 sg13g2_nand2_1 _36187_ (.Y(_10416_),
    .A(net4708),
    .B(_10415_));
 sg13g2_o21ai_1 _36188_ (.B1(_10416_),
    .Y(_10417_),
    .A1(net4708),
    .A2(_10408_));
 sg13g2_o21ai_1 _36189_ (.B1(net5603),
    .Y(_10418_),
    .A1(net4418),
    .A2(_10397_));
 sg13g2_a21oi_1 _36190_ (.A1(net4418),
    .A2(_10417_),
    .Y(_10419_),
    .B1(_10418_));
 sg13g2_a21o_1 _36191_ (.A2(net4210),
    .A1(net2926),
    .B1(_10419_),
    .X(_00823_));
 sg13g2_o21ai_1 _36192_ (.B1(_09241_),
    .Y(_10420_),
    .A1(_09237_),
    .A2(_10361_));
 sg13g2_a21oi_1 _36193_ (.A1(_09047_),
    .A2(_10420_),
    .Y(_10421_),
    .B1(_08997_));
 sg13g2_and3_1 _36194_ (.X(_10422_),
    .A(_08997_),
    .B(_09047_),
    .C(_10420_));
 sg13g2_nor3_1 _36195_ (.A(net5369),
    .B(_10421_),
    .C(_10422_),
    .Y(_10423_));
 sg13g2_a21o_2 _36196_ (.A2(_08995_),
    .A1(net5369),
    .B1(_10423_),
    .X(_10424_));
 sg13g2_nand3_1 _36197_ (.B(net4641),
    .C(_10424_),
    .A(net4633),
    .Y(_10425_));
 sg13g2_a21o_1 _36198_ (.A2(net4641),
    .A1(net4633),
    .B1(_10424_),
    .X(_10426_));
 sg13g2_nand2_1 _36199_ (.Y(_10427_),
    .A(_10425_),
    .B(_10426_));
 sg13g2_o21ai_1 _36200_ (.B1(_10409_),
    .Y(_10428_),
    .A1(_10411_),
    .A2(_10414_));
 sg13g2_a21oi_1 _36201_ (.A1(_10427_),
    .A2(_10428_),
    .Y(_10429_),
    .B1(net4671));
 sg13g2_o21ai_1 _36202_ (.B1(_10429_),
    .Y(_10430_),
    .A1(_10427_),
    .A2(_10428_));
 sg13g2_o21ai_1 _36203_ (.B1(_10430_),
    .Y(_10431_),
    .A1(net4708),
    .A2(_10424_));
 sg13g2_o21ai_1 _36204_ (.B1(net5603),
    .Y(_10432_),
    .A1(net4418),
    .A2(_10408_));
 sg13g2_a21oi_1 _36205_ (.A1(net4418),
    .A2(_10431_),
    .Y(_10433_),
    .B1(_10432_));
 sg13g2_a21o_1 _36206_ (.A2(net4210),
    .A1(net3304),
    .B1(_10433_),
    .X(_00824_));
 sg13g2_nor2_1 _36207_ (.A(_08996_),
    .B(_10421_),
    .Y(_10434_));
 sg13g2_xnor2_1 _36208_ (.Y(_10435_),
    .A(_09008_),
    .B(_10434_));
 sg13g2_nor2_1 _36209_ (.A(net5372),
    .B(_10435_),
    .Y(_10436_));
 sg13g2_a21oi_2 _36210_ (.B1(_10436_),
    .Y(_10437_),
    .A2(_09005_),
    .A1(net5369));
 sg13g2_xnor2_1 _36211_ (.Y(_10438_),
    .A(net4558),
    .B(_10437_));
 sg13g2_xnor2_1 _36212_ (.Y(_10439_),
    .A(net4606),
    .B(_10437_));
 sg13g2_nand4_1 _36213_ (.B(_10410_),
    .C(_10425_),
    .A(_10409_),
    .Y(_10440_),
    .D(_10426_));
 sg13g2_and2_1 _36214_ (.A(_10409_),
    .B(_10425_),
    .X(_10441_));
 sg13g2_o21ai_1 _36215_ (.B1(_10441_),
    .Y(_10442_),
    .A1(_10412_),
    .A2(_10440_));
 sg13g2_nor3_1 _36216_ (.A(_10376_),
    .B(_10399_),
    .C(_10440_),
    .Y(_10443_));
 sg13g2_a21oi_1 _36217_ (.A1(_10386_),
    .A2(_10443_),
    .Y(_10444_),
    .B1(_10442_));
 sg13g2_nor2_1 _36218_ (.A(_10439_),
    .B(_10444_),
    .Y(_10445_));
 sg13g2_and2_1 _36219_ (.A(_10439_),
    .B(_10444_),
    .X(_10446_));
 sg13g2_o21ai_1 _36220_ (.B1(net4708),
    .Y(_10447_),
    .A1(_10445_),
    .A2(_10446_));
 sg13g2_o21ai_1 _36221_ (.B1(_10447_),
    .Y(_10448_),
    .A1(net4709),
    .A2(_10437_));
 sg13g2_o21ai_1 _36222_ (.B1(net5603),
    .Y(_10449_),
    .A1(net4418),
    .A2(_10424_));
 sg13g2_a21oi_1 _36223_ (.A1(net4419),
    .A2(_10448_),
    .Y(_10450_),
    .B1(_10449_));
 sg13g2_a21o_1 _36224_ (.A2(net4210),
    .A1(net2645),
    .B1(_10450_),
    .X(_00825_));
 sg13g2_nand2_1 _36225_ (.Y(_10451_),
    .A(net5373),
    .B(_08986_));
 sg13g2_o21ai_1 _36226_ (.B1(_09007_),
    .Y(_10452_),
    .A1(_09050_),
    .A2(_10421_));
 sg13g2_nor2_1 _36227_ (.A(_08988_),
    .B(_10452_),
    .Y(_10453_));
 sg13g2_a21o_1 _36228_ (.A2(_10452_),
    .A1(_08988_),
    .B1(net5373),
    .X(_10454_));
 sg13g2_o21ai_1 _36229_ (.B1(_10451_),
    .Y(_10455_),
    .A1(_10453_),
    .A2(_10454_));
 sg13g2_and2_1 _36230_ (.A(net4606),
    .B(_10455_),
    .X(_10456_));
 sg13g2_nand2b_1 _36231_ (.Y(_10457_),
    .B(net4558),
    .A_N(_10455_));
 sg13g2_xnor2_1 _36232_ (.Y(_10458_),
    .A(net4558),
    .B(_10455_));
 sg13g2_a21oi_1 _36233_ (.A1(net4606),
    .A2(_10437_),
    .Y(_10459_),
    .B1(_10445_));
 sg13g2_a21oi_1 _36234_ (.A1(_10458_),
    .A2(_10459_),
    .Y(_10460_),
    .B1(net4671));
 sg13g2_o21ai_1 _36235_ (.B1(_10460_),
    .Y(_10461_),
    .A1(_10458_),
    .A2(_10459_));
 sg13g2_o21ai_1 _36236_ (.B1(_10461_),
    .Y(_10462_),
    .A1(net4709),
    .A2(_10455_));
 sg13g2_o21ai_1 _36237_ (.B1(net5603),
    .Y(_10463_),
    .A1(net4419),
    .A2(_10437_));
 sg13g2_a21oi_1 _36238_ (.A1(net4419),
    .A2(_10462_),
    .Y(_10464_),
    .B1(_10463_));
 sg13g2_a21o_1 _36239_ (.A2(net4210),
    .A1(net2740),
    .B1(_10464_),
    .X(_00826_));
 sg13g2_nand2_1 _36240_ (.Y(_10465_),
    .A(net5373),
    .B(_08979_));
 sg13g2_nor2_1 _36241_ (.A(_08987_),
    .B(_10453_),
    .Y(_10466_));
 sg13g2_xor2_1 _36242_ (.B(_10466_),
    .A(_08981_),
    .X(_10467_));
 sg13g2_o21ai_1 _36243_ (.B1(_10465_),
    .Y(_10468_),
    .A1(net5373),
    .A2(_10467_));
 sg13g2_or2_1 _36244_ (.X(_10469_),
    .B(_10468_),
    .A(net4558));
 sg13g2_xnor2_1 _36245_ (.Y(_10470_),
    .A(net4606),
    .B(_10468_));
 sg13g2_a21o_1 _36246_ (.A2(_10437_),
    .A1(net4605),
    .B1(_10456_),
    .X(_10471_));
 sg13g2_or2_1 _36247_ (.X(_10472_),
    .B(_10471_),
    .A(_10445_));
 sg13g2_nand3_1 _36248_ (.B(_10470_),
    .C(_10472_),
    .A(_10457_),
    .Y(_10473_));
 sg13g2_a21oi_1 _36249_ (.A1(_10457_),
    .A2(_10472_),
    .Y(_10474_),
    .B1(_10470_));
 sg13g2_nor2_1 _36250_ (.A(net4671),
    .B(_10474_),
    .Y(_10475_));
 sg13g2_nor2_1 _36251_ (.A(net4709),
    .B(_10468_),
    .Y(_10476_));
 sg13g2_a21oi_1 _36252_ (.A1(_10473_),
    .A2(_10475_),
    .Y(_10477_),
    .B1(_10476_));
 sg13g2_o21ai_1 _36253_ (.B1(net5603),
    .Y(_10478_),
    .A1(net4419),
    .A2(_10455_));
 sg13g2_a21oi_1 _36254_ (.A1(net4419),
    .A2(_10477_),
    .Y(_10479_),
    .B1(_10478_));
 sg13g2_a21o_1 _36255_ (.A2(net4210),
    .A1(net2438),
    .B1(_10479_),
    .X(_00827_));
 sg13g2_nand2_1 _36256_ (.Y(_10480_),
    .A(net5373),
    .B(_08953_));
 sg13g2_o21ai_1 _36257_ (.B1(_09243_),
    .Y(_10481_),
    .A1(_09237_),
    .A2(_10361_));
 sg13g2_a21o_2 _36258_ (.A2(_10481_),
    .A1(_09052_),
    .B1(_08963_),
    .X(_10482_));
 sg13g2_nand3_1 _36259_ (.B(_09052_),
    .C(_10481_),
    .A(_08963_),
    .Y(_10483_));
 sg13g2_nand3_1 _36260_ (.B(_10482_),
    .C(_10483_),
    .A(net5414),
    .Y(_10484_));
 sg13g2_nand2_2 _36261_ (.Y(_10485_),
    .A(_10480_),
    .B(_10484_));
 sg13g2_nand2_1 _36262_ (.Y(_10486_),
    .A(net4606),
    .B(_10485_));
 sg13g2_xnor2_1 _36263_ (.Y(_10487_),
    .A(net4558),
    .B(_10485_));
 sg13g2_nand2_1 _36264_ (.Y(_10488_),
    .A(_10469_),
    .B(_10473_));
 sg13g2_o21ai_1 _36265_ (.B1(net4709),
    .Y(_10489_),
    .A1(_10487_),
    .A2(_10488_));
 sg13g2_a21o_1 _36266_ (.A2(_10488_),
    .A1(_10487_),
    .B1(_10489_),
    .X(_10490_));
 sg13g2_nand2_1 _36267_ (.Y(_10491_),
    .A(net4671),
    .B(_10485_));
 sg13g2_nand3_1 _36268_ (.B(_10490_),
    .C(_10491_),
    .A(net4419),
    .Y(_10492_));
 sg13g2_a21oi_1 _36269_ (.A1(net4365),
    .A2(_10468_),
    .Y(_10493_),
    .B1(net5564));
 sg13g2_a22oi_1 _36270_ (.Y(_10494_),
    .B1(_10492_),
    .B2(_10493_),
    .A2(net4210),
    .A1(net1726));
 sg13g2_inv_1 _36271_ (.Y(_00828_),
    .A(_10494_));
 sg13g2_nand2_1 _36272_ (.Y(_10495_),
    .A(net5373),
    .B(_08946_));
 sg13g2_nor2b_1 _36273_ (.A(_08954_),
    .B_N(_10482_),
    .Y(_10496_));
 sg13g2_xnor2_1 _36274_ (.Y(_10497_),
    .A(_08962_),
    .B(_10496_));
 sg13g2_o21ai_1 _36275_ (.B1(_10495_),
    .Y(_10498_),
    .A1(net5373),
    .A2(_10497_));
 sg13g2_xnor2_1 _36276_ (.Y(_10499_),
    .A(net4560),
    .B(_10498_));
 sg13g2_xnor2_1 _36277_ (.Y(_10500_),
    .A(net4612),
    .B(_10498_));
 sg13g2_and2_1 _36278_ (.A(_10470_),
    .B(_10487_),
    .X(_10501_));
 sg13g2_and4_1 _36279_ (.A(_10438_),
    .B(_10458_),
    .C(_10470_),
    .D(_10487_),
    .X(_10502_));
 sg13g2_nand2_1 _36280_ (.Y(_10503_),
    .A(_10469_),
    .B(_10486_));
 sg13g2_a221oi_1 _36281_ (.B2(_10442_),
    .C1(_10503_),
    .B1(_10502_),
    .A1(_10471_),
    .Y(_10504_),
    .A2(_10501_));
 sg13g2_nand2_1 _36282_ (.Y(_10505_),
    .A(_10443_),
    .B(_10502_));
 sg13g2_o21ai_1 _36283_ (.B1(_10504_),
    .Y(_10506_),
    .A1(_10385_),
    .A2(_10505_));
 sg13g2_and2_1 _36284_ (.A(_10499_),
    .B(_10506_),
    .X(_10507_));
 sg13g2_nor2_1 _36285_ (.A(_10499_),
    .B(_10506_),
    .Y(_10508_));
 sg13g2_o21ai_1 _36286_ (.B1(net4714),
    .Y(_10509_),
    .A1(_10507_),
    .A2(_10508_));
 sg13g2_o21ai_1 _36287_ (.B1(_10509_),
    .Y(_10510_),
    .A1(net4714),
    .A2(_10498_));
 sg13g2_o21ai_1 _36288_ (.B1(net5604),
    .Y(_10511_),
    .A1(net4426),
    .A2(_10485_));
 sg13g2_a21oi_1 _36289_ (.A1(net4426),
    .A2(_10510_),
    .Y(_10512_),
    .B1(_10511_));
 sg13g2_a21o_1 _36290_ (.A2(net4211),
    .A1(net2590),
    .B1(_10512_),
    .X(_00829_));
 sg13g2_nand2_1 _36291_ (.Y(_10513_),
    .A(net5373),
    .B(_08925_));
 sg13g2_a22oi_1 _36292_ (.Y(_10514_),
    .B1(_08955_),
    .B2(_10482_),
    .A2(_08947_),
    .A1(net4817));
 sg13g2_a221oi_1 _36293_ (.B2(_10482_),
    .C1(_08927_),
    .B1(_08955_),
    .A1(net4817),
    .Y(_10515_),
    .A2(_08947_));
 sg13g2_xor2_1 _36294_ (.B(_10514_),
    .A(_08927_),
    .X(_10516_));
 sg13g2_o21ai_1 _36295_ (.B1(_10513_),
    .Y(_10517_),
    .A1(net5375),
    .A2(_10516_));
 sg13g2_a21oi_1 _36296_ (.A1(net4612),
    .A2(_10498_),
    .Y(_10518_),
    .B1(_10507_));
 sg13g2_xnor2_1 _36297_ (.Y(_10519_),
    .A(net4612),
    .B(_10517_));
 sg13g2_nor2_1 _36298_ (.A(_10518_),
    .B(_10519_),
    .Y(_10520_));
 sg13g2_nand2_1 _36299_ (.Y(_10521_),
    .A(_10518_),
    .B(_10519_));
 sg13g2_nand3b_1 _36300_ (.B(_10521_),
    .C(net4714),
    .Y(_10522_),
    .A_N(_10520_));
 sg13g2_a21oi_1 _36301_ (.A1(net4673),
    .A2(_10517_),
    .Y(_10523_),
    .B1(net4366));
 sg13g2_o21ai_1 _36302_ (.B1(net5604),
    .Y(_10524_),
    .A1(net4426),
    .A2(_10498_));
 sg13g2_a21oi_1 _36303_ (.A1(_10522_),
    .A2(_10523_),
    .Y(_10525_),
    .B1(_10524_));
 sg13g2_a21o_1 _36304_ (.A2(net4211),
    .A1(net2177),
    .B1(_10525_),
    .X(_00830_));
 sg13g2_nor2_1 _36305_ (.A(net5414),
    .B(_08935_),
    .Y(_10526_));
 sg13g2_nor2_1 _36306_ (.A(_08926_),
    .B(_10515_),
    .Y(_10527_));
 sg13g2_xor2_1 _36307_ (.B(_10527_),
    .A(_08936_),
    .X(_10528_));
 sg13g2_a21o_2 _36308_ (.A2(_10528_),
    .A1(net5414),
    .B1(_10526_),
    .X(_10529_));
 sg13g2_nand2_1 _36309_ (.Y(_10530_),
    .A(net4673),
    .B(_10529_));
 sg13g2_nand3b_1 _36310_ (.B(net4633),
    .C(net4641),
    .Y(_10531_),
    .A_N(_10529_));
 sg13g2_o21ai_1 _36311_ (.B1(_10529_),
    .Y(_10532_),
    .A1(_09669_),
    .A2(_09672_));
 sg13g2_nand2_1 _36312_ (.Y(_10533_),
    .A(_10531_),
    .B(_10532_));
 sg13g2_o21ai_1 _36313_ (.B1(net4612),
    .Y(_10534_),
    .A1(_10498_),
    .A2(_10517_));
 sg13g2_nand2b_1 _36314_ (.Y(_10535_),
    .B(_10534_),
    .A_N(_10507_));
 sg13g2_o21ai_1 _36315_ (.B1(_10535_),
    .Y(_10536_),
    .A1(net4612),
    .A2(_10517_));
 sg13g2_xor2_1 _36316_ (.B(_10536_),
    .A(_10533_),
    .X(_10537_));
 sg13g2_o21ai_1 _36317_ (.B1(_10530_),
    .Y(_10538_),
    .A1(net4673),
    .A2(_10537_));
 sg13g2_o21ai_1 _36318_ (.B1(net5604),
    .Y(_10539_),
    .A1(net4426),
    .A2(_10517_));
 sg13g2_a21oi_1 _36319_ (.A1(net4426),
    .A2(_10538_),
    .Y(_10540_),
    .B1(_10539_));
 sg13g2_a21o_1 _36320_ (.A2(net4211),
    .A1(net2624),
    .B1(_10540_),
    .X(_00831_));
 sg13g2_nand2_1 _36321_ (.Y(_10541_),
    .A(net5376),
    .B(_08913_));
 sg13g2_a21oi_1 _36322_ (.A1(_09052_),
    .A2(_10481_),
    .Y(_10542_),
    .B1(_08964_));
 sg13g2_o21ai_1 _36323_ (.B1(_08915_),
    .Y(_10543_),
    .A1(_08957_),
    .A2(_10542_));
 sg13g2_or3_1 _36324_ (.A(_08915_),
    .B(_08957_),
    .C(_10542_),
    .X(_10544_));
 sg13g2_nand2_1 _36325_ (.Y(_10545_),
    .A(_10543_),
    .B(_10544_));
 sg13g2_o21ai_1 _36326_ (.B1(_10541_),
    .Y(_10546_),
    .A1(net5375),
    .A2(_10545_));
 sg13g2_nand3_1 _36327_ (.B(net4641),
    .C(_10546_),
    .A(net4633),
    .Y(_10547_));
 sg13g2_a21o_1 _36328_ (.A2(net4641),
    .A1(net4633),
    .B1(_10546_),
    .X(_10548_));
 sg13g2_nand2_1 _36329_ (.Y(_10549_),
    .A(_10547_),
    .B(_10548_));
 sg13g2_o21ai_1 _36330_ (.B1(_10531_),
    .Y(_10550_),
    .A1(_10533_),
    .A2(_10536_));
 sg13g2_xnor2_1 _36331_ (.Y(_10551_),
    .A(_10549_),
    .B(_10550_));
 sg13g2_nand2_1 _36332_ (.Y(_10552_),
    .A(net4714),
    .B(_10551_));
 sg13g2_nand2_1 _36333_ (.Y(_10553_),
    .A(net4673),
    .B(_10546_));
 sg13g2_nand3_1 _36334_ (.B(_10552_),
    .C(_10553_),
    .A(net4426),
    .Y(_10554_));
 sg13g2_a21oi_1 _36335_ (.A1(net4366),
    .A2(_10529_),
    .Y(_10555_),
    .B1(net5569));
 sg13g2_a22oi_1 _36336_ (.Y(_10556_),
    .B1(_10554_),
    .B2(_10555_),
    .A2(net4211),
    .A1(net2606));
 sg13g2_inv_1 _36337_ (.Y(_00832_),
    .A(_10556_));
 sg13g2_a21oi_1 _36338_ (.A1(_08897_),
    .A2(_08902_),
    .Y(_10557_),
    .B1(net5419));
 sg13g2_nand2_1 _36339_ (.Y(_10558_),
    .A(_08914_),
    .B(_10543_));
 sg13g2_xnor2_1 _36340_ (.Y(_10559_),
    .A(_08906_),
    .B(_10558_));
 sg13g2_a21oi_2 _36341_ (.B1(_10557_),
    .Y(_10560_),
    .A2(_10559_),
    .A1(net5419));
 sg13g2_nand2_1 _36342_ (.Y(_10561_),
    .A(net4613),
    .B(_10560_));
 sg13g2_xnor2_1 _36343_ (.Y(_10562_),
    .A(net4562),
    .B(_10560_));
 sg13g2_xnor2_1 _36344_ (.Y(_10563_),
    .A(net4613),
    .B(_10560_));
 sg13g2_nand4_1 _36345_ (.B(_10532_),
    .C(_10547_),
    .A(_10531_),
    .Y(_10564_),
    .D(_10548_));
 sg13g2_and2_1 _36346_ (.A(_10531_),
    .B(_10547_),
    .X(_10565_));
 sg13g2_o21ai_1 _36347_ (.B1(_10565_),
    .Y(_10566_),
    .A1(_10534_),
    .A2(_10564_));
 sg13g2_or3_1 _36348_ (.A(_10500_),
    .B(_10519_),
    .C(_10564_),
    .X(_10567_));
 sg13g2_nor2b_1 _36349_ (.A(_10567_),
    .B_N(_10506_),
    .Y(_10568_));
 sg13g2_nor2_2 _36350_ (.A(_10566_),
    .B(_10568_),
    .Y(_10569_));
 sg13g2_nor2_1 _36351_ (.A(_10563_),
    .B(_10569_),
    .Y(_10570_));
 sg13g2_xnor2_1 _36352_ (.Y(_10571_),
    .A(_10563_),
    .B(_10569_));
 sg13g2_nand2_1 _36353_ (.Y(_10572_),
    .A(net4715),
    .B(_10571_));
 sg13g2_o21ai_1 _36354_ (.B1(_10572_),
    .Y(_10573_),
    .A1(net4715),
    .A2(_10560_));
 sg13g2_o21ai_1 _36355_ (.B1(net5604),
    .Y(_10574_),
    .A1(net4426),
    .A2(_10546_));
 sg13g2_a21oi_1 _36356_ (.A1(net4426),
    .A2(_10573_),
    .Y(_10575_),
    .B1(_10574_));
 sg13g2_a21o_1 _36357_ (.A2(net4211),
    .A1(net2117),
    .B1(_10575_),
    .X(_00833_));
 sg13g2_o21ai_1 _36358_ (.B1(_10561_),
    .Y(_10576_),
    .A1(_10563_),
    .A2(_10569_));
 sg13g2_a21o_1 _36359_ (.A2(_10543_),
    .A1(_08958_),
    .B1(_08904_),
    .X(_10577_));
 sg13g2_xnor2_1 _36360_ (.Y(_10578_),
    .A(_08878_),
    .B(_10577_));
 sg13g2_mux2_1 _36361_ (.A0(_08876_),
    .A1(_10578_),
    .S(net5419),
    .X(_10579_));
 sg13g2_nand2_1 _36362_ (.Y(_10580_),
    .A(net4562),
    .B(_10579_));
 sg13g2_xnor2_1 _36363_ (.Y(_10581_),
    .A(net4613),
    .B(_10579_));
 sg13g2_nand2_1 _36364_ (.Y(_10582_),
    .A(net4675),
    .B(_10579_));
 sg13g2_xor2_1 _36365_ (.B(_10581_),
    .A(_10576_),
    .X(_10583_));
 sg13g2_o21ai_1 _36366_ (.B1(_10582_),
    .Y(_10584_),
    .A1(net4675),
    .A2(_10583_));
 sg13g2_o21ai_1 _36367_ (.B1(net5606),
    .Y(_10585_),
    .A1(net4428),
    .A2(_10560_));
 sg13g2_a21oi_1 _36368_ (.A1(net4428),
    .A2(_10584_),
    .Y(_10586_),
    .B1(_10585_));
 sg13g2_a21o_1 _36369_ (.A2(net4225),
    .A1(net2347),
    .B1(_10586_),
    .X(_00834_));
 sg13g2_a21oi_1 _36370_ (.A1(_08881_),
    .A2(_08886_),
    .Y(_10587_),
    .B1(net5419));
 sg13g2_o21ai_1 _36371_ (.B1(_08877_),
    .Y(_10588_),
    .A1(_08878_),
    .A2(_10577_));
 sg13g2_xnor2_1 _36372_ (.Y(_10589_),
    .A(_08890_),
    .B(_10588_));
 sg13g2_a21oi_2 _36373_ (.B1(_10587_),
    .Y(_10590_),
    .A2(_10589_),
    .A1(net5419));
 sg13g2_and2_1 _36374_ (.A(net4613),
    .B(_10590_),
    .X(_10591_));
 sg13g2_xnor2_1 _36375_ (.Y(_10592_),
    .A(net4562),
    .B(_10590_));
 sg13g2_o21ai_1 _36376_ (.B1(_10561_),
    .Y(_10593_),
    .A1(net4562),
    .A2(_10579_));
 sg13g2_or2_1 _36377_ (.X(_10594_),
    .B(_10593_),
    .A(_10570_));
 sg13g2_a21o_1 _36378_ (.A2(_10594_),
    .A1(_10580_),
    .B1(_10592_),
    .X(_10595_));
 sg13g2_nand3_1 _36379_ (.B(_10592_),
    .C(_10594_),
    .A(_10580_),
    .Y(_10596_));
 sg13g2_nand3_1 _36380_ (.B(_10595_),
    .C(_10596_),
    .A(net4715),
    .Y(_10597_));
 sg13g2_nand2_1 _36381_ (.Y(_10598_),
    .A(net4675),
    .B(_10590_));
 sg13g2_nand3_1 _36382_ (.B(_10597_),
    .C(_10598_),
    .A(net4428),
    .Y(_10599_));
 sg13g2_a21oi_1 _36383_ (.A1(net4369),
    .A2(_10579_),
    .Y(_10600_),
    .B1(net5572));
 sg13g2_a22oi_1 _36384_ (.Y(_10601_),
    .B1(_10599_),
    .B2(_10600_),
    .A2(net4225),
    .A1(net2600));
 sg13g2_inv_1 _36385_ (.Y(_00835_),
    .A(_10601_));
 sg13g2_o21ai_1 _36386_ (.B1(net5419),
    .Y(_10602_),
    .A1(_09602_),
    .A2(_09606_));
 sg13g2_a21oi_1 _36387_ (.A1(_09602_),
    .A2(_09606_),
    .Y(_10603_),
    .B1(_10602_));
 sg13g2_a21oi_2 _36388_ (.B1(_10603_),
    .Y(_10604_),
    .A2(_08816_),
    .A1(net5376));
 sg13g2_nand2_1 _36389_ (.Y(_10605_),
    .A(net4675),
    .B(_10604_));
 sg13g2_nor2_1 _36390_ (.A(net4562),
    .B(_10604_),
    .Y(_10606_));
 sg13g2_xnor2_1 _36391_ (.Y(_10607_),
    .A(net4613),
    .B(_10604_));
 sg13g2_nor2b_1 _36392_ (.A(_10591_),
    .B_N(_10596_),
    .Y(_10608_));
 sg13g2_xnor2_1 _36393_ (.Y(_10609_),
    .A(_10607_),
    .B(_10608_));
 sg13g2_o21ai_1 _36394_ (.B1(_10605_),
    .Y(_10610_),
    .A1(net4675),
    .A2(_10609_));
 sg13g2_o21ai_1 _36395_ (.B1(net5606),
    .Y(_10611_),
    .A1(net4428),
    .A2(_10590_));
 sg13g2_a21oi_1 _36396_ (.A1(net4428),
    .A2(_10610_),
    .Y(_10612_),
    .B1(_10611_));
 sg13g2_a21o_1 _36397_ (.A2(net4225),
    .A1(net1582),
    .B1(_10612_),
    .X(_00836_));
 sg13g2_nand2_1 _36398_ (.Y(_10613_),
    .A(net4369),
    .B(_10604_));
 sg13g2_o21ai_1 _36399_ (.B1(_08817_),
    .Y(_10614_),
    .A1(_09602_),
    .A2(_09606_));
 sg13g2_o21ai_1 _36400_ (.B1(net5419),
    .Y(_10615_),
    .A1(_09604_),
    .A2(_10614_));
 sg13g2_a21o_1 _36401_ (.A2(_10614_),
    .A1(_09604_),
    .B1(_10615_),
    .X(_10616_));
 sg13g2_o21ai_1 _36402_ (.B1(_10616_),
    .Y(_10617_),
    .A1(net5419),
    .A2(_08811_));
 sg13g2_nand2_1 _36403_ (.Y(_10618_),
    .A(net4613),
    .B(_10617_));
 sg13g2_xnor2_1 _36404_ (.Y(_10619_),
    .A(net4562),
    .B(_10617_));
 sg13g2_and2_1 _36405_ (.A(_10592_),
    .B(_10607_),
    .X(_10620_));
 sg13g2_and4_1 _36406_ (.A(_10562_),
    .B(_10581_),
    .C(_10592_),
    .D(_10607_),
    .X(_10621_));
 sg13g2_nand2b_2 _36407_ (.Y(_10622_),
    .B(_10621_),
    .A_N(_10567_));
 sg13g2_nor2_1 _36408_ (.A(_10505_),
    .B(_10622_),
    .Y(_10623_));
 sg13g2_nand2b_1 _36409_ (.Y(_10624_),
    .B(_10623_),
    .A_N(_10383_));
 sg13g2_or2_1 _36410_ (.X(_10625_),
    .B(_10606_),
    .A(_10591_));
 sg13g2_a221oi_1 _36411_ (.B2(_10566_),
    .C1(_10625_),
    .B1(_10621_),
    .A1(_10593_),
    .Y(_10626_),
    .A2(_10620_));
 sg13g2_o21ai_1 _36412_ (.B1(_10626_),
    .Y(_10627_),
    .A1(_10504_),
    .A2(_10622_));
 sg13g2_a21oi_1 _36413_ (.A1(_10382_),
    .A2(_10623_),
    .Y(_10628_),
    .B1(_10627_));
 sg13g2_o21ai_1 _36414_ (.B1(_10628_),
    .Y(_10629_),
    .A1(_10136_),
    .A2(_10624_));
 sg13g2_nand2_1 _36415_ (.Y(_10630_),
    .A(_10619_),
    .B(_10629_));
 sg13g2_or2_1 _36416_ (.X(_10631_),
    .B(_10629_),
    .A(_10619_));
 sg13g2_a21o_1 _36417_ (.A2(_10631_),
    .A1(_10630_),
    .B1(net4675),
    .X(_10632_));
 sg13g2_o21ai_1 _36418_ (.B1(_10632_),
    .Y(_10633_),
    .A1(net4715),
    .A2(_10617_));
 sg13g2_a21oi_1 _36419_ (.A1(net4428),
    .A2(_10633_),
    .Y(_10634_),
    .B1(net5572));
 sg13g2_a22oi_1 _36420_ (.Y(_10635_),
    .B1(_10613_),
    .B2(_10634_),
    .A2(net4225),
    .A1(net2678));
 sg13g2_inv_1 _36421_ (.Y(_00837_),
    .A(_10635_));
 sg13g2_nand2_1 _36422_ (.Y(_10636_),
    .A(net2641),
    .B(net4225));
 sg13g2_nor2_1 _36423_ (.A(net5422),
    .B(_08790_),
    .Y(_10637_));
 sg13g2_o21ai_1 _36424_ (.B1(_08818_),
    .Y(_10638_),
    .A1(_09602_),
    .A2(_09606_));
 sg13g2_nand3_1 _36425_ (.B(_09603_),
    .C(_10638_),
    .A(_08792_),
    .Y(_10639_));
 sg13g2_a21o_1 _36426_ (.A2(_10638_),
    .A1(_09603_),
    .B1(_08792_),
    .X(_10640_));
 sg13g2_and2_1 _36427_ (.A(_10639_),
    .B(_10640_),
    .X(_10641_));
 sg13g2_a21oi_2 _36428_ (.B1(_10637_),
    .Y(_10642_),
    .A2(_10641_),
    .A1(net5422));
 sg13g2_inv_1 _36429_ (.Y(_10643_),
    .A(_10642_));
 sg13g2_nand2_1 _36430_ (.Y(_10644_),
    .A(_10618_),
    .B(_10630_));
 sg13g2_xnor2_1 _36431_ (.Y(_10645_),
    .A(net4613),
    .B(_10642_));
 sg13g2_xor2_1 _36432_ (.B(_10645_),
    .A(_10644_),
    .X(_10646_));
 sg13g2_o21ai_1 _36433_ (.B1(net4429),
    .Y(_10647_),
    .A1(net4715),
    .A2(_10642_));
 sg13g2_a21oi_1 _36434_ (.A1(net4715),
    .A2(_10646_),
    .Y(_10648_),
    .B1(_10647_));
 sg13g2_o21ai_1 _36435_ (.B1(net5606),
    .Y(_10649_),
    .A1(net4429),
    .A2(_10617_));
 sg13g2_o21ai_1 _36436_ (.B1(_10636_),
    .Y(_00838_),
    .A1(_10648_),
    .A2(_10649_));
 sg13g2_and2_1 _36437_ (.A(net5378),
    .B(_08800_),
    .X(_10650_));
 sg13g2_nor2b_1 _36438_ (.A(_08791_),
    .B_N(_10639_),
    .Y(_10651_));
 sg13g2_xor2_1 _36439_ (.B(_10651_),
    .A(_08801_),
    .X(_10652_));
 sg13g2_a21oi_2 _36440_ (.B1(_10650_),
    .Y(_10653_),
    .A2(_10652_),
    .A1(net5422));
 sg13g2_nand3_1 _36441_ (.B(net4639),
    .C(_10653_),
    .A(net4631),
    .Y(_10654_));
 sg13g2_inv_1 _36442_ (.Y(_10655_),
    .A(_10654_));
 sg13g2_a21o_1 _36443_ (.A2(net4639),
    .A1(net4631),
    .B1(_10653_),
    .X(_10656_));
 sg13g2_and2_1 _36444_ (.A(_10654_),
    .B(_10656_),
    .X(_10657_));
 sg13g2_o21ai_1 _36445_ (.B1(net4613),
    .Y(_10658_),
    .A1(_10617_),
    .A2(_10643_));
 sg13g2_a22oi_1 _36446_ (.Y(_10659_),
    .B1(_10658_),
    .B2(_10630_),
    .A2(_10642_),
    .A1(net4562));
 sg13g2_xnor2_1 _36447_ (.Y(_10660_),
    .A(_10657_),
    .B(_10659_));
 sg13g2_nand2_1 _36448_ (.Y(_10661_),
    .A(net4717),
    .B(_10660_));
 sg13g2_o21ai_1 _36449_ (.B1(_10661_),
    .Y(_10662_),
    .A1(net4715),
    .A2(_10653_));
 sg13g2_nand2_1 _36450_ (.Y(_10663_),
    .A(net4429),
    .B(_10662_));
 sg13g2_a21oi_1 _36451_ (.A1(net4369),
    .A2(_10642_),
    .Y(_10664_),
    .B1(net5572));
 sg13g2_a22oi_1 _36452_ (.Y(_10665_),
    .B1(_10663_),
    .B2(_10664_),
    .A2(net4227),
    .A1(net2334));
 sg13g2_inv_1 _36453_ (.Y(_00839_),
    .A(_10665_));
 sg13g2_nand2_1 _36454_ (.Y(_10666_),
    .A(net5378),
    .B(_08779_));
 sg13g2_o21ai_1 _36455_ (.B1(_09607_),
    .Y(_10667_),
    .A1(_09245_),
    .A2(net1064));
 sg13g2_nand2b_1 _36456_ (.Y(_10668_),
    .B(_10667_),
    .A_N(_08820_));
 sg13g2_and2_1 _36457_ (.A(_08782_),
    .B(_10668_),
    .X(_10669_));
 sg13g2_xnor2_1 _36458_ (.Y(_10670_),
    .A(_08782_),
    .B(_10668_));
 sg13g2_o21ai_1 _36459_ (.B1(_10666_),
    .Y(_10671_),
    .A1(net5378),
    .A2(_10670_));
 sg13g2_nand3_1 _36460_ (.B(net4639),
    .C(_10671_),
    .A(net4631),
    .Y(_10672_));
 sg13g2_a21o_1 _36461_ (.A2(net4639),
    .A1(net4631),
    .B1(_10671_),
    .X(_10673_));
 sg13g2_nand2_1 _36462_ (.Y(_10674_),
    .A(_10672_),
    .B(_10673_));
 sg13g2_a21oi_1 _36463_ (.A1(_10657_),
    .A2(_10659_),
    .Y(_10675_),
    .B1(_10655_));
 sg13g2_xnor2_1 _36464_ (.Y(_10676_),
    .A(_10674_),
    .B(_10675_));
 sg13g2_nand2_1 _36465_ (.Y(_10677_),
    .A(net4717),
    .B(_10676_));
 sg13g2_o21ai_1 _36466_ (.B1(_10677_),
    .Y(_10678_),
    .A1(net4717),
    .A2(_10671_));
 sg13g2_o21ai_1 _36467_ (.B1(net5606),
    .Y(_10679_),
    .A1(net4429),
    .A2(_10653_));
 sg13g2_a21oi_1 _36468_ (.A1(net4429),
    .A2(_10678_),
    .Y(_10680_),
    .B1(_10679_));
 sg13g2_a21o_1 _36469_ (.A2(net4227),
    .A1(net5880),
    .B1(_10680_),
    .X(_00840_));
 sg13g2_nor2_1 _36470_ (.A(_08780_),
    .B(_10669_),
    .Y(_10681_));
 sg13g2_xnor2_1 _36471_ (.Y(_10682_),
    .A(_08774_),
    .B(_10681_));
 sg13g2_nand2_1 _36472_ (.Y(_10683_),
    .A(net5422),
    .B(_10682_));
 sg13g2_o21ai_1 _36473_ (.B1(_10683_),
    .Y(_10684_),
    .A1(net5422),
    .A2(_08772_));
 sg13g2_and2_1 _36474_ (.A(net4617),
    .B(_10684_),
    .X(_10685_));
 sg13g2_xnor2_1 _36475_ (.Y(_10686_),
    .A(net4617),
    .B(_10684_));
 sg13g2_nand4_1 _36476_ (.B(_10656_),
    .C(_10672_),
    .A(_10654_),
    .Y(_10687_),
    .D(_10673_));
 sg13g2_and2_1 _36477_ (.A(_10654_),
    .B(_10672_),
    .X(_10688_));
 sg13g2_o21ai_1 _36478_ (.B1(_10688_),
    .Y(_10689_),
    .A1(_10658_),
    .A2(_10687_));
 sg13g2_nand2_1 _36479_ (.Y(_10690_),
    .A(_10619_),
    .B(_10645_));
 sg13g2_nor2_2 _36480_ (.A(_10687_),
    .B(_10690_),
    .Y(_10691_));
 sg13g2_a21oi_1 _36481_ (.A1(_10629_),
    .A2(_10691_),
    .Y(_10692_),
    .B1(_10689_));
 sg13g2_nor2_1 _36482_ (.A(_10686_),
    .B(_10692_),
    .Y(_10693_));
 sg13g2_xnor2_1 _36483_ (.Y(_10694_),
    .A(_10686_),
    .B(_10692_));
 sg13g2_nand2_1 _36484_ (.Y(_10695_),
    .A(net4717),
    .B(_10694_));
 sg13g2_o21ai_1 _36485_ (.B1(_10695_),
    .Y(_10696_),
    .A1(net4717),
    .A2(_10684_));
 sg13g2_o21ai_1 _36486_ (.B1(net5607),
    .Y(_10697_),
    .A1(net4432),
    .A2(_10671_));
 sg13g2_a21oi_1 _36487_ (.A1(net4432),
    .A2(_10696_),
    .Y(_10698_),
    .B1(_10697_));
 sg13g2_a21o_1 _36488_ (.A2(net4227),
    .A1(net2879),
    .B1(_10698_),
    .X(_00841_));
 sg13g2_nand2_1 _36489_ (.Y(_10699_),
    .A(net2871),
    .B(net4228));
 sg13g2_nor2_1 _36490_ (.A(net5422),
    .B(_08750_),
    .Y(_10700_));
 sg13g2_o21ai_1 _36491_ (.B1(_08773_),
    .Y(_10701_),
    .A1(_08822_),
    .A2(_10669_));
 sg13g2_xnor2_1 _36492_ (.Y(_10702_),
    .A(_08753_),
    .B(_10701_));
 sg13g2_a21oi_2 _36493_ (.B1(_10700_),
    .Y(_10703_),
    .A2(_10702_),
    .A1(net5422));
 sg13g2_nor2_1 _36494_ (.A(_10685_),
    .B(_10693_),
    .Y(_10704_));
 sg13g2_nand2_1 _36495_ (.Y(_10705_),
    .A(net4566),
    .B(_10703_));
 sg13g2_nor2_1 _36496_ (.A(net4566),
    .B(_10703_),
    .Y(_10706_));
 sg13g2_xnor2_1 _36497_ (.Y(_10707_),
    .A(net4566),
    .B(_10703_));
 sg13g2_xor2_1 _36498_ (.B(_10707_),
    .A(_10704_),
    .X(_10708_));
 sg13g2_o21ai_1 _36499_ (.B1(net4432),
    .Y(_10709_),
    .A1(net4717),
    .A2(_10703_));
 sg13g2_a21oi_1 _36500_ (.A1(net4717),
    .A2(_10708_),
    .Y(_10710_),
    .B1(_10709_));
 sg13g2_o21ai_1 _36501_ (.B1(net5608),
    .Y(_10711_),
    .A1(net4432),
    .A2(_10684_));
 sg13g2_o21ai_1 _36502_ (.B1(_10699_),
    .Y(_00842_),
    .A1(_10710_),
    .A2(_10711_));
 sg13g2_nand2_1 _36503_ (.Y(_10712_),
    .A(net5378),
    .B(_08761_));
 sg13g2_o21ai_1 _36504_ (.B1(_08751_),
    .Y(_10713_),
    .A1(_08752_),
    .A2(_10701_));
 sg13g2_xor2_1 _36505_ (.B(_10713_),
    .A(_08762_),
    .X(_10714_));
 sg13g2_o21ai_1 _36506_ (.B1(_10712_),
    .Y(_10715_),
    .A1(net5378),
    .A2(_10714_));
 sg13g2_nand2_1 _36507_ (.Y(_10716_),
    .A(net4678),
    .B(_10715_));
 sg13g2_or2_1 _36508_ (.X(_10717_),
    .B(_10715_),
    .A(net4566));
 sg13g2_xnor2_1 _36509_ (.Y(_10718_),
    .A(net4566),
    .B(_10715_));
 sg13g2_or2_1 _36510_ (.X(_10719_),
    .B(_10706_),
    .A(_10685_));
 sg13g2_o21ai_1 _36511_ (.B1(_10705_),
    .Y(_10720_),
    .A1(_10693_),
    .A2(_10719_));
 sg13g2_xor2_1 _36512_ (.B(_10720_),
    .A(_10718_),
    .X(_10721_));
 sg13g2_o21ai_1 _36513_ (.B1(_10716_),
    .Y(_10722_),
    .A1(net4678),
    .A2(_10721_));
 sg13g2_nand2_1 _36514_ (.Y(_10723_),
    .A(net4432),
    .B(_10722_));
 sg13g2_a21oi_1 _36515_ (.A1(net4368),
    .A2(_10703_),
    .Y(_10724_),
    .B1(net5571));
 sg13g2_a22oi_1 _36516_ (.Y(_10725_),
    .B1(_10723_),
    .B2(_10724_),
    .A2(net4228),
    .A1(net2952));
 sg13g2_inv_1 _36517_ (.Y(_00843_),
    .A(_10725_));
 sg13g2_nand2_1 _36518_ (.Y(_10726_),
    .A(net5378),
    .B(_08721_));
 sg13g2_o21ai_1 _36519_ (.B1(_09608_),
    .Y(_10727_),
    .A1(_09245_),
    .A2(net1064));
 sg13g2_a21o_2 _36520_ (.A2(_10727_),
    .A1(_08823_),
    .B1(_08723_),
    .X(_10728_));
 sg13g2_nand3_1 _36521_ (.B(_08823_),
    .C(_10727_),
    .A(_08723_),
    .Y(_10729_));
 sg13g2_nand2_1 _36522_ (.Y(_10730_),
    .A(_10728_),
    .B(_10729_));
 sg13g2_o21ai_1 _36523_ (.B1(_10726_),
    .Y(_10731_),
    .A1(net5378),
    .A2(_10730_));
 sg13g2_nand2_1 _36524_ (.Y(_10732_),
    .A(net4617),
    .B(_10731_));
 sg13g2_xnor2_1 _36525_ (.Y(_10733_),
    .A(net4617),
    .B(_10731_));
 sg13g2_o21ai_1 _36526_ (.B1(_10717_),
    .Y(_10734_),
    .A1(_10718_),
    .A2(_10720_));
 sg13g2_o21ai_1 _36527_ (.B1(net4718),
    .Y(_10735_),
    .A1(_10733_),
    .A2(_10734_));
 sg13g2_a21o_1 _36528_ (.A2(_10734_),
    .A1(_10733_),
    .B1(_10735_),
    .X(_10736_));
 sg13g2_o21ai_1 _36529_ (.B1(_10736_),
    .Y(_10737_),
    .A1(net4718),
    .A2(_10731_));
 sg13g2_nand2_1 _36530_ (.Y(_10738_),
    .A(net4432),
    .B(_10737_));
 sg13g2_a21oi_1 _36531_ (.A1(net4368),
    .A2(_10715_),
    .Y(_10739_),
    .B1(net5571));
 sg13g2_a22oi_1 _36532_ (.Y(_10740_),
    .B1(_10738_),
    .B2(_10739_),
    .A2(net4228),
    .A1(net5879));
 sg13g2_inv_1 _36533_ (.Y(_00844_),
    .A(_10740_));
 sg13g2_nand2_1 _36534_ (.Y(_10741_),
    .A(_08722_),
    .B(_10728_));
 sg13g2_xnor2_1 _36535_ (.Y(_10742_),
    .A(_08733_),
    .B(_10741_));
 sg13g2_nor2_1 _36536_ (.A(net5378),
    .B(_10742_),
    .Y(_10743_));
 sg13g2_a21oi_2 _36537_ (.B1(_10743_),
    .Y(_10744_),
    .A2(_08732_),
    .A1(net5382));
 sg13g2_xnor2_1 _36538_ (.Y(_10745_),
    .A(net4617),
    .B(_10744_));
 sg13g2_nor2_1 _36539_ (.A(_10718_),
    .B(_10733_),
    .Y(_10746_));
 sg13g2_nor4_1 _36540_ (.A(_10686_),
    .B(_10707_),
    .C(_10718_),
    .D(_10733_),
    .Y(_10747_));
 sg13g2_nand2_1 _36541_ (.Y(_10748_),
    .A(_10717_),
    .B(_10732_));
 sg13g2_a221oi_1 _36542_ (.B2(_10689_),
    .C1(_10748_),
    .B1(_10747_),
    .A1(_10719_),
    .Y(_10749_),
    .A2(_10746_));
 sg13g2_nand3_1 _36543_ (.B(_10691_),
    .C(_10747_),
    .A(_10629_),
    .Y(_10750_));
 sg13g2_and2_1 _36544_ (.A(_10749_),
    .B(_10750_),
    .X(_10751_));
 sg13g2_nor2_1 _36545_ (.A(_10745_),
    .B(_10751_),
    .Y(_10752_));
 sg13g2_and2_1 _36546_ (.A(_10745_),
    .B(_10751_),
    .X(_10753_));
 sg13g2_o21ai_1 _36547_ (.B1(net4718),
    .Y(_10754_),
    .A1(_10752_),
    .A2(_10753_));
 sg13g2_o21ai_1 _36548_ (.B1(_10754_),
    .Y(_10755_),
    .A1(net4718),
    .A2(_10744_));
 sg13g2_o21ai_1 _36549_ (.B1(net5608),
    .Y(_10756_),
    .A1(net4432),
    .A2(_10731_));
 sg13g2_a21oi_1 _36550_ (.A1(net4432),
    .A2(_10755_),
    .Y(_10757_),
    .B1(_10756_));
 sg13g2_a21o_1 _36551_ (.A2(net4228),
    .A1(net2536),
    .B1(_10757_),
    .X(_00845_));
 sg13g2_nand2_1 _36552_ (.Y(_10758_),
    .A(net5382),
    .B(_08706_));
 sg13g2_nand2_1 _36553_ (.Y(_10759_),
    .A(_08828_),
    .B(_10728_));
 sg13g2_o21ai_1 _36554_ (.B1(_10759_),
    .Y(_10760_),
    .A1(net4777),
    .A2(_08731_));
 sg13g2_a221oi_1 _36555_ (.B2(_10728_),
    .C1(_08708_),
    .B1(_08828_),
    .A1(net4825),
    .Y(_10761_),
    .A2(_08732_));
 sg13g2_a21o_1 _36556_ (.A2(_10760_),
    .A1(_08708_),
    .B1(net5382),
    .X(_10762_));
 sg13g2_o21ai_1 _36557_ (.B1(_10758_),
    .Y(_10763_),
    .A1(_10761_),
    .A2(_10762_));
 sg13g2_xnor2_1 _36558_ (.Y(_10764_),
    .A(net4617),
    .B(_10763_));
 sg13g2_a21oi_1 _36559_ (.A1(net4617),
    .A2(_10744_),
    .Y(_10765_),
    .B1(_10752_));
 sg13g2_xnor2_1 _36560_ (.Y(_10766_),
    .A(_10764_),
    .B(_10765_));
 sg13g2_nand2_1 _36561_ (.Y(_10767_),
    .A(net4718),
    .B(_10766_));
 sg13g2_o21ai_1 _36562_ (.B1(_10767_),
    .Y(_10768_),
    .A1(net4718),
    .A2(_10763_));
 sg13g2_o21ai_1 _36563_ (.B1(net5608),
    .Y(_10769_),
    .A1(net4433),
    .A2(_10744_));
 sg13g2_a21oi_1 _36564_ (.A1(net4433),
    .A2(_10768_),
    .Y(_10770_),
    .B1(_10769_));
 sg13g2_a21o_1 _36565_ (.A2(net4228),
    .A1(net5878),
    .B1(_10770_),
    .X(_00846_));
 sg13g2_nor2_1 _36566_ (.A(net5424),
    .B(_08714_),
    .Y(_10771_));
 sg13g2_nor2_1 _36567_ (.A(_08707_),
    .B(_10761_),
    .Y(_10772_));
 sg13g2_xor2_1 _36568_ (.B(_10772_),
    .A(_08715_),
    .X(_10773_));
 sg13g2_a21oi_2 _36569_ (.B1(_10771_),
    .Y(_10774_),
    .A2(_10773_),
    .A1(net5424));
 sg13g2_nand3_1 _36570_ (.B(net4639),
    .C(_10774_),
    .A(net4631),
    .Y(_10775_));
 sg13g2_a21o_1 _36571_ (.A2(net4639),
    .A1(net4631),
    .B1(_10774_),
    .X(_10776_));
 sg13g2_nand2_1 _36572_ (.Y(_10777_),
    .A(_10775_),
    .B(_10776_));
 sg13g2_o21ai_1 _36573_ (.B1(net4622),
    .Y(_10778_),
    .A1(_10744_),
    .A2(_10763_));
 sg13g2_o21ai_1 _36574_ (.B1(_10778_),
    .Y(_10779_),
    .A1(_10745_),
    .A2(_10751_));
 sg13g2_o21ai_1 _36575_ (.B1(_10779_),
    .Y(_10780_),
    .A1(net4622),
    .A2(_10763_));
 sg13g2_xnor2_1 _36576_ (.Y(_10781_),
    .A(_10777_),
    .B(_10780_));
 sg13g2_nand2_1 _36577_ (.Y(_10782_),
    .A(net4722),
    .B(_10781_));
 sg13g2_o21ai_1 _36578_ (.B1(_10782_),
    .Y(_10783_),
    .A1(net4717),
    .A2(_10774_));
 sg13g2_o21ai_1 _36579_ (.B1(net5608),
    .Y(_10784_),
    .A1(net4433),
    .A2(_10763_));
 sg13g2_a21oi_1 _36580_ (.A1(net4433),
    .A2(_10783_),
    .Y(_10785_),
    .B1(_10784_));
 sg13g2_a21o_1 _36581_ (.A2(net4228),
    .A1(net2963),
    .B1(_10785_),
    .X(_00847_));
 sg13g2_a21oi_1 _36582_ (.A1(_08823_),
    .A2(_10727_),
    .Y(_10786_),
    .B1(_08735_));
 sg13g2_o21ai_1 _36583_ (.B1(_08699_),
    .Y(_10787_),
    .A1(_08830_),
    .A2(_10786_));
 sg13g2_or3_1 _36584_ (.A(_08699_),
    .B(_08830_),
    .C(_10786_),
    .X(_10788_));
 sg13g2_and2_1 _36585_ (.A(_10787_),
    .B(_10788_),
    .X(_10789_));
 sg13g2_mux2_1 _36586_ (.A0(_08697_),
    .A1(_10789_),
    .S(net5424),
    .X(_10790_));
 sg13g2_nand3_1 _36587_ (.B(net4639),
    .C(_10790_),
    .A(net4631),
    .Y(_10791_));
 sg13g2_a21o_1 _36588_ (.A2(net4639),
    .A1(net4631),
    .B1(_10790_),
    .X(_10792_));
 sg13g2_nand2_1 _36589_ (.Y(_10793_),
    .A(_10791_),
    .B(_10792_));
 sg13g2_o21ai_1 _36590_ (.B1(_10775_),
    .Y(_10794_),
    .A1(_10777_),
    .A2(_10780_));
 sg13g2_o21ai_1 _36591_ (.B1(net4722),
    .Y(_10795_),
    .A1(_10793_),
    .A2(_10794_));
 sg13g2_a21o_1 _36592_ (.A2(_10794_),
    .A1(_10793_),
    .B1(_10795_),
    .X(_10796_));
 sg13g2_o21ai_1 _36593_ (.B1(_10796_),
    .Y(_10797_),
    .A1(net4722),
    .A2(_10790_));
 sg13g2_o21ai_1 _36594_ (.B1(net5608),
    .Y(_10798_),
    .A1(net4433),
    .A2(_10774_));
 sg13g2_a21oi_1 _36595_ (.A1(net4433),
    .A2(_10797_),
    .Y(_10799_),
    .B1(_10798_));
 sg13g2_a21o_1 _36596_ (.A2(net4228),
    .A1(net5877),
    .B1(_10799_),
    .X(_00848_));
 sg13g2_nand2_1 _36597_ (.Y(_10800_),
    .A(_08698_),
    .B(_10787_));
 sg13g2_xor2_1 _36598_ (.B(_10800_),
    .A(_08691_),
    .X(_10801_));
 sg13g2_nor2_1 _36599_ (.A(net5424),
    .B(_08689_),
    .Y(_10802_));
 sg13g2_a21oi_2 _36600_ (.B1(_10802_),
    .Y(_10803_),
    .A2(_10801_),
    .A1(net5424));
 sg13g2_nand2_1 _36601_ (.Y(_10804_),
    .A(net4681),
    .B(_10803_));
 sg13g2_nor2_1 _36602_ (.A(net4568),
    .B(_10803_),
    .Y(_10805_));
 sg13g2_xnor2_1 _36603_ (.Y(_10806_),
    .A(net4622),
    .B(_10803_));
 sg13g2_nand4_1 _36604_ (.B(_10776_),
    .C(_10791_),
    .A(_10775_),
    .Y(_10807_),
    .D(_10792_));
 sg13g2_and2_1 _36605_ (.A(_10775_),
    .B(_10791_),
    .X(_10808_));
 sg13g2_o21ai_1 _36606_ (.B1(_10808_),
    .Y(_10809_),
    .A1(_10778_),
    .A2(_10807_));
 sg13g2_or3_1 _36607_ (.A(_10745_),
    .B(_10764_),
    .C(_10807_),
    .X(_10810_));
 sg13g2_nor2_1 _36608_ (.A(_10751_),
    .B(_10810_),
    .Y(_10811_));
 sg13g2_nor2_1 _36609_ (.A(_10809_),
    .B(_10811_),
    .Y(_10812_));
 sg13g2_nor2b_1 _36610_ (.A(_10812_),
    .B_N(_10806_),
    .Y(_10813_));
 sg13g2_xnor2_1 _36611_ (.Y(_10814_),
    .A(_10806_),
    .B(_10812_));
 sg13g2_o21ai_1 _36612_ (.B1(_10804_),
    .Y(_10815_),
    .A1(net4681),
    .A2(_10814_));
 sg13g2_o21ai_1 _36613_ (.B1(net5610),
    .Y(_10816_),
    .A1(net4440),
    .A2(_10790_));
 sg13g2_a21oi_1 _36614_ (.A1(net4440),
    .A2(_10815_),
    .Y(_10817_),
    .B1(_10816_));
 sg13g2_a21o_1 _36615_ (.A2(net4228),
    .A1(net1954),
    .B1(_10817_),
    .X(_00849_));
 sg13g2_nor2_1 _36616_ (.A(net5424),
    .B(_08665_),
    .Y(_10818_));
 sg13g2_a22oi_1 _36617_ (.Y(_10819_),
    .B1(_08825_),
    .B2(_10787_),
    .A2(_08689_),
    .A1(net4825));
 sg13g2_xnor2_1 _36618_ (.Y(_10820_),
    .A(_08668_),
    .B(_10819_));
 sg13g2_a21oi_2 _36619_ (.B1(_10818_),
    .Y(_10821_),
    .A2(_10820_),
    .A1(net5424));
 sg13g2_nand2_1 _36620_ (.Y(_10822_),
    .A(net4568),
    .B(_10821_));
 sg13g2_xnor2_1 _36621_ (.Y(_10823_),
    .A(net4622),
    .B(_10821_));
 sg13g2_nor2_1 _36622_ (.A(_10805_),
    .B(_10813_),
    .Y(_10824_));
 sg13g2_nand2_1 _36623_ (.Y(_10825_),
    .A(net4681),
    .B(_10821_));
 sg13g2_xnor2_1 _36624_ (.Y(_10826_),
    .A(_10823_),
    .B(_10824_));
 sg13g2_o21ai_1 _36625_ (.B1(_10825_),
    .Y(_10827_),
    .A1(net4681),
    .A2(_10826_));
 sg13g2_nand2_1 _36626_ (.Y(_10828_),
    .A(net4440),
    .B(_10827_));
 sg13g2_a21oi_1 _36627_ (.A1(net4370),
    .A2(_10803_),
    .Y(_10829_),
    .B1(net5578));
 sg13g2_a22oi_1 _36628_ (.Y(_10830_),
    .B1(_10828_),
    .B2(_10829_),
    .A2(net4242),
    .A1(net2974));
 sg13g2_inv_1 _36629_ (.Y(_00850_),
    .A(_10830_));
 sg13g2_a21oi_1 _36630_ (.A1(_08671_),
    .A2(_08676_),
    .Y(_10831_),
    .B1(net5424));
 sg13g2_a21oi_1 _36631_ (.A1(_08667_),
    .A2(_10819_),
    .Y(_10832_),
    .B1(_08666_));
 sg13g2_xor2_1 _36632_ (.B(_10832_),
    .A(_08679_),
    .X(_10833_));
 sg13g2_a21oi_2 _36633_ (.B1(_10831_),
    .Y(_10834_),
    .A2(_10833_),
    .A1(net5430));
 sg13g2_nand2_1 _36634_ (.Y(_10835_),
    .A(net4622),
    .B(_10834_));
 sg13g2_xnor2_1 _36635_ (.Y(_10836_),
    .A(net4568),
    .B(_10834_));
 sg13g2_a21o_1 _36636_ (.A2(_10821_),
    .A1(_10803_),
    .B1(net4568),
    .X(_10837_));
 sg13g2_nand2b_1 _36637_ (.Y(_10838_),
    .B(_10837_),
    .A_N(_10813_));
 sg13g2_nand3_1 _36638_ (.B(_10836_),
    .C(_10838_),
    .A(_10822_),
    .Y(_10839_));
 sg13g2_a21o_1 _36639_ (.A2(_10838_),
    .A1(_10822_),
    .B1(_10836_),
    .X(_10840_));
 sg13g2_nand3_1 _36640_ (.B(_10839_),
    .C(_10840_),
    .A(net4725),
    .Y(_10841_));
 sg13g2_nand2_1 _36641_ (.Y(_10842_),
    .A(net4681),
    .B(_10834_));
 sg13g2_nand3_1 _36642_ (.B(_10841_),
    .C(_10842_),
    .A(net4439),
    .Y(_10843_));
 sg13g2_a21oi_1 _36643_ (.A1(net4370),
    .A2(_10821_),
    .Y(_10844_),
    .B1(net5578));
 sg13g2_a22oi_1 _36644_ (.Y(_10845_),
    .B1(_10843_),
    .B2(_10844_),
    .A2(net4242),
    .A1(net3087));
 sg13g2_inv_1 _36645_ (.Y(_00851_),
    .A(_10845_));
 sg13g2_nand2_1 _36646_ (.Y(_10846_),
    .A(net5383),
    .B(_08608_));
 sg13g2_o21ai_1 _36647_ (.B1(_09609_),
    .Y(_10847_),
    .A1(_09245_),
    .A2(net1064));
 sg13g2_a21o_2 _36648_ (.A2(_10847_),
    .A1(_08833_),
    .B1(_08610_),
    .X(_10848_));
 sg13g2_nand3_1 _36649_ (.B(_08833_),
    .C(_10847_),
    .A(_08610_),
    .Y(_10849_));
 sg13g2_nand3_1 _36650_ (.B(_10848_),
    .C(_10849_),
    .A(net5427),
    .Y(_10850_));
 sg13g2_nand2_2 _36651_ (.Y(_10851_),
    .A(_10846_),
    .B(_10850_));
 sg13g2_xnor2_1 _36652_ (.Y(_10852_),
    .A(net4568),
    .B(_10851_));
 sg13g2_nand2_1 _36653_ (.Y(_10853_),
    .A(_10835_),
    .B(_10839_));
 sg13g2_xnor2_1 _36654_ (.Y(_10854_),
    .A(_10852_),
    .B(_10853_));
 sg13g2_nand2_1 _36655_ (.Y(_10855_),
    .A(net4725),
    .B(_10854_));
 sg13g2_o21ai_1 _36656_ (.B1(_10855_),
    .Y(_10856_),
    .A1(net4725),
    .A2(_10851_));
 sg13g2_o21ai_1 _36657_ (.B1(net5610),
    .Y(_10857_),
    .A1(net4439),
    .A2(_10834_));
 sg13g2_a21oi_1 _36658_ (.A1(net4439),
    .A2(_10856_),
    .Y(_10858_),
    .B1(_10857_));
 sg13g2_a21o_1 _36659_ (.A2(net4242),
    .A1(net2306),
    .B1(_10858_),
    .X(_00852_));
 sg13g2_nor2_1 _36660_ (.A(net5427),
    .B(_08639_),
    .Y(_10859_));
 sg13g2_nand2b_1 _36661_ (.Y(_10860_),
    .B(_10848_),
    .A_N(_08609_));
 sg13g2_xnor2_1 _36662_ (.Y(_10861_),
    .A(_08641_),
    .B(_10860_));
 sg13g2_a21oi_2 _36663_ (.B1(_10859_),
    .Y(_10862_),
    .A2(_10861_),
    .A1(net5427));
 sg13g2_inv_1 _36664_ (.Y(_10863_),
    .A(_10862_));
 sg13g2_xnor2_1 _36665_ (.Y(_10864_),
    .A(net4623),
    .B(_10862_));
 sg13g2_nand2_1 _36666_ (.Y(_10865_),
    .A(_10836_),
    .B(_10852_));
 sg13g2_and4_1 _36667_ (.A(_10806_),
    .B(_10823_),
    .C(_10836_),
    .D(_10852_),
    .X(_10866_));
 sg13g2_nor2b_1 _36668_ (.A(_10810_),
    .B_N(_10866_),
    .Y(_10867_));
 sg13g2_nor2b_1 _36669_ (.A(_10749_),
    .B_N(_10867_),
    .Y(_10868_));
 sg13g2_o21ai_1 _36670_ (.B1(net4622),
    .Y(_10869_),
    .A1(_10834_),
    .A2(_10851_));
 sg13g2_o21ai_1 _36671_ (.B1(_10869_),
    .Y(_10870_),
    .A1(_10837_),
    .A2(_10865_));
 sg13g2_and2_1 _36672_ (.A(_10809_),
    .B(_10866_),
    .X(_10871_));
 sg13g2_nor3_1 _36673_ (.A(_10868_),
    .B(_10870_),
    .C(_10871_),
    .Y(_10872_));
 sg13g2_nand3_1 _36674_ (.B(_10747_),
    .C(_10867_),
    .A(_10691_),
    .Y(_10873_));
 sg13g2_nand2b_1 _36675_ (.Y(_10874_),
    .B(_10629_),
    .A_N(_10873_));
 sg13g2_and2_1 _36676_ (.A(_10872_),
    .B(_10874_),
    .X(_10875_));
 sg13g2_nor2_1 _36677_ (.A(_10864_),
    .B(_10875_),
    .Y(_10876_));
 sg13g2_and2_1 _36678_ (.A(_10864_),
    .B(_10875_),
    .X(_10877_));
 sg13g2_o21ai_1 _36679_ (.B1(net4722),
    .Y(_10878_),
    .A1(_10876_),
    .A2(_10877_));
 sg13g2_o21ai_1 _36680_ (.B1(_10878_),
    .Y(_10879_),
    .A1(net4722),
    .A2(_10862_));
 sg13g2_o21ai_1 _36681_ (.B1(net5610),
    .Y(_10880_),
    .A1(net4439),
    .A2(_10851_));
 sg13g2_a21oi_1 _36682_ (.A1(net4439),
    .A2(_10879_),
    .Y(_10881_),
    .B1(_10880_));
 sg13g2_a21o_1 _36683_ (.A2(net4243),
    .A1(net3027),
    .B1(_10881_),
    .X(_00853_));
 sg13g2_nor2_1 _36684_ (.A(net5427),
    .B(_08619_),
    .Y(_10882_));
 sg13g2_a22oi_1 _36685_ (.Y(_10883_),
    .B1(_08835_),
    .B2(_10848_),
    .A2(_08640_),
    .A1(net4826));
 sg13g2_a221oi_1 _36686_ (.B2(_10848_),
    .C1(_08621_),
    .B1(_08835_),
    .A1(net4826),
    .Y(_10884_),
    .A2(_08640_));
 sg13g2_xnor2_1 _36687_ (.Y(_10885_),
    .A(_08621_),
    .B(_10883_));
 sg13g2_a21oi_2 _36688_ (.B1(_10882_),
    .Y(_10886_),
    .A2(_10885_),
    .A1(net5427));
 sg13g2_nand2_1 _36689_ (.Y(_10887_),
    .A(net4682),
    .B(_10886_));
 sg13g2_a21oi_1 _36690_ (.A1(net4623),
    .A2(_10862_),
    .Y(_10888_),
    .B1(_10876_));
 sg13g2_nand2_1 _36691_ (.Y(_10889_),
    .A(net4569),
    .B(_10886_));
 sg13g2_xnor2_1 _36692_ (.Y(_10890_),
    .A(net4623),
    .B(_10886_));
 sg13g2_xnor2_1 _36693_ (.Y(_10891_),
    .A(_10888_),
    .B(_10890_));
 sg13g2_o21ai_1 _36694_ (.B1(_10887_),
    .Y(_10892_),
    .A1(net4682),
    .A2(_10891_));
 sg13g2_o21ai_1 _36695_ (.B1(net5610),
    .Y(_10893_),
    .A1(net4439),
    .A2(_10862_));
 sg13g2_a21oi_1 _36696_ (.A1(net4439),
    .A2(_10892_),
    .Y(_10894_),
    .B1(_10893_));
 sg13g2_a21o_1 _36697_ (.A2(net4242),
    .A1(net2849),
    .B1(_10894_),
    .X(_00854_));
 sg13g2_or3_1 _36698_ (.A(_08620_),
    .B(_08631_),
    .C(_10884_),
    .X(_10895_));
 sg13g2_o21ai_1 _36699_ (.B1(_08631_),
    .Y(_10896_),
    .A1(_08620_),
    .A2(_10884_));
 sg13g2_a21oi_1 _36700_ (.A1(_10895_),
    .A2(_10896_),
    .Y(_10897_),
    .B1(net5383));
 sg13g2_a21oi_2 _36701_ (.B1(_10897_),
    .Y(_10898_),
    .A2(_08630_),
    .A1(net5383));
 sg13g2_nand3_1 _36702_ (.B(net4640),
    .C(_10898_),
    .A(net4632),
    .Y(_10899_));
 sg13g2_a21o_1 _36703_ (.A2(net4640),
    .A1(net4632),
    .B1(_10898_),
    .X(_10900_));
 sg13g2_nand2_1 _36704_ (.Y(_10901_),
    .A(_10899_),
    .B(_10900_));
 sg13g2_a21o_1 _36705_ (.A2(_10886_),
    .A1(_10863_),
    .B1(net4569),
    .X(_10902_));
 sg13g2_o21ai_1 _36706_ (.B1(_10902_),
    .Y(_10903_),
    .A1(_10864_),
    .A2(_10875_));
 sg13g2_nand2_1 _36707_ (.Y(_10904_),
    .A(_10889_),
    .B(_10903_));
 sg13g2_xnor2_1 _36708_ (.Y(_10905_),
    .A(_10901_),
    .B(_10904_));
 sg13g2_nand2_1 _36709_ (.Y(_10906_),
    .A(net4726),
    .B(_10905_));
 sg13g2_o21ai_1 _36710_ (.B1(_10906_),
    .Y(_10907_),
    .A1(net4726),
    .A2(_10898_));
 sg13g2_nand2_1 _36711_ (.Y(_10908_),
    .A(net4439),
    .B(_10907_));
 sg13g2_a21oi_1 _36712_ (.A1(net4370),
    .A2(_10886_),
    .Y(_10909_),
    .B1(net5578));
 sg13g2_a22oi_1 _36713_ (.Y(_10910_),
    .B1(_10908_),
    .B2(_10909_),
    .A2(net4242),
    .A1(net2928));
 sg13g2_inv_1 _36714_ (.Y(_00855_),
    .A(_10910_));
 sg13g2_a21oi_1 _36715_ (.A1(_08833_),
    .A2(_10847_),
    .Y(_10911_),
    .B1(_08643_));
 sg13g2_o21ai_1 _36716_ (.B1(_08601_),
    .Y(_10912_),
    .A1(_08837_),
    .A2(_10911_));
 sg13g2_or3_1 _36717_ (.A(_08601_),
    .B(_08837_),
    .C(_10911_),
    .X(_10913_));
 sg13g2_and2_1 _36718_ (.A(_10912_),
    .B(_10913_),
    .X(_10914_));
 sg13g2_mux2_1 _36719_ (.A0(_08599_),
    .A1(_10914_),
    .S(net5428),
    .X(_10915_));
 sg13g2_nand3_1 _36720_ (.B(net4640),
    .C(_10915_),
    .A(net4632),
    .Y(_10916_));
 sg13g2_a21o_1 _36721_ (.A2(net4640),
    .A1(net4632),
    .B1(_10915_),
    .X(_10917_));
 sg13g2_nand2_1 _36722_ (.Y(_10918_),
    .A(_10916_),
    .B(_10917_));
 sg13g2_o21ai_1 _36723_ (.B1(_10899_),
    .Y(_10919_),
    .A1(_10901_),
    .A2(_10904_));
 sg13g2_o21ai_1 _36724_ (.B1(net4726),
    .Y(_10920_),
    .A1(_10918_),
    .A2(_10919_));
 sg13g2_a21o_1 _36725_ (.A2(_10919_),
    .A1(_10918_),
    .B1(_10920_),
    .X(_10921_));
 sg13g2_o21ai_1 _36726_ (.B1(_10921_),
    .Y(_10922_),
    .A1(net4726),
    .A2(_10915_));
 sg13g2_o21ai_1 _36727_ (.B1(net5612),
    .Y(_10923_),
    .A1(net4444),
    .A2(_10898_));
 sg13g2_a21oi_1 _36728_ (.A1(net4444),
    .A2(_10922_),
    .Y(_10924_),
    .B1(_10923_));
 sg13g2_a21o_1 _36729_ (.A2(net4246),
    .A1(net2448),
    .B1(_10924_),
    .X(_00856_));
 sg13g2_nand2_1 _36730_ (.Y(_10925_),
    .A(_08600_),
    .B(_10912_));
 sg13g2_xnor2_1 _36731_ (.Y(_10926_),
    .A(_08594_),
    .B(_10925_));
 sg13g2_mux2_1 _36732_ (.A0(_08593_),
    .A1(_10926_),
    .S(net5428),
    .X(_10927_));
 sg13g2_nand2_1 _36733_ (.Y(_10928_),
    .A(net4683),
    .B(_10927_));
 sg13g2_nor2_1 _36734_ (.A(net4569),
    .B(_10927_),
    .Y(_10929_));
 sg13g2_xnor2_1 _36735_ (.Y(_10930_),
    .A(net4569),
    .B(_10927_));
 sg13g2_nand4_1 _36736_ (.B(_10900_),
    .C(_10916_),
    .A(_10899_),
    .Y(_10931_),
    .D(_10917_));
 sg13g2_and2_1 _36737_ (.A(_10899_),
    .B(_10916_),
    .X(_10932_));
 sg13g2_o21ai_1 _36738_ (.B1(_10932_),
    .Y(_10933_),
    .A1(_10902_),
    .A2(_10931_));
 sg13g2_nor2_1 _36739_ (.A(_10864_),
    .B(_10931_),
    .Y(_10934_));
 sg13g2_nand3b_1 _36740_ (.B(_10890_),
    .C(_10934_),
    .Y(_10935_),
    .A_N(_10875_));
 sg13g2_nor2b_1 _36741_ (.A(_10933_),
    .B_N(_10935_),
    .Y(_10936_));
 sg13g2_nor2_1 _36742_ (.A(_10930_),
    .B(_10936_),
    .Y(_10937_));
 sg13g2_xor2_1 _36743_ (.B(_10936_),
    .A(_10930_),
    .X(_10938_));
 sg13g2_o21ai_1 _36744_ (.B1(_10928_),
    .Y(_10939_),
    .A1(net4683),
    .A2(_10938_));
 sg13g2_o21ai_1 _36745_ (.B1(net5612),
    .Y(_10940_),
    .A1(net4444),
    .A2(_10915_));
 sg13g2_a21oi_1 _36746_ (.A1(net4444),
    .A2(_10939_),
    .Y(_10941_),
    .B1(_10940_));
 sg13g2_a21o_1 _36747_ (.A2(net4246),
    .A1(net2636),
    .B1(_10941_),
    .X(_00857_));
 sg13g2_nand2_1 _36748_ (.Y(_10942_),
    .A(net5383),
    .B(_08569_));
 sg13g2_a22oi_1 _36749_ (.Y(_10943_),
    .B1(_08839_),
    .B2(_10912_),
    .A2(_08593_),
    .A1(net4828));
 sg13g2_xor2_1 _36750_ (.B(_10943_),
    .A(_08572_),
    .X(_10944_));
 sg13g2_o21ai_1 _36751_ (.B1(_10942_),
    .Y(_10945_),
    .A1(net5383),
    .A2(_10944_));
 sg13g2_nor2_1 _36752_ (.A(_10929_),
    .B(_10937_),
    .Y(_10946_));
 sg13g2_nand2b_1 _36753_ (.Y(_10947_),
    .B(net4570),
    .A_N(_10945_));
 sg13g2_xnor2_1 _36754_ (.Y(_10948_),
    .A(net4624),
    .B(_10945_));
 sg13g2_xor2_1 _36755_ (.B(_10948_),
    .A(_10946_),
    .X(_10949_));
 sg13g2_nand2_1 _36756_ (.Y(_10950_),
    .A(net4726),
    .B(_10949_));
 sg13g2_a21oi_1 _36757_ (.A1(net4682),
    .A2(_10945_),
    .Y(_10951_),
    .B1(net4371));
 sg13g2_a221oi_1 _36758_ (.B2(_10951_),
    .C1(net5579),
    .B1(_10950_),
    .A1(net4371),
    .Y(_10952_),
    .A2(_10927_));
 sg13g2_a21o_1 _36759_ (.A2(net4246),
    .A1(net2810),
    .B1(_10952_),
    .X(_00858_));
 sg13g2_nor2_1 _36760_ (.A(net5428),
    .B(_08580_),
    .Y(_10953_));
 sg13g2_a21oi_1 _36761_ (.A1(_08571_),
    .A2(_10943_),
    .Y(_10954_),
    .B1(_08570_));
 sg13g2_xnor2_1 _36762_ (.Y(_10955_),
    .A(_08581_),
    .B(_10954_));
 sg13g2_a21oi_2 _36763_ (.B1(_10953_),
    .Y(_10956_),
    .A2(_10955_),
    .A1(net5428));
 sg13g2_and2_1 _36764_ (.A(net4624),
    .B(_10956_),
    .X(_10957_));
 sg13g2_xnor2_1 _36765_ (.Y(_10958_),
    .A(net4624),
    .B(_10956_));
 sg13g2_a21o_1 _36766_ (.A2(_10945_),
    .A1(net4624),
    .B1(_10929_),
    .X(_10959_));
 sg13g2_o21ai_1 _36767_ (.B1(_10947_),
    .Y(_10960_),
    .A1(_10937_),
    .A2(_10959_));
 sg13g2_nor2_1 _36768_ (.A(_10958_),
    .B(_10960_),
    .Y(_10961_));
 sg13g2_and2_1 _36769_ (.A(_10958_),
    .B(_10960_),
    .X(_10962_));
 sg13g2_o21ai_1 _36770_ (.B1(net4726),
    .Y(_10963_),
    .A1(_10961_),
    .A2(_10962_));
 sg13g2_o21ai_1 _36771_ (.B1(_10963_),
    .Y(_10964_),
    .A1(net4727),
    .A2(_10956_));
 sg13g2_o21ai_1 _36772_ (.B1(net5612),
    .Y(_10965_),
    .A1(net4445),
    .A2(_10945_));
 sg13g2_a21oi_1 _36773_ (.A1(net4445),
    .A2(_10964_),
    .Y(_10966_),
    .B1(_10965_));
 sg13g2_a21o_1 _36774_ (.A2(net4246),
    .A1(net2468),
    .B1(_10966_),
    .X(_00859_));
 sg13g2_nand2_1 _36775_ (.Y(_10967_),
    .A(net5383),
    .B(_08545_));
 sg13g2_a21oi_2 _36776_ (.B1(_08645_),
    .Y(_10968_),
    .A2(_10847_),
    .A1(_08833_));
 sg13g2_nor3_1 _36777_ (.A(_08547_),
    .B(_08842_),
    .C(_10968_),
    .Y(_10969_));
 sg13g2_o21ai_1 _36778_ (.B1(_08547_),
    .Y(_10970_),
    .A1(_08842_),
    .A2(_10968_));
 sg13g2_nand2_1 _36779_ (.Y(_10971_),
    .A(net5429),
    .B(_10970_));
 sg13g2_o21ai_1 _36780_ (.B1(_10967_),
    .Y(_10972_),
    .A1(_10969_),
    .A2(_10971_));
 sg13g2_xnor2_1 _36781_ (.Y(_10973_),
    .A(net4624),
    .B(_10972_));
 sg13g2_nor2_1 _36782_ (.A(_10957_),
    .B(_10961_),
    .Y(_10974_));
 sg13g2_xnor2_1 _36783_ (.Y(_10975_),
    .A(_10973_),
    .B(_10974_));
 sg13g2_nand2_1 _36784_ (.Y(_10976_),
    .A(net4727),
    .B(_10975_));
 sg13g2_o21ai_1 _36785_ (.B1(_10976_),
    .Y(_10977_),
    .A1(net4727),
    .A2(_10972_));
 sg13g2_o21ai_1 _36786_ (.B1(net5612),
    .Y(_10978_),
    .A1(net4445),
    .A2(_10956_));
 sg13g2_a21oi_1 _36787_ (.A1(net4445),
    .A2(_10977_),
    .Y(_10979_),
    .B1(_10978_));
 sg13g2_a21o_1 _36788_ (.A2(net4246),
    .A1(net2276),
    .B1(_10979_),
    .X(_00860_));
 sg13g2_nand2_1 _36789_ (.Y(_10980_),
    .A(net1524),
    .B(net4246));
 sg13g2_nand2_1 _36790_ (.Y(_10981_),
    .A(net5384),
    .B(_08537_));
 sg13g2_nand2_1 _36791_ (.Y(_10982_),
    .A(_08546_),
    .B(_10970_));
 sg13g2_xor2_1 _36792_ (.B(_10982_),
    .A(_08539_),
    .X(_10983_));
 sg13g2_o21ai_1 _36793_ (.B1(_10981_),
    .Y(_10984_),
    .A1(net5384),
    .A2(_10983_));
 sg13g2_nor2_1 _36794_ (.A(net4570),
    .B(_10984_),
    .Y(_10985_));
 sg13g2_xnor2_1 _36795_ (.Y(_10986_),
    .A(net4625),
    .B(_10984_));
 sg13g2_nor2_1 _36796_ (.A(_10958_),
    .B(_10973_),
    .Y(_10987_));
 sg13g2_nor4_1 _36797_ (.A(_10930_),
    .B(_10948_),
    .C(_10958_),
    .D(_10973_),
    .Y(_10988_));
 sg13g2_a21o_1 _36798_ (.A2(_10972_),
    .A1(net4624),
    .B1(_10957_),
    .X(_10989_));
 sg13g2_a221oi_1 _36799_ (.B2(_10933_),
    .C1(_10989_),
    .B1(_10988_),
    .A1(_10959_),
    .Y(_10990_),
    .A2(_10987_));
 sg13g2_nand3_1 _36800_ (.B(_10934_),
    .C(_10988_),
    .A(_10890_),
    .Y(_10991_));
 sg13g2_o21ai_1 _36801_ (.B1(_10990_),
    .Y(_10992_),
    .A1(_10875_),
    .A2(_10991_));
 sg13g2_and2_1 _36802_ (.A(_10986_),
    .B(_10992_),
    .X(_10993_));
 sg13g2_o21ai_1 _36803_ (.B1(net4727),
    .Y(_10994_),
    .A1(_10986_),
    .A2(_10992_));
 sg13g2_nor2_1 _36804_ (.A(_10993_),
    .B(_10994_),
    .Y(_10995_));
 sg13g2_o21ai_1 _36805_ (.B1(net4447),
    .Y(_10996_),
    .A1(net4728),
    .A2(_10984_));
 sg13g2_nor2_1 _36806_ (.A(_10995_),
    .B(_10996_),
    .Y(_10997_));
 sg13g2_o21ai_1 _36807_ (.B1(net5612),
    .Y(_10998_),
    .A1(net4444),
    .A2(_10972_));
 sg13g2_o21ai_1 _36808_ (.B1(_10980_),
    .Y(_00861_),
    .A1(_10997_),
    .A2(_10998_));
 sg13g2_nor2_1 _36809_ (.A(net5429),
    .B(_08525_),
    .Y(_10999_));
 sg13g2_a22oi_1 _36810_ (.Y(_11000_),
    .B1(_08844_),
    .B2(_10970_),
    .A2(_08537_),
    .A1(net4827));
 sg13g2_xor2_1 _36811_ (.B(_11000_),
    .A(_08527_),
    .X(_11001_));
 sg13g2_a21oi_2 _36812_ (.B1(_10999_),
    .Y(_11002_),
    .A2(_11001_),
    .A1(net5429));
 sg13g2_nor2_1 _36813_ (.A(_10985_),
    .B(_10993_),
    .Y(_11003_));
 sg13g2_nand2_1 _36814_ (.Y(_11004_),
    .A(net4570),
    .B(_11002_));
 sg13g2_xnor2_1 _36815_ (.Y(_11005_),
    .A(net4625),
    .B(_11002_));
 sg13g2_xnor2_1 _36816_ (.Y(_11006_),
    .A(_11003_),
    .B(_11005_));
 sg13g2_o21ai_1 _36817_ (.B1(net4447),
    .Y(_11007_),
    .A1(net4727),
    .A2(_11002_));
 sg13g2_a21oi_1 _36818_ (.A1(net4727),
    .A2(_11006_),
    .Y(_11008_),
    .B1(_11007_));
 sg13g2_a21oi_1 _36819_ (.A1(net4371),
    .A2(_10984_),
    .Y(_11009_),
    .B1(net5579));
 sg13g2_nor2b_1 _36820_ (.A(_11008_),
    .B_N(_11009_),
    .Y(_11010_));
 sg13g2_a21o_1 _36821_ (.A2(net4244),
    .A1(net3270),
    .B1(_11010_),
    .X(_00862_));
 sg13g2_nand2b_1 _36822_ (.Y(_11011_),
    .B(net5384),
    .A_N(_08518_));
 sg13g2_a21oi_1 _36823_ (.A1(_08527_),
    .A2(_11000_),
    .Y(_11012_),
    .B1(_08526_));
 sg13g2_xor2_1 _36824_ (.B(_11012_),
    .A(_08519_),
    .X(_11013_));
 sg13g2_o21ai_1 _36825_ (.B1(_11011_),
    .Y(_11014_),
    .A1(net5384),
    .A2(_11013_));
 sg13g2_nor2_1 _36826_ (.A(net4727),
    .B(_11014_),
    .Y(_11015_));
 sg13g2_nand2_1 _36827_ (.Y(_11016_),
    .A(net4625),
    .B(_11014_));
 sg13g2_xnor2_1 _36828_ (.Y(_11017_),
    .A(net4570),
    .B(_11014_));
 sg13g2_a21oi_1 _36829_ (.A1(_10984_),
    .A2(_11002_),
    .Y(_11018_),
    .B1(net4570));
 sg13g2_or2_1 _36830_ (.X(_11019_),
    .B(_11018_),
    .A(_10993_));
 sg13g2_nand3_1 _36831_ (.B(_11017_),
    .C(_11019_),
    .A(_11004_),
    .Y(_11020_));
 sg13g2_a21o_1 _36832_ (.A2(_11019_),
    .A1(_11004_),
    .B1(_11017_),
    .X(_11021_));
 sg13g2_a21oi_1 _36833_ (.A1(_11020_),
    .A2(_11021_),
    .Y(_11022_),
    .B1(net4683));
 sg13g2_o21ai_1 _36834_ (.B1(net4446),
    .Y(_11023_),
    .A1(_11015_),
    .A2(_11022_));
 sg13g2_a21oi_1 _36835_ (.A1(net4371),
    .A2(_11002_),
    .Y(_11024_),
    .B1(net5579));
 sg13g2_a22oi_1 _36836_ (.Y(_11025_),
    .B1(_11023_),
    .B2(_11024_),
    .A2(net4244),
    .A1(net3047));
 sg13g2_inv_1 _36837_ (.Y(_00863_),
    .A(_11025_));
 sg13g2_nand2_1 _36838_ (.Y(_11026_),
    .A(net2853),
    .B(net4244));
 sg13g2_o21ai_1 _36839_ (.B1(_08548_),
    .Y(_11027_),
    .A1(_08842_),
    .A2(_10968_));
 sg13g2_nand3_1 _36840_ (.B(_08847_),
    .C(_11027_),
    .A(_08505_),
    .Y(_11028_));
 sg13g2_a21oi_1 _36841_ (.A1(_08847_),
    .A2(_11027_),
    .Y(_11029_),
    .B1(_08505_));
 sg13g2_a21o_1 _36842_ (.A2(_11027_),
    .A1(_08847_),
    .B1(_08505_),
    .X(_11030_));
 sg13g2_nand3_1 _36843_ (.B(_11028_),
    .C(_11030_),
    .A(net5429),
    .Y(_11031_));
 sg13g2_o21ai_1 _36844_ (.B1(_11031_),
    .Y(_11032_),
    .A1(net5429),
    .A2(_08503_));
 sg13g2_xnor2_1 _36845_ (.Y(_11033_),
    .A(net4571),
    .B(_11032_));
 sg13g2_nand2_1 _36846_ (.Y(_11034_),
    .A(_11016_),
    .B(_11020_));
 sg13g2_xnor2_1 _36847_ (.Y(_11035_),
    .A(_11033_),
    .B(_11034_));
 sg13g2_a21oi_1 _36848_ (.A1(net4683),
    .A2(_11032_),
    .Y(_11036_),
    .B1(net4371));
 sg13g2_o21ai_1 _36849_ (.B1(_11036_),
    .Y(_11037_),
    .A1(net4683),
    .A2(_11035_));
 sg13g2_o21ai_1 _36850_ (.B1(_11037_),
    .Y(_11038_),
    .A1(net4446),
    .A2(_11014_));
 sg13g2_o21ai_1 _36851_ (.B1(_11026_),
    .Y(_00864_),
    .A1(net5579),
    .A2(_11038_));
 sg13g2_nor2_1 _36852_ (.A(net5428),
    .B(_08496_),
    .Y(_11039_));
 sg13g2_nand2_1 _36853_ (.Y(_11040_),
    .A(_08504_),
    .B(_11030_));
 sg13g2_xnor2_1 _36854_ (.Y(_11041_),
    .A(_08498_),
    .B(_11040_));
 sg13g2_a21oi_2 _36855_ (.B1(_11039_),
    .Y(_11042_),
    .A2(_11041_),
    .A1(net5427));
 sg13g2_nand2_1 _36856_ (.Y(_11043_),
    .A(net4623),
    .B(_11042_));
 sg13g2_xnor2_1 _36857_ (.Y(_11044_),
    .A(net4623),
    .B(_11042_));
 sg13g2_nand3_1 _36858_ (.B(_11018_),
    .C(_11033_),
    .A(_11017_),
    .Y(_11045_));
 sg13g2_o21ai_1 _36859_ (.B1(net4625),
    .Y(_11046_),
    .A1(_11014_),
    .A2(_11032_));
 sg13g2_nand2_1 _36860_ (.Y(_11047_),
    .A(_11045_),
    .B(_11046_));
 sg13g2_and4_1 _36861_ (.A(_10986_),
    .B(_11005_),
    .C(_11017_),
    .D(_11033_),
    .X(_11048_));
 sg13g2_a21oi_1 _36862_ (.A1(_10992_),
    .A2(_11048_),
    .Y(_11049_),
    .B1(_11047_));
 sg13g2_nor2_1 _36863_ (.A(_11044_),
    .B(_11049_),
    .Y(_11050_));
 sg13g2_and2_1 _36864_ (.A(_11044_),
    .B(_11049_),
    .X(_11051_));
 sg13g2_o21ai_1 _36865_ (.B1(net4726),
    .Y(_11052_),
    .A1(_11050_),
    .A2(_11051_));
 sg13g2_o21ai_1 _36866_ (.B1(_11052_),
    .Y(_11053_),
    .A1(net4726),
    .A2(_11042_));
 sg13g2_o21ai_1 _36867_ (.B1(net5612),
    .Y(_11054_),
    .A1(net4446),
    .A2(_11032_));
 sg13g2_a21oi_1 _36868_ (.A1(net4446),
    .A2(_11053_),
    .Y(_11055_),
    .B1(_11054_));
 sg13g2_a21o_1 _36869_ (.A2(net4245),
    .A1(net2667),
    .B1(_11055_),
    .X(_00865_));
 sg13g2_nor2_1 _36870_ (.A(net5427),
    .B(_08486_),
    .Y(_11056_));
 sg13g2_a21oi_1 _36871_ (.A1(_08498_),
    .A2(_11029_),
    .Y(_11057_),
    .B1(_08849_));
 sg13g2_xor2_1 _36872_ (.B(_11057_),
    .A(_08488_),
    .X(_11058_));
 sg13g2_a21oi_2 _36873_ (.B1(_11056_),
    .Y(_11059_),
    .A2(_11058_),
    .A1(net5427));
 sg13g2_nand2_1 _36874_ (.Y(_11060_),
    .A(net4682),
    .B(_11059_));
 sg13g2_o21ai_1 _36875_ (.B1(_11043_),
    .Y(_11061_),
    .A1(_11044_),
    .A2(_11049_));
 sg13g2_nand2_1 _36876_ (.Y(_11062_),
    .A(net4569),
    .B(_11059_));
 sg13g2_xnor2_1 _36877_ (.Y(_11063_),
    .A(net4623),
    .B(_11059_));
 sg13g2_xor2_1 _36878_ (.B(_11063_),
    .A(_11061_),
    .X(_11064_));
 sg13g2_o21ai_1 _36879_ (.B1(_11060_),
    .Y(_11065_),
    .A1(net4682),
    .A2(_11064_));
 sg13g2_o21ai_1 _36880_ (.B1(net5612),
    .Y(_11066_),
    .A1(net4444),
    .A2(_11042_));
 sg13g2_a21oi_1 _36881_ (.A1(net4444),
    .A2(_11065_),
    .Y(_11067_),
    .B1(_11066_));
 sg13g2_a21o_1 _36882_ (.A2(net4245),
    .A1(net2388),
    .B1(_11067_),
    .X(_00866_));
 sg13g2_nor2_1 _36883_ (.A(net5428),
    .B(_08479_),
    .Y(_11068_));
 sg13g2_o21ai_1 _36884_ (.B1(_08487_),
    .Y(_11069_),
    .A1(_08488_),
    .A2(_11057_));
 sg13g2_xor2_1 _36885_ (.B(_11069_),
    .A(_08480_),
    .X(_11070_));
 sg13g2_a21oi_2 _36886_ (.B1(_11068_),
    .Y(_11071_),
    .A2(_11070_),
    .A1(net5428));
 sg13g2_nor2_1 _36887_ (.A(net4722),
    .B(_11071_),
    .Y(_11072_));
 sg13g2_nand2_1 _36888_ (.Y(_11073_),
    .A(net4623),
    .B(_11071_));
 sg13g2_xnor2_1 _36889_ (.Y(_11074_),
    .A(net4569),
    .B(_11071_));
 sg13g2_xnor2_1 _36890_ (.Y(_11075_),
    .A(net4624),
    .B(_11071_));
 sg13g2_o21ai_1 _36891_ (.B1(_11043_),
    .Y(_11076_),
    .A1(net4569),
    .A2(_11059_));
 sg13g2_o21ai_1 _36892_ (.B1(_11062_),
    .Y(_11077_),
    .A1(_11050_),
    .A2(_11076_));
 sg13g2_xnor2_1 _36893_ (.Y(_11078_),
    .A(_11074_),
    .B(_11077_));
 sg13g2_nor2_1 _36894_ (.A(net4682),
    .B(_11078_),
    .Y(_11079_));
 sg13g2_o21ai_1 _36895_ (.B1(net4440),
    .Y(_11080_),
    .A1(_11072_),
    .A2(_11079_));
 sg13g2_a21oi_1 _36896_ (.A1(net4370),
    .A2(_11059_),
    .Y(_11081_),
    .B1(net5578));
 sg13g2_a22oi_1 _36897_ (.Y(_11082_),
    .B1(_11080_),
    .B2(_11081_),
    .A2(net4242),
    .A1(net3315));
 sg13g2_inv_1 _36898_ (.Y(_00867_),
    .A(_11082_));
 sg13g2_nand2_1 _36899_ (.Y(_11083_),
    .A(net5380),
    .B(_08428_));
 sg13g2_nand2_1 _36900_ (.Y(_11084_),
    .A(_08430_),
    .B(_09612_));
 sg13g2_xnor2_1 _36901_ (.Y(_11085_),
    .A(_08430_),
    .B(_09612_));
 sg13g2_o21ai_1 _36902_ (.B1(_11083_),
    .Y(_11086_),
    .A1(net5380),
    .A2(_11085_));
 sg13g2_nand2_1 _36903_ (.Y(_11087_),
    .A(net4623),
    .B(_11086_));
 sg13g2_xnor2_1 _36904_ (.Y(_11088_),
    .A(net4569),
    .B(_11086_));
 sg13g2_o21ai_1 _36905_ (.B1(_11073_),
    .Y(_11089_),
    .A1(_11075_),
    .A2(_11077_));
 sg13g2_xnor2_1 _36906_ (.Y(_11090_),
    .A(_11088_),
    .B(_11089_));
 sg13g2_a21oi_1 _36907_ (.A1(net4682),
    .A2(_11086_),
    .Y(_11091_),
    .B1(net4370));
 sg13g2_o21ai_1 _36908_ (.B1(_11091_),
    .Y(_11092_),
    .A1(net4682),
    .A2(_11090_));
 sg13g2_nor2_1 _36909_ (.A(net4444),
    .B(_11071_),
    .Y(_11093_));
 sg13g2_nor2_1 _36910_ (.A(net5579),
    .B(_11093_),
    .Y(_11094_));
 sg13g2_a22oi_1 _36911_ (.Y(_11095_),
    .B1(_11092_),
    .B2(_11094_),
    .A2(net4246),
    .A1(net2626));
 sg13g2_inv_1 _36912_ (.Y(_00868_),
    .A(_11095_));
 sg13g2_nor2_1 _36913_ (.A(net5425),
    .B(_08420_),
    .Y(_11096_));
 sg13g2_a21oi_1 _36914_ (.A1(_08430_),
    .A2(_09612_),
    .Y(_11097_),
    .B1(_08429_));
 sg13g2_xor2_1 _36915_ (.B(_11097_),
    .A(_08422_),
    .X(_11098_));
 sg13g2_a21oi_2 _36916_ (.B1(_11096_),
    .Y(_11099_),
    .A2(_11098_),
    .A1(net5425));
 sg13g2_and2_1 _36917_ (.A(net4620),
    .B(_11099_),
    .X(_11100_));
 sg13g2_xnor2_1 _36918_ (.Y(_11101_),
    .A(net4621),
    .B(_11099_));
 sg13g2_nor2b_1 _36919_ (.A(_11044_),
    .B_N(_11063_),
    .Y(_11102_));
 sg13g2_nand4_1 _36920_ (.B(_11074_),
    .C(_11088_),
    .A(_11048_),
    .Y(_11103_),
    .D(_11102_));
 sg13g2_or2_1 _36921_ (.X(_11104_),
    .B(_11103_),
    .A(_10991_));
 sg13g2_nor2_1 _36922_ (.A(_10873_),
    .B(_11104_),
    .Y(_11105_));
 sg13g2_nor2_1 _36923_ (.A(_10990_),
    .B(_11103_),
    .Y(_11106_));
 sg13g2_and4_1 _36924_ (.A(_11047_),
    .B(_11074_),
    .C(_11088_),
    .D(_11102_),
    .X(_11107_));
 sg13g2_nand3_1 _36925_ (.B(_11076_),
    .C(_11088_),
    .A(_11074_),
    .Y(_11108_));
 sg13g2_nand3_1 _36926_ (.B(_11087_),
    .C(_11108_),
    .A(_11073_),
    .Y(_11109_));
 sg13g2_nor3_2 _36927_ (.A(_11106_),
    .B(_11107_),
    .C(_11109_),
    .Y(_11110_));
 sg13g2_o21ai_1 _36928_ (.B1(_11110_),
    .Y(_11111_),
    .A1(_10872_),
    .A2(_11104_));
 sg13g2_a21oi_2 _36929_ (.B1(_11111_),
    .Y(_11112_),
    .A2(_11105_),
    .A1(_10629_));
 sg13g2_nor2_1 _36930_ (.A(_11101_),
    .B(_11112_),
    .Y(_11113_));
 sg13g2_xnor2_1 _36931_ (.Y(_11114_),
    .A(_11101_),
    .B(_11112_));
 sg13g2_nand2_1 _36932_ (.Y(_11115_),
    .A(net4722),
    .B(_11114_));
 sg13g2_o21ai_1 _36933_ (.B1(_11115_),
    .Y(_11116_),
    .A1(net4722),
    .A2(_11099_));
 sg13g2_o21ai_1 _36934_ (.B1(net5610),
    .Y(_11117_),
    .A1(net4440),
    .A2(_11086_));
 sg13g2_a21oi_1 _36935_ (.A1(net4440),
    .A2(_11116_),
    .Y(_11118_),
    .B1(_11117_));
 sg13g2_a21o_1 _36936_ (.A2(net4243),
    .A1(net2944),
    .B1(_11118_),
    .X(_00869_));
 sg13g2_nor2_1 _36937_ (.A(net5429),
    .B(_08397_),
    .Y(_11119_));
 sg13g2_a22oi_1 _36938_ (.Y(_11120_),
    .B1(_09615_),
    .B2(_11084_),
    .A2(_08421_),
    .A1(net4823));
 sg13g2_xnor2_1 _36939_ (.Y(_11121_),
    .A(_08401_),
    .B(_11120_));
 sg13g2_a21oi_2 _36940_ (.B1(_11119_),
    .Y(_11122_),
    .A2(_11121_),
    .A1(net5429));
 sg13g2_nand2_1 _36941_ (.Y(_11123_),
    .A(net4683),
    .B(_11122_));
 sg13g2_nor2_1 _36942_ (.A(_11100_),
    .B(_11113_),
    .Y(_11124_));
 sg13g2_nor2_1 _36943_ (.A(net4567),
    .B(_11122_),
    .Y(_11125_));
 sg13g2_nand2_1 _36944_ (.Y(_11126_),
    .A(net4567),
    .B(_11122_));
 sg13g2_nor2b_2 _36945_ (.A(_11125_),
    .B_N(_11126_),
    .Y(_11127_));
 sg13g2_xnor2_1 _36946_ (.Y(_11128_),
    .A(_11124_),
    .B(_11127_));
 sg13g2_o21ai_1 _36947_ (.B1(_11123_),
    .Y(_11129_),
    .A1(net4680),
    .A2(_11128_));
 sg13g2_o21ai_1 _36948_ (.B1(net5610),
    .Y(_11130_),
    .A1(net4443),
    .A2(_11099_));
 sg13g2_a21oi_1 _36949_ (.A1(net4443),
    .A2(_11129_),
    .Y(_11131_),
    .B1(_11130_));
 sg13g2_a21o_1 _36950_ (.A2(net4242),
    .A1(net3044),
    .B1(_11131_),
    .X(_00870_));
 sg13g2_a21oi_1 _36951_ (.A1(_08400_),
    .A2(_11120_),
    .Y(_11132_),
    .B1(_08399_));
 sg13g2_nand2_1 _36952_ (.Y(_11133_),
    .A(net5383),
    .B(_08409_));
 sg13g2_xnor2_1 _36953_ (.Y(_11134_),
    .A(_08410_),
    .B(_11132_));
 sg13g2_o21ai_1 _36954_ (.B1(_11133_),
    .Y(_11135_),
    .A1(net5383),
    .A2(_11134_));
 sg13g2_nor2_1 _36955_ (.A(net4570),
    .B(_11135_),
    .Y(_11136_));
 sg13g2_xnor2_1 _36956_ (.Y(_11137_),
    .A(net4570),
    .B(_11135_));
 sg13g2_nor2_1 _36957_ (.A(_11100_),
    .B(_11125_),
    .Y(_11138_));
 sg13g2_o21ai_1 _36958_ (.B1(_11138_),
    .Y(_11139_),
    .A1(_11101_),
    .A2(_11112_));
 sg13g2_nand2_1 _36959_ (.Y(_11140_),
    .A(_11126_),
    .B(_11139_));
 sg13g2_or2_1 _36960_ (.X(_11141_),
    .B(_11140_),
    .A(_11137_));
 sg13g2_nand2_1 _36961_ (.Y(_11142_),
    .A(net4724),
    .B(_11141_));
 sg13g2_a21oi_1 _36962_ (.A1(_11137_),
    .A2(_11140_),
    .Y(_11143_),
    .B1(_11142_));
 sg13g2_nor2_1 _36963_ (.A(net4724),
    .B(_11135_),
    .Y(_11144_));
 sg13g2_or3_1 _36964_ (.A(net4370),
    .B(_11143_),
    .C(_11144_),
    .X(_11145_));
 sg13g2_a21oi_1 _36965_ (.A1(net4370),
    .A2(_11122_),
    .Y(_11146_),
    .B1(net5578));
 sg13g2_a22oi_1 _36966_ (.Y(_11147_),
    .B1(_11145_),
    .B2(_11146_),
    .A2(net4242),
    .A1(net3104));
 sg13g2_inv_1 _36967_ (.Y(_00871_),
    .A(_11147_));
 sg13g2_nand2_1 _36968_ (.Y(_11148_),
    .A(net5380),
    .B(_08438_));
 sg13g2_a21oi_1 _36969_ (.A1(_08851_),
    .A2(_09611_),
    .Y(_11149_),
    .B1(_08432_));
 sg13g2_nor2_1 _36970_ (.A(_09618_),
    .B(_11149_),
    .Y(_11150_));
 sg13g2_o21ai_1 _36971_ (.B1(_08440_),
    .Y(_11151_),
    .A1(_09618_),
    .A2(_11149_));
 sg13g2_xor2_1 _36972_ (.B(_11150_),
    .A(_08440_),
    .X(_11152_));
 sg13g2_o21ai_1 _36973_ (.B1(_11148_),
    .Y(_11153_),
    .A1(net5380),
    .A2(_11152_));
 sg13g2_xnor2_1 _36974_ (.Y(_11154_),
    .A(net4621),
    .B(_11153_));
 sg13g2_nor2b_1 _36975_ (.A(_11136_),
    .B_N(_11141_),
    .Y(_11155_));
 sg13g2_xnor2_1 _36976_ (.Y(_11156_),
    .A(_11154_),
    .B(_11155_));
 sg13g2_nand2_1 _36977_ (.Y(_11157_),
    .A(net4724),
    .B(_11156_));
 sg13g2_o21ai_1 _36978_ (.B1(_11157_),
    .Y(_11158_),
    .A1(net4724),
    .A2(_11153_));
 sg13g2_nand2_1 _36979_ (.Y(_11159_),
    .A(net4443),
    .B(_11158_));
 sg13g2_a21oi_1 _36980_ (.A1(net4371),
    .A2(_11135_),
    .Y(_11160_),
    .B1(net5578));
 sg13g2_a22oi_1 _36981_ (.Y(_11161_),
    .B1(_11159_),
    .B2(_11160_),
    .A2(net4247),
    .A1(net3381));
 sg13g2_inv_1 _36982_ (.Y(_00872_),
    .A(_11161_));
 sg13g2_nor2_1 _36983_ (.A(net5425),
    .B(_08448_),
    .Y(_11162_));
 sg13g2_nand2_1 _36984_ (.Y(_11163_),
    .A(_08439_),
    .B(_11151_));
 sg13g2_xnor2_1 _36985_ (.Y(_11164_),
    .A(_08450_),
    .B(_11163_));
 sg13g2_a21oi_2 _36986_ (.B1(_11162_),
    .Y(_11165_),
    .A2(_11164_),
    .A1(net5425));
 sg13g2_nand2_1 _36987_ (.Y(_11166_),
    .A(net4620),
    .B(_11165_));
 sg13g2_xnor2_1 _36988_ (.Y(_11167_),
    .A(net4571),
    .B(_11165_));
 sg13g2_or2_1 _36989_ (.X(_11168_),
    .B(_11154_),
    .A(_11137_));
 sg13g2_a21oi_1 _36990_ (.A1(net4621),
    .A2(_11153_),
    .Y(_11169_),
    .B1(_11136_));
 sg13g2_o21ai_1 _36991_ (.B1(_11169_),
    .Y(_11170_),
    .A1(_11138_),
    .A2(_11168_));
 sg13g2_nor2_1 _36992_ (.A(_11101_),
    .B(_11168_),
    .Y(_11171_));
 sg13g2_nand2_1 _36993_ (.Y(_11172_),
    .A(_11127_),
    .B(_11171_));
 sg13g2_nor2_1 _36994_ (.A(_11112_),
    .B(_11172_),
    .Y(_11173_));
 sg13g2_nor3_1 _36995_ (.A(_11167_),
    .B(_11170_),
    .C(_11173_),
    .Y(_11174_));
 sg13g2_o21ai_1 _36996_ (.B1(_11167_),
    .Y(_11175_),
    .A1(_11170_),
    .A2(_11173_));
 sg13g2_nor2_1 _36997_ (.A(net4680),
    .B(_11174_),
    .Y(_11176_));
 sg13g2_a22oi_1 _36998_ (.Y(_11177_),
    .B1(_11175_),
    .B2(_11176_),
    .A2(_11165_),
    .A1(net4680));
 sg13g2_o21ai_1 _36999_ (.B1(net5611),
    .Y(_11178_),
    .A1(net4443),
    .A2(_11153_));
 sg13g2_a21oi_1 _37000_ (.A1(net4443),
    .A2(_11177_),
    .Y(_11179_),
    .B1(_11178_));
 sg13g2_a21o_1 _37001_ (.A2(net4247),
    .A1(net2420),
    .B1(_11179_),
    .X(_00873_));
 sg13g2_nor2_1 _37002_ (.A(net5425),
    .B(_08375_),
    .Y(_11180_));
 sg13g2_a21oi_1 _37003_ (.A1(_09614_),
    .A2(_11151_),
    .Y(_11181_),
    .B1(_08449_));
 sg13g2_xor2_1 _37004_ (.B(_11181_),
    .A(_08378_),
    .X(_11182_));
 sg13g2_a21oi_2 _37005_ (.B1(_11180_),
    .Y(_11183_),
    .A2(_11182_),
    .A1(net5425));
 sg13g2_nand2_1 _37006_ (.Y(_11184_),
    .A(net4680),
    .B(_11183_));
 sg13g2_nor2_1 _37007_ (.A(net4568),
    .B(_11183_),
    .Y(_11185_));
 sg13g2_xnor2_1 _37008_ (.Y(_11186_),
    .A(net4620),
    .B(_11183_));
 sg13g2_nand2_1 _37009_ (.Y(_11187_),
    .A(_11166_),
    .B(_11175_));
 sg13g2_xor2_1 _37010_ (.B(_11187_),
    .A(_11186_),
    .X(_11188_));
 sg13g2_o21ai_1 _37011_ (.B1(_11184_),
    .Y(_11189_),
    .A1(net4680),
    .A2(_11188_));
 sg13g2_o21ai_1 _37012_ (.B1(net5611),
    .Y(_11190_),
    .A1(net4443),
    .A2(_11165_));
 sg13g2_a21oi_1 _37013_ (.A1(net4443),
    .A2(_11189_),
    .Y(_11191_),
    .B1(_11190_));
 sg13g2_a21o_1 _37014_ (.A2(net4243),
    .A1(net2337),
    .B1(_11191_),
    .X(_00874_));
 sg13g2_and2_1 _37015_ (.A(net5381),
    .B(_08386_),
    .X(_11192_));
 sg13g2_a21oi_1 _37016_ (.A1(_08378_),
    .A2(_11181_),
    .Y(_11193_),
    .B1(_08377_));
 sg13g2_xor2_1 _37017_ (.B(_11193_),
    .A(_08387_),
    .X(_11194_));
 sg13g2_a21oi_2 _37018_ (.B1(_11192_),
    .Y(_11195_),
    .A2(_11194_),
    .A1(net5426));
 sg13g2_xnor2_1 _37019_ (.Y(_11196_),
    .A(net4620),
    .B(_11195_));
 sg13g2_a21oi_1 _37020_ (.A1(net4620),
    .A2(_11165_),
    .Y(_11197_),
    .B1(_11185_));
 sg13g2_a22oi_1 _37021_ (.Y(_11198_),
    .B1(_11197_),
    .B2(_11175_),
    .A2(_11183_),
    .A1(net4568));
 sg13g2_nor2b_1 _37022_ (.A(_11196_),
    .B_N(_11198_),
    .Y(_11199_));
 sg13g2_xor2_1 _37023_ (.B(_11198_),
    .A(_11196_),
    .X(_11200_));
 sg13g2_nand2_1 _37024_ (.Y(_11201_),
    .A(net4724),
    .B(_11200_));
 sg13g2_o21ai_1 _37025_ (.B1(_11201_),
    .Y(_11202_),
    .A1(net4724),
    .A2(_11195_));
 sg13g2_nand2_1 _37026_ (.Y(_11203_),
    .A(net4442),
    .B(_11202_));
 sg13g2_a21oi_1 _37027_ (.A1(net4370),
    .A2(_11183_),
    .Y(_11204_),
    .B1(net5578));
 sg13g2_a22oi_1 _37028_ (.Y(_11205_),
    .B1(_11203_),
    .B2(_11204_),
    .A2(net4247),
    .A1(net2612));
 sg13g2_inv_1 _37029_ (.Y(_00875_),
    .A(_11205_));
 sg13g2_and2_1 _37030_ (.A(net5381),
    .B(_08349_),
    .X(_11206_));
 sg13g2_a21oi_1 _37031_ (.A1(_08851_),
    .A2(_09611_),
    .Y(_11207_),
    .B1(_08453_));
 sg13g2_nor2_1 _37032_ (.A(_09622_),
    .B(_11207_),
    .Y(_11208_));
 sg13g2_or2_1 _37033_ (.X(_11209_),
    .B(_11208_),
    .A(_08351_));
 sg13g2_a21oi_1 _37034_ (.A1(_08351_),
    .A2(_11208_),
    .Y(_11210_),
    .B1(net5380));
 sg13g2_a21o_2 _37035_ (.A2(_11210_),
    .A1(_11209_),
    .B1(_11206_),
    .X(_11211_));
 sg13g2_xnor2_1 _37036_ (.Y(_11212_),
    .A(net4620),
    .B(_11211_));
 sg13g2_a21oi_1 _37037_ (.A1(net4620),
    .A2(_11195_),
    .Y(_11213_),
    .B1(_11199_));
 sg13g2_xnor2_1 _37038_ (.Y(_11214_),
    .A(_11212_),
    .B(_11213_));
 sg13g2_nand2_1 _37039_ (.Y(_11215_),
    .A(net4724),
    .B(_11214_));
 sg13g2_o21ai_1 _37040_ (.B1(_11215_),
    .Y(_11216_),
    .A1(net4724),
    .A2(_11211_));
 sg13g2_o21ai_1 _37041_ (.B1(net5611),
    .Y(_11217_),
    .A1(net4442),
    .A2(_11195_));
 sg13g2_a21oi_1 _37042_ (.A1(net4441),
    .A2(_11216_),
    .Y(_11218_),
    .B1(_11217_));
 sg13g2_a21o_1 _37043_ (.A2(net4243),
    .A1(net2327),
    .B1(_11218_),
    .X(_00876_));
 sg13g2_nand2b_1 _37044_ (.Y(_11219_),
    .B(_11209_),
    .A_N(_08350_));
 sg13g2_xnor2_1 _37045_ (.Y(_11220_),
    .A(_08361_),
    .B(_11219_));
 sg13g2_nor2_1 _37046_ (.A(net5380),
    .B(_11220_),
    .Y(_11221_));
 sg13g2_a21oi_2 _37047_ (.B1(_11221_),
    .Y(_11222_),
    .A2(_08359_),
    .A1(net5380));
 sg13g2_nand2_1 _37048_ (.Y(_11223_),
    .A(net4619),
    .B(_11222_));
 sg13g2_xnor2_1 _37049_ (.Y(_11224_),
    .A(net4619),
    .B(_11222_));
 sg13g2_or2_1 _37050_ (.X(_11225_),
    .B(_11212_),
    .A(_11196_));
 sg13g2_nand2_1 _37051_ (.Y(_11226_),
    .A(_11167_),
    .B(_11186_));
 sg13g2_nor2_1 _37052_ (.A(_11225_),
    .B(_11226_),
    .Y(_11227_));
 sg13g2_o21ai_1 _37053_ (.B1(net4620),
    .Y(_11228_),
    .A1(_11195_),
    .A2(_11211_));
 sg13g2_o21ai_1 _37054_ (.B1(_11228_),
    .Y(_11229_),
    .A1(_11197_),
    .A2(_11225_));
 sg13g2_a21o_2 _37055_ (.A2(_11227_),
    .A1(_11170_),
    .B1(_11229_),
    .X(_11230_));
 sg13g2_nand3_1 _37056_ (.B(_11171_),
    .C(_11227_),
    .A(_11127_),
    .Y(_11231_));
 sg13g2_nor2_1 _37057_ (.A(_11112_),
    .B(_11231_),
    .Y(_11232_));
 sg13g2_or2_1 _37058_ (.X(_11233_),
    .B(_11232_),
    .A(_11230_));
 sg13g2_nand2b_1 _37059_ (.Y(_11234_),
    .B(_11233_),
    .A_N(_11224_));
 sg13g2_nand2b_1 _37060_ (.Y(_11235_),
    .B(_11224_),
    .A_N(_11233_));
 sg13g2_a21o_1 _37061_ (.A2(_11235_),
    .A1(_11234_),
    .B1(net4679),
    .X(_11236_));
 sg13g2_o21ai_1 _37062_ (.B1(_11236_),
    .Y(_11237_),
    .A1(net4723),
    .A2(_11222_));
 sg13g2_o21ai_1 _37063_ (.B1(net5611),
    .Y(_11238_),
    .A1(net4442),
    .A2(_11211_));
 sg13g2_a21oi_1 _37064_ (.A1(net4441),
    .A2(_11237_),
    .Y(_11239_),
    .B1(_11238_));
 sg13g2_a21o_1 _37065_ (.A2(net4243),
    .A1(net1640),
    .B1(_11239_),
    .X(_00877_));
 sg13g2_nand2_1 _37066_ (.Y(_11240_),
    .A(_11223_),
    .B(_11234_));
 sg13g2_nand2_1 _37067_ (.Y(_11241_),
    .A(net5380),
    .B(_08340_));
 sg13g2_a22oi_1 _37068_ (.Y(_11242_),
    .B1(_09624_),
    .B2(_11209_),
    .A2(_08359_),
    .A1(net4824));
 sg13g2_xnor2_1 _37069_ (.Y(_11243_),
    .A(_08343_),
    .B(_11242_));
 sg13g2_o21ai_1 _37070_ (.B1(_11241_),
    .Y(_11244_),
    .A1(net5381),
    .A2(_11243_));
 sg13g2_nor2_1 _37071_ (.A(net4618),
    .B(_11244_),
    .Y(_11245_));
 sg13g2_xnor2_1 _37072_ (.Y(_11246_),
    .A(net4567),
    .B(_11244_));
 sg13g2_inv_1 _37073_ (.Y(_11247_),
    .A(_11246_));
 sg13g2_o21ai_1 _37074_ (.B1(net4723),
    .Y(_11248_),
    .A1(_11240_),
    .A2(_11246_));
 sg13g2_a21oi_1 _37075_ (.A1(_11240_),
    .A2(_11246_),
    .Y(_11249_),
    .B1(_11248_));
 sg13g2_a21oi_1 _37076_ (.A1(net4679),
    .A2(_11244_),
    .Y(_11250_),
    .B1(_11249_));
 sg13g2_o21ai_1 _37077_ (.B1(net5611),
    .Y(_11251_),
    .A1(net4441),
    .A2(_11222_));
 sg13g2_a21oi_1 _37078_ (.A1(net4441),
    .A2(_11250_),
    .Y(_11252_),
    .B1(_11251_));
 sg13g2_a21o_1 _37079_ (.A2(net4243),
    .A1(net2321),
    .B1(_11252_),
    .X(_00878_));
 sg13g2_nor2_1 _37080_ (.A(net5425),
    .B(_08333_),
    .Y(_11253_));
 sg13g2_a21oi_1 _37081_ (.A1(_08343_),
    .A2(_11242_),
    .Y(_11254_),
    .B1(_08342_));
 sg13g2_xor2_1 _37082_ (.B(_11254_),
    .A(_08334_),
    .X(_11255_));
 sg13g2_a21oi_2 _37083_ (.B1(_11253_),
    .Y(_11256_),
    .A2(_11255_),
    .A1(net5425));
 sg13g2_and2_1 _37084_ (.A(net4619),
    .B(_11256_),
    .X(_11257_));
 sg13g2_xnor2_1 _37085_ (.Y(_11258_),
    .A(net4618),
    .B(_11256_));
 sg13g2_o21ai_1 _37086_ (.B1(net4618),
    .Y(_11259_),
    .A1(_11222_),
    .A2(_11244_));
 sg13g2_a21oi_1 _37087_ (.A1(_11234_),
    .A2(_11259_),
    .Y(_11260_),
    .B1(_11245_));
 sg13g2_nor2b_1 _37088_ (.A(_11258_),
    .B_N(_11260_),
    .Y(_11261_));
 sg13g2_xor2_1 _37089_ (.B(_11260_),
    .A(_11258_),
    .X(_11262_));
 sg13g2_nand2_1 _37090_ (.Y(_11263_),
    .A(net4723),
    .B(_11262_));
 sg13g2_o21ai_1 _37091_ (.B1(_11263_),
    .Y(_11264_),
    .A1(net4723),
    .A2(_11256_));
 sg13g2_o21ai_1 _37092_ (.B1(net5610),
    .Y(_11265_),
    .A1(net4441),
    .A2(_11244_));
 sg13g2_a21oi_1 _37093_ (.A1(net4441),
    .A2(_11264_),
    .Y(_11266_),
    .B1(_11265_));
 sg13g2_a21o_1 _37094_ (.A2(net4243),
    .A1(net2514),
    .B1(_11266_),
    .X(_00879_));
 sg13g2_nor2_1 _37095_ (.A(net5426),
    .B(_08320_),
    .Y(_11267_));
 sg13g2_o21ai_1 _37096_ (.B1(_08363_),
    .Y(_11268_),
    .A1(_09622_),
    .A2(_11207_));
 sg13g2_nand2_1 _37097_ (.Y(_11269_),
    .A(_09627_),
    .B(_11268_));
 sg13g2_xor2_1 _37098_ (.B(_11269_),
    .A(_08322_),
    .X(_11270_));
 sg13g2_a21oi_2 _37099_ (.B1(_11267_),
    .Y(_11271_),
    .A2(_11270_),
    .A1(net5426));
 sg13g2_nand2_1 _37100_ (.Y(_11272_),
    .A(net4679),
    .B(_11271_));
 sg13g2_nor2_1 _37101_ (.A(net4567),
    .B(_11271_),
    .Y(_11273_));
 sg13g2_xnor2_1 _37102_ (.Y(_11274_),
    .A(net4567),
    .B(_11271_));
 sg13g2_nor2_1 _37103_ (.A(_11257_),
    .B(_11261_),
    .Y(_11275_));
 sg13g2_xor2_1 _37104_ (.B(_11275_),
    .A(_11274_),
    .X(_11276_));
 sg13g2_o21ai_1 _37105_ (.B1(_11272_),
    .Y(_11277_),
    .A1(net4679),
    .A2(_11276_));
 sg13g2_o21ai_1 _37106_ (.B1(net5610),
    .Y(_11278_),
    .A1(net4441),
    .A2(_11256_));
 sg13g2_a21oi_1 _37107_ (.A1(net4441),
    .A2(_11277_),
    .Y(_11279_),
    .B1(_11278_));
 sg13g2_a21o_1 _37108_ (.A2(net4258),
    .A1(net3097),
    .B1(_11279_),
    .X(_00880_));
 sg13g2_a21oi_1 _37109_ (.A1(_08322_),
    .A2(_11269_),
    .Y(_11280_),
    .B1(_08321_));
 sg13g2_xnor2_1 _37110_ (.Y(_11281_),
    .A(_08314_),
    .B(_11280_));
 sg13g2_mux2_1 _37111_ (.A0(_08313_),
    .A1(_11281_),
    .S(net5426),
    .X(_11282_));
 sg13g2_nand2_1 _37112_ (.Y(_11283_),
    .A(net4619),
    .B(_11282_));
 sg13g2_xnor2_1 _37113_ (.Y(_11284_),
    .A(net4619),
    .B(_11282_));
 sg13g2_nor3_1 _37114_ (.A(_11258_),
    .B(_11259_),
    .C(_11274_),
    .Y(_11285_));
 sg13g2_or3_1 _37115_ (.A(_11257_),
    .B(_11273_),
    .C(_11285_),
    .X(_11286_));
 sg13g2_nor4_1 _37116_ (.A(_11224_),
    .B(_11247_),
    .C(_11258_),
    .D(_11274_),
    .Y(_11287_));
 sg13g2_a21oi_1 _37117_ (.A1(_11233_),
    .A2(_11287_),
    .Y(_11288_),
    .B1(_11286_));
 sg13g2_nor2_1 _37118_ (.A(_11284_),
    .B(_11288_),
    .Y(_11289_));
 sg13g2_a21oi_1 _37119_ (.A1(_11284_),
    .A2(_11288_),
    .Y(_11290_),
    .B1(net4679));
 sg13g2_nand2b_1 _37120_ (.Y(_11291_),
    .B(_11290_),
    .A_N(_11289_));
 sg13g2_nand2_1 _37121_ (.Y(_11292_),
    .A(net4679),
    .B(_11282_));
 sg13g2_nand3_1 _37122_ (.B(_11291_),
    .C(_11292_),
    .A(net4442),
    .Y(_11293_));
 sg13g2_a21oi_1 _37123_ (.A1(net4371),
    .A2(_11271_),
    .Y(_11294_),
    .B1(net5578));
 sg13g2_a22oi_1 _37124_ (.Y(_11295_),
    .B1(_11293_),
    .B2(_11294_),
    .A2(net4229),
    .A1(net3231));
 sg13g2_inv_1 _37125_ (.Y(_00881_),
    .A(_11295_));
 sg13g2_nor2_1 _37126_ (.A(net5426),
    .B(_08291_),
    .Y(_11296_));
 sg13g2_a21oi_1 _37127_ (.A1(_09627_),
    .A2(_11268_),
    .Y(_11297_),
    .B1(_08323_));
 sg13g2_o21ai_1 _37128_ (.B1(_08294_),
    .Y(_11298_),
    .A1(_09629_),
    .A2(_11297_));
 sg13g2_nor3_1 _37129_ (.A(_08294_),
    .B(_09629_),
    .C(_11297_),
    .Y(_11299_));
 sg13g2_nor2_1 _37130_ (.A(net5381),
    .B(_11299_),
    .Y(_11300_));
 sg13g2_a21o_2 _37131_ (.A2(_11300_),
    .A1(_11298_),
    .B1(_11296_),
    .X(_11301_));
 sg13g2_o21ai_1 _37132_ (.B1(_11283_),
    .Y(_11302_),
    .A1(_11284_),
    .A2(_11288_));
 sg13g2_nand2_1 _37133_ (.Y(_11303_),
    .A(net4618),
    .B(_11301_));
 sg13g2_nand2b_1 _37134_ (.Y(_11304_),
    .B(net4567),
    .A_N(_11301_));
 sg13g2_nand2_1 _37135_ (.Y(_11305_),
    .A(_11303_),
    .B(_11304_));
 sg13g2_xor2_1 _37136_ (.B(_11305_),
    .A(_11302_),
    .X(_11306_));
 sg13g2_nand2_1 _37137_ (.Y(_11307_),
    .A(net4723),
    .B(_11306_));
 sg13g2_o21ai_1 _37138_ (.B1(_11307_),
    .Y(_11308_),
    .A1(net4723),
    .A2(_11301_));
 sg13g2_o21ai_1 _37139_ (.B1(net5608),
    .Y(_11309_),
    .A1(net4436),
    .A2(_11282_));
 sg13g2_a21oi_1 _37140_ (.A1(net4435),
    .A2(_11308_),
    .Y(_11310_),
    .B1(_11309_));
 sg13g2_a21o_1 _37141_ (.A2(net4229),
    .A1(net2516),
    .B1(_11310_),
    .X(_00882_));
 sg13g2_nor2_1 _37142_ (.A(net5426),
    .B(_08302_),
    .Y(_11311_));
 sg13g2_nand2_1 _37143_ (.Y(_11312_),
    .A(_08292_),
    .B(_11298_));
 sg13g2_xor2_1 _37144_ (.B(_11312_),
    .A(_08303_),
    .X(_11313_));
 sg13g2_a21oi_2 _37145_ (.B1(_11311_),
    .Y(_11314_),
    .A2(_11313_),
    .A1(net5426));
 sg13g2_nand2_1 _37146_ (.Y(_11315_),
    .A(net4618),
    .B(_11314_));
 sg13g2_xnor2_1 _37147_ (.Y(_11316_),
    .A(net4618),
    .B(_11314_));
 sg13g2_nand2_1 _37148_ (.Y(_11317_),
    .A(_11283_),
    .B(_11303_));
 sg13g2_o21ai_1 _37149_ (.B1(_11304_),
    .Y(_11318_),
    .A1(_11289_),
    .A2(_11317_));
 sg13g2_xnor2_1 _37150_ (.Y(_11319_),
    .A(_11316_),
    .B(_11318_));
 sg13g2_nand2_1 _37151_ (.Y(_11320_),
    .A(net4723),
    .B(_11319_));
 sg13g2_o21ai_1 _37152_ (.B1(_11320_),
    .Y(_11321_),
    .A1(net4723),
    .A2(_11314_));
 sg13g2_o21ai_1 _37153_ (.B1(net5609),
    .Y(_11322_),
    .A1(net4436),
    .A2(_11301_));
 sg13g2_a21oi_1 _37154_ (.A1(net4435),
    .A2(_11321_),
    .Y(_11323_),
    .B1(_11322_));
 sg13g2_a21o_1 _37155_ (.A2(net4235),
    .A1(net1421),
    .B1(_11323_),
    .X(_00883_));
 sg13g2_nand2_1 _37156_ (.Y(_11324_),
    .A(net1534),
    .B(net4229));
 sg13g2_nand2_1 _37157_ (.Y(_11325_),
    .A(net5377),
    .B(_08270_));
 sg13g2_a21oi_1 _37158_ (.A1(_08851_),
    .A2(_09611_),
    .Y(_11326_),
    .B1(_08454_));
 sg13g2_nor2_1 _37159_ (.A(_09631_),
    .B(_11326_),
    .Y(_11327_));
 sg13g2_o21ai_1 _37160_ (.B1(_08272_),
    .Y(_11328_),
    .A1(_09631_),
    .A2(_11326_));
 sg13g2_xor2_1 _37161_ (.B(_11327_),
    .A(_08272_),
    .X(_11329_));
 sg13g2_o21ai_1 _37162_ (.B1(_11325_),
    .Y(_11330_),
    .A1(net5377),
    .A2(_11329_));
 sg13g2_xnor2_1 _37163_ (.Y(_11331_),
    .A(net4567),
    .B(_11330_));
 sg13g2_inv_1 _37164_ (.Y(_11332_),
    .A(_11331_));
 sg13g2_o21ai_1 _37165_ (.B1(_11315_),
    .Y(_11333_),
    .A1(_11316_),
    .A2(_11318_));
 sg13g2_xnor2_1 _37166_ (.Y(_11334_),
    .A(_11331_),
    .B(_11333_));
 sg13g2_nand2_1 _37167_ (.Y(_11335_),
    .A(net4720),
    .B(_11334_));
 sg13g2_o21ai_1 _37168_ (.B1(_11335_),
    .Y(_11336_),
    .A1(net4720),
    .A2(_11330_));
 sg13g2_a21oi_1 _37169_ (.A1(net4436),
    .A2(_11336_),
    .Y(_11337_),
    .B1(net5571));
 sg13g2_o21ai_1 _37170_ (.B1(_11337_),
    .Y(_11338_),
    .A1(net4435),
    .A2(_11314_));
 sg13g2_nand2_1 _37171_ (.Y(_00884_),
    .A(_11324_),
    .B(_11338_));
 sg13g2_nor2_1 _37172_ (.A(net5420),
    .B(_08263_),
    .Y(_11339_));
 sg13g2_nand2_1 _37173_ (.Y(_11340_),
    .A(_08271_),
    .B(_11328_));
 sg13g2_xnor2_1 _37174_ (.Y(_11341_),
    .A(_08265_),
    .B(_11340_));
 sg13g2_a21oi_2 _37175_ (.B1(_11339_),
    .Y(_11342_),
    .A2(_11341_),
    .A1(net5420));
 sg13g2_nand2_1 _37176_ (.Y(_11343_),
    .A(net4618),
    .B(_11342_));
 sg13g2_xnor2_1 _37177_ (.Y(_11344_),
    .A(net4615),
    .B(_11342_));
 sg13g2_nor4_1 _37178_ (.A(_11284_),
    .B(_11305_),
    .C(_11316_),
    .D(_11332_),
    .Y(_11345_));
 sg13g2_and2_1 _37179_ (.A(_11287_),
    .B(_11345_),
    .X(_11346_));
 sg13g2_nand3b_1 _37180_ (.B(_11317_),
    .C(_11331_),
    .Y(_11347_),
    .A_N(_11316_));
 sg13g2_o21ai_1 _37181_ (.B1(net4618),
    .Y(_11348_),
    .A1(_11314_),
    .A2(_11330_));
 sg13g2_nand2_1 _37182_ (.Y(_11349_),
    .A(_11347_),
    .B(_11348_));
 sg13g2_a221oi_1 _37183_ (.B2(_11230_),
    .C1(_11349_),
    .B1(_11346_),
    .A1(_11286_),
    .Y(_11350_),
    .A2(_11345_));
 sg13g2_nand2b_2 _37184_ (.Y(_11351_),
    .B(_11346_),
    .A_N(_11231_));
 sg13g2_o21ai_1 _37185_ (.B1(_11350_),
    .Y(_11352_),
    .A1(_11112_),
    .A2(_11351_));
 sg13g2_nand2b_1 _37186_ (.Y(_11353_),
    .B(_11352_),
    .A_N(_11344_));
 sg13g2_nand2b_1 _37187_ (.Y(_11354_),
    .B(_11344_),
    .A_N(_11352_));
 sg13g2_a21o_1 _37188_ (.A2(_11354_),
    .A1(_11353_),
    .B1(net4679),
    .X(_11355_));
 sg13g2_o21ai_1 _37189_ (.B1(_11355_),
    .Y(_11356_),
    .A1(net4720),
    .A2(_11342_));
 sg13g2_o21ai_1 _37190_ (.B1(net5608),
    .Y(_11357_),
    .A1(net4435),
    .A2(_11330_));
 sg13g2_a21oi_1 _37191_ (.A1(net4436),
    .A2(_11356_),
    .Y(_11358_),
    .B1(_11357_));
 sg13g2_a21o_1 _37192_ (.A2(net4229),
    .A1(net2919),
    .B1(_11358_),
    .X(_00885_));
 sg13g2_nand2_1 _37193_ (.Y(_11359_),
    .A(net2437),
    .B(net4229));
 sg13g2_a21oi_1 _37194_ (.A1(_09632_),
    .A2(_11328_),
    .Y(_11360_),
    .B1(_08264_));
 sg13g2_o21ai_1 _37195_ (.B1(net5420),
    .Y(_11361_),
    .A1(_08254_),
    .A2(_11360_));
 sg13g2_a21o_1 _37196_ (.A2(_11360_),
    .A1(_08254_),
    .B1(_11361_),
    .X(_11362_));
 sg13g2_o21ai_1 _37197_ (.B1(_11362_),
    .Y(_11363_),
    .A1(net5420),
    .A2(_08252_));
 sg13g2_nor2_1 _37198_ (.A(net4720),
    .B(_11363_),
    .Y(_11364_));
 sg13g2_nand2_1 _37199_ (.Y(_11365_),
    .A(_11343_),
    .B(_11353_));
 sg13g2_nor2_1 _37200_ (.A(net4615),
    .B(_11363_),
    .Y(_11366_));
 sg13g2_xnor2_1 _37201_ (.Y(_11367_),
    .A(net4615),
    .B(_11363_));
 sg13g2_o21ai_1 _37202_ (.B1(net4720),
    .Y(_11368_),
    .A1(_11365_),
    .A2(_11367_));
 sg13g2_a21oi_1 _37203_ (.A1(_11365_),
    .A2(_11367_),
    .Y(_11369_),
    .B1(_11368_));
 sg13g2_o21ai_1 _37204_ (.B1(net4435),
    .Y(_11370_),
    .A1(_11364_),
    .A2(_11369_));
 sg13g2_o21ai_1 _37205_ (.B1(_11370_),
    .Y(_11371_),
    .A1(net4435),
    .A2(_11342_));
 sg13g2_o21ai_1 _37206_ (.B1(_11359_),
    .Y(_00886_),
    .A1(net5571),
    .A2(_11371_));
 sg13g2_or2_1 _37207_ (.X(_11372_),
    .B(_08245_),
    .A(net5421));
 sg13g2_a21oi_1 _37208_ (.A1(_08254_),
    .A2(_11360_),
    .Y(_11373_),
    .B1(_08253_));
 sg13g2_xnor2_1 _37209_ (.Y(_11374_),
    .A(_08246_),
    .B(_11373_));
 sg13g2_o21ai_1 _37210_ (.B1(_11372_),
    .Y(_11375_),
    .A1(net5379),
    .A2(_11374_));
 sg13g2_nand2_1 _37211_ (.Y(_11376_),
    .A(net4679),
    .B(_11375_));
 sg13g2_nor2_1 _37212_ (.A(net4564),
    .B(_11375_),
    .Y(_11377_));
 sg13g2_nand2_1 _37213_ (.Y(_11378_),
    .A(net4567),
    .B(_11375_));
 sg13g2_xnor2_1 _37214_ (.Y(_11379_),
    .A(net4565),
    .B(_11375_));
 sg13g2_o21ai_1 _37215_ (.B1(net4616),
    .Y(_11380_),
    .A1(_11342_),
    .A2(_11363_));
 sg13g2_a21oi_1 _37216_ (.A1(_11353_),
    .A2(_11380_),
    .Y(_11381_),
    .B1(_11366_));
 sg13g2_xnor2_1 _37217_ (.Y(_11382_),
    .A(_11379_),
    .B(_11381_));
 sg13g2_o21ai_1 _37218_ (.B1(_11376_),
    .Y(_11383_),
    .A1(net4677),
    .A2(_11382_));
 sg13g2_o21ai_1 _37219_ (.B1(net5608),
    .Y(_11384_),
    .A1(net4435),
    .A2(_11363_));
 sg13g2_a21oi_1 _37220_ (.A1(net4435),
    .A2(_11383_),
    .Y(_11385_),
    .B1(_11384_));
 sg13g2_a21o_1 _37221_ (.A2(net4235),
    .A1(net2569),
    .B1(_11385_),
    .X(_00887_));
 sg13g2_and2_1 _37222_ (.A(net5379),
    .B(_08233_),
    .X(_11386_));
 sg13g2_or2_1 _37223_ (.X(_11387_),
    .B(_11327_),
    .A(_08273_));
 sg13g2_a21oi_1 _37224_ (.A1(_09635_),
    .A2(_11387_),
    .Y(_11388_),
    .B1(_08235_));
 sg13g2_nand3_1 _37225_ (.B(_09635_),
    .C(_11387_),
    .A(_08235_),
    .Y(_11389_));
 sg13g2_nor2b_1 _37226_ (.A(_11388_),
    .B_N(_11389_),
    .Y(_11390_));
 sg13g2_a21oi_2 _37227_ (.B1(_11386_),
    .Y(_11391_),
    .A2(_11390_),
    .A1(net5420));
 sg13g2_xnor2_1 _37228_ (.Y(_11392_),
    .A(net4565),
    .B(_11391_));
 sg13g2_a21oi_1 _37229_ (.A1(_11378_),
    .A2(_11381_),
    .Y(_11393_),
    .B1(_11377_));
 sg13g2_xnor2_1 _37230_ (.Y(_11394_),
    .A(_11392_),
    .B(_11393_));
 sg13g2_nor2_1 _37231_ (.A(net4720),
    .B(_11391_),
    .Y(_11395_));
 sg13g2_nor2_1 _37232_ (.A(net4368),
    .B(_11395_),
    .Y(_11396_));
 sg13g2_o21ai_1 _37233_ (.B1(_11396_),
    .Y(_11397_),
    .A1(net4677),
    .A2(_11394_));
 sg13g2_a21oi_1 _37234_ (.A1(net4368),
    .A2(_11375_),
    .Y(_11398_),
    .B1(net5571));
 sg13g2_a22oi_1 _37235_ (.Y(_11399_),
    .B1(_11397_),
    .B2(_11398_),
    .A2(net4229),
    .A1(net2372));
 sg13g2_inv_1 _37236_ (.Y(_00888_),
    .A(_11399_));
 sg13g2_nor2_1 _37237_ (.A(_08234_),
    .B(_11388_),
    .Y(_11400_));
 sg13g2_xnor2_1 _37238_ (.Y(_11401_),
    .A(_08227_),
    .B(_11400_));
 sg13g2_mux2_1 _37239_ (.A0(_08226_),
    .A1(_11401_),
    .S(net5420),
    .X(_11402_));
 sg13g2_xnor2_1 _37240_ (.Y(_11403_),
    .A(net4565),
    .B(_11402_));
 sg13g2_or2_1 _37241_ (.X(_11404_),
    .B(_11392_),
    .A(_11379_));
 sg13g2_a21o_1 _37242_ (.A2(_11391_),
    .A1(_11375_),
    .B1(net4565),
    .X(_11405_));
 sg13g2_o21ai_1 _37243_ (.B1(_11405_),
    .Y(_11406_),
    .A1(_11380_),
    .A2(_11404_));
 sg13g2_nor3_1 _37244_ (.A(_11344_),
    .B(_11367_),
    .C(_11404_),
    .Y(_11407_));
 sg13g2_a21oi_1 _37245_ (.A1(_11352_),
    .A2(_11407_),
    .Y(_11408_),
    .B1(_11406_));
 sg13g2_nor2b_1 _37246_ (.A(_11408_),
    .B_N(_11403_),
    .Y(_11409_));
 sg13g2_xor2_1 _37247_ (.B(_11408_),
    .A(_11403_),
    .X(_11410_));
 sg13g2_nor2_1 _37248_ (.A(net4677),
    .B(_11410_),
    .Y(_11411_));
 sg13g2_a21oi_1 _37249_ (.A1(net4677),
    .A2(_11402_),
    .Y(_11412_),
    .B1(_11411_));
 sg13g2_nand2_1 _37250_ (.Y(_11413_),
    .A(net4434),
    .B(_11412_));
 sg13g2_a21oi_1 _37251_ (.A1(net4368),
    .A2(_11391_),
    .Y(_11414_),
    .B1(net5572));
 sg13g2_a22oi_1 _37252_ (.Y(_11415_),
    .B1(_11413_),
    .B2(_11414_),
    .A2(net4229),
    .A1(net2370));
 sg13g2_inv_1 _37253_ (.Y(_00889_),
    .A(_11415_));
 sg13g2_nor2_1 _37254_ (.A(net5421),
    .B(_08214_),
    .Y(_11416_));
 sg13g2_a21oi_1 _37255_ (.A1(_08227_),
    .A2(_11388_),
    .Y(_11417_),
    .B1(_09637_));
 sg13g2_xnor2_1 _37256_ (.Y(_11418_),
    .A(_08216_),
    .B(_11417_));
 sg13g2_a21oi_2 _37257_ (.B1(_11416_),
    .Y(_11419_),
    .A2(_11418_),
    .A1(net5420));
 sg13g2_inv_1 _37258_ (.Y(_11420_),
    .A(_11419_));
 sg13g2_nand2_1 _37259_ (.Y(_11421_),
    .A(net4678),
    .B(_11419_));
 sg13g2_a21oi_1 _37260_ (.A1(net4615),
    .A2(_11402_),
    .Y(_11422_),
    .B1(_11409_));
 sg13g2_nand2_1 _37261_ (.Y(_11423_),
    .A(net4565),
    .B(_11419_));
 sg13g2_xnor2_1 _37262_ (.Y(_11424_),
    .A(net4615),
    .B(_11419_));
 sg13g2_xnor2_1 _37263_ (.Y(_11425_),
    .A(_11422_),
    .B(_11424_));
 sg13g2_o21ai_1 _37264_ (.B1(_11421_),
    .Y(_11426_),
    .A1(net4678),
    .A2(_11425_));
 sg13g2_o21ai_1 _37265_ (.B1(net5609),
    .Y(_11427_),
    .A1(net4434),
    .A2(_11402_));
 sg13g2_a21oi_1 _37266_ (.A1(net4434),
    .A2(_11426_),
    .Y(_11428_),
    .B1(_11427_));
 sg13g2_a21o_1 _37267_ (.A2(net4234),
    .A1(net2906),
    .B1(_11428_),
    .X(_00890_));
 sg13g2_and3_1 _37268_ (.X(_11429_),
    .A(net5377),
    .B(_08193_),
    .C(_08205_));
 sg13g2_o21ai_1 _37269_ (.B1(_08215_),
    .Y(_11430_),
    .A1(_08217_),
    .A2(_11417_));
 sg13g2_xor2_1 _37270_ (.B(_11430_),
    .A(_08208_),
    .X(_11431_));
 sg13g2_a21oi_2 _37271_ (.B1(_11429_),
    .Y(_11432_),
    .A2(_11431_),
    .A1(net5420));
 sg13g2_nand2b_1 _37272_ (.Y(_11433_),
    .B(net4615),
    .A_N(_11432_));
 sg13g2_xnor2_1 _37273_ (.Y(_11434_),
    .A(net4615),
    .B(_11432_));
 sg13g2_o21ai_1 _37274_ (.B1(net4615),
    .Y(_11435_),
    .A1(_11402_),
    .A2(_11420_));
 sg13g2_nand2b_1 _37275_ (.Y(_11436_),
    .B(_11435_),
    .A_N(_11409_));
 sg13g2_a21o_1 _37276_ (.A2(_11436_),
    .A1(_11423_),
    .B1(_11434_),
    .X(_11437_));
 sg13g2_nand3_1 _37277_ (.B(_11434_),
    .C(_11436_),
    .A(_11423_),
    .Y(_11438_));
 sg13g2_a21oi_1 _37278_ (.A1(_11437_),
    .A2(_11438_),
    .Y(_11439_),
    .B1(net4677));
 sg13g2_a21oi_1 _37279_ (.A1(net4678),
    .A2(_11432_),
    .Y(_11440_),
    .B1(_11439_));
 sg13g2_o21ai_1 _37280_ (.B1(net5609),
    .Y(_11441_),
    .A1(net4368),
    .A2(_11440_));
 sg13g2_a21oi_1 _37281_ (.A1(net4368),
    .A2(_11419_),
    .Y(_11442_),
    .B1(_11441_));
 sg13g2_a21o_1 _37282_ (.A2(net4234),
    .A1(net3066),
    .B1(_11442_),
    .X(_00891_));
 sg13g2_nand2_1 _37283_ (.Y(_11443_),
    .A(net5377),
    .B(_08181_));
 sg13g2_o21ai_1 _37284_ (.B1(_08274_),
    .Y(_11444_),
    .A1(_09631_),
    .A2(_11326_));
 sg13g2_a21oi_1 _37285_ (.A1(_09640_),
    .A2(_11444_),
    .Y(_11445_),
    .B1(_08183_));
 sg13g2_nand3_1 _37286_ (.B(_09640_),
    .C(_11444_),
    .A(_08183_),
    .Y(_11446_));
 sg13g2_nand2_1 _37287_ (.Y(_11447_),
    .A(net5421),
    .B(_11446_));
 sg13g2_o21ai_1 _37288_ (.B1(_11443_),
    .Y(_11448_),
    .A1(_11445_),
    .A2(_11447_));
 sg13g2_nand2_1 _37289_ (.Y(_11449_),
    .A(net4616),
    .B(_11448_));
 sg13g2_xnor2_1 _37290_ (.Y(_11450_),
    .A(net4564),
    .B(_11448_));
 sg13g2_nand2_1 _37291_ (.Y(_11451_),
    .A(_11433_),
    .B(_11438_));
 sg13g2_xor2_1 _37292_ (.B(_11451_),
    .A(_11450_),
    .X(_11452_));
 sg13g2_nand2_1 _37293_ (.Y(_11453_),
    .A(net4719),
    .B(_11452_));
 sg13g2_a21oi_1 _37294_ (.A1(net4677),
    .A2(_11448_),
    .Y(_11454_),
    .B1(net4373));
 sg13g2_a221oi_1 _37295_ (.B2(_11454_),
    .C1(net5571),
    .B1(_11453_),
    .A1(net4369),
    .Y(_11455_),
    .A2(_11432_));
 sg13g2_a21o_1 _37296_ (.A2(net4226),
    .A1(net2638),
    .B1(_11455_),
    .X(_00892_));
 sg13g2_a21oi_1 _37297_ (.A1(net4775),
    .A2(_08181_),
    .Y(_11456_),
    .B1(_11445_));
 sg13g2_xnor2_1 _37298_ (.Y(_11457_),
    .A(_08176_),
    .B(_11456_));
 sg13g2_nor2_1 _37299_ (.A(net5377),
    .B(_11457_),
    .Y(_11458_));
 sg13g2_a21oi_2 _37300_ (.B1(_11458_),
    .Y(_11459_),
    .A2(_08175_),
    .A1(net5377));
 sg13g2_nand2_1 _37301_ (.Y(_11460_),
    .A(net4616),
    .B(_11459_));
 sg13g2_xnor2_1 _37302_ (.Y(_11461_),
    .A(net4616),
    .B(_11459_));
 sg13g2_and2_1 _37303_ (.A(_11403_),
    .B(_11424_),
    .X(_11462_));
 sg13g2_nand4_1 _37304_ (.B(_11434_),
    .C(_11450_),
    .A(_11406_),
    .Y(_11463_),
    .D(_11462_));
 sg13g2_nand3b_1 _37305_ (.B(_11450_),
    .C(_11434_),
    .Y(_11464_),
    .A_N(_11435_));
 sg13g2_nand4_1 _37306_ (.B(_11449_),
    .C(_11463_),
    .A(_11433_),
    .Y(_11465_),
    .D(_11464_));
 sg13g2_nand4_1 _37307_ (.B(_11434_),
    .C(_11450_),
    .A(_11407_),
    .Y(_11466_),
    .D(_11462_));
 sg13g2_inv_1 _37308_ (.Y(_11467_),
    .A(_11466_));
 sg13g2_a21oi_2 _37309_ (.B1(_11465_),
    .Y(_11468_),
    .A2(_11467_),
    .A1(_11352_));
 sg13g2_nor2_1 _37310_ (.A(_11461_),
    .B(_11468_),
    .Y(_11469_));
 sg13g2_xnor2_1 _37311_ (.Y(_11470_),
    .A(_11461_),
    .B(_11468_));
 sg13g2_nand2_1 _37312_ (.Y(_11471_),
    .A(net4719),
    .B(_11470_));
 sg13g2_o21ai_1 _37313_ (.B1(_11471_),
    .Y(_11472_),
    .A1(net4720),
    .A2(_11459_));
 sg13g2_o21ai_1 _37314_ (.B1(net5609),
    .Y(_11473_),
    .A1(net4437),
    .A2(_11448_));
 sg13g2_a21oi_1 _37315_ (.A1(net4437),
    .A2(_11472_),
    .Y(_11474_),
    .B1(_11473_));
 sg13g2_a21o_1 _37316_ (.A2(net4226),
    .A1(net2883),
    .B1(_11474_),
    .X(_00893_));
 sg13g2_nor2_1 _37317_ (.A(net4434),
    .B(_11459_),
    .Y(_11475_));
 sg13g2_nor2_1 _37318_ (.A(net5421),
    .B(_08153_),
    .Y(_11476_));
 sg13g2_a21oi_1 _37319_ (.A1(_08176_),
    .A2(_11445_),
    .Y(_11477_),
    .B1(_09641_));
 sg13g2_xnor2_1 _37320_ (.Y(_11478_),
    .A(_08156_),
    .B(_11477_));
 sg13g2_a21oi_2 _37321_ (.B1(_11476_),
    .Y(_11479_),
    .A2(_11478_),
    .A1(net5421));
 sg13g2_o21ai_1 _37322_ (.B1(_11460_),
    .Y(_11480_),
    .A1(_11461_),
    .A2(_11468_));
 sg13g2_nand2_1 _37323_ (.Y(_11481_),
    .A(net4564),
    .B(_11479_));
 sg13g2_xnor2_1 _37324_ (.Y(_11482_),
    .A(net4564),
    .B(_11479_));
 sg13g2_xnor2_1 _37325_ (.Y(_11483_),
    .A(_11480_),
    .B(_11482_));
 sg13g2_o21ai_1 _37326_ (.B1(net4434),
    .Y(_11484_),
    .A1(net4719),
    .A2(_11479_));
 sg13g2_a21oi_1 _37327_ (.A1(net4719),
    .A2(_11483_),
    .Y(_11485_),
    .B1(_11484_));
 sg13g2_nor3_1 _37328_ (.A(net5571),
    .B(_11475_),
    .C(_11485_),
    .Y(_11486_));
 sg13g2_a21o_1 _37329_ (.A2(net4226),
    .A1(net3068),
    .B1(_11486_),
    .X(_00894_));
 sg13g2_nand2_1 _37330_ (.Y(_11487_),
    .A(net5377),
    .B(_08164_));
 sg13g2_o21ai_1 _37331_ (.B1(_08154_),
    .Y(_11488_),
    .A1(_08155_),
    .A2(_11477_));
 sg13g2_xnor2_1 _37332_ (.Y(_11489_),
    .A(_08166_),
    .B(_11488_));
 sg13g2_o21ai_1 _37333_ (.B1(_11487_),
    .Y(_11490_),
    .A1(net5377),
    .A2(_11489_));
 sg13g2_nand2_1 _37334_ (.Y(_11491_),
    .A(net4616),
    .B(_11490_));
 sg13g2_xnor2_1 _37335_ (.Y(_11492_),
    .A(net4564),
    .B(_11490_));
 sg13g2_o21ai_1 _37336_ (.B1(_11460_),
    .Y(_11493_),
    .A1(net4564),
    .A2(_11479_));
 sg13g2_or2_1 _37337_ (.X(_11494_),
    .B(_11493_),
    .A(_11469_));
 sg13g2_nand3_1 _37338_ (.B(_11492_),
    .C(_11494_),
    .A(_11481_),
    .Y(_11495_));
 sg13g2_a21o_1 _37339_ (.A2(_11494_),
    .A1(_11481_),
    .B1(_11492_),
    .X(_11496_));
 sg13g2_nand3_1 _37340_ (.B(_11495_),
    .C(_11496_),
    .A(net4719),
    .Y(_11497_));
 sg13g2_nand2_1 _37341_ (.Y(_11498_),
    .A(net4677),
    .B(_11490_));
 sg13g2_nand3_1 _37342_ (.B(_11497_),
    .C(_11498_),
    .A(net4434),
    .Y(_11499_));
 sg13g2_a21oi_1 _37343_ (.A1(net4368),
    .A2(_11479_),
    .Y(_11500_),
    .B1(net5571));
 sg13g2_a22oi_1 _37344_ (.Y(_11501_),
    .B1(_11499_),
    .B2(_11500_),
    .A2(net4229),
    .A1(net3287));
 sg13g2_inv_1 _37345_ (.Y(_00895_),
    .A(_11501_));
 sg13g2_nand2_1 _37346_ (.Y(_11502_),
    .A(net2137),
    .B(net4226));
 sg13g2_nand2_1 _37347_ (.Y(_11503_),
    .A(net5376),
    .B(_08143_));
 sg13g2_a21oi_2 _37348_ (.B1(_08185_),
    .Y(_11504_),
    .A2(_11444_),
    .A1(_09640_));
 sg13g2_nor3_1 _37349_ (.A(_08145_),
    .B(_09643_),
    .C(_11504_),
    .Y(_11505_));
 sg13g2_o21ai_1 _37350_ (.B1(_08145_),
    .Y(_11506_),
    .A1(_09643_),
    .A2(_11504_));
 sg13g2_nand2_1 _37351_ (.Y(_11507_),
    .A(net5421),
    .B(_11506_));
 sg13g2_o21ai_1 _37352_ (.B1(_11503_),
    .Y(_11508_),
    .A1(_11505_),
    .A2(_11507_));
 sg13g2_nand2_1 _37353_ (.Y(_11509_),
    .A(net4616),
    .B(_11508_));
 sg13g2_xnor2_1 _37354_ (.Y(_11510_),
    .A(net4564),
    .B(_11508_));
 sg13g2_nand2_1 _37355_ (.Y(_11511_),
    .A(_11491_),
    .B(_11495_));
 sg13g2_o21ai_1 _37356_ (.B1(net4719),
    .Y(_11512_),
    .A1(_11510_),
    .A2(_11511_));
 sg13g2_a21oi_1 _37357_ (.A1(_11510_),
    .A2(_11511_),
    .Y(_11513_),
    .B1(_11512_));
 sg13g2_a21oi_1 _37358_ (.A1(net4677),
    .A2(_11508_),
    .Y(_11514_),
    .B1(_11513_));
 sg13g2_a21oi_1 _37359_ (.A1(net4434),
    .A2(_11514_),
    .Y(_11515_),
    .B1(net5572));
 sg13g2_o21ai_1 _37360_ (.B1(_11515_),
    .Y(_11516_),
    .A1(net4434),
    .A2(_11490_));
 sg13g2_nand2_1 _37361_ (.Y(_00896_),
    .A(_11502_),
    .B(_11516_));
 sg13g2_nand2_1 _37362_ (.Y(_11517_),
    .A(net2621),
    .B(net4226));
 sg13g2_nand3_1 _37363_ (.B(_11493_),
    .C(_11510_),
    .A(_11492_),
    .Y(_11518_));
 sg13g2_nand3_1 _37364_ (.B(_11509_),
    .C(_11518_),
    .A(_11491_),
    .Y(_11519_));
 sg13g2_nor2_1 _37365_ (.A(_11461_),
    .B(_11482_),
    .Y(_11520_));
 sg13g2_nand3_1 _37366_ (.B(_11510_),
    .C(_11520_),
    .A(_11492_),
    .Y(_11521_));
 sg13g2_nor2_1 _37367_ (.A(_11468_),
    .B(_11521_),
    .Y(_11522_));
 sg13g2_nand2b_1 _37368_ (.Y(_11523_),
    .B(_11506_),
    .A_N(_08144_));
 sg13g2_xnor2_1 _37369_ (.Y(_11524_),
    .A(_08138_),
    .B(_11523_));
 sg13g2_nand2_1 _37370_ (.Y(_11525_),
    .A(net5421),
    .B(_11524_));
 sg13g2_o21ai_1 _37371_ (.B1(_11525_),
    .Y(_11526_),
    .A1(net5417),
    .A2(_08137_));
 sg13g2_nor2_1 _37372_ (.A(net4564),
    .B(_11526_),
    .Y(_11527_));
 sg13g2_xnor2_1 _37373_ (.Y(_11528_),
    .A(net4616),
    .B(_11526_));
 sg13g2_o21ai_1 _37374_ (.B1(_11528_),
    .Y(_11529_),
    .A1(_11519_),
    .A2(_11522_));
 sg13g2_or3_1 _37375_ (.A(_11519_),
    .B(_11522_),
    .C(_11528_),
    .X(_11530_));
 sg13g2_and2_1 _37376_ (.A(net4719),
    .B(_11530_),
    .X(_11531_));
 sg13g2_o21ai_1 _37377_ (.B1(net4430),
    .Y(_11532_),
    .A1(net4719),
    .A2(_11526_));
 sg13g2_a21oi_1 _37378_ (.A1(_11529_),
    .A2(_11531_),
    .Y(_11533_),
    .B1(_11532_));
 sg13g2_o21ai_1 _37379_ (.B1(net5607),
    .Y(_11534_),
    .A1(net4430),
    .A2(_11508_));
 sg13g2_o21ai_1 _37380_ (.B1(_11517_),
    .Y(_00897_),
    .A1(_11533_),
    .A2(_11534_));
 sg13g2_nand2_1 _37381_ (.Y(_11535_),
    .A(net4369),
    .B(_11526_));
 sg13g2_nand2_1 _37382_ (.Y(_11536_),
    .A(net5376),
    .B(_08116_));
 sg13g2_o21ai_1 _37383_ (.B1(_08146_),
    .Y(_11537_),
    .A1(_09643_),
    .A2(_11504_));
 sg13g2_a21oi_1 _37384_ (.A1(_09646_),
    .A2(_11537_),
    .Y(_11538_),
    .B1(_08118_));
 sg13g2_nand3_1 _37385_ (.B(_09646_),
    .C(_11537_),
    .A(_08118_),
    .Y(_11539_));
 sg13g2_nand2_1 _37386_ (.Y(_11540_),
    .A(net5417),
    .B(_11539_));
 sg13g2_o21ai_1 _37387_ (.B1(_11536_),
    .Y(_11541_),
    .A1(_11538_),
    .A2(_11540_));
 sg13g2_inv_1 _37388_ (.Y(_11542_),
    .A(_11541_));
 sg13g2_xnor2_1 _37389_ (.Y(_11543_),
    .A(net4561),
    .B(_11541_));
 sg13g2_nor2b_1 _37390_ (.A(_11527_),
    .B_N(_11529_),
    .Y(_11544_));
 sg13g2_a21oi_1 _37391_ (.A1(_11543_),
    .A2(_11544_),
    .Y(_11545_),
    .B1(net4676));
 sg13g2_o21ai_1 _37392_ (.B1(_11545_),
    .Y(_11546_),
    .A1(_11543_),
    .A2(_11544_));
 sg13g2_o21ai_1 _37393_ (.B1(_11546_),
    .Y(_11547_),
    .A1(net4716),
    .A2(_11541_));
 sg13g2_a21oi_1 _37394_ (.A1(net4431),
    .A2(_11547_),
    .Y(_11548_),
    .B1(net5572));
 sg13g2_a22oi_1 _37395_ (.Y(_11549_),
    .B1(_11535_),
    .B2(_11548_),
    .A2(net4226),
    .A1(net2697));
 sg13g2_inv_1 _37396_ (.Y(_00898_),
    .A(_11549_));
 sg13g2_or3_1 _37397_ (.A(_08117_),
    .B(_08129_),
    .C(_11538_),
    .X(_11550_));
 sg13g2_o21ai_1 _37398_ (.B1(_08129_),
    .Y(_11551_),
    .A1(_08117_),
    .A2(_11538_));
 sg13g2_nand3_1 _37399_ (.B(_11550_),
    .C(_11551_),
    .A(net5418),
    .Y(_11552_));
 sg13g2_o21ai_1 _37400_ (.B1(_11552_),
    .Y(_11553_),
    .A1(net5418),
    .A2(_08127_));
 sg13g2_nand2_1 _37401_ (.Y(_11554_),
    .A(net4676),
    .B(_11553_));
 sg13g2_nor2_1 _37402_ (.A(net4563),
    .B(_11553_),
    .Y(_11555_));
 sg13g2_nand2_1 _37403_ (.Y(_11556_),
    .A(net4561),
    .B(_11553_));
 sg13g2_xnor2_1 _37404_ (.Y(_11557_),
    .A(net4561),
    .B(_11553_));
 sg13g2_a21o_1 _37405_ (.A2(_11542_),
    .A1(_11526_),
    .B1(net4561),
    .X(_11558_));
 sg13g2_a22oi_1 _37406_ (.Y(_11559_),
    .B1(_11558_),
    .B2(_11529_),
    .A2(_11542_),
    .A1(net4563));
 sg13g2_xnor2_1 _37407_ (.Y(_11560_),
    .A(_11557_),
    .B(_11559_));
 sg13g2_o21ai_1 _37408_ (.B1(_11554_),
    .Y(_11561_),
    .A1(net4676),
    .A2(_11560_));
 sg13g2_o21ai_1 _37409_ (.B1(net5607),
    .Y(_11562_),
    .A1(net4431),
    .A2(_11541_));
 sg13g2_a21oi_1 _37410_ (.A1(net4431),
    .A2(_11561_),
    .Y(_11563_),
    .B1(_11562_));
 sg13g2_a21o_1 _37411_ (.A2(net4226),
    .A1(net3222),
    .B1(_11563_),
    .X(_00899_));
 sg13g2_nand2_1 _37412_ (.Y(_11564_),
    .A(net5376),
    .B(_07659_));
 sg13g2_nand3_1 _37413_ (.B(_09649_),
    .C(_09651_),
    .A(_09613_),
    .Y(_11565_));
 sg13g2_a21o_1 _37414_ (.A2(_09649_),
    .A1(_09613_),
    .B1(_09651_),
    .X(_11566_));
 sg13g2_nand3_1 _37415_ (.B(_11565_),
    .C(_11566_),
    .A(net5418),
    .Y(_11567_));
 sg13g2_nand2_2 _37416_ (.Y(_11568_),
    .A(_11564_),
    .B(_11567_));
 sg13g2_xnor2_1 _37417_ (.Y(_11569_),
    .A(net4563),
    .B(_11568_));
 sg13g2_a21oi_1 _37418_ (.A1(_11556_),
    .A2(_11559_),
    .Y(_11570_),
    .B1(_11555_));
 sg13g2_xnor2_1 _37419_ (.Y(_11571_),
    .A(_11569_),
    .B(_11570_));
 sg13g2_nand2_1 _37420_ (.Y(_11572_),
    .A(net4716),
    .B(_11571_));
 sg13g2_nand2_1 _37421_ (.Y(_11573_),
    .A(net4676),
    .B(_11568_));
 sg13g2_nand3_1 _37422_ (.B(_11572_),
    .C(_11573_),
    .A(net4430),
    .Y(_11574_));
 sg13g2_a21oi_1 _37423_ (.A1(net4369),
    .A2(_11553_),
    .Y(_11575_),
    .B1(net5572));
 sg13g2_a22oi_1 _37424_ (.Y(_11576_),
    .B1(_11574_),
    .B2(_11575_),
    .A2(net4227),
    .A1(net2443));
 sg13g2_inv_1 _37425_ (.Y(_00900_),
    .A(_11576_));
 sg13g2_nand2b_1 _37426_ (.Y(_11577_),
    .B(_11566_),
    .A_N(_07660_));
 sg13g2_xnor2_1 _37427_ (.Y(_11578_),
    .A(_09650_),
    .B(_11577_));
 sg13g2_nand2_1 _37428_ (.Y(_11579_),
    .A(net5418),
    .B(_11578_));
 sg13g2_o21ai_1 _37429_ (.B1(_11579_),
    .Y(_11580_),
    .A1(net5418),
    .A2(_07653_));
 sg13g2_nand2_1 _37430_ (.Y(_11581_),
    .A(net4614),
    .B(_11580_));
 sg13g2_xnor2_1 _37431_ (.Y(_11582_),
    .A(net4561),
    .B(_11580_));
 sg13g2_nor2b_1 _37432_ (.A(_11557_),
    .B_N(_11569_),
    .Y(_11583_));
 sg13g2_nand2b_2 _37433_ (.Y(_11584_),
    .B(_11569_),
    .A_N(_11557_));
 sg13g2_nand2_1 _37434_ (.Y(_11585_),
    .A(_11528_),
    .B(_11543_));
 sg13g2_nor3_1 _37435_ (.A(_11521_),
    .B(_11584_),
    .C(_11585_),
    .Y(_11586_));
 sg13g2_nor4_1 _37436_ (.A(_11466_),
    .B(_11521_),
    .C(_11584_),
    .D(_11585_),
    .Y(_11587_));
 sg13g2_nor2b_1 _37437_ (.A(_11350_),
    .B_N(_11587_),
    .Y(_11588_));
 sg13g2_and2_1 _37438_ (.A(_11465_),
    .B(_11586_),
    .X(_11589_));
 sg13g2_and4_1 _37439_ (.A(_11519_),
    .B(_11528_),
    .C(_11543_),
    .D(_11583_),
    .X(_11590_));
 sg13g2_a21oi_1 _37440_ (.A1(net4614),
    .A2(_11568_),
    .Y(_11591_),
    .B1(_11555_));
 sg13g2_o21ai_1 _37441_ (.B1(_11591_),
    .Y(_11592_),
    .A1(_11558_),
    .A2(_11584_));
 sg13g2_nor4_1 _37442_ (.A(_11588_),
    .B(_11589_),
    .C(_11590_),
    .D(_11592_),
    .Y(_11593_));
 sg13g2_nand2b_1 _37443_ (.Y(_11594_),
    .B(_11587_),
    .A_N(_11351_));
 sg13g2_o21ai_1 _37444_ (.B1(_11593_),
    .Y(_11595_),
    .A1(_11594_),
    .A2(_11112_));
 sg13g2_nor2_1 _37445_ (.A(_11582_),
    .B(net1067),
    .Y(_11596_));
 sg13g2_nand2_1 _37446_ (.Y(_11597_),
    .A(_11582_),
    .B(net1067));
 sg13g2_nor2_1 _37447_ (.A(net4676),
    .B(_11596_),
    .Y(_11598_));
 sg13g2_a22oi_1 _37448_ (.Y(_11599_),
    .B1(_11597_),
    .B2(_11598_),
    .A2(_11580_),
    .A1(net4676));
 sg13g2_o21ai_1 _37449_ (.B1(net5606),
    .Y(_11600_),
    .A1(net4430),
    .A2(_11568_));
 sg13g2_a21oi_1 _37450_ (.A1(net4430),
    .A2(_11599_),
    .Y(_11601_),
    .B1(_11600_));
 sg13g2_a21o_1 _37451_ (.A2(net4226),
    .A1(net2092),
    .B1(_11601_),
    .X(_00901_));
 sg13g2_nand2_1 _37452_ (.Y(_11602_),
    .A(net2976),
    .B(net4225));
 sg13g2_a22oi_1 _37453_ (.Y(_11603_),
    .B1(_07661_),
    .B2(_11566_),
    .A2(_07653_),
    .A1(net4819));
 sg13g2_xnor2_1 _37454_ (.Y(_11604_),
    .A(_07633_),
    .B(_11603_));
 sg13g2_mux2_1 _37455_ (.A0(_07630_),
    .A1(_11604_),
    .S(net5417),
    .X(_11605_));
 sg13g2_nand2_1 _37456_ (.Y(_11606_),
    .A(_11581_),
    .B(_11597_));
 sg13g2_nand2b_1 _37457_ (.Y(_11607_),
    .B(net4562),
    .A_N(_11605_));
 sg13g2_xnor2_1 _37458_ (.Y(_11608_),
    .A(net4561),
    .B(_11605_));
 sg13g2_xor2_1 _37459_ (.B(_11608_),
    .A(_11606_),
    .X(_11609_));
 sg13g2_a21o_1 _37460_ (.A2(_11605_),
    .A1(net4675),
    .B1(net4369),
    .X(_11610_));
 sg13g2_a21oi_1 _37461_ (.A1(net4716),
    .A2(_11609_),
    .Y(_11611_),
    .B1(_11610_));
 sg13g2_o21ai_1 _37462_ (.B1(net5606),
    .Y(_11612_),
    .A1(net4428),
    .A2(_11580_));
 sg13g2_o21ai_1 _37463_ (.B1(_11602_),
    .Y(_00902_),
    .A1(_11611_),
    .A2(_11612_));
 sg13g2_and2_1 _37464_ (.A(net5376),
    .B(_07642_),
    .X(_11613_));
 sg13g2_a21oi_1 _37465_ (.A1(_07632_),
    .A2(_11603_),
    .Y(_11614_),
    .B1(_07631_));
 sg13g2_xor2_1 _37466_ (.B(_11614_),
    .A(_07644_),
    .X(_11615_));
 sg13g2_a21oi_2 _37467_ (.B1(_11613_),
    .Y(_11616_),
    .A2(_11615_),
    .A1(net5417));
 sg13g2_nand2_1 _37468_ (.Y(_11617_),
    .A(net4614),
    .B(_11616_));
 sg13g2_xnor2_1 _37469_ (.Y(_11618_),
    .A(net4561),
    .B(_11616_));
 sg13g2_o21ai_1 _37470_ (.B1(net4614),
    .Y(_11619_),
    .A1(_11580_),
    .A2(_11605_));
 sg13g2_nand2_1 _37471_ (.Y(_11620_),
    .A(_11597_),
    .B(_11619_));
 sg13g2_a21o_1 _37472_ (.A2(_11620_),
    .A1(_11607_),
    .B1(_11618_),
    .X(_11621_));
 sg13g2_nand3_1 _37473_ (.B(_11618_),
    .C(_11620_),
    .A(_11607_),
    .Y(_11622_));
 sg13g2_and2_1 _37474_ (.A(net4715),
    .B(_11622_),
    .X(_11623_));
 sg13g2_a22oi_1 _37475_ (.Y(_11624_),
    .B1(_11621_),
    .B2(_11623_),
    .A2(_11616_),
    .A1(net4675));
 sg13g2_o21ai_1 _37476_ (.B1(net5606),
    .Y(_11625_),
    .A1(net4428),
    .A2(_11605_));
 sg13g2_a21oi_1 _37477_ (.A1(net4429),
    .A2(_11624_),
    .Y(_11626_),
    .B1(_11625_));
 sg13g2_a21o_1 _37478_ (.A2(net4225),
    .A1(net2610),
    .B1(_11626_),
    .X(_00903_));
 sg13g2_nand2_1 _37479_ (.Y(_11627_),
    .A(net5376),
    .B(_07619_));
 sg13g2_a21oi_1 _37480_ (.A1(_09613_),
    .A2(_09649_),
    .Y(_11628_),
    .B1(_09653_));
 sg13g2_nor2_1 _37481_ (.A(_07663_),
    .B(_11628_),
    .Y(_11629_));
 sg13g2_o21ai_1 _37482_ (.B1(_07621_),
    .Y(_11630_),
    .A1(_07663_),
    .A2(_11628_));
 sg13g2_xor2_1 _37483_ (.B(_11629_),
    .A(_07621_),
    .X(_11631_));
 sg13g2_o21ai_1 _37484_ (.B1(_11627_),
    .Y(_11632_),
    .A1(net5376),
    .A2(_11631_));
 sg13g2_xnor2_1 _37485_ (.Y(_11633_),
    .A(net4561),
    .B(_11632_));
 sg13g2_nand2_1 _37486_ (.Y(_11634_),
    .A(_11617_),
    .B(_11622_));
 sg13g2_a21oi_1 _37487_ (.A1(_11633_),
    .A2(_11634_),
    .Y(_11635_),
    .B1(net4676));
 sg13g2_or2_1 _37488_ (.X(_11636_),
    .B(_11634_),
    .A(_11633_));
 sg13g2_a22oi_1 _37489_ (.Y(_11637_),
    .B1(_11635_),
    .B2(_11636_),
    .A2(_11632_),
    .A1(net4676));
 sg13g2_o21ai_1 _37490_ (.B1(net5606),
    .Y(_11638_),
    .A1(net4430),
    .A2(_11616_));
 sg13g2_a21oi_1 _37491_ (.A1(net4430),
    .A2(_11637_),
    .Y(_11639_),
    .B1(_11638_));
 sg13g2_a21o_1 _37492_ (.A2(net4225),
    .A1(net2317),
    .B1(_11639_),
    .X(_00904_));
 sg13g2_nor2_1 _37493_ (.A(net5417),
    .B(_07610_),
    .Y(_11640_));
 sg13g2_nand2_1 _37494_ (.Y(_11641_),
    .A(_07620_),
    .B(_11630_));
 sg13g2_xnor2_1 _37495_ (.Y(_11642_),
    .A(_07614_),
    .B(_11641_));
 sg13g2_a21oi_2 _37496_ (.B1(_11640_),
    .Y(_11643_),
    .A2(_11642_),
    .A1(net5417));
 sg13g2_nand2_1 _37497_ (.Y(_11644_),
    .A(net4614),
    .B(_11643_));
 sg13g2_xnor2_1 _37498_ (.Y(_11645_),
    .A(net4614),
    .B(_11643_));
 sg13g2_nand2_1 _37499_ (.Y(_11646_),
    .A(_11618_),
    .B(_11633_));
 sg13g2_o21ai_1 _37500_ (.B1(net4614),
    .Y(_11647_),
    .A1(_11616_),
    .A2(_11632_));
 sg13g2_o21ai_1 _37501_ (.B1(_11647_),
    .Y(_11648_),
    .A1(_11619_),
    .A2(_11646_));
 sg13g2_nand4_1 _37502_ (.B(_11608_),
    .C(_11618_),
    .A(_11582_),
    .Y(_11649_),
    .D(_11633_));
 sg13g2_inv_1 _37503_ (.Y(_11650_),
    .A(_11649_));
 sg13g2_a21oi_1 _37504_ (.A1(net1067),
    .A2(_11650_),
    .Y(_11651_),
    .B1(_11648_));
 sg13g2_xnor2_1 _37505_ (.Y(_11652_),
    .A(_11645_),
    .B(_11651_));
 sg13g2_nand2_1 _37506_ (.Y(_11653_),
    .A(net4716),
    .B(_11652_));
 sg13g2_o21ai_1 _37507_ (.B1(_11653_),
    .Y(_11654_),
    .A1(net4716),
    .A2(_11643_));
 sg13g2_o21ai_1 _37508_ (.B1(net5604),
    .Y(_11655_),
    .A1(net4430),
    .A2(_11632_));
 sg13g2_a21oi_1 _37509_ (.A1(net4424),
    .A2(_11654_),
    .Y(_11656_),
    .B1(_11655_));
 sg13g2_a21o_1 _37510_ (.A2(net4211),
    .A1(net2693),
    .B1(_11656_),
    .X(_00905_));
 sg13g2_nand2_1 _37511_ (.Y(_11657_),
    .A(net2470),
    .B(net4211));
 sg13g2_nor2_1 _37512_ (.A(net4424),
    .B(_11643_),
    .Y(_11658_));
 sg13g2_nand2_1 _37513_ (.Y(_11659_),
    .A(net5379),
    .B(_07597_));
 sg13g2_a22oi_1 _37514_ (.Y(_11660_),
    .B1(_07664_),
    .B2(_11630_),
    .A2(_07611_),
    .A1(net4819));
 sg13g2_xor2_1 _37515_ (.B(_11660_),
    .A(_07600_),
    .X(_11661_));
 sg13g2_o21ai_1 _37516_ (.B1(_11659_),
    .Y(_11662_),
    .A1(net5379),
    .A2(_11661_));
 sg13g2_o21ai_1 _37517_ (.B1(_11644_),
    .Y(_11663_),
    .A1(_11645_),
    .A2(_11651_));
 sg13g2_nand2b_1 _37518_ (.Y(_11664_),
    .B(net4560),
    .A_N(_11662_));
 sg13g2_xnor2_1 _37519_ (.Y(_11665_),
    .A(net4611),
    .B(_11662_));
 sg13g2_xnor2_1 _37520_ (.Y(_11666_),
    .A(_11663_),
    .B(_11665_));
 sg13g2_mux2_1 _37521_ (.A0(_11662_),
    .A1(_11666_),
    .S(net4714),
    .X(_11667_));
 sg13g2_o21ai_1 _37522_ (.B1(net5604),
    .Y(_11668_),
    .A1(net4365),
    .A2(_11667_));
 sg13g2_o21ai_1 _37523_ (.B1(_11657_),
    .Y(_00906_),
    .A1(_11658_),
    .A2(_11668_));
 sg13g2_a21oi_1 _37524_ (.A1(_07576_),
    .A2(_07587_),
    .Y(_11669_),
    .B1(net5417));
 sg13g2_a21oi_1 _37525_ (.A1(_07599_),
    .A2(_11660_),
    .Y(_11670_),
    .B1(_07598_));
 sg13g2_xnor2_1 _37526_ (.Y(_11671_),
    .A(_07590_),
    .B(_11670_));
 sg13g2_a21oi_2 _37527_ (.B1(_11669_),
    .Y(_11672_),
    .A2(_11671_),
    .A1(net5417));
 sg13g2_nand2_1 _37528_ (.Y(_11673_),
    .A(net4611),
    .B(_11672_));
 sg13g2_xnor2_1 _37529_ (.Y(_11674_),
    .A(net4560),
    .B(_11672_));
 sg13g2_o21ai_1 _37530_ (.B1(net4611),
    .Y(_11675_),
    .A1(_11643_),
    .A2(_11662_));
 sg13g2_o21ai_1 _37531_ (.B1(_11675_),
    .Y(_11676_),
    .A1(_11645_),
    .A2(_11651_));
 sg13g2_a21o_1 _37532_ (.A2(_11676_),
    .A1(_11664_),
    .B1(_11674_),
    .X(_11677_));
 sg13g2_nand3_1 _37533_ (.B(_11674_),
    .C(_11676_),
    .A(_11664_),
    .Y(_11678_));
 sg13g2_and2_1 _37534_ (.A(net4713),
    .B(_11678_),
    .X(_11679_));
 sg13g2_a22oi_1 _37535_ (.Y(_11680_),
    .B1(_11677_),
    .B2(_11679_),
    .A2(_11672_),
    .A1(net4673));
 sg13g2_o21ai_1 _37536_ (.B1(net5604),
    .Y(_11681_),
    .A1(net4425),
    .A2(_11662_));
 sg13g2_a21oi_1 _37537_ (.A1(net4425),
    .A2(_11680_),
    .Y(_11682_),
    .B1(_11681_));
 sg13g2_a21o_1 _37538_ (.A2(net4211),
    .A1(net3074),
    .B1(_11682_),
    .X(_00907_));
 sg13g2_nand2_1 _37539_ (.Y(_11683_),
    .A(net2632),
    .B(net4212));
 sg13g2_nand2_1 _37540_ (.Y(_11684_),
    .A(net5374),
    .B(_07552_));
 sg13g2_a21o_1 _37541_ (.A2(_09649_),
    .A1(_09613_),
    .B1(_09654_),
    .X(_11685_));
 sg13g2_nand2_1 _37542_ (.Y(_11686_),
    .A(_07667_),
    .B(_11685_));
 sg13g2_a21o_1 _37543_ (.A2(_11685_),
    .A1(_07667_),
    .B1(_07555_),
    .X(_11687_));
 sg13g2_xnor2_1 _37544_ (.Y(_11688_),
    .A(_07554_),
    .B(_11686_));
 sg13g2_o21ai_1 _37545_ (.B1(_11684_),
    .Y(_11689_),
    .A1(net5374),
    .A2(_11688_));
 sg13g2_nand2_1 _37546_ (.Y(_11690_),
    .A(net4611),
    .B(_11689_));
 sg13g2_xnor2_1 _37547_ (.Y(_11691_),
    .A(net4559),
    .B(_11689_));
 sg13g2_nand2_1 _37548_ (.Y(_11692_),
    .A(_11673_),
    .B(_11678_));
 sg13g2_o21ai_1 _37549_ (.B1(net4714),
    .Y(_11693_),
    .A1(_11691_),
    .A2(_11692_));
 sg13g2_a21oi_1 _37550_ (.A1(_11691_),
    .A2(_11692_),
    .Y(_11694_),
    .B1(_11693_));
 sg13g2_a21oi_1 _37551_ (.A1(net4673),
    .A2(_11689_),
    .Y(_11695_),
    .B1(_11694_));
 sg13g2_a21oi_1 _37552_ (.A1(net4425),
    .A2(_11695_),
    .Y(_11696_),
    .B1(net5564));
 sg13g2_o21ai_1 _37553_ (.B1(_11696_),
    .Y(_11697_),
    .A1(net4425),
    .A2(_11672_));
 sg13g2_nand2_1 _37554_ (.Y(_00908_),
    .A(_11683_),
    .B(_11697_));
 sg13g2_nand2_1 _37555_ (.Y(_11698_),
    .A(net5374),
    .B(_07564_));
 sg13g2_nand2b_1 _37556_ (.Y(_11699_),
    .B(_11687_),
    .A_N(_07553_));
 sg13g2_xor2_1 _37557_ (.B(_11699_),
    .A(_07566_),
    .X(_11700_));
 sg13g2_o21ai_1 _37558_ (.B1(_11698_),
    .Y(_11701_),
    .A1(net5374),
    .A2(_11700_));
 sg13g2_nand2_1 _37559_ (.Y(_11702_),
    .A(net4672),
    .B(_11701_));
 sg13g2_or2_1 _37560_ (.X(_11703_),
    .B(_11701_),
    .A(net4559));
 sg13g2_xnor2_1 _37561_ (.Y(_11704_),
    .A(net4559),
    .B(_11701_));
 sg13g2_nor2_1 _37562_ (.A(_11645_),
    .B(_11665_),
    .Y(_11705_));
 sg13g2_nand3_1 _37563_ (.B(_11691_),
    .C(_11705_),
    .A(_11674_),
    .Y(_11706_));
 sg13g2_nand2b_1 _37564_ (.Y(_11707_),
    .B(_11648_),
    .A_N(_11706_));
 sg13g2_nand3b_1 _37565_ (.B(_11691_),
    .C(_11674_),
    .Y(_11708_),
    .A_N(_11675_));
 sg13g2_nand4_1 _37566_ (.B(_11690_),
    .C(_11707_),
    .A(_11673_),
    .Y(_11709_),
    .D(_11708_));
 sg13g2_nor2_2 _37567_ (.A(_11649_),
    .B(_11706_),
    .Y(_11710_));
 sg13g2_a21oi_2 _37568_ (.B1(_11709_),
    .Y(_11711_),
    .A2(_11710_),
    .A1(net1067));
 sg13g2_xor2_1 _37569_ (.B(_11711_),
    .A(_11704_),
    .X(_11712_));
 sg13g2_o21ai_1 _37570_ (.B1(_11702_),
    .Y(_11713_),
    .A1(net4673),
    .A2(_11712_));
 sg13g2_o21ai_1 _37571_ (.B1(net5605),
    .Y(_11714_),
    .A1(net4425),
    .A2(_11689_));
 sg13g2_a21oi_1 _37572_ (.A1(net4425),
    .A2(_11713_),
    .Y(_11715_),
    .B1(_11714_));
 sg13g2_a21o_1 _37573_ (.A2(net4212),
    .A1(net2996),
    .B1(_11715_),
    .X(_00909_));
 sg13g2_nor2_1 _37574_ (.A(net5414),
    .B(_07542_),
    .Y(_11716_));
 sg13g2_nand2_1 _37575_ (.Y(_11717_),
    .A(_07669_),
    .B(_11687_));
 sg13g2_a221oi_1 _37576_ (.B2(_11687_),
    .C1(_07545_),
    .B1(_07669_),
    .A1(net4816),
    .Y(_11718_),
    .A2(_07564_));
 sg13g2_a21oi_1 _37577_ (.A1(_07565_),
    .A2(_11717_),
    .Y(_11719_),
    .B1(_07544_));
 sg13g2_nor2_1 _37578_ (.A(_11718_),
    .B(_11719_),
    .Y(_11720_));
 sg13g2_a21oi_2 _37579_ (.B1(_11716_),
    .Y(_11721_),
    .A2(_11720_),
    .A1(net5414));
 sg13g2_and2_1 _37580_ (.A(net4672),
    .B(_11721_),
    .X(_11722_));
 sg13g2_o21ai_1 _37581_ (.B1(_11703_),
    .Y(_11723_),
    .A1(_11704_),
    .A2(_11711_));
 sg13g2_nand2_1 _37582_ (.Y(_11724_),
    .A(net4559),
    .B(_11721_));
 sg13g2_xnor2_1 _37583_ (.Y(_11725_),
    .A(net4610),
    .B(_11721_));
 sg13g2_xnor2_1 _37584_ (.Y(_11726_),
    .A(_11723_),
    .B(_11725_));
 sg13g2_a21oi_1 _37585_ (.A1(net4713),
    .A2(_11726_),
    .Y(_11727_),
    .B1(_11722_));
 sg13g2_o21ai_1 _37586_ (.B1(net5604),
    .Y(_11728_),
    .A1(net4365),
    .A2(_11727_));
 sg13g2_a21oi_1 _37587_ (.A1(net4366),
    .A2(_11701_),
    .Y(_11729_),
    .B1(_11728_));
 sg13g2_a21o_1 _37588_ (.A2(net4212),
    .A1(net2145),
    .B1(_11729_),
    .X(_00910_));
 sg13g2_or3_1 _37589_ (.A(_07537_),
    .B(_07543_),
    .C(_11718_),
    .X(_11730_));
 sg13g2_o21ai_1 _37590_ (.B1(_07537_),
    .Y(_11731_),
    .A1(_07543_),
    .A2(_11718_));
 sg13g2_a21oi_1 _37591_ (.A1(_11730_),
    .A2(_11731_),
    .Y(_11732_),
    .B1(net5374));
 sg13g2_a21oi_2 _37592_ (.B1(_11732_),
    .Y(_11733_),
    .A2(_07536_),
    .A1(net5375));
 sg13g2_nor2_1 _37593_ (.A(net4713),
    .B(_11733_),
    .Y(_11734_));
 sg13g2_nand2_1 _37594_ (.Y(_11735_),
    .A(net4611),
    .B(_11733_));
 sg13g2_xnor2_1 _37595_ (.Y(_11736_),
    .A(net4559),
    .B(_11733_));
 sg13g2_a21o_1 _37596_ (.A2(_11721_),
    .A1(_11701_),
    .B1(net4560),
    .X(_11737_));
 sg13g2_o21ai_1 _37597_ (.B1(_11737_),
    .Y(_11738_),
    .A1(_11704_),
    .A2(_11711_));
 sg13g2_a21o_1 _37598_ (.A2(_11738_),
    .A1(_11724_),
    .B1(_11736_),
    .X(_11739_));
 sg13g2_nand3_1 _37599_ (.B(_11736_),
    .C(_11738_),
    .A(_11724_),
    .Y(_11740_));
 sg13g2_a21oi_1 _37600_ (.A1(_11739_),
    .A2(_11740_),
    .Y(_11741_),
    .B1(net4672));
 sg13g2_o21ai_1 _37601_ (.B1(net4424),
    .Y(_11742_),
    .A1(_11734_),
    .A2(_11741_));
 sg13g2_a21oi_1 _37602_ (.A1(net4366),
    .A2(_11721_),
    .Y(_11743_),
    .B1(net5564));
 sg13g2_a22oi_1 _37603_ (.Y(_11744_),
    .B1(_11742_),
    .B2(_11743_),
    .A2(net4212),
    .A1(net3235));
 sg13g2_inv_1 _37604_ (.Y(_00911_),
    .A(_11744_));
 sg13g2_nand2_1 _37605_ (.Y(_11745_),
    .A(net1969),
    .B(net4212));
 sg13g2_nand2_1 _37606_ (.Y(_11746_),
    .A(net5374),
    .B(_07524_));
 sg13g2_a21oi_1 _37607_ (.A1(_07667_),
    .A2(_11685_),
    .Y(_11747_),
    .B1(_07567_));
 sg13g2_nor3_1 _37608_ (.A(_07526_),
    .B(_07671_),
    .C(_11747_),
    .Y(_11748_));
 sg13g2_o21ai_1 _37609_ (.B1(_07526_),
    .Y(_11749_),
    .A1(_07671_),
    .A2(_11747_));
 sg13g2_nand2_1 _37610_ (.Y(_11750_),
    .A(net5414),
    .B(_11749_));
 sg13g2_o21ai_1 _37611_ (.B1(_11746_),
    .Y(_11751_),
    .A1(_11748_),
    .A2(_11750_));
 sg13g2_xnor2_1 _37612_ (.Y(_11752_),
    .A(net4559),
    .B(_11751_));
 sg13g2_nand2_1 _37613_ (.Y(_11753_),
    .A(_11735_),
    .B(_11740_));
 sg13g2_o21ai_1 _37614_ (.B1(net4713),
    .Y(_11754_),
    .A1(_11752_),
    .A2(_11753_));
 sg13g2_a21oi_1 _37615_ (.A1(_11752_),
    .A2(_11753_),
    .Y(_11755_),
    .B1(_11754_));
 sg13g2_a21oi_1 _37616_ (.A1(net4672),
    .A2(_11751_),
    .Y(_11756_),
    .B1(_11755_));
 sg13g2_a21oi_1 _37617_ (.A1(net4424),
    .A2(_11756_),
    .Y(_11757_),
    .B1(net5564));
 sg13g2_o21ai_1 _37618_ (.B1(_11757_),
    .Y(_11758_),
    .A1(net4424),
    .A2(_11733_));
 sg13g2_nand2_1 _37619_ (.Y(_00912_),
    .A(_11745_),
    .B(_11758_));
 sg13g2_nand2_1 _37620_ (.Y(_11759_),
    .A(_07525_),
    .B(_11749_));
 sg13g2_xor2_1 _37621_ (.B(_11759_),
    .A(_07519_),
    .X(_11760_));
 sg13g2_nor2_1 _37622_ (.A(net5374),
    .B(_11760_),
    .Y(_11761_));
 sg13g2_a21oi_2 _37623_ (.B1(_11761_),
    .Y(_11762_),
    .A2(_07516_),
    .A1(net5374));
 sg13g2_xnor2_1 _37624_ (.Y(_11763_),
    .A(net4610),
    .B(_11762_));
 sg13g2_nand2_1 _37625_ (.Y(_11764_),
    .A(_11736_),
    .B(_11752_));
 sg13g2_o21ai_1 _37626_ (.B1(_11735_),
    .Y(_11765_),
    .A1(_11737_),
    .A2(_11764_));
 sg13g2_a21o_1 _37627_ (.A2(_11751_),
    .A1(net4610),
    .B1(_11765_),
    .X(_11766_));
 sg13g2_nand2b_1 _37628_ (.Y(_11767_),
    .B(_11725_),
    .A_N(_11704_));
 sg13g2_nor2_1 _37629_ (.A(_11764_),
    .B(_11767_),
    .Y(_11768_));
 sg13g2_nor2b_1 _37630_ (.A(_11711_),
    .B_N(_11768_),
    .Y(_11769_));
 sg13g2_nor2_1 _37631_ (.A(_11766_),
    .B(_11769_),
    .Y(_11770_));
 sg13g2_nor2_1 _37632_ (.A(_11763_),
    .B(_11770_),
    .Y(_11771_));
 sg13g2_and2_1 _37633_ (.A(_11763_),
    .B(_11770_),
    .X(_11772_));
 sg13g2_o21ai_1 _37634_ (.B1(net4713),
    .Y(_11773_),
    .A1(_11771_),
    .A2(_11772_));
 sg13g2_o21ai_1 _37635_ (.B1(_11773_),
    .Y(_11774_),
    .A1(net4713),
    .A2(_11762_));
 sg13g2_o21ai_1 _37636_ (.B1(net5605),
    .Y(_11775_),
    .A1(net4424),
    .A2(_11751_));
 sg13g2_a21oi_1 _37637_ (.A1(net4424),
    .A2(_11774_),
    .Y(_11776_),
    .B1(_11775_));
 sg13g2_a21o_1 _37638_ (.A2(net4212),
    .A1(net2814),
    .B1(_11776_),
    .X(_00913_));
 sg13g2_nand2_1 _37639_ (.Y(_11777_),
    .A(net2739),
    .B(net4215));
 sg13g2_nor2_1 _37640_ (.A(net5414),
    .B(_07492_),
    .Y(_11778_));
 sg13g2_a22oi_1 _37641_ (.Y(_11779_),
    .B1(_07673_),
    .B2(_11749_),
    .A2(_07516_),
    .A1(net4816));
 sg13g2_xnor2_1 _37642_ (.Y(_11780_),
    .A(_07496_),
    .B(_11779_));
 sg13g2_a21oi_2 _37643_ (.B1(_11778_),
    .Y(_11781_),
    .A2(_11780_),
    .A1(net5415));
 sg13g2_nand2_1 _37644_ (.Y(_11782_),
    .A(net4672),
    .B(_11781_));
 sg13g2_nor2_1 _37645_ (.A(net4559),
    .B(_11781_),
    .Y(_11783_));
 sg13g2_nand2_1 _37646_ (.Y(_11784_),
    .A(net4559),
    .B(_11781_));
 sg13g2_nand2b_1 _37647_ (.Y(_11785_),
    .B(_11784_),
    .A_N(_11783_));
 sg13g2_a21oi_1 _37648_ (.A1(net4610),
    .A2(_11762_),
    .Y(_11786_),
    .B1(_11771_));
 sg13g2_xor2_1 _37649_ (.B(_11786_),
    .A(_11785_),
    .X(_11787_));
 sg13g2_o21ai_1 _37650_ (.B1(_11782_),
    .Y(_11788_),
    .A1(net4672),
    .A2(_11787_));
 sg13g2_a21oi_1 _37651_ (.A1(net4424),
    .A2(_11788_),
    .Y(_11789_),
    .B1(net5569));
 sg13g2_o21ai_1 _37652_ (.B1(_11789_),
    .Y(_11790_),
    .A1(net4421),
    .A2(_11762_));
 sg13g2_nand2_1 _37653_ (.Y(_00914_),
    .A(_11777_),
    .B(_11790_));
 sg13g2_a21oi_1 _37654_ (.A1(_07499_),
    .A2(_07503_),
    .Y(_11791_),
    .B1(net5415));
 sg13g2_a21oi_1 _37655_ (.A1(_07495_),
    .A2(_11779_),
    .Y(_11792_),
    .B1(_07494_));
 sg13g2_xor2_1 _37656_ (.B(_11792_),
    .A(_07506_),
    .X(_11793_));
 sg13g2_a21oi_2 _37657_ (.B1(_11791_),
    .Y(_11794_),
    .A2(_11793_),
    .A1(net5414));
 sg13g2_nor2_1 _37658_ (.A(net4713),
    .B(_11794_),
    .Y(_11795_));
 sg13g2_nand2_1 _37659_ (.Y(_11796_),
    .A(net4610),
    .B(_11794_));
 sg13g2_xnor2_1 _37660_ (.Y(_11797_),
    .A(net4610),
    .B(_11794_));
 sg13g2_a21oi_1 _37661_ (.A1(net4611),
    .A2(_11762_),
    .Y(_11798_),
    .B1(_11783_));
 sg13g2_inv_1 _37662_ (.Y(_11799_),
    .A(_11798_));
 sg13g2_o21ai_1 _37663_ (.B1(_11784_),
    .Y(_11800_),
    .A1(_11771_),
    .A2(_11799_));
 sg13g2_xor2_1 _37664_ (.B(_11800_),
    .A(_11797_),
    .X(_11801_));
 sg13g2_nor2_1 _37665_ (.A(net4672),
    .B(_11801_),
    .Y(_11802_));
 sg13g2_o21ai_1 _37666_ (.B1(net4421),
    .Y(_11803_),
    .A1(_11795_),
    .A2(_11802_));
 sg13g2_a21oi_1 _37667_ (.A1(net4366),
    .A2(_11781_),
    .Y(_11804_),
    .B1(net5564));
 sg13g2_a22oi_1 _37668_ (.Y(_11805_),
    .B1(_11803_),
    .B2(_11804_),
    .A2(net4208),
    .A1(net2519));
 sg13g2_inv_1 _37669_ (.Y(_00915_),
    .A(_11805_));
 sg13g2_a21o_2 _37670_ (.A2(_09649_),
    .A1(_09613_),
    .B1(_09655_),
    .X(_11806_));
 sg13g2_a21o_1 _37671_ (.A2(_11806_),
    .A1(_07675_),
    .B1(_07676_),
    .X(_11807_));
 sg13g2_nand3_1 _37672_ (.B(_07676_),
    .C(_11806_),
    .A(_07675_),
    .Y(_11808_));
 sg13g2_nand2_1 _37673_ (.Y(_11809_),
    .A(net5370),
    .B(_07456_));
 sg13g2_nand3_1 _37674_ (.B(_11807_),
    .C(_11808_),
    .A(net5412),
    .Y(_11810_));
 sg13g2_nand2_2 _37675_ (.Y(_11811_),
    .A(_11809_),
    .B(_11810_));
 sg13g2_nand2_1 _37676_ (.Y(_11812_),
    .A(net4610),
    .B(_11811_));
 sg13g2_xnor2_1 _37677_ (.Y(_11813_),
    .A(net4610),
    .B(_11811_));
 sg13g2_o21ai_1 _37678_ (.B1(_11796_),
    .Y(_11814_),
    .A1(_11797_),
    .A2(_11800_));
 sg13g2_a21oi_1 _37679_ (.A1(_11813_),
    .A2(_11814_),
    .Y(_11815_),
    .B1(net4672));
 sg13g2_o21ai_1 _37680_ (.B1(_11815_),
    .Y(_11816_),
    .A1(_11813_),
    .A2(_11814_));
 sg13g2_o21ai_1 _37681_ (.B1(_11816_),
    .Y(_11817_),
    .A1(net4713),
    .A2(_11811_));
 sg13g2_o21ai_1 _37682_ (.B1(net5605),
    .Y(_11818_),
    .A1(net4421),
    .A2(_11794_));
 sg13g2_a21oi_1 _37683_ (.A1(net4422),
    .A2(_11817_),
    .Y(_11819_),
    .B1(_11818_));
 sg13g2_a21o_1 _37684_ (.A2(net4209),
    .A1(net2552),
    .B1(_11819_),
    .X(_00916_));
 sg13g2_nand2_1 _37685_ (.Y(_11820_),
    .A(_07457_),
    .B(_11807_));
 sg13g2_nor2_1 _37686_ (.A(net5412),
    .B(_07465_),
    .Y(_11821_));
 sg13g2_xor2_1 _37687_ (.B(_11820_),
    .A(_07677_),
    .X(_11822_));
 sg13g2_a21oi_2 _37688_ (.B1(_11821_),
    .Y(_11823_),
    .A2(_11822_),
    .A1(net5412));
 sg13g2_nand2_1 _37689_ (.Y(_11824_),
    .A(net4608),
    .B(_11823_));
 sg13g2_xnor2_1 _37690_ (.Y(_11825_),
    .A(net4608),
    .B(_11823_));
 sg13g2_nor4_1 _37691_ (.A(_11763_),
    .B(_11785_),
    .C(_11797_),
    .D(_11813_),
    .Y(_11826_));
 sg13g2_and2_1 _37692_ (.A(_11768_),
    .B(_11826_),
    .X(_11827_));
 sg13g2_or3_1 _37693_ (.A(_11797_),
    .B(_11798_),
    .C(_11813_),
    .X(_11828_));
 sg13g2_nand3_1 _37694_ (.B(_11812_),
    .C(_11828_),
    .A(_11796_),
    .Y(_11829_));
 sg13g2_a21o_1 _37695_ (.A2(_11826_),
    .A1(_11766_),
    .B1(_11829_),
    .X(_11830_));
 sg13g2_a221oi_1 _37696_ (.B2(_11709_),
    .C1(_11829_),
    .B1(_11827_),
    .A1(_11766_),
    .Y(_11831_),
    .A2(_11826_));
 sg13g2_and2_1 _37697_ (.A(_11710_),
    .B(_11827_),
    .X(_11832_));
 sg13g2_a221oi_1 _37698_ (.B2(net1067),
    .C1(_11830_),
    .B1(_11832_),
    .A1(_11709_),
    .Y(_11833_),
    .A2(_11827_));
 sg13g2_xnor2_1 _37699_ (.Y(_11834_),
    .A(_11825_),
    .B(_11833_));
 sg13g2_nand2_1 _37700_ (.Y(_11835_),
    .A(net4710),
    .B(_11834_));
 sg13g2_o21ai_1 _37701_ (.B1(_11835_),
    .Y(_11836_),
    .A1(net4710),
    .A2(_11823_));
 sg13g2_o21ai_1 _37702_ (.B1(net5602),
    .Y(_11837_),
    .A1(net4421),
    .A2(_11811_));
 sg13g2_a21oi_1 _37703_ (.A1(net4421),
    .A2(_11836_),
    .Y(_11838_),
    .B1(_11837_));
 sg13g2_a21o_1 _37704_ (.A2(net4209),
    .A1(net2249),
    .B1(_11838_),
    .X(_00917_));
 sg13g2_nand2_1 _37705_ (.Y(_11839_),
    .A(net5371),
    .B(_07438_));
 sg13g2_a22oi_1 _37706_ (.Y(_11840_),
    .B1(_07467_),
    .B2(_11807_),
    .A2(_07466_),
    .A1(net4815));
 sg13g2_xnor2_1 _37707_ (.Y(_11841_),
    .A(_07440_),
    .B(_11840_));
 sg13g2_o21ai_1 _37708_ (.B1(_11839_),
    .Y(_11842_),
    .A1(net5371),
    .A2(_11841_));
 sg13g2_o21ai_1 _37709_ (.B1(_11824_),
    .Y(_11843_),
    .A1(_11825_),
    .A2(_11833_));
 sg13g2_nand2b_1 _37710_ (.Y(_11844_),
    .B(net4557),
    .A_N(_11842_));
 sg13g2_xnor2_1 _37711_ (.Y(_11845_),
    .A(net4557),
    .B(_11842_));
 sg13g2_xnor2_1 _37712_ (.Y(_11846_),
    .A(_11843_),
    .B(_11845_));
 sg13g2_nand2_1 _37713_ (.Y(_11847_),
    .A(net4711),
    .B(_11846_));
 sg13g2_o21ai_1 _37714_ (.B1(_11847_),
    .Y(_11848_),
    .A1(net4711),
    .A2(_11842_));
 sg13g2_o21ai_1 _37715_ (.B1(net5602),
    .Y(_11849_),
    .A1(net4421),
    .A2(_11823_));
 sg13g2_a21oi_1 _37716_ (.A1(net4421),
    .A2(_11848_),
    .Y(_11850_),
    .B1(_11849_));
 sg13g2_a21o_1 _37717_ (.A2(net4209),
    .A1(net2682),
    .B1(_11850_),
    .X(_00918_));
 sg13g2_nor2_1 _37718_ (.A(net5412),
    .B(_07448_),
    .Y(_11851_));
 sg13g2_a21oi_1 _37719_ (.A1(_07440_),
    .A2(_11840_),
    .Y(_11852_),
    .B1(_07439_));
 sg13g2_xor2_1 _37720_ (.B(_11852_),
    .A(_07449_),
    .X(_11853_));
 sg13g2_a21oi_2 _37721_ (.B1(_11851_),
    .Y(_11854_),
    .A2(_11853_),
    .A1(net5412));
 sg13g2_and2_1 _37722_ (.A(net4608),
    .B(_11854_),
    .X(_11855_));
 sg13g2_xnor2_1 _37723_ (.Y(_11856_),
    .A(net4557),
    .B(_11854_));
 sg13g2_o21ai_1 _37724_ (.B1(net4608),
    .Y(_11857_),
    .A1(_11823_),
    .A2(_11842_));
 sg13g2_inv_1 _37725_ (.Y(_11858_),
    .A(_11857_));
 sg13g2_o21ai_1 _37726_ (.B1(_11857_),
    .Y(_11859_),
    .A1(_11825_),
    .A2(_11833_));
 sg13g2_a21o_1 _37727_ (.A2(_11859_),
    .A1(_11844_),
    .B1(_11856_),
    .X(_11860_));
 sg13g2_nand3_1 _37728_ (.B(_11856_),
    .C(_11859_),
    .A(_11844_),
    .Y(_11861_));
 sg13g2_and2_1 _37729_ (.A(net4710),
    .B(_11861_),
    .X(_11862_));
 sg13g2_a22oi_1 _37730_ (.Y(_11863_),
    .B1(_11860_),
    .B2(_11862_),
    .A2(_11854_),
    .A1(net4674));
 sg13g2_o21ai_1 _37731_ (.B1(net5602),
    .Y(_11864_),
    .A1(net4421),
    .A2(_11842_));
 sg13g2_a21oi_1 _37732_ (.A1(net4422),
    .A2(_11863_),
    .Y(_11865_),
    .B1(_11864_));
 sg13g2_a21o_1 _37733_ (.A2(net4208),
    .A1(net5876),
    .B1(_11865_),
    .X(_00919_));
 sg13g2_nand2_1 _37734_ (.Y(_11866_),
    .A(net5371),
    .B(_07429_));
 sg13g2_a21oi_1 _37735_ (.A1(_07675_),
    .A2(_11806_),
    .Y(_11867_),
    .B1(_07679_));
 sg13g2_nor3_1 _37736_ (.A(_07431_),
    .B(_07469_),
    .C(_11867_),
    .Y(_11868_));
 sg13g2_o21ai_1 _37737_ (.B1(_07431_),
    .Y(_11869_),
    .A1(_07469_),
    .A2(_11867_));
 sg13g2_nand2_1 _37738_ (.Y(_11870_),
    .A(net5411),
    .B(_11869_));
 sg13g2_o21ai_1 _37739_ (.B1(_11866_),
    .Y(_11871_),
    .A1(_11868_),
    .A2(_11870_));
 sg13g2_xnor2_1 _37740_ (.Y(_11872_),
    .A(net4557),
    .B(_11871_));
 sg13g2_nor2b_1 _37741_ (.A(_11855_),
    .B_N(_11861_),
    .Y(_11873_));
 sg13g2_a21oi_1 _37742_ (.A1(_11872_),
    .A2(_11873_),
    .Y(_11874_),
    .B1(net4674));
 sg13g2_o21ai_1 _37743_ (.B1(_11874_),
    .Y(_11875_),
    .A1(_11872_),
    .A2(_11873_));
 sg13g2_o21ai_1 _37744_ (.B1(_11875_),
    .Y(_11876_),
    .A1(net4711),
    .A2(_11871_));
 sg13g2_o21ai_1 _37745_ (.B1(net5602),
    .Y(_11877_),
    .A1(net4422),
    .A2(_11854_));
 sg13g2_a21oi_1 _37746_ (.A1(net4422),
    .A2(_11876_),
    .Y(_11878_),
    .B1(_11877_));
 sg13g2_a21o_1 _37747_ (.A2(net4209),
    .A1(net2756),
    .B1(_11878_),
    .X(_00920_));
 sg13g2_nand2_1 _37748_ (.Y(_11879_),
    .A(net2973),
    .B(net4208));
 sg13g2_and2_1 _37749_ (.A(_11856_),
    .B(_11872_),
    .X(_11880_));
 sg13g2_a221oi_1 _37750_ (.B2(_11858_),
    .C1(_11855_),
    .B1(_11880_),
    .A1(net4608),
    .Y(_11881_),
    .A2(_11871_));
 sg13g2_nand3b_1 _37751_ (.B(_11845_),
    .C(_11880_),
    .Y(_11882_),
    .A_N(_11825_));
 sg13g2_nor2_1 _37752_ (.A(_11833_),
    .B(_11882_),
    .Y(_11883_));
 sg13g2_inv_1 _37753_ (.Y(_11884_),
    .A(_11883_));
 sg13g2_nand3_1 _37754_ (.B(_07430_),
    .C(_11869_),
    .A(_07423_),
    .Y(_11885_));
 sg13g2_a21o_1 _37755_ (.A2(_11869_),
    .A1(_07430_),
    .B1(_07423_),
    .X(_11886_));
 sg13g2_nand3_1 _37756_ (.B(_11885_),
    .C(_11886_),
    .A(net5412),
    .Y(_11887_));
 sg13g2_o21ai_1 _37757_ (.B1(_11887_),
    .Y(_11888_),
    .A1(net5412),
    .A2(_07421_));
 sg13g2_nor2_1 _37758_ (.A(net4557),
    .B(_11888_),
    .Y(_11889_));
 sg13g2_xnor2_1 _37759_ (.Y(_11890_),
    .A(net4557),
    .B(_11888_));
 sg13g2_a21oi_1 _37760_ (.A1(_11881_),
    .A2(_11884_),
    .Y(_11891_),
    .B1(_11890_));
 sg13g2_nand3_1 _37761_ (.B(_11884_),
    .C(_11890_),
    .A(_11881_),
    .Y(_11892_));
 sg13g2_nor2b_1 _37762_ (.A(_11891_),
    .B_N(_11892_),
    .Y(_11893_));
 sg13g2_o21ai_1 _37763_ (.B1(net4420),
    .Y(_11894_),
    .A1(net4711),
    .A2(_11888_));
 sg13g2_a21oi_1 _37764_ (.A1(net4711),
    .A2(_11893_),
    .Y(_11895_),
    .B1(_11894_));
 sg13g2_o21ai_1 _37765_ (.B1(net5602),
    .Y(_11896_),
    .A1(net4422),
    .A2(_11871_));
 sg13g2_o21ai_1 _37766_ (.B1(_11879_),
    .Y(_00921_),
    .A1(_11895_),
    .A2(_11896_));
 sg13g2_nand2_1 _37767_ (.Y(_11897_),
    .A(net5371),
    .B(_07400_));
 sg13g2_a22oi_1 _37768_ (.Y(_11898_),
    .B1(_07471_),
    .B2(_11869_),
    .A2(_07422_),
    .A1(net4815));
 sg13g2_xnor2_1 _37769_ (.Y(_11899_),
    .A(_07403_),
    .B(_11898_));
 sg13g2_o21ai_1 _37770_ (.B1(_11897_),
    .Y(_11900_),
    .A1(net5371),
    .A2(_11899_));
 sg13g2_nor2_1 _37771_ (.A(net4710),
    .B(_11900_),
    .Y(_11901_));
 sg13g2_nor2_1 _37772_ (.A(_11889_),
    .B(_11891_),
    .Y(_11902_));
 sg13g2_nand2b_1 _37773_ (.Y(_11903_),
    .B(net4556),
    .A_N(_11900_));
 sg13g2_xnor2_1 _37774_ (.Y(_11904_),
    .A(net4557),
    .B(_11900_));
 sg13g2_xnor2_1 _37775_ (.Y(_11905_),
    .A(_11902_),
    .B(_11904_));
 sg13g2_nor2_1 _37776_ (.A(net4674),
    .B(_11905_),
    .Y(_11906_));
 sg13g2_o21ai_1 _37777_ (.B1(net4420),
    .Y(_11907_),
    .A1(_11901_),
    .A2(_11906_));
 sg13g2_a21oi_1 _37778_ (.A1(net4365),
    .A2(_11888_),
    .Y(_11908_),
    .B1(net5564));
 sg13g2_a22oi_1 _37779_ (.Y(_11909_),
    .B1(_11907_),
    .B2(_11908_),
    .A2(net4208),
    .A1(net2942));
 sg13g2_inv_1 _37780_ (.Y(_00922_),
    .A(_11909_));
 sg13g2_nand2_1 _37781_ (.Y(_11910_),
    .A(net2932),
    .B(net4208));
 sg13g2_a21oi_1 _37782_ (.A1(_07403_),
    .A2(_11898_),
    .Y(_11911_),
    .B1(_07401_));
 sg13g2_xor2_1 _37783_ (.B(_11911_),
    .A(_07412_),
    .X(_11912_));
 sg13g2_nand2_1 _37784_ (.Y(_11913_),
    .A(net5370),
    .B(_07411_));
 sg13g2_o21ai_1 _37785_ (.B1(_11913_),
    .Y(_11914_),
    .A1(net5370),
    .A2(_11912_));
 sg13g2_nand2_1 _37786_ (.Y(_11915_),
    .A(net4607),
    .B(_11914_));
 sg13g2_xnor2_1 _37787_ (.Y(_11916_),
    .A(net4556),
    .B(_11914_));
 sg13g2_inv_1 _37788_ (.Y(_11917_),
    .A(_11916_));
 sg13g2_a21o_1 _37789_ (.A2(_11900_),
    .A1(net4608),
    .B1(_11889_),
    .X(_11918_));
 sg13g2_o21ai_1 _37790_ (.B1(_11903_),
    .Y(_11919_),
    .A1(_11891_),
    .A2(_11918_));
 sg13g2_or2_1 _37791_ (.X(_11920_),
    .B(_11919_),
    .A(_11917_));
 sg13g2_a21oi_1 _37792_ (.A1(_11917_),
    .A2(_11919_),
    .Y(_11921_),
    .B1(net4670));
 sg13g2_a221oi_1 _37793_ (.B2(_11921_),
    .C1(net4365),
    .B1(_11920_),
    .A1(net4670),
    .Y(_11922_),
    .A2(_11914_));
 sg13g2_o21ai_1 _37794_ (.B1(net5602),
    .Y(_11923_),
    .A1(net4420),
    .A2(_11900_));
 sg13g2_o21ai_1 _37795_ (.B1(_11910_),
    .Y(_00923_),
    .A1(_11922_),
    .A2(_11923_));
 sg13g2_nand2_1 _37796_ (.Y(_11924_),
    .A(net5370),
    .B(_07372_));
 sg13g2_a21oi_1 _37797_ (.A1(_07675_),
    .A2(_11806_),
    .Y(_11925_),
    .B1(_07680_));
 sg13g2_o21ai_1 _37798_ (.B1(_07383_),
    .Y(_11926_),
    .A1(_07475_),
    .A2(_11925_));
 sg13g2_or3_1 _37799_ (.A(_07383_),
    .B(_07475_),
    .C(_11925_),
    .X(_11927_));
 sg13g2_nand3_1 _37800_ (.B(_11926_),
    .C(_11927_),
    .A(net5411),
    .Y(_11928_));
 sg13g2_nand2_2 _37801_ (.Y(_11929_),
    .A(_11924_),
    .B(_11928_));
 sg13g2_nand2_1 _37802_ (.Y(_11930_),
    .A(net4607),
    .B(_11929_));
 sg13g2_xnor2_1 _37803_ (.Y(_11931_),
    .A(net4556),
    .B(_11929_));
 sg13g2_nand2_1 _37804_ (.Y(_11932_),
    .A(_11915_),
    .B(_11920_));
 sg13g2_xnor2_1 _37805_ (.Y(_11933_),
    .A(_11931_),
    .B(_11932_));
 sg13g2_a21oi_1 _37806_ (.A1(net4670),
    .A2(_11929_),
    .Y(_11934_),
    .B1(net4365));
 sg13g2_o21ai_1 _37807_ (.B1(_11934_),
    .Y(_11935_),
    .A1(net4670),
    .A2(_11933_));
 sg13g2_o21ai_1 _37808_ (.B1(net5602),
    .Y(_11936_),
    .A1(net4420),
    .A2(_11914_));
 sg13g2_inv_1 _37809_ (.Y(_11937_),
    .A(_11936_));
 sg13g2_a22oi_1 _37810_ (.Y(_11938_),
    .B1(_11935_),
    .B2(_11937_),
    .A2(net4208),
    .A1(net3003));
 sg13g2_inv_1 _37811_ (.Y(_00924_),
    .A(_11938_));
 sg13g2_nand2_1 _37812_ (.Y(_11939_),
    .A(_07373_),
    .B(_11926_));
 sg13g2_nor2_1 _37813_ (.A(net5411),
    .B(_07366_),
    .Y(_11940_));
 sg13g2_xor2_1 _37814_ (.B(_11939_),
    .A(_07381_),
    .X(_11941_));
 sg13g2_a21oi_2 _37815_ (.B1(_11940_),
    .Y(_11942_),
    .A2(_11941_),
    .A1(net5411));
 sg13g2_and2_1 _37816_ (.A(net4607),
    .B(_11942_),
    .X(_11943_));
 sg13g2_xnor2_1 _37817_ (.Y(_11944_),
    .A(net4556),
    .B(_11942_));
 sg13g2_inv_1 _37818_ (.Y(_11945_),
    .A(_11944_));
 sg13g2_nor2b_1 _37819_ (.A(_11890_),
    .B_N(_11904_),
    .Y(_11946_));
 sg13g2_nand3_1 _37820_ (.B(_11931_),
    .C(_11946_),
    .A(_11916_),
    .Y(_11947_));
 sg13g2_nor2_1 _37821_ (.A(_11881_),
    .B(_11947_),
    .Y(_11948_));
 sg13g2_nand3_1 _37822_ (.B(_11918_),
    .C(_11931_),
    .A(_11916_),
    .Y(_11949_));
 sg13g2_nand3_1 _37823_ (.B(_11930_),
    .C(_11949_),
    .A(_11915_),
    .Y(_11950_));
 sg13g2_nor2_1 _37824_ (.A(_11948_),
    .B(_11950_),
    .Y(_11951_));
 sg13g2_or2_1 _37825_ (.X(_11952_),
    .B(_11947_),
    .A(_11882_));
 sg13g2_o21ai_1 _37826_ (.B1(_11951_),
    .Y(_11953_),
    .A1(_11833_),
    .A2(_11952_));
 sg13g2_and2_1 _37827_ (.A(_11944_),
    .B(_11953_),
    .X(_11954_));
 sg13g2_nor2_1 _37828_ (.A(_11944_),
    .B(_11953_),
    .Y(_11955_));
 sg13g2_o21ai_1 _37829_ (.B1(net4710),
    .Y(_11956_),
    .A1(_11954_),
    .A2(_11955_));
 sg13g2_o21ai_1 _37830_ (.B1(_11956_),
    .Y(_11957_),
    .A1(net4710),
    .A2(_11942_));
 sg13g2_o21ai_1 _37831_ (.B1(net5602),
    .Y(_11958_),
    .A1(net4423),
    .A2(_11929_));
 sg13g2_a21oi_1 _37832_ (.A1(net4423),
    .A2(_11957_),
    .Y(_11959_),
    .B1(_11958_));
 sg13g2_a21o_1 _37833_ (.A2(net4208),
    .A1(net3220),
    .B1(_11959_),
    .X(_00925_));
 sg13g2_nand2_1 _37834_ (.Y(_11960_),
    .A(net2381),
    .B(net4193));
 sg13g2_nand2_1 _37835_ (.Y(_11961_),
    .A(net5368),
    .B(_07345_));
 sg13g2_a22oi_1 _37836_ (.Y(_11962_),
    .B1(_07374_),
    .B2(_11926_),
    .A2(_07367_),
    .A1(net4814));
 sg13g2_xnor2_1 _37837_ (.Y(_11963_),
    .A(_07347_),
    .B(_11962_));
 sg13g2_o21ai_1 _37838_ (.B1(_11961_),
    .Y(_11964_),
    .A1(net5368),
    .A2(_11963_));
 sg13g2_nand2b_1 _37839_ (.Y(_11965_),
    .B(net4555),
    .A_N(_11964_));
 sg13g2_xnor2_1 _37840_ (.Y(_11966_),
    .A(net4603),
    .B(_11964_));
 sg13g2_nor2_1 _37841_ (.A(_11943_),
    .B(_11954_),
    .Y(_11967_));
 sg13g2_xnor2_1 _37842_ (.Y(_11968_),
    .A(_11966_),
    .B(_11967_));
 sg13g2_nand2_1 _37843_ (.Y(_11969_),
    .A(net4706),
    .B(_11968_));
 sg13g2_o21ai_1 _37844_ (.B1(_11969_),
    .Y(_11970_),
    .A1(net4707),
    .A2(_11964_));
 sg13g2_a21oi_1 _37845_ (.A1(net4416),
    .A2(_11970_),
    .Y(_11971_),
    .B1(net5558));
 sg13g2_o21ai_1 _37846_ (.B1(_11971_),
    .Y(_11972_),
    .A1(net4416),
    .A2(_11942_));
 sg13g2_nand2_1 _37847_ (.Y(_00926_),
    .A(_11960_),
    .B(_11972_));
 sg13g2_nand2_1 _37848_ (.Y(_11973_),
    .A(net2433),
    .B(net4193));
 sg13g2_nor2_1 _37849_ (.A(net5410),
    .B(_07355_),
    .Y(_11974_));
 sg13g2_a21oi_1 _37850_ (.A1(_07347_),
    .A2(_11962_),
    .Y(_11975_),
    .B1(_07346_));
 sg13g2_xor2_1 _37851_ (.B(_11975_),
    .A(_07356_),
    .X(_11976_));
 sg13g2_a21oi_2 _37852_ (.B1(_11974_),
    .Y(_11977_),
    .A2(_11976_),
    .A1(net5416));
 sg13g2_nand2_1 _37853_ (.Y(_11978_),
    .A(net4603),
    .B(_11977_));
 sg13g2_xnor2_1 _37854_ (.Y(_11979_),
    .A(net4604),
    .B(_11977_));
 sg13g2_a21o_1 _37855_ (.A2(_11964_),
    .A1(net4604),
    .B1(_11943_),
    .X(_11980_));
 sg13g2_o21ai_1 _37856_ (.B1(_11965_),
    .Y(_11981_),
    .A1(_11954_),
    .A2(_11980_));
 sg13g2_or2_1 _37857_ (.X(_11982_),
    .B(_11981_),
    .A(_11979_));
 sg13g2_a21oi_1 _37858_ (.A1(_11979_),
    .A2(_11981_),
    .Y(_11983_),
    .B1(net4669));
 sg13g2_a221oi_1 _37859_ (.B2(_11983_),
    .C1(net4364),
    .B1(_11982_),
    .A1(net4669),
    .Y(_11984_),
    .A2(_11977_));
 sg13g2_o21ai_1 _37860_ (.B1(net5600),
    .Y(_11985_),
    .A1(net4416),
    .A2(_11964_));
 sg13g2_o21ai_1 _37861_ (.B1(_11973_),
    .Y(_00927_),
    .A1(_11984_),
    .A2(_11985_));
 sg13g2_nand2_1 _37862_ (.Y(_11986_),
    .A(net2406),
    .B(net4193));
 sg13g2_nand2_1 _37863_ (.Y(_11987_),
    .A(_11978_),
    .B(_11982_));
 sg13g2_nand2_1 _37864_ (.Y(_11988_),
    .A(net5370),
    .B(_07336_));
 sg13g2_o21ai_1 _37865_ (.B1(_07384_),
    .Y(_11989_),
    .A1(_07475_),
    .A2(_11925_));
 sg13g2_nor2b_2 _37866_ (.A(_07376_),
    .B_N(_11989_),
    .Y(_11990_));
 sg13g2_nor2b_1 _37867_ (.A(_11990_),
    .B_N(_07338_),
    .Y(_11991_));
 sg13g2_xor2_1 _37868_ (.B(_11990_),
    .A(_07338_),
    .X(_11992_));
 sg13g2_o21ai_1 _37869_ (.B1(_11988_),
    .Y(_11993_),
    .A1(net5370),
    .A2(_11992_));
 sg13g2_xnor2_1 _37870_ (.Y(_11994_),
    .A(net4555),
    .B(_11993_));
 sg13g2_inv_1 _37871_ (.Y(_11995_),
    .A(_11994_));
 sg13g2_xnor2_1 _37872_ (.Y(_11996_),
    .A(_11987_),
    .B(_11995_));
 sg13g2_a21o_1 _37873_ (.A2(_11993_),
    .A1(net4669),
    .B1(net4364),
    .X(_11997_));
 sg13g2_a21oi_1 _37874_ (.A1(net4707),
    .A2(_11996_),
    .Y(_11998_),
    .B1(_11997_));
 sg13g2_o21ai_1 _37875_ (.B1(net5600),
    .Y(_11999_),
    .A1(net4416),
    .A2(_11977_));
 sg13g2_o21ai_1 _37876_ (.B1(_11986_),
    .Y(_00928_),
    .A1(_11998_),
    .A2(_11999_));
 sg13g2_and2_1 _37877_ (.A(net5370),
    .B(_07330_),
    .X(_12000_));
 sg13g2_a21oi_1 _37878_ (.A1(net4760),
    .A2(_07336_),
    .Y(_12001_),
    .B1(_11991_));
 sg13g2_xor2_1 _37879_ (.B(_12001_),
    .A(_07331_),
    .X(_12002_));
 sg13g2_a21oi_2 _37880_ (.B1(_12000_),
    .Y(_12003_),
    .A2(_12002_),
    .A1(net5411));
 sg13g2_and2_1 _37881_ (.A(net4607),
    .B(_12003_),
    .X(_12004_));
 sg13g2_xnor2_1 _37882_ (.Y(_12005_),
    .A(net4556),
    .B(_12003_));
 sg13g2_xnor2_1 _37883_ (.Y(_12006_),
    .A(net4607),
    .B(_12003_));
 sg13g2_nand3b_1 _37884_ (.B(_11980_),
    .C(_11994_),
    .Y(_12007_),
    .A_N(_11979_));
 sg13g2_o21ai_1 _37885_ (.B1(net4604),
    .Y(_12008_),
    .A1(_11977_),
    .A2(_11993_));
 sg13g2_nand2_1 _37886_ (.Y(_12009_),
    .A(_12007_),
    .B(_12008_));
 sg13g2_nor4_1 _37887_ (.A(_11945_),
    .B(_11966_),
    .C(_11979_),
    .D(_11995_),
    .Y(_12010_));
 sg13g2_inv_1 _37888_ (.Y(_12011_),
    .A(_12010_));
 sg13g2_a21oi_1 _37889_ (.A1(_11953_),
    .A2(_12010_),
    .Y(_12012_),
    .B1(_12009_));
 sg13g2_nor2_1 _37890_ (.A(_12006_),
    .B(_12012_),
    .Y(_12013_));
 sg13g2_a21oi_1 _37891_ (.A1(_12006_),
    .A2(_12012_),
    .Y(_12014_),
    .B1(net4670));
 sg13g2_nor2b_1 _37892_ (.A(_12013_),
    .B_N(_12014_),
    .Y(_12015_));
 sg13g2_a21oi_1 _37893_ (.A1(net4670),
    .A2(_12003_),
    .Y(_12016_),
    .B1(_12015_));
 sg13g2_o21ai_1 _37894_ (.B1(net5601),
    .Y(_12017_),
    .A1(net4417),
    .A2(_11993_));
 sg13g2_a21oi_1 _37895_ (.A1(net4417),
    .A2(_12016_),
    .Y(_12018_),
    .B1(_12017_));
 sg13g2_a21o_1 _37896_ (.A2(net4193),
    .A1(net2062),
    .B1(_12018_),
    .X(_00929_));
 sg13g2_nand2_1 _37897_ (.Y(_12019_),
    .A(net2383),
    .B(net4193));
 sg13g2_nor2_1 _37898_ (.A(_12004_),
    .B(_12013_),
    .Y(_12020_));
 sg13g2_o21ai_1 _37899_ (.B1(_07378_),
    .Y(_12021_),
    .A1(_07339_),
    .A2(_11990_));
 sg13g2_o21ai_1 _37900_ (.B1(net5411),
    .Y(_12022_),
    .A1(_07308_),
    .A2(_12021_));
 sg13g2_a21o_1 _37901_ (.A2(_12021_),
    .A1(_07308_),
    .B1(_12022_),
    .X(_12023_));
 sg13g2_o21ai_1 _37902_ (.B1(_12023_),
    .Y(_12024_),
    .A1(net5411),
    .A2(_07304_));
 sg13g2_nand2b_1 _37903_ (.Y(_12025_),
    .B(net4556),
    .A_N(_12024_));
 sg13g2_xnor2_1 _37904_ (.Y(_12026_),
    .A(net4556),
    .B(_12024_));
 sg13g2_a21oi_1 _37905_ (.A1(_12020_),
    .A2(_12026_),
    .Y(_12027_),
    .B1(net4670));
 sg13g2_o21ai_1 _37906_ (.B1(_12027_),
    .Y(_12028_),
    .A1(_12020_),
    .A2(_12026_));
 sg13g2_o21ai_1 _37907_ (.B1(_12028_),
    .Y(_12029_),
    .A1(net4710),
    .A2(_12024_));
 sg13g2_a21oi_1 _37908_ (.A1(net4420),
    .A2(_12029_),
    .Y(_12030_),
    .B1(net5564));
 sg13g2_o21ai_1 _37909_ (.B1(_12030_),
    .Y(_12031_),
    .A1(net4420),
    .A2(_12003_));
 sg13g2_nand2_1 _37910_ (.Y(_00930_),
    .A(_12019_),
    .B(_12031_));
 sg13g2_nand2_1 _37911_ (.Y(_12032_),
    .A(net3029),
    .B(net4208));
 sg13g2_a21oi_1 _37912_ (.A1(_07308_),
    .A2(_12021_),
    .Y(_12033_),
    .B1(_07306_));
 sg13g2_xnor2_1 _37913_ (.Y(_12034_),
    .A(_07320_),
    .B(_12033_));
 sg13g2_and3_1 _37914_ (.X(_12035_),
    .A(net5370),
    .B(_07311_),
    .C(_07316_));
 sg13g2_a21oi_2 _37915_ (.B1(_12035_),
    .Y(_12036_),
    .A2(_12034_),
    .A1(net5411));
 sg13g2_nand2b_1 _37916_ (.Y(_12037_),
    .B(net4607),
    .A_N(_12036_));
 sg13g2_xnor2_1 _37917_ (.Y(_12038_),
    .A(net4607),
    .B(_12036_));
 sg13g2_xnor2_1 _37918_ (.Y(_12039_),
    .A(net4556),
    .B(_12036_));
 sg13g2_a21o_1 _37919_ (.A2(_12024_),
    .A1(net4607),
    .B1(_12004_),
    .X(_12040_));
 sg13g2_o21ai_1 _37920_ (.B1(_12025_),
    .Y(_12041_),
    .A1(_12013_),
    .A2(_12040_));
 sg13g2_or2_1 _37921_ (.X(_12042_),
    .B(_12041_),
    .A(_12039_));
 sg13g2_a21oi_1 _37922_ (.A1(_12039_),
    .A2(_12041_),
    .Y(_12043_),
    .B1(net4670));
 sg13g2_o21ai_1 _37923_ (.B1(net4420),
    .Y(_12044_),
    .A1(net4710),
    .A2(_12036_));
 sg13g2_a21oi_1 _37924_ (.A1(_12042_),
    .A2(_12043_),
    .Y(_12045_),
    .B1(_12044_));
 sg13g2_o21ai_1 _37925_ (.B1(net5603),
    .Y(_12046_),
    .A1(net4420),
    .A2(_12024_));
 sg13g2_o21ai_1 _37926_ (.B1(_12032_),
    .Y(_00931_),
    .A1(_12045_),
    .A2(_12046_));
 sg13g2_nor3_1 _37927_ (.A(_07683_),
    .B(_08041_),
    .C(_09657_),
    .Y(_12047_));
 sg13g2_o21ai_1 _37928_ (.B1(_08041_),
    .Y(_12048_),
    .A1(_07683_),
    .A2(_09657_));
 sg13g2_nand2_1 _37929_ (.Y(_12049_),
    .A(net5367),
    .B(_08039_));
 sg13g2_nand2_1 _37930_ (.Y(_12050_),
    .A(net5413),
    .B(_12048_));
 sg13g2_o21ai_1 _37931_ (.B1(_12049_),
    .Y(_12051_),
    .A1(_12047_),
    .A2(_12050_));
 sg13g2_nand2_1 _37932_ (.Y(_12052_),
    .A(net4605),
    .B(_12051_));
 sg13g2_xnor2_1 _37933_ (.Y(_12053_),
    .A(net4605),
    .B(_12051_));
 sg13g2_inv_2 _37934_ (.Y(_12054_),
    .A(_12053_));
 sg13g2_nand2_1 _37935_ (.Y(_12055_),
    .A(_12037_),
    .B(_12042_));
 sg13g2_xnor2_1 _37936_ (.Y(_12056_),
    .A(_12054_),
    .B(_12055_));
 sg13g2_a21oi_1 _37937_ (.A1(net4671),
    .A2(_12051_),
    .Y(_12057_),
    .B1(net4365));
 sg13g2_o21ai_1 _37938_ (.B1(_12057_),
    .Y(_12058_),
    .A1(net4671),
    .A2(_12056_));
 sg13g2_a21oi_1 _37939_ (.A1(net4365),
    .A2(_12036_),
    .Y(_12059_),
    .B1(net5564));
 sg13g2_a22oi_1 _37940_ (.Y(_12060_),
    .B1(_12058_),
    .B2(_12059_),
    .A2(net4193),
    .A1(net3254));
 sg13g2_inv_1 _37941_ (.Y(_00932_),
    .A(_12060_));
 sg13g2_nand2_1 _37942_ (.Y(_12061_),
    .A(_08040_),
    .B(_12048_));
 sg13g2_and2_1 _37943_ (.A(net5367),
    .B(_08032_),
    .X(_12062_));
 sg13g2_xnor2_1 _37944_ (.Y(_12063_),
    .A(_08034_),
    .B(_12061_));
 sg13g2_a21oi_2 _37945_ (.B1(_12062_),
    .Y(_12064_),
    .A2(_12063_),
    .A1(net5410));
 sg13g2_and2_1 _37946_ (.A(net4603),
    .B(_12064_),
    .X(_12065_));
 sg13g2_xnor2_1 _37947_ (.Y(_12066_),
    .A(net4603),
    .B(_12064_));
 sg13g2_nand4_1 _37948_ (.B(_12026_),
    .C(_12038_),
    .A(_12005_),
    .Y(_12067_),
    .D(_12054_));
 sg13g2_nor3_1 _37949_ (.A(_11952_),
    .B(_12011_),
    .C(_12067_),
    .Y(_12068_));
 sg13g2_and2_1 _37950_ (.A(_11832_),
    .B(_12068_),
    .X(_12069_));
 sg13g2_nor2b_1 _37951_ (.A(_11831_),
    .B_N(_12068_),
    .Y(_12070_));
 sg13g2_nor3_1 _37952_ (.A(_11951_),
    .B(_12011_),
    .C(_12067_),
    .Y(_12071_));
 sg13g2_nand2b_1 _37953_ (.Y(_12072_),
    .B(_12009_),
    .A_N(_12067_));
 sg13g2_nand3_1 _37954_ (.B(_12040_),
    .C(_12054_),
    .A(_12038_),
    .Y(_12073_));
 sg13g2_nand4_1 _37955_ (.B(_12052_),
    .C(_12072_),
    .A(_12037_),
    .Y(_12074_),
    .D(_12073_));
 sg13g2_or3_1 _37956_ (.A(_12070_),
    .B(_12071_),
    .C(_12074_),
    .X(_12075_));
 sg13g2_a21oi_2 _37957_ (.B1(_12075_),
    .Y(_12076_),
    .A2(_12069_),
    .A1(net1067));
 sg13g2_nor2_1 _37958_ (.A(_12066_),
    .B(_12076_),
    .Y(_12077_));
 sg13g2_or2_1 _37959_ (.X(_12078_),
    .B(_12076_),
    .A(_12066_));
 sg13g2_a21oi_1 _37960_ (.A1(_12066_),
    .A2(_12076_),
    .Y(_12079_),
    .B1(net4668));
 sg13g2_a22oi_1 _37961_ (.Y(_12080_),
    .B1(_12078_),
    .B2(_12079_),
    .A2(_12064_),
    .A1(net4671));
 sg13g2_o21ai_1 _37962_ (.B1(net5600),
    .Y(_12081_),
    .A1(net4415),
    .A2(_12051_));
 sg13g2_a21oi_1 _37963_ (.A1(net4415),
    .A2(_12080_),
    .Y(_12082_),
    .B1(_12081_));
 sg13g2_a21o_1 _37964_ (.A2(net4192),
    .A1(net3400),
    .B1(_12082_),
    .X(_00933_));
 sg13g2_nand2_1 _37965_ (.Y(_12083_),
    .A(net2732),
    .B(net4192));
 sg13g2_nor2_1 _37966_ (.A(net5410),
    .B(_08021_),
    .Y(_12084_));
 sg13g2_a22oi_1 _37967_ (.Y(_12085_),
    .B1(_08064_),
    .B2(_12048_),
    .A2(_08032_),
    .A1(net4811));
 sg13g2_xor2_1 _37968_ (.B(_12085_),
    .A(_08023_),
    .X(_12086_));
 sg13g2_a21oi_2 _37969_ (.B1(_12084_),
    .Y(_12087_),
    .A2(_12086_),
    .A1(net5410));
 sg13g2_nor2_1 _37970_ (.A(_12065_),
    .B(_12077_),
    .Y(_12088_));
 sg13g2_nor2_1 _37971_ (.A(net4553),
    .B(_12087_),
    .Y(_12089_));
 sg13g2_nand2_1 _37972_ (.Y(_12090_),
    .A(net4553),
    .B(_12087_));
 sg13g2_nand2b_1 _37973_ (.Y(_12091_),
    .B(_12090_),
    .A_N(_12089_));
 sg13g2_xor2_1 _37974_ (.B(_12091_),
    .A(_12088_),
    .X(_12092_));
 sg13g2_o21ai_1 _37975_ (.B1(net4415),
    .Y(_12093_),
    .A1(net4706),
    .A2(_12087_));
 sg13g2_a21oi_1 _37976_ (.A1(net4706),
    .A2(_12092_),
    .Y(_12094_),
    .B1(_12093_));
 sg13g2_nor2_1 _37977_ (.A(net5558),
    .B(_12094_),
    .Y(_12095_));
 sg13g2_o21ai_1 _37978_ (.B1(_12095_),
    .Y(_12096_),
    .A1(net4415),
    .A2(_12064_));
 sg13g2_nand2_1 _37979_ (.Y(_00934_),
    .A(_12083_),
    .B(_12096_));
 sg13g2_nand2_1 _37980_ (.Y(_12097_),
    .A(net5367),
    .B(_08013_));
 sg13g2_a21oi_1 _37981_ (.A1(_08023_),
    .A2(_12085_),
    .Y(_12098_),
    .B1(_08022_));
 sg13g2_xnor2_1 _37982_ (.Y(_12099_),
    .A(_08014_),
    .B(_12098_));
 sg13g2_o21ai_1 _37983_ (.B1(_12097_),
    .Y(_12100_),
    .A1(net5367),
    .A2(_12099_));
 sg13g2_nand2_1 _37984_ (.Y(_12101_),
    .A(net4668),
    .B(_12100_));
 sg13g2_or2_1 _37985_ (.X(_12102_),
    .B(_12100_),
    .A(net4553));
 sg13g2_xnor2_1 _37986_ (.Y(_12103_),
    .A(net4554),
    .B(_12100_));
 sg13g2_or2_1 _37987_ (.X(_12104_),
    .B(_12089_),
    .A(_12065_));
 sg13g2_o21ai_1 _37988_ (.B1(_12090_),
    .Y(_12105_),
    .A1(_12077_),
    .A2(_12104_));
 sg13g2_xor2_1 _37989_ (.B(_12105_),
    .A(_12103_),
    .X(_12106_));
 sg13g2_o21ai_1 _37990_ (.B1(_12101_),
    .Y(_12107_),
    .A1(net4668),
    .A2(_12106_));
 sg13g2_nand2_1 _37991_ (.Y(_12108_),
    .A(net4416),
    .B(_12107_));
 sg13g2_a21oi_1 _37992_ (.A1(net4363),
    .A2(_12087_),
    .Y(_12109_),
    .B1(net5558));
 sg13g2_a22oi_1 _37993_ (.Y(_12110_),
    .B1(_12108_),
    .B2(_12109_),
    .A2(net4192),
    .A1(net2722));
 sg13g2_inv_1 _37994_ (.Y(_00935_),
    .A(_12110_));
 sg13g2_nand2_1 _37995_ (.Y(_12111_),
    .A(net5367),
    .B(_07988_));
 sg13g2_a21oi_1 _37996_ (.A1(_07682_),
    .A2(_09658_),
    .Y(_12112_),
    .B1(_08042_));
 sg13g2_o21ai_1 _37997_ (.B1(_07990_),
    .Y(_12113_),
    .A1(_08067_),
    .A2(_12112_));
 sg13g2_or3_1 _37998_ (.A(_07990_),
    .B(_08067_),
    .C(_12112_),
    .X(_12114_));
 sg13g2_nand2_1 _37999_ (.Y(_12115_),
    .A(_12113_),
    .B(_12114_));
 sg13g2_o21ai_1 _38000_ (.B1(_12111_),
    .Y(_12116_),
    .A1(net5367),
    .A2(_12115_));
 sg13g2_nand2_1 _38001_ (.Y(_12117_),
    .A(net4603),
    .B(_12116_));
 sg13g2_xnor2_1 _38002_ (.Y(_12118_),
    .A(net4554),
    .B(_12116_));
 sg13g2_o21ai_1 _38003_ (.B1(_12102_),
    .Y(_12119_),
    .A1(_12103_),
    .A2(_12105_));
 sg13g2_xor2_1 _38004_ (.B(_12119_),
    .A(_12118_),
    .X(_12120_));
 sg13g2_nand2_1 _38005_ (.Y(_12121_),
    .A(net4706),
    .B(_12120_));
 sg13g2_a21oi_1 _38006_ (.A1(net4668),
    .A2(_12116_),
    .Y(_12122_),
    .B1(net4363));
 sg13g2_a22oi_1 _38007_ (.Y(_12123_),
    .B1(_12121_),
    .B2(_12122_),
    .A2(_12100_),
    .A1(net4364));
 sg13g2_a22oi_1 _38008_ (.Y(_12124_),
    .B1(_12123_),
    .B2(net5600),
    .A2(net4192),
    .A1(net3082));
 sg13g2_inv_1 _38009_ (.Y(_00936_),
    .A(_12124_));
 sg13g2_nand2_1 _38010_ (.Y(_12125_),
    .A(net2908),
    .B(net4193));
 sg13g2_nand2_1 _38011_ (.Y(_12126_),
    .A(net5367),
    .B(_07998_));
 sg13g2_nor2b_1 _38012_ (.A(_07989_),
    .B_N(_12113_),
    .Y(_12127_));
 sg13g2_xnor2_1 _38013_ (.Y(_12128_),
    .A(_08000_),
    .B(_12127_));
 sg13g2_o21ai_1 _38014_ (.B1(_12126_),
    .Y(_12129_),
    .A1(net5367),
    .A2(_12128_));
 sg13g2_nor2_1 _38015_ (.A(net4553),
    .B(_12129_),
    .Y(_12130_));
 sg13g2_xnor2_1 _38016_ (.Y(_12131_),
    .A(net4603),
    .B(_12129_));
 sg13g2_inv_1 _38017_ (.Y(_12132_),
    .A(_12131_));
 sg13g2_nand3b_1 _38018_ (.B(_12104_),
    .C(_12118_),
    .Y(_12133_),
    .A_N(_12103_));
 sg13g2_nand3_1 _38019_ (.B(_12117_),
    .C(_12133_),
    .A(_12102_),
    .Y(_12134_));
 sg13g2_nor2_1 _38020_ (.A(_12066_),
    .B(_12091_),
    .Y(_12135_));
 sg13g2_nand3b_1 _38021_ (.B(_12118_),
    .C(_12135_),
    .Y(_12136_),
    .A_N(_12103_));
 sg13g2_inv_1 _38022_ (.Y(_12137_),
    .A(_12136_));
 sg13g2_nor2_1 _38023_ (.A(_12076_),
    .B(_12136_),
    .Y(_12138_));
 sg13g2_o21ai_1 _38024_ (.B1(_12131_),
    .Y(_12139_),
    .A1(_12134_),
    .A2(_12138_));
 sg13g2_nor3_1 _38025_ (.A(_12131_),
    .B(_12134_),
    .C(_12138_),
    .Y(_12140_));
 sg13g2_nor2_1 _38026_ (.A(net4668),
    .B(_12140_),
    .Y(_12141_));
 sg13g2_o21ai_1 _38027_ (.B1(net4416),
    .Y(_12142_),
    .A1(net4706),
    .A2(_12129_));
 sg13g2_a21oi_1 _38028_ (.A1(_12139_),
    .A2(_12141_),
    .Y(_12143_),
    .B1(_12142_));
 sg13g2_o21ai_1 _38029_ (.B1(net5600),
    .Y(_12144_),
    .A1(net4416),
    .A2(_12116_));
 sg13g2_o21ai_1 _38030_ (.B1(_12125_),
    .Y(_00937_),
    .A1(_12143_),
    .A2(_12144_));
 sg13g2_nor2_1 _38031_ (.A(net5410),
    .B(_07980_),
    .Y(_12145_));
 sg13g2_a22oi_1 _38032_ (.Y(_12146_),
    .B1(_08063_),
    .B2(_12113_),
    .A2(_07998_),
    .A1(net4811));
 sg13g2_nand2_1 _38033_ (.Y(_12147_),
    .A(_07981_),
    .B(_12146_));
 sg13g2_xor2_1 _38034_ (.B(_12146_),
    .A(_07981_),
    .X(_12148_));
 sg13g2_a21oi_2 _38035_ (.B1(_12145_),
    .Y(_12149_),
    .A2(_12148_),
    .A1(net5410));
 sg13g2_nand2_1 _38036_ (.Y(_12150_),
    .A(net4553),
    .B(_12149_));
 sg13g2_xnor2_1 _38037_ (.Y(_12151_),
    .A(net4553),
    .B(_12149_));
 sg13g2_nor2b_1 _38038_ (.A(_12130_),
    .B_N(_12139_),
    .Y(_12152_));
 sg13g2_a21oi_1 _38039_ (.A1(_12151_),
    .A2(_12152_),
    .Y(_12153_),
    .B1(net4668));
 sg13g2_o21ai_1 _38040_ (.B1(_12153_),
    .Y(_12154_),
    .A1(_12151_),
    .A2(_12152_));
 sg13g2_o21ai_1 _38041_ (.B1(_12154_),
    .Y(_12155_),
    .A1(net4706),
    .A2(_12149_));
 sg13g2_o21ai_1 _38042_ (.B1(net5600),
    .Y(_12156_),
    .A1(net4364),
    .A2(_12155_));
 sg13g2_a21oi_1 _38043_ (.A1(net4364),
    .A2(_12129_),
    .Y(_12157_),
    .B1(_12156_));
 sg13g2_a21o_1 _38044_ (.A2(net4192),
    .A1(net3384),
    .B1(_12157_),
    .X(_00938_));
 sg13g2_a21oi_1 _38045_ (.A1(_07966_),
    .A2(_07972_),
    .Y(_12158_),
    .B1(net5410));
 sg13g2_o21ai_1 _38046_ (.B1(_12147_),
    .Y(_12159_),
    .A1(net4812),
    .A2(_07980_));
 sg13g2_xnor2_1 _38047_ (.Y(_12160_),
    .A(_07974_),
    .B(_12159_));
 sg13g2_a21oi_2 _38048_ (.B1(_12158_),
    .Y(_12161_),
    .A2(_12160_),
    .A1(net5410));
 sg13g2_nor2_1 _38049_ (.A(net4706),
    .B(_12161_),
    .Y(_12162_));
 sg13g2_nand2_1 _38050_ (.Y(_12163_),
    .A(net4603),
    .B(_12161_));
 sg13g2_xnor2_1 _38051_ (.Y(_12164_),
    .A(net4553),
    .B(_12161_));
 sg13g2_a21o_1 _38052_ (.A2(_12149_),
    .A1(_12129_),
    .B1(net4553),
    .X(_12165_));
 sg13g2_nand2_1 _38053_ (.Y(_12166_),
    .A(_12139_),
    .B(_12165_));
 sg13g2_nand3_1 _38054_ (.B(_12164_),
    .C(_12166_),
    .A(_12150_),
    .Y(_12167_));
 sg13g2_a21o_1 _38055_ (.A2(_12166_),
    .A1(_12150_),
    .B1(_12164_),
    .X(_12168_));
 sg13g2_a21oi_1 _38056_ (.A1(_12167_),
    .A2(_12168_),
    .Y(_12169_),
    .B1(net4668));
 sg13g2_o21ai_1 _38057_ (.B1(net4415),
    .Y(_12170_),
    .A1(_12162_),
    .A2(_12169_));
 sg13g2_a21oi_1 _38058_ (.A1(net4364),
    .A2(_12149_),
    .Y(_12171_),
    .B1(net5558));
 sg13g2_a22oi_1 _38059_ (.Y(_12172_),
    .B1(_12170_),
    .B2(_12171_),
    .A2(net4192),
    .A1(net3130));
 sg13g2_inv_1 _38060_ (.Y(_00939_),
    .A(_12172_));
 sg13g2_and2_1 _38061_ (.A(net5366),
    .B(_07956_),
    .X(_12173_));
 sg13g2_a21oi_1 _38062_ (.A1(_07682_),
    .A2(_09658_),
    .Y(_12174_),
    .B1(_08044_));
 sg13g2_o21ai_1 _38063_ (.B1(_07958_),
    .Y(_12175_),
    .A1(_08071_),
    .A2(_12174_));
 sg13g2_nor3_1 _38064_ (.A(_07958_),
    .B(_08071_),
    .C(_12174_),
    .Y(_12176_));
 sg13g2_nor2_1 _38065_ (.A(net5366),
    .B(_12176_),
    .Y(_12177_));
 sg13g2_a21o_2 _38066_ (.A2(_12177_),
    .A1(_12175_),
    .B1(_12173_),
    .X(_12178_));
 sg13g2_nand2_1 _38067_ (.Y(_12179_),
    .A(net4603),
    .B(_12178_));
 sg13g2_xnor2_1 _38068_ (.Y(_12180_),
    .A(net4554),
    .B(_12178_));
 sg13g2_nand2_1 _38069_ (.Y(_12181_),
    .A(_12163_),
    .B(_12167_));
 sg13g2_o21ai_1 _38070_ (.B1(net4706),
    .Y(_12182_),
    .A1(_12180_),
    .A2(_12181_));
 sg13g2_a21oi_1 _38071_ (.A1(_12180_),
    .A2(_12181_),
    .Y(_12183_),
    .B1(_12182_));
 sg13g2_a21oi_1 _38072_ (.A1(net4668),
    .A2(_12178_),
    .Y(_12184_),
    .B1(_12183_));
 sg13g2_o21ai_1 _38073_ (.B1(net5600),
    .Y(_12185_),
    .A1(net4415),
    .A2(_12161_));
 sg13g2_a21oi_1 _38074_ (.A1(net4415),
    .A2(_12184_),
    .Y(_12186_),
    .B1(_12185_));
 sg13g2_a21o_1 _38075_ (.A2(net4192),
    .A1(net2875),
    .B1(_12186_),
    .X(_00940_));
 sg13g2_nand2_1 _38076_ (.Y(_12187_),
    .A(net5366),
    .B(_07949_));
 sg13g2_nand2_1 _38077_ (.Y(_12188_),
    .A(_07957_),
    .B(_12175_));
 sg13g2_xnor2_1 _38078_ (.Y(_12189_),
    .A(_07951_),
    .B(_12188_));
 sg13g2_o21ai_1 _38079_ (.B1(_12187_),
    .Y(_12190_),
    .A1(net5366),
    .A2(_12189_));
 sg13g2_nand2_1 _38080_ (.Y(_12191_),
    .A(net4600),
    .B(_12190_));
 sg13g2_xnor2_1 _38081_ (.Y(_12192_),
    .A(net4550),
    .B(_12190_));
 sg13g2_inv_1 _38082_ (.Y(_12193_),
    .A(_12192_));
 sg13g2_nor2_1 _38083_ (.A(_12132_),
    .B(_12151_),
    .Y(_12194_));
 sg13g2_nand4_1 _38084_ (.B(_12164_),
    .C(_12180_),
    .A(_12134_),
    .Y(_12195_),
    .D(_12194_));
 sg13g2_nand3b_1 _38085_ (.B(_12180_),
    .C(_12164_),
    .Y(_12196_),
    .A_N(_12165_));
 sg13g2_and4_1 _38086_ (.A(_12163_),
    .B(_12179_),
    .C(_12195_),
    .D(_12196_),
    .X(_12197_));
 sg13g2_nand4_1 _38087_ (.B(_12164_),
    .C(_12180_),
    .A(_12137_),
    .Y(_12198_),
    .D(_12194_));
 sg13g2_o21ai_1 _38088_ (.B1(_12197_),
    .Y(_12199_),
    .A1(_12076_),
    .A2(_12198_));
 sg13g2_nand2_1 _38089_ (.Y(_12200_),
    .A(_12192_),
    .B(_12199_));
 sg13g2_nor2_1 _38090_ (.A(_12192_),
    .B(_12199_),
    .Y(_12201_));
 sg13g2_nor2_1 _38091_ (.A(net4665),
    .B(_12201_),
    .Y(_12202_));
 sg13g2_a22oi_1 _38092_ (.Y(_12203_),
    .B1(_12200_),
    .B2(_12202_),
    .A2(_12190_),
    .A1(net4665));
 sg13g2_o21ai_1 _38093_ (.B1(net5601),
    .Y(_12204_),
    .A1(net4410),
    .A2(_12178_));
 sg13g2_a21oi_1 _38094_ (.A1(net4410),
    .A2(_12203_),
    .Y(_12205_),
    .B1(_12204_));
 sg13g2_a21o_1 _38095_ (.A2(net4190),
    .A1(net2936),
    .B1(_12205_),
    .X(_00941_));
 sg13g2_nand2_1 _38096_ (.Y(_12206_),
    .A(net2561),
    .B(net4190));
 sg13g2_nand2_1 _38097_ (.Y(_12207_),
    .A(net5366),
    .B(_07929_));
 sg13g2_a22oi_1 _38098_ (.Y(_12208_),
    .B1(_08073_),
    .B2(_12175_),
    .A2(_07950_),
    .A1(net4808));
 sg13g2_a221oi_1 _38099_ (.B2(_12175_),
    .C1(_07931_),
    .B1(_08073_),
    .A1(net4808),
    .Y(_12209_),
    .A2(_07950_));
 sg13g2_o21ai_1 _38100_ (.B1(net5408),
    .Y(_12210_),
    .A1(_07930_),
    .A2(_12208_));
 sg13g2_o21ai_1 _38101_ (.B1(_12207_),
    .Y(_12211_),
    .A1(_12209_),
    .A2(_12210_));
 sg13g2_nor2_1 _38102_ (.A(net4600),
    .B(_12211_),
    .Y(_12212_));
 sg13g2_xnor2_1 _38103_ (.Y(_12213_),
    .A(net4600),
    .B(_12211_));
 sg13g2_nand2_1 _38104_ (.Y(_12214_),
    .A(_12191_),
    .B(_12200_));
 sg13g2_o21ai_1 _38105_ (.B1(net4704),
    .Y(_12215_),
    .A1(_12213_),
    .A2(_12214_));
 sg13g2_a21o_1 _38106_ (.A2(_12214_),
    .A1(_12213_),
    .B1(_12215_),
    .X(_12216_));
 sg13g2_o21ai_1 _38107_ (.B1(_12216_),
    .Y(_12217_),
    .A1(net4704),
    .A2(_12211_));
 sg13g2_a21oi_1 _38108_ (.A1(net4411),
    .A2(_12217_),
    .Y(_12218_),
    .B1(net5557));
 sg13g2_o21ai_1 _38109_ (.B1(_12218_),
    .Y(_12219_),
    .A1(net4411),
    .A2(_12190_));
 sg13g2_nand2_1 _38110_ (.Y(_00942_),
    .A(_12206_),
    .B(_12219_));
 sg13g2_nor2_1 _38111_ (.A(net5408),
    .B(_07939_),
    .Y(_12220_));
 sg13g2_a21oi_1 _38112_ (.A1(net4757),
    .A2(_07929_),
    .Y(_12221_),
    .B1(_12209_));
 sg13g2_xor2_1 _38113_ (.B(_12221_),
    .A(_07940_),
    .X(_12222_));
 sg13g2_a21oi_2 _38114_ (.B1(_12220_),
    .Y(_12223_),
    .A2(_12222_),
    .A1(net5408));
 sg13g2_nand2_1 _38115_ (.Y(_12224_),
    .A(net4600),
    .B(_12223_));
 sg13g2_xnor2_1 _38116_ (.Y(_12225_),
    .A(net4600),
    .B(_12223_));
 sg13g2_o21ai_1 _38117_ (.B1(net4600),
    .Y(_12226_),
    .A1(_12190_),
    .A2(_12211_));
 sg13g2_a21oi_1 _38118_ (.A1(_12200_),
    .A2(_12226_),
    .Y(_12227_),
    .B1(_12212_));
 sg13g2_inv_1 _38119_ (.Y(_12228_),
    .A(_12227_));
 sg13g2_xor2_1 _38120_ (.B(_12227_),
    .A(_12225_),
    .X(_12229_));
 sg13g2_nand2_1 _38121_ (.Y(_12230_),
    .A(net4705),
    .B(_12229_));
 sg13g2_o21ai_1 _38122_ (.B1(_12230_),
    .Y(_12231_),
    .A1(net4705),
    .A2(_12223_));
 sg13g2_o21ai_1 _38123_ (.B1(net5601),
    .Y(_12232_),
    .A1(net4411),
    .A2(_12211_));
 sg13g2_a21oi_1 _38124_ (.A1(net4411),
    .A2(_12231_),
    .Y(_12233_),
    .B1(_12232_));
 sg13g2_a21o_1 _38125_ (.A2(net4191),
    .A1(net2587),
    .B1(_12233_),
    .X(_00943_));
 sg13g2_nand2_1 _38126_ (.Y(_12234_),
    .A(net2284),
    .B(net4190));
 sg13g2_o21ai_1 _38127_ (.B1(_07959_),
    .Y(_12235_),
    .A1(_08071_),
    .A2(_12174_));
 sg13g2_a21oi_1 _38128_ (.A1(_08076_),
    .A2(_12235_),
    .Y(_12236_),
    .B1(_07913_));
 sg13g2_nand3_1 _38129_ (.B(_08076_),
    .C(_12235_),
    .A(_07913_),
    .Y(_12237_));
 sg13g2_nand3b_1 _38130_ (.B(_12237_),
    .C(net5408),
    .Y(_12238_),
    .A_N(_12236_));
 sg13g2_o21ai_1 _38131_ (.B1(_12238_),
    .Y(_12239_),
    .A1(net5408),
    .A2(_07910_));
 sg13g2_xnor2_1 _38132_ (.Y(_12240_),
    .A(net4600),
    .B(_12239_));
 sg13g2_o21ai_1 _38133_ (.B1(_12224_),
    .Y(_12241_),
    .A1(_12225_),
    .A2(_12228_));
 sg13g2_xor2_1 _38134_ (.B(_12241_),
    .A(_12240_),
    .X(_12242_));
 sg13g2_a21oi_1 _38135_ (.A1(net4666),
    .A2(_12239_),
    .Y(_12243_),
    .B1(net4363));
 sg13g2_o21ai_1 _38136_ (.B1(_12243_),
    .Y(_12244_),
    .A1(net4666),
    .A2(_12242_));
 sg13g2_o21ai_1 _38137_ (.B1(_12244_),
    .Y(_12245_),
    .A1(net4410),
    .A2(_12223_));
 sg13g2_o21ai_1 _38138_ (.B1(_12234_),
    .Y(_00944_),
    .A1(net5557),
    .A2(_12245_));
 sg13g2_nand2_1 _38139_ (.Y(_12246_),
    .A(net1581),
    .B(net4191));
 sg13g2_nor2_1 _38140_ (.A(net5409),
    .B(_07921_),
    .Y(_12247_));
 sg13g2_nor2_1 _38141_ (.A(_07911_),
    .B(_12236_),
    .Y(_12248_));
 sg13g2_xor2_1 _38142_ (.B(_12248_),
    .A(_07922_),
    .X(_12249_));
 sg13g2_a21oi_2 _38143_ (.B1(_12247_),
    .Y(_12250_),
    .A2(_12249_),
    .A1(net5408));
 sg13g2_nand2_1 _38144_ (.Y(_12251_),
    .A(net4601),
    .B(_12250_));
 sg13g2_xnor2_1 _38145_ (.Y(_12252_),
    .A(net4601),
    .B(_12250_));
 sg13g2_or2_1 _38146_ (.X(_12253_),
    .B(_12240_),
    .A(_12225_));
 sg13g2_o21ai_1 _38147_ (.B1(_12224_),
    .Y(_12254_),
    .A1(_12226_),
    .A2(_12253_));
 sg13g2_a21o_1 _38148_ (.A2(_12239_),
    .A1(net4600),
    .B1(_12254_),
    .X(_12255_));
 sg13g2_nor3_1 _38149_ (.A(_12193_),
    .B(_12213_),
    .C(_12253_),
    .Y(_12256_));
 sg13g2_a21oi_1 _38150_ (.A1(_12199_),
    .A2(_12256_),
    .Y(_12257_),
    .B1(_12255_));
 sg13g2_nor2_1 _38151_ (.A(_12252_),
    .B(_12257_),
    .Y(_12258_));
 sg13g2_xnor2_1 _38152_ (.Y(_12259_),
    .A(_12252_),
    .B(_12257_));
 sg13g2_nand2_1 _38153_ (.Y(_12260_),
    .A(net4704),
    .B(_12259_));
 sg13g2_o21ai_1 _38154_ (.B1(_12260_),
    .Y(_12261_),
    .A1(net4704),
    .A2(_12250_));
 sg13g2_a21oi_1 _38155_ (.A1(net4410),
    .A2(_12261_),
    .Y(_12262_),
    .B1(net5557));
 sg13g2_o21ai_1 _38156_ (.B1(_12262_),
    .Y(_12263_),
    .A1(net4411),
    .A2(_12239_));
 sg13g2_nand2_1 _38157_ (.Y(_00945_),
    .A(_12246_),
    .B(_12263_));
 sg13g2_nand2_1 _38158_ (.Y(_12264_),
    .A(net2246),
    .B(net4190));
 sg13g2_o21ai_1 _38159_ (.B1(_12251_),
    .Y(_12265_),
    .A1(_12252_),
    .A2(_12257_));
 sg13g2_nor2_1 _38160_ (.A(net5408),
    .B(_07893_),
    .Y(_12266_));
 sg13g2_a21oi_1 _38161_ (.A1(_07922_),
    .A2(_12236_),
    .Y(_12267_),
    .B1(_08078_));
 sg13g2_xor2_1 _38162_ (.B(_12267_),
    .A(_07895_),
    .X(_12268_));
 sg13g2_a21oi_2 _38163_ (.B1(_12266_),
    .Y(_12269_),
    .A2(_12268_),
    .A1(net5408));
 sg13g2_nand2_1 _38164_ (.Y(_12270_),
    .A(net4550),
    .B(_12269_));
 sg13g2_xnor2_1 _38165_ (.Y(_12271_),
    .A(net4550),
    .B(_12269_));
 sg13g2_xnor2_1 _38166_ (.Y(_12272_),
    .A(_12265_),
    .B(_12271_));
 sg13g2_o21ai_1 _38167_ (.B1(net4410),
    .Y(_12273_),
    .A1(net4704),
    .A2(_12269_));
 sg13g2_a21oi_1 _38168_ (.A1(net4704),
    .A2(_12272_),
    .Y(_12274_),
    .B1(_12273_));
 sg13g2_o21ai_1 _38169_ (.B1(net5601),
    .Y(_12275_),
    .A1(net4410),
    .A2(_12250_));
 sg13g2_o21ai_1 _38170_ (.B1(_12264_),
    .Y(_00946_),
    .A1(_12274_),
    .A2(_12275_));
 sg13g2_nand2_1 _38171_ (.Y(_12276_),
    .A(net5366),
    .B(_07903_));
 sg13g2_o21ai_1 _38172_ (.B1(_07894_),
    .Y(_12277_),
    .A1(_07895_),
    .A2(_12267_));
 sg13g2_xnor2_1 _38173_ (.Y(_12278_),
    .A(_07904_),
    .B(_12277_));
 sg13g2_o21ai_1 _38174_ (.B1(_12276_),
    .Y(_12279_),
    .A1(net5366),
    .A2(_12278_));
 sg13g2_or2_1 _38175_ (.X(_12280_),
    .B(_12279_),
    .A(net4550));
 sg13g2_xnor2_1 _38176_ (.Y(_12281_),
    .A(net4550),
    .B(_12279_));
 sg13g2_o21ai_1 _38177_ (.B1(_12251_),
    .Y(_12282_),
    .A1(net4552),
    .A2(_12269_));
 sg13g2_o21ai_1 _38178_ (.B1(_12270_),
    .Y(_12283_),
    .A1(_12258_),
    .A2(_12282_));
 sg13g2_or2_1 _38179_ (.X(_12284_),
    .B(_12283_),
    .A(_12281_));
 sg13g2_a21oi_1 _38180_ (.A1(_12281_),
    .A2(_12283_),
    .Y(_12285_),
    .B1(net4665));
 sg13g2_nor2_1 _38181_ (.A(net4704),
    .B(_12279_),
    .Y(_12286_));
 sg13g2_a21oi_1 _38182_ (.A1(_12284_),
    .A2(_12285_),
    .Y(_12287_),
    .B1(_12286_));
 sg13g2_nand2_1 _38183_ (.Y(_12288_),
    .A(net4363),
    .B(_12269_));
 sg13g2_a21oi_1 _38184_ (.A1(net4410),
    .A2(_12287_),
    .Y(_12289_),
    .B1(net5557));
 sg13g2_a22oi_1 _38185_ (.Y(_12290_),
    .B1(_12288_),
    .B2(_12289_),
    .A2(net4190),
    .A1(net2538));
 sg13g2_inv_1 _38186_ (.Y(_00947_),
    .A(_12290_));
 sg13g2_a21oi_2 _38187_ (.B1(_08084_),
    .Y(_12291_),
    .A2(_09658_),
    .A1(_07682_));
 sg13g2_nor2_1 _38188_ (.A(_08081_),
    .B(_12291_),
    .Y(_12292_));
 sg13g2_o21ai_1 _38189_ (.B1(_07873_),
    .Y(_12293_),
    .A1(_08081_),
    .A2(_12291_));
 sg13g2_xnor2_1 _38190_ (.Y(_12294_),
    .A(_07873_),
    .B(_12292_));
 sg13g2_mux2_1 _38191_ (.A0(_07870_),
    .A1(_12294_),
    .S(net5409),
    .X(_12295_));
 sg13g2_xnor2_1 _38192_ (.Y(_12296_),
    .A(net4552),
    .B(_12295_));
 sg13g2_inv_1 _38193_ (.Y(_12297_),
    .A(_12296_));
 sg13g2_nand2_1 _38194_ (.Y(_12298_),
    .A(_12280_),
    .B(_12284_));
 sg13g2_xnor2_1 _38195_ (.Y(_12299_),
    .A(_12296_),
    .B(_12298_));
 sg13g2_a21oi_1 _38196_ (.A1(net4665),
    .A2(_12295_),
    .Y(_12300_),
    .B1(net4363));
 sg13g2_o21ai_1 _38197_ (.B1(_12300_),
    .Y(_12301_),
    .A1(net4666),
    .A2(_12299_));
 sg13g2_a21oi_1 _38198_ (.A1(net4363),
    .A2(_12279_),
    .Y(_12302_),
    .B1(net5557));
 sg13g2_a22oi_1 _38199_ (.Y(_12303_),
    .B1(_12301_),
    .B2(_12302_),
    .A2(net4190),
    .A1(net2707));
 sg13g2_inv_1 _38200_ (.Y(_00948_),
    .A(_12303_));
 sg13g2_nand2_1 _38201_ (.Y(_12304_),
    .A(net5365),
    .B(_07863_));
 sg13g2_nand2_1 _38202_ (.Y(_12305_),
    .A(_07871_),
    .B(_12293_));
 sg13g2_xnor2_1 _38203_ (.Y(_12306_),
    .A(_07865_),
    .B(_12305_));
 sg13g2_o21ai_1 _38204_ (.B1(_12304_),
    .Y(_12307_),
    .A1(net5365),
    .A2(_12306_));
 sg13g2_xnor2_1 _38205_ (.Y(_12308_),
    .A(net4551),
    .B(_12307_));
 sg13g2_nor2_1 _38206_ (.A(_12281_),
    .B(_12297_),
    .Y(_12309_));
 sg13g2_nor4_1 _38207_ (.A(_12252_),
    .B(_12271_),
    .C(_12281_),
    .D(_12297_),
    .Y(_12310_));
 sg13g2_nand2_1 _38208_ (.Y(_12311_),
    .A(_12256_),
    .B(_12310_));
 sg13g2_nor2_1 _38209_ (.A(_12197_),
    .B(_12311_),
    .Y(_12312_));
 sg13g2_a22oi_1 _38210_ (.Y(_12313_),
    .B1(_12309_),
    .B2(_12282_),
    .A2(_12295_),
    .A1(net4601));
 sg13g2_nand2_1 _38211_ (.Y(_12314_),
    .A(_12280_),
    .B(_12313_));
 sg13g2_and2_1 _38212_ (.A(_12255_),
    .B(_12310_),
    .X(_12315_));
 sg13g2_nor3_1 _38213_ (.A(_12312_),
    .B(_12314_),
    .C(_12315_),
    .Y(_12316_));
 sg13g2_or3_1 _38214_ (.A(_12312_),
    .B(_12314_),
    .C(_12315_),
    .X(_12317_));
 sg13g2_nor2_2 _38215_ (.A(_12198_),
    .B(_12311_),
    .Y(_12318_));
 sg13g2_inv_1 _38216_ (.Y(_12319_),
    .A(_12318_));
 sg13g2_o21ai_1 _38217_ (.B1(_12316_),
    .Y(_12320_),
    .A1(_12076_),
    .A2(_12319_));
 sg13g2_and2_1 _38218_ (.A(_12308_),
    .B(_12320_),
    .X(_12321_));
 sg13g2_nor2_1 _38219_ (.A(_12308_),
    .B(_12320_),
    .Y(_12322_));
 sg13g2_o21ai_1 _38220_ (.B1(net4705),
    .Y(_12323_),
    .A1(_12321_),
    .A2(_12322_));
 sg13g2_o21ai_1 _38221_ (.B1(_12323_),
    .Y(_12324_),
    .A1(net4705),
    .A2(_12307_));
 sg13g2_o21ai_1 _38222_ (.B1(net5601),
    .Y(_12325_),
    .A1(net4413),
    .A2(_12295_));
 sg13g2_a21oi_1 _38223_ (.A1(net4412),
    .A2(_12324_),
    .Y(_12326_),
    .B1(_12325_));
 sg13g2_a21o_1 _38224_ (.A2(net4191),
    .A1(net1423),
    .B1(_12326_),
    .X(_00949_));
 sg13g2_nand2_1 _38225_ (.Y(_12327_),
    .A(net2140),
    .B(net4191));
 sg13g2_nand2_1 _38226_ (.Y(_12328_),
    .A(net5365),
    .B(_07852_));
 sg13g2_a22oi_1 _38227_ (.Y(_12329_),
    .B1(_08046_),
    .B2(_12293_),
    .A2(_07864_),
    .A1(net4813));
 sg13g2_xnor2_1 _38228_ (.Y(_12330_),
    .A(_07854_),
    .B(_12329_));
 sg13g2_o21ai_1 _38229_ (.B1(_12328_),
    .Y(_12331_),
    .A1(net5368),
    .A2(_12330_));
 sg13g2_nand2b_1 _38230_ (.Y(_12332_),
    .B(net4551),
    .A_N(_12331_));
 sg13g2_xnor2_1 _38231_ (.Y(_12333_),
    .A(net4551),
    .B(_12331_));
 sg13g2_a21oi_1 _38232_ (.A1(net4602),
    .A2(_12307_),
    .Y(_12334_),
    .B1(_12321_));
 sg13g2_a21oi_1 _38233_ (.A1(_12333_),
    .A2(_12334_),
    .Y(_12335_),
    .B1(net4666));
 sg13g2_o21ai_1 _38234_ (.B1(_12335_),
    .Y(_12336_),
    .A1(_12333_),
    .A2(_12334_));
 sg13g2_o21ai_1 _38235_ (.B1(_12336_),
    .Y(_12337_),
    .A1(net4705),
    .A2(_12331_));
 sg13g2_a21oi_1 _38236_ (.A1(net4412),
    .A2(_12337_),
    .Y(_12338_),
    .B1(net5558));
 sg13g2_o21ai_1 _38237_ (.B1(_12338_),
    .Y(_12339_),
    .A1(net4413),
    .A2(_12307_));
 sg13g2_nand2_1 _38238_ (.Y(_00950_),
    .A(_12327_),
    .B(_12339_));
 sg13g2_a21oi_1 _38239_ (.A1(_07854_),
    .A2(_12329_),
    .Y(_12340_),
    .B1(_07853_));
 sg13g2_xnor2_1 _38240_ (.Y(_12341_),
    .A(_07847_),
    .B(_12340_));
 sg13g2_and2_1 _38241_ (.A(net5368),
    .B(_07846_),
    .X(_12342_));
 sg13g2_a21oi_2 _38242_ (.B1(_12342_),
    .Y(_12343_),
    .A2(_12341_),
    .A1(net5409));
 sg13g2_xnor2_1 _38243_ (.Y(_12344_),
    .A(net4602),
    .B(_12343_));
 sg13g2_o21ai_1 _38244_ (.B1(net4602),
    .Y(_12345_),
    .A1(_12307_),
    .A2(_12331_));
 sg13g2_nand2b_1 _38245_ (.Y(_12346_),
    .B(_12345_),
    .A_N(_12321_));
 sg13g2_nand3_1 _38246_ (.B(_12344_),
    .C(_12346_),
    .A(_12332_),
    .Y(_12347_));
 sg13g2_a21o_1 _38247_ (.A2(_12346_),
    .A1(_12332_),
    .B1(_12344_),
    .X(_12348_));
 sg13g2_nand2_1 _38248_ (.Y(_12349_),
    .A(_12347_),
    .B(_12348_));
 sg13g2_mux2_1 _38249_ (.A0(_12343_),
    .A1(_12349_),
    .S(net4705),
    .X(_12350_));
 sg13g2_o21ai_1 _38250_ (.B1(net5601),
    .Y(_12351_),
    .A1(net4413),
    .A2(_12331_));
 sg13g2_a21oi_1 _38251_ (.A1(net4413),
    .A2(_12350_),
    .Y(_12352_),
    .B1(_12351_));
 sg13g2_a21o_1 _38252_ (.A2(net4191),
    .A1(net1982),
    .B1(_12352_),
    .X(_00951_));
 sg13g2_or2_1 _38253_ (.X(_12353_),
    .B(_07833_),
    .A(net5409));
 sg13g2_o21ai_1 _38254_ (.B1(_07874_),
    .Y(_12354_),
    .A1(_08081_),
    .A2(_12291_));
 sg13g2_nand2_1 _38255_ (.Y(_12355_),
    .A(_08049_),
    .B(_12354_));
 sg13g2_xnor2_1 _38256_ (.Y(_12356_),
    .A(_07835_),
    .B(_12355_));
 sg13g2_o21ai_1 _38257_ (.B1(_12353_),
    .Y(_12357_),
    .A1(net5365),
    .A2(_12356_));
 sg13g2_nand2_1 _38258_ (.Y(_12358_),
    .A(net4604),
    .B(_12357_));
 sg13g2_xnor2_1 _38259_ (.Y(_12359_),
    .A(net4552),
    .B(_12357_));
 sg13g2_o21ai_1 _38260_ (.B1(_12347_),
    .Y(_12360_),
    .A1(net4552),
    .A2(_12343_));
 sg13g2_or2_1 _38261_ (.X(_12361_),
    .B(_12360_),
    .A(_12359_));
 sg13g2_a21oi_1 _38262_ (.A1(_12359_),
    .A2(_12360_),
    .Y(_12362_),
    .B1(net4666));
 sg13g2_a22oi_1 _38263_ (.Y(_12363_),
    .B1(_12361_),
    .B2(_12362_),
    .A2(_12357_),
    .A1(net4666));
 sg13g2_nand2_1 _38264_ (.Y(_12364_),
    .A(net4412),
    .B(_12363_));
 sg13g2_a21oi_1 _38265_ (.A1(net4363),
    .A2(_12343_),
    .Y(_12365_),
    .B1(net5558));
 sg13g2_a22oi_1 _38266_ (.Y(_12366_),
    .B1(_12364_),
    .B2(_12365_),
    .A2(net4191),
    .A1(net2418));
 sg13g2_inv_1 _38267_ (.Y(_00952_),
    .A(_12366_));
 sg13g2_nand2_1 _38268_ (.Y(_12367_),
    .A(net1661),
    .B(net4194));
 sg13g2_a21oi_1 _38269_ (.A1(_07835_),
    .A2(_12355_),
    .Y(_12368_),
    .B1(_07834_));
 sg13g2_xnor2_1 _38270_ (.Y(_12369_),
    .A(_07828_),
    .B(_12368_));
 sg13g2_nor2_1 _38271_ (.A(net5365),
    .B(_12369_),
    .Y(_12370_));
 sg13g2_a21oi_2 _38272_ (.B1(_12370_),
    .Y(_12371_),
    .A2(_07823_),
    .A1(net5365));
 sg13g2_and2_1 _38273_ (.A(net4602),
    .B(_12371_),
    .X(_12372_));
 sg13g2_xnor2_1 _38274_ (.Y(_12373_),
    .A(net4602),
    .B(_12371_));
 sg13g2_and2_1 _38275_ (.A(_12344_),
    .B(_12359_),
    .X(_12374_));
 sg13g2_nor2b_1 _38276_ (.A(_12345_),
    .B_N(_12374_),
    .Y(_12375_));
 sg13g2_o21ai_1 _38277_ (.B1(_12358_),
    .Y(_12376_),
    .A1(net4552),
    .A2(_12343_));
 sg13g2_nor2_1 _38278_ (.A(_12375_),
    .B(_12376_),
    .Y(_12377_));
 sg13g2_and3_1 _38279_ (.X(_12378_),
    .A(_12308_),
    .B(_12333_),
    .C(_12374_));
 sg13g2_nand2_1 _38280_ (.Y(_12379_),
    .A(_12320_),
    .B(_12378_));
 sg13g2_a21oi_1 _38281_ (.A1(_12377_),
    .A2(_12379_),
    .Y(_12380_),
    .B1(_12373_));
 sg13g2_nand3_1 _38282_ (.B(_12377_),
    .C(_12379_),
    .A(_12373_),
    .Y(_12381_));
 sg13g2_nand2b_1 _38283_ (.Y(_12382_),
    .B(_12381_),
    .A_N(_12380_));
 sg13g2_nand2_1 _38284_ (.Y(_12383_),
    .A(net4705),
    .B(_12382_));
 sg13g2_o21ai_1 _38285_ (.B1(_12383_),
    .Y(_12384_),
    .A1(net4707),
    .A2(_12371_));
 sg13g2_a21oi_1 _38286_ (.A1(net4412),
    .A2(_12384_),
    .Y(_12385_),
    .B1(net5557));
 sg13g2_o21ai_1 _38287_ (.B1(_12385_),
    .Y(_12386_),
    .A1(net4412),
    .A2(_12357_));
 sg13g2_nand2_1 _38288_ (.Y(_00953_),
    .A(_12367_),
    .B(_12386_));
 sg13g2_nand2_1 _38289_ (.Y(_12387_),
    .A(net2836),
    .B(net4191));
 sg13g2_nor2_1 _38290_ (.A(_12372_),
    .B(_12380_),
    .Y(_12388_));
 sg13g2_a221oi_1 _38291_ (.B2(_12354_),
    .C1(_07836_),
    .B1(_08049_),
    .A1(_07826_),
    .Y(_12389_),
    .A2(_07827_));
 sg13g2_o21ai_1 _38292_ (.B1(_07812_),
    .Y(_12390_),
    .A1(_08051_),
    .A2(_12389_));
 sg13g2_or3_1 _38293_ (.A(_07812_),
    .B(_08051_),
    .C(_12389_),
    .X(_12391_));
 sg13g2_a21oi_1 _38294_ (.A1(_12390_),
    .A2(_12391_),
    .Y(_12392_),
    .B1(net5365));
 sg13g2_a21o_2 _38295_ (.A2(_07810_),
    .A1(net5365),
    .B1(_12392_),
    .X(_12393_));
 sg13g2_nand2_1 _38296_ (.Y(_12394_),
    .A(net4551),
    .B(_12393_));
 sg13g2_nor2_1 _38297_ (.A(net4551),
    .B(_12393_),
    .Y(_12395_));
 sg13g2_xnor2_1 _38298_ (.Y(_12396_),
    .A(net4602),
    .B(_12393_));
 sg13g2_xnor2_1 _38299_ (.Y(_12397_),
    .A(_12388_),
    .B(_12396_));
 sg13g2_nand2_1 _38300_ (.Y(_12398_),
    .A(net4666),
    .B(_12393_));
 sg13g2_o21ai_1 _38301_ (.B1(_12398_),
    .Y(_12399_),
    .A1(net4667),
    .A2(_12397_));
 sg13g2_a21oi_1 _38302_ (.A1(net4412),
    .A2(_12399_),
    .Y(_12400_),
    .B1(net5557));
 sg13g2_o21ai_1 _38303_ (.B1(_12400_),
    .Y(_12401_),
    .A1(net4412),
    .A2(_12371_));
 sg13g2_nand2_1 _38304_ (.Y(_00954_),
    .A(_12387_),
    .B(_12401_));
 sg13g2_nand2_1 _38305_ (.Y(_12402_),
    .A(_07811_),
    .B(_12390_));
 sg13g2_xnor2_1 _38306_ (.Y(_12403_),
    .A(_07804_),
    .B(_12402_));
 sg13g2_mux2_1 _38307_ (.A0(_07801_),
    .A1(_12403_),
    .S(net5409),
    .X(_12404_));
 sg13g2_nor2_1 _38308_ (.A(net4551),
    .B(_12404_),
    .Y(_12405_));
 sg13g2_xnor2_1 _38309_ (.Y(_12406_),
    .A(net4551),
    .B(_12404_));
 sg13g2_or2_1 _38310_ (.X(_12407_),
    .B(_12395_),
    .A(_12372_));
 sg13g2_o21ai_1 _38311_ (.B1(_12394_),
    .Y(_12408_),
    .A1(_12380_),
    .A2(_12407_));
 sg13g2_or2_1 _38312_ (.X(_12409_),
    .B(_12408_),
    .A(_12406_));
 sg13g2_a21oi_1 _38313_ (.A1(_12406_),
    .A2(_12408_),
    .Y(_12410_),
    .B1(net4667));
 sg13g2_o21ai_1 _38314_ (.B1(net4412),
    .Y(_12411_),
    .A1(net4707),
    .A2(_12404_));
 sg13g2_a21oi_1 _38315_ (.A1(_12409_),
    .A2(_12410_),
    .Y(_12412_),
    .B1(_12411_));
 sg13g2_a21oi_1 _38316_ (.A1(net4363),
    .A2(_12393_),
    .Y(_12413_),
    .B1(_12412_));
 sg13g2_a22oi_1 _38317_ (.Y(_12414_),
    .B1(_12413_),
    .B2(net5601),
    .A2(net4190),
    .A1(net2663));
 sg13g2_inv_1 _38318_ (.Y(_00955_),
    .A(_12414_));
 sg13g2_nand2_1 _38319_ (.Y(_12415_),
    .A(net2385),
    .B(net4172));
 sg13g2_nand2_1 _38320_ (.Y(_12416_),
    .A(net5363),
    .B(_07777_));
 sg13g2_o21ai_1 _38321_ (.B1(_07875_),
    .Y(_12417_),
    .A1(_08081_),
    .A2(_12291_));
 sg13g2_a21o_1 _38322_ (.A2(_12417_),
    .A1(_08052_),
    .B1(_07780_),
    .X(_12418_));
 sg13g2_nand3b_1 _38323_ (.B(_08052_),
    .C(_12417_),
    .Y(_12419_),
    .A_N(_07779_));
 sg13g2_nand3_1 _38324_ (.B(_12418_),
    .C(_12419_),
    .A(net5403),
    .Y(_12420_));
 sg13g2_nand2_2 _38325_ (.Y(_12421_),
    .A(_12416_),
    .B(_12420_));
 sg13g2_xnor2_1 _38326_ (.Y(_12422_),
    .A(net4551),
    .B(_12421_));
 sg13g2_xnor2_1 _38327_ (.Y(_12423_),
    .A(net4602),
    .B(_12421_));
 sg13g2_nand2b_1 _38328_ (.Y(_12424_),
    .B(_12409_),
    .A_N(_12405_));
 sg13g2_nand2b_1 _38329_ (.Y(_12425_),
    .B(_12423_),
    .A_N(_12424_));
 sg13g2_a21oi_1 _38330_ (.A1(_12422_),
    .A2(_12424_),
    .Y(_12426_),
    .B1(net4667));
 sg13g2_a221oi_1 _38331_ (.B2(_12426_),
    .C1(net4360),
    .B1(_12425_),
    .A1(net4667),
    .Y(_12427_),
    .A2(_12421_));
 sg13g2_a21o_1 _38332_ (.A2(_12404_),
    .A1(net4360),
    .B1(net5549),
    .X(_12428_));
 sg13g2_o21ai_1 _38333_ (.B1(_12415_),
    .Y(_00956_),
    .A1(_12427_),
    .A2(_12428_));
 sg13g2_nand2_1 _38334_ (.Y(_12429_),
    .A(net2802),
    .B(net4194));
 sg13g2_nor2_1 _38335_ (.A(net5403),
    .B(_07769_),
    .Y(_12430_));
 sg13g2_nand2_1 _38336_ (.Y(_12431_),
    .A(_07778_),
    .B(_12418_));
 sg13g2_xnor2_1 _38337_ (.Y(_12432_),
    .A(_07771_),
    .B(_12431_));
 sg13g2_a21oi_2 _38338_ (.B1(_12430_),
    .Y(_12433_),
    .A2(_12432_),
    .A1(net5404));
 sg13g2_nand2_1 _38339_ (.Y(_12434_),
    .A(net4596),
    .B(_12433_));
 sg13g2_inv_1 _38340_ (.Y(_12435_),
    .A(_12434_));
 sg13g2_xnor2_1 _38341_ (.Y(_12436_),
    .A(net4597),
    .B(_12433_));
 sg13g2_nor2_1 _38342_ (.A(_12406_),
    .B(_12423_),
    .Y(_12437_));
 sg13g2_nor2b_1 _38343_ (.A(_12373_),
    .B_N(_12437_),
    .Y(_12438_));
 sg13g2_nand2_1 _38344_ (.Y(_12439_),
    .A(_12396_),
    .B(_12438_));
 sg13g2_a221oi_1 _38345_ (.B2(_12407_),
    .C1(_12405_),
    .B1(_12437_),
    .A1(net4602),
    .Y(_12440_),
    .A2(_12421_));
 sg13g2_o21ai_1 _38346_ (.B1(_12440_),
    .Y(_12441_),
    .A1(_12377_),
    .A2(_12439_));
 sg13g2_nand3_1 _38347_ (.B(_12396_),
    .C(_12438_),
    .A(_12378_),
    .Y(_12442_));
 sg13g2_inv_1 _38348_ (.Y(_12443_),
    .A(_12442_));
 sg13g2_a21oi_2 _38349_ (.B1(_12441_),
    .Y(_12444_),
    .A2(_12443_),
    .A1(_12320_));
 sg13g2_nor2_1 _38350_ (.A(_12436_),
    .B(_12444_),
    .Y(_12445_));
 sg13g2_xnor2_1 _38351_ (.Y(_12446_),
    .A(_12436_),
    .B(_12444_));
 sg13g2_nand2_1 _38352_ (.Y(_12447_),
    .A(net4702),
    .B(_12446_));
 sg13g2_o21ai_1 _38353_ (.B1(_12447_),
    .Y(_12448_),
    .A1(net4702),
    .A2(_12433_));
 sg13g2_a21oi_1 _38354_ (.A1(net4406),
    .A2(_12448_),
    .Y(_12449_),
    .B1(net5549));
 sg13g2_o21ai_1 _38355_ (.B1(_12449_),
    .Y(_12450_),
    .A1(net4406),
    .A2(_12421_));
 sg13g2_nand2_1 _38356_ (.Y(_00957_),
    .A(_12429_),
    .B(_12450_));
 sg13g2_nand2_1 _38357_ (.Y(_12451_),
    .A(net5363),
    .B(_07749_));
 sg13g2_o21ai_1 _38358_ (.B1(_08055_),
    .Y(_12452_),
    .A1(_07772_),
    .A2(_12418_));
 sg13g2_xnor2_1 _38359_ (.Y(_12453_),
    .A(_07752_),
    .B(_12452_));
 sg13g2_o21ai_1 _38360_ (.B1(_12451_),
    .Y(_12454_),
    .A1(net5363),
    .A2(_12453_));
 sg13g2_nor2_1 _38361_ (.A(_12435_),
    .B(_12445_),
    .Y(_12455_));
 sg13g2_nand2b_1 _38362_ (.Y(_12456_),
    .B(net4547),
    .A_N(_12454_));
 sg13g2_xnor2_1 _38363_ (.Y(_12457_),
    .A(net4547),
    .B(_12454_));
 sg13g2_xor2_1 _38364_ (.B(_12457_),
    .A(_12455_),
    .X(_12458_));
 sg13g2_nor2_1 _38365_ (.A(net4663),
    .B(_12458_),
    .Y(_12459_));
 sg13g2_a21oi_1 _38366_ (.A1(net4662),
    .A2(_12454_),
    .Y(_12460_),
    .B1(_12459_));
 sg13g2_o21ai_1 _38367_ (.B1(net5597),
    .Y(_12461_),
    .A1(net4406),
    .A2(_12433_));
 sg13g2_a21oi_1 _38368_ (.A1(net4406),
    .A2(_12460_),
    .Y(_12462_),
    .B1(_12461_));
 sg13g2_a21o_1 _38369_ (.A2(net4173),
    .A1(net2909),
    .B1(_12462_),
    .X(_00958_));
 sg13g2_nand2_1 _38370_ (.Y(_12463_),
    .A(net1999),
    .B(net4173));
 sg13g2_nor2_1 _38371_ (.A(net5404),
    .B(_07760_),
    .Y(_12464_));
 sg13g2_a21oi_1 _38372_ (.A1(_07752_),
    .A2(_12452_),
    .Y(_12465_),
    .B1(_07751_));
 sg13g2_xor2_1 _38373_ (.B(_12465_),
    .A(_07761_),
    .X(_12466_));
 sg13g2_a21oi_2 _38374_ (.B1(_12464_),
    .Y(_12467_),
    .A2(_12466_),
    .A1(net5404));
 sg13g2_nand2_1 _38375_ (.Y(_12468_),
    .A(net4596),
    .B(_12467_));
 sg13g2_xnor2_1 _38376_ (.Y(_12469_),
    .A(net4596),
    .B(_12467_));
 sg13g2_a21o_1 _38377_ (.A2(_12454_),
    .A1(net4597),
    .B1(_12435_),
    .X(_12470_));
 sg13g2_o21ai_1 _38378_ (.B1(_12456_),
    .Y(_12471_),
    .A1(_12445_),
    .A2(_12470_));
 sg13g2_or2_1 _38379_ (.X(_12472_),
    .B(_12471_),
    .A(_12469_));
 sg13g2_a21oi_1 _38380_ (.A1(_12469_),
    .A2(_12471_),
    .Y(_12473_),
    .B1(net4661));
 sg13g2_a221oi_1 _38381_ (.B2(_12473_),
    .C1(net4360),
    .B1(_12472_),
    .A1(net4661),
    .Y(_12474_),
    .A2(_12467_));
 sg13g2_o21ai_1 _38382_ (.B1(net5597),
    .Y(_12475_),
    .A1(net4407),
    .A2(_12454_));
 sg13g2_o21ai_1 _38383_ (.B1(_12463_),
    .Y(_00959_),
    .A1(_12474_),
    .A2(_12475_));
 sg13g2_nand2_1 _38384_ (.Y(_12476_),
    .A(net2205),
    .B(net4173));
 sg13g2_a21oi_1 _38385_ (.A1(_08052_),
    .A2(_12417_),
    .Y(_12477_),
    .B1(_07781_));
 sg13g2_nor3_1 _38386_ (.A(_07729_),
    .B(_08058_),
    .C(_12477_),
    .Y(_12478_));
 sg13g2_o21ai_1 _38387_ (.B1(_07729_),
    .Y(_12479_),
    .A1(_08058_),
    .A2(_12477_));
 sg13g2_nand2b_1 _38388_ (.Y(_12480_),
    .B(_12479_),
    .A_N(_12478_));
 sg13g2_mux2_1 _38389_ (.A0(_07727_),
    .A1(_12480_),
    .S(net5403),
    .X(_12481_));
 sg13g2_nor2_1 _38390_ (.A(net4547),
    .B(_12481_),
    .Y(_12482_));
 sg13g2_xnor2_1 _38391_ (.Y(_12483_),
    .A(net4547),
    .B(_12481_));
 sg13g2_nand2_1 _38392_ (.Y(_12484_),
    .A(_12468_),
    .B(_12472_));
 sg13g2_xnor2_1 _38393_ (.Y(_12485_),
    .A(_12483_),
    .B(_12484_));
 sg13g2_o21ai_1 _38394_ (.B1(net4407),
    .Y(_12486_),
    .A1(net4701),
    .A2(_12481_));
 sg13g2_a21oi_1 _38395_ (.A1(net4701),
    .A2(_12485_),
    .Y(_12487_),
    .B1(_12486_));
 sg13g2_o21ai_1 _38396_ (.B1(net5598),
    .Y(_12488_),
    .A1(net4407),
    .A2(_12467_));
 sg13g2_o21ai_1 _38397_ (.B1(_12476_),
    .Y(_00960_),
    .A1(_12487_),
    .A2(_12488_));
 sg13g2_nor2_1 _38398_ (.A(net5403),
    .B(_07737_),
    .Y(_12489_));
 sg13g2_nand2_1 _38399_ (.Y(_12490_),
    .A(_07728_),
    .B(_12479_));
 sg13g2_xnor2_1 _38400_ (.Y(_12491_),
    .A(_07739_),
    .B(_12490_));
 sg13g2_a21oi_2 _38401_ (.B1(_12489_),
    .Y(_12492_),
    .A2(_12491_),
    .A1(net5403));
 sg13g2_nand2_1 _38402_ (.Y(_12493_),
    .A(net4596),
    .B(_12492_));
 sg13g2_xnor2_1 _38403_ (.Y(_12494_),
    .A(net4548),
    .B(_12492_));
 sg13g2_nor2_1 _38404_ (.A(_12469_),
    .B(_12483_),
    .Y(_12495_));
 sg13g2_a221oi_1 _38405_ (.B2(_12495_),
    .C1(_12482_),
    .B1(_12470_),
    .A1(net4598),
    .Y(_12496_),
    .A2(_12467_));
 sg13g2_nand3b_1 _38406_ (.B(_12457_),
    .C(_12495_),
    .Y(_12497_),
    .A_N(_12436_));
 sg13g2_o21ai_1 _38407_ (.B1(_12496_),
    .Y(_12498_),
    .A1(_12444_),
    .A2(_12497_));
 sg13g2_nand2_1 _38408_ (.Y(_12499_),
    .A(_12494_),
    .B(_12498_));
 sg13g2_or2_1 _38409_ (.X(_12500_),
    .B(_12498_),
    .A(_12494_));
 sg13g2_a21o_1 _38410_ (.A2(_12500_),
    .A1(_12499_),
    .B1(net4663),
    .X(_12501_));
 sg13g2_o21ai_1 _38411_ (.B1(_12501_),
    .Y(_12502_),
    .A1(net4701),
    .A2(_12492_));
 sg13g2_nand2_1 _38412_ (.Y(_12503_),
    .A(net4360),
    .B(_12481_));
 sg13g2_a21oi_1 _38413_ (.A1(net4406),
    .A2(_12502_),
    .Y(_12504_),
    .B1(net5549));
 sg13g2_a22oi_1 _38414_ (.Y(_12505_),
    .B1(_12503_),
    .B2(_12504_),
    .A2(net4173),
    .A1(net3076));
 sg13g2_inv_1 _38415_ (.Y(_00961_),
    .A(_12505_));
 sg13g2_o21ai_1 _38416_ (.B1(_07741_),
    .Y(_12506_),
    .A1(_08058_),
    .A2(_12477_));
 sg13g2_a21o_1 _38417_ (.A2(_12506_),
    .A1(_08059_),
    .B1(_07712_),
    .X(_12507_));
 sg13g2_nand3_1 _38418_ (.B(_08059_),
    .C(_12506_),
    .A(_07712_),
    .Y(_12508_));
 sg13g2_nand3_1 _38419_ (.B(_12507_),
    .C(_12508_),
    .A(net5403),
    .Y(_12509_));
 sg13g2_o21ai_1 _38420_ (.B1(_12509_),
    .Y(_12510_),
    .A1(net5403),
    .A2(_07710_));
 sg13g2_nor2_1 _38421_ (.A(net4596),
    .B(_12510_),
    .Y(_12511_));
 sg13g2_xnor2_1 _38422_ (.Y(_12512_),
    .A(net4548),
    .B(_12510_));
 sg13g2_nand2_1 _38423_ (.Y(_12513_),
    .A(_12493_),
    .B(_12499_));
 sg13g2_xnor2_1 _38424_ (.Y(_12514_),
    .A(_12512_),
    .B(_12513_));
 sg13g2_a21oi_1 _38425_ (.A1(net4661),
    .A2(_12510_),
    .Y(_12515_),
    .B1(net4361));
 sg13g2_o21ai_1 _38426_ (.B1(_12515_),
    .Y(_12516_),
    .A1(net4661),
    .A2(_12514_));
 sg13g2_o21ai_1 _38427_ (.B1(net5597),
    .Y(_12517_),
    .A1(net4406),
    .A2(_12492_));
 sg13g2_inv_1 _38428_ (.Y(_12518_),
    .A(_12517_));
 sg13g2_a22oi_1 _38429_ (.Y(_12519_),
    .B1(_12516_),
    .B2(_12518_),
    .A2(net4173),
    .A1(net2341));
 sg13g2_inv_1 _38430_ (.Y(_00962_),
    .A(_12519_));
 sg13g2_a21oi_1 _38431_ (.A1(_07711_),
    .A2(_12507_),
    .Y(_12520_),
    .B1(_07722_));
 sg13g2_and3_1 _38432_ (.X(_12521_),
    .A(_07711_),
    .B(_07722_),
    .C(_12507_));
 sg13g2_o21ai_1 _38433_ (.B1(net5403),
    .Y(_12522_),
    .A1(_12520_),
    .A2(_12521_));
 sg13g2_o21ai_1 _38434_ (.B1(_12522_),
    .Y(_12523_),
    .A1(net5405),
    .A2(_07720_));
 sg13g2_nor2_1 _38435_ (.A(net4548),
    .B(_12523_),
    .Y(_12524_));
 sg13g2_xnor2_1 _38436_ (.Y(_12525_),
    .A(net4596),
    .B(_12523_));
 sg13g2_o21ai_1 _38437_ (.B1(net4596),
    .Y(_12526_),
    .A1(_12492_),
    .A2(_12510_));
 sg13g2_a21oi_1 _38438_ (.A1(_12499_),
    .A2(_12526_),
    .Y(_12527_),
    .B1(_12511_));
 sg13g2_xor2_1 _38439_ (.B(_12527_),
    .A(_12525_),
    .X(_12528_));
 sg13g2_nand2_1 _38440_ (.Y(_12529_),
    .A(net4661),
    .B(_12523_));
 sg13g2_o21ai_1 _38441_ (.B1(_12529_),
    .Y(_12530_),
    .A1(net4661),
    .A2(_12528_));
 sg13g2_o21ai_1 _38442_ (.B1(net5597),
    .Y(_12531_),
    .A1(net4406),
    .A2(_12510_));
 sg13g2_a21oi_1 _38443_ (.A1(net4406),
    .A2(_12530_),
    .Y(_12532_),
    .B1(_12531_));
 sg13g2_a21o_1 _38444_ (.A2(net4173),
    .A1(net2021),
    .B1(_12532_),
    .X(_00963_));
 sg13g2_nand2_1 _38445_ (.Y(_12533_),
    .A(net2292),
    .B(net4173));
 sg13g2_a21oi_1 _38446_ (.A1(_12525_),
    .A2(_12527_),
    .Y(_12534_),
    .B1(_12524_));
 sg13g2_nand2_1 _38447_ (.Y(_12535_),
    .A(net5359),
    .B(_07198_));
 sg13g2_xnor2_1 _38448_ (.Y(_12536_),
    .A(_07275_),
    .B(_09659_));
 sg13g2_o21ai_1 _38449_ (.B1(_12535_),
    .Y(_12537_),
    .A1(net5359),
    .A2(_12536_));
 sg13g2_nand2_1 _38450_ (.Y(_12538_),
    .A(net4596),
    .B(_12537_));
 sg13g2_xnor2_1 _38451_ (.Y(_12539_),
    .A(net4548),
    .B(_12537_));
 sg13g2_inv_1 _38452_ (.Y(_12540_),
    .A(_12539_));
 sg13g2_nand2b_1 _38453_ (.Y(_12541_),
    .B(_12539_),
    .A_N(_12534_));
 sg13g2_a21oi_1 _38454_ (.A1(_12534_),
    .A2(_12540_),
    .Y(_12542_),
    .B1(net4661));
 sg13g2_a221oi_1 _38455_ (.B2(_12542_),
    .C1(net4361),
    .B1(_12541_),
    .A1(net4661),
    .Y(_12543_),
    .A2(_12537_));
 sg13g2_a21o_1 _38456_ (.A2(_12523_),
    .A1(net4361),
    .B1(net5556),
    .X(_12544_));
 sg13g2_o21ai_1 _38457_ (.B1(_12533_),
    .Y(_00964_),
    .A1(_12543_),
    .A2(_12544_));
 sg13g2_nand2_1 _38458_ (.Y(_12545_),
    .A(net1343),
    .B(net4171));
 sg13g2_nor2_1 _38459_ (.A(net5402),
    .B(_07192_),
    .Y(_12546_));
 sg13g2_o21ai_1 _38460_ (.B1(_07199_),
    .Y(_12547_),
    .A1(_07275_),
    .A2(_09659_));
 sg13g2_xnor2_1 _38461_ (.Y(_12548_),
    .A(_07273_),
    .B(_12547_));
 sg13g2_a21oi_2 _38462_ (.B1(_12546_),
    .Y(_12549_),
    .A2(_12548_),
    .A1(net5406));
 sg13g2_inv_1 _38463_ (.Y(_12550_),
    .A(_12549_));
 sg13g2_xnor2_1 _38464_ (.Y(_12551_),
    .A(net4594),
    .B(_12549_));
 sg13g2_nand2_1 _38465_ (.Y(_12552_),
    .A(_12525_),
    .B(_12539_));
 sg13g2_nand4_1 _38466_ (.B(_12512_),
    .C(_12525_),
    .A(_12494_),
    .Y(_12553_),
    .D(_12539_));
 sg13g2_nor2_1 _38467_ (.A(_12497_),
    .B(_12553_),
    .Y(_12554_));
 sg13g2_nor2b_2 _38468_ (.A(_12442_),
    .B_N(_12554_),
    .Y(_12555_));
 sg13g2_nor2_1 _38469_ (.A(_12496_),
    .B(_12553_),
    .Y(_12556_));
 sg13g2_o21ai_1 _38470_ (.B1(_12538_),
    .Y(_12557_),
    .A1(_12526_),
    .A2(_12552_));
 sg13g2_or3_1 _38471_ (.A(_12524_),
    .B(_12556_),
    .C(_12557_),
    .X(_12558_));
 sg13g2_a221oi_1 _38472_ (.B2(_12317_),
    .C1(_12558_),
    .B1(_12555_),
    .A1(_12441_),
    .Y(_12559_),
    .A2(_12554_));
 sg13g2_nand3_1 _38473_ (.B(_12318_),
    .C(_12555_),
    .A(_12075_),
    .Y(_12560_));
 sg13g2_nand4_1 _38474_ (.B(_12069_),
    .C(_12318_),
    .A(net1067),
    .Y(_12561_),
    .D(_12555_));
 sg13g2_and3_2 _38475_ (.X(_12562_),
    .A(_12559_),
    .B(_12560_),
    .C(_12561_));
 sg13g2_nand3_1 _38476_ (.B(_12560_),
    .C(_12561_),
    .A(_12559_),
    .Y(_12563_));
 sg13g2_nor2_1 _38477_ (.A(_12551_),
    .B(_12562_),
    .Y(_12564_));
 sg13g2_xnor2_1 _38478_ (.Y(_12565_),
    .A(_12551_),
    .B(_12562_));
 sg13g2_nand2_1 _38479_ (.Y(_12566_),
    .A(net4658),
    .B(_12549_));
 sg13g2_o21ai_1 _38480_ (.B1(_12566_),
    .Y(_12567_),
    .A1(net4658),
    .A2(_12565_));
 sg13g2_nor2_1 _38481_ (.A(net4404),
    .B(_12537_),
    .Y(_12568_));
 sg13g2_o21ai_1 _38482_ (.B1(net5598),
    .Y(_12569_),
    .A1(net4358),
    .A2(_12567_));
 sg13g2_o21ai_1 _38483_ (.B1(_12545_),
    .Y(_00965_),
    .A1(_12568_),
    .A2(_12569_));
 sg13g2_nand2_1 _38484_ (.Y(_12570_),
    .A(net1725),
    .B(net4171));
 sg13g2_nor2_1 _38485_ (.A(net5402),
    .B(_07171_),
    .Y(_12571_));
 sg13g2_o21ai_1 _38486_ (.B1(_07200_),
    .Y(_12572_),
    .A1(_07275_),
    .A2(_09659_));
 sg13g2_nand3_1 _38487_ (.B(_07272_),
    .C(_12572_),
    .A(_07173_),
    .Y(_12573_));
 sg13g2_a21oi_1 _38488_ (.A1(_07272_),
    .A2(_12572_),
    .Y(_12574_),
    .B1(_07173_));
 sg13g2_nor2_1 _38489_ (.A(net5359),
    .B(_12574_),
    .Y(_12575_));
 sg13g2_a21oi_2 _38490_ (.B1(_12571_),
    .Y(_12576_),
    .A2(_12575_),
    .A1(_12573_));
 sg13g2_nand2_1 _38491_ (.Y(_12577_),
    .A(net4659),
    .B(_12576_));
 sg13g2_nand2_1 _38492_ (.Y(_12578_),
    .A(net4546),
    .B(_12576_));
 sg13g2_xnor2_1 _38493_ (.Y(_12579_),
    .A(net4594),
    .B(_12576_));
 sg13g2_a21oi_1 _38494_ (.A1(net4594),
    .A2(_12549_),
    .Y(_12580_),
    .B1(_12564_));
 sg13g2_xnor2_1 _38495_ (.Y(_12581_),
    .A(_12579_),
    .B(_12580_));
 sg13g2_o21ai_1 _38496_ (.B1(_12577_),
    .Y(_12582_),
    .A1(net4659),
    .A2(_12581_));
 sg13g2_a21oi_1 _38497_ (.A1(net4404),
    .A2(_12582_),
    .Y(_12583_),
    .B1(net5547));
 sg13g2_o21ai_1 _38498_ (.B1(_12583_),
    .Y(_12584_),
    .A1(net4404),
    .A2(_12549_));
 sg13g2_nand2_1 _38499_ (.Y(_00966_),
    .A(_12570_),
    .B(_12584_));
 sg13g2_a21o_1 _38500_ (.A2(_12573_),
    .A1(_07172_),
    .B1(_07183_),
    .X(_12585_));
 sg13g2_nand3_1 _38501_ (.B(_07183_),
    .C(_12573_),
    .A(_07172_),
    .Y(_12586_));
 sg13g2_a21oi_1 _38502_ (.A1(_12585_),
    .A2(_12586_),
    .Y(_12587_),
    .B1(net5360));
 sg13g2_and3_1 _38503_ (.X(_12588_),
    .A(net5360),
    .B(_07177_),
    .C(_07180_));
 sg13g2_nor2_1 _38504_ (.A(_12587_),
    .B(_12588_),
    .Y(_12589_));
 sg13g2_o21ai_1 _38505_ (.B1(net4594),
    .Y(_12590_),
    .A1(_12587_),
    .A2(_12588_));
 sg13g2_or3_1 _38506_ (.A(net4598),
    .B(_12587_),
    .C(_12588_),
    .X(_12591_));
 sg13g2_nand2_1 _38507_ (.Y(_12592_),
    .A(_12590_),
    .B(_12591_));
 sg13g2_a21oi_1 _38508_ (.A1(_12550_),
    .A2(_12576_),
    .Y(_12593_),
    .B1(net4546));
 sg13g2_o21ai_1 _38509_ (.B1(_12578_),
    .Y(_12594_),
    .A1(_12564_),
    .A2(_12593_));
 sg13g2_or2_1 _38510_ (.X(_12595_),
    .B(_12594_),
    .A(_12592_));
 sg13g2_a21oi_1 _38511_ (.A1(_12592_),
    .A2(_12594_),
    .Y(_12596_),
    .B1(net4659));
 sg13g2_a21oi_1 _38512_ (.A1(_12595_),
    .A2(_12596_),
    .Y(_12597_),
    .B1(net4359));
 sg13g2_o21ai_1 _38513_ (.B1(_12597_),
    .Y(_12598_),
    .A1(net4700),
    .A2(_12589_));
 sg13g2_a21oi_1 _38514_ (.A1(net4359),
    .A2(_12576_),
    .Y(_12599_),
    .B1(net5548));
 sg13g2_a22oi_1 _38515_ (.Y(_12600_),
    .B1(_12598_),
    .B2(_12599_),
    .A2(net4171),
    .A1(net2462));
 sg13g2_inv_1 _38516_ (.Y(_00967_),
    .A(_12600_));
 sg13g2_nand2_1 _38517_ (.Y(_12601_),
    .A(net5360),
    .B(_07146_));
 sg13g2_a21o_1 _38518_ (.A2(_09660_),
    .A1(_07276_),
    .B1(_07204_),
    .X(_12602_));
 sg13g2_nand2_1 _38519_ (.Y(_12603_),
    .A(_07159_),
    .B(_12602_));
 sg13g2_xnor2_1 _38520_ (.Y(_12604_),
    .A(_07159_),
    .B(_12602_));
 sg13g2_o21ai_1 _38521_ (.B1(_12601_),
    .Y(_12605_),
    .A1(net5360),
    .A2(_12604_));
 sg13g2_and2_1 _38522_ (.A(net4598),
    .B(_12605_),
    .X(_12606_));
 sg13g2_inv_1 _38523_ (.Y(_12607_),
    .A(_12606_));
 sg13g2_xnor2_1 _38524_ (.Y(_12608_),
    .A(net4546),
    .B(_12605_));
 sg13g2_and3_1 _38525_ (.X(_12609_),
    .A(_12590_),
    .B(_12595_),
    .C(_12608_));
 sg13g2_a21oi_1 _38526_ (.A1(_12590_),
    .A2(_12595_),
    .Y(_12610_),
    .B1(_12608_));
 sg13g2_nor2_1 _38527_ (.A(_12609_),
    .B(_12610_),
    .Y(_12611_));
 sg13g2_a21oi_1 _38528_ (.A1(net4659),
    .A2(_12605_),
    .Y(_12612_),
    .B1(net4359));
 sg13g2_o21ai_1 _38529_ (.B1(_12612_),
    .Y(_12613_),
    .A1(net4659),
    .A2(_12611_));
 sg13g2_a21oi_1 _38530_ (.A1(net4359),
    .A2(_12589_),
    .Y(_12614_),
    .B1(net5548));
 sg13g2_a22oi_1 _38531_ (.Y(_12615_),
    .B1(_12613_),
    .B2(_12614_),
    .A2(net4171),
    .A1(net2279));
 sg13g2_inv_1 _38532_ (.Y(_00968_),
    .A(_12615_));
 sg13g2_nand2_1 _38533_ (.Y(_12616_),
    .A(net2305),
    .B(net4171));
 sg13g2_nor2_1 _38534_ (.A(net5402),
    .B(_07156_),
    .Y(_12617_));
 sg13g2_a21oi_1 _38535_ (.A1(_07159_),
    .A2(_12602_),
    .Y(_12618_),
    .B1(_07147_));
 sg13g2_xnor2_1 _38536_ (.Y(_12619_),
    .A(_07161_),
    .B(_12618_));
 sg13g2_a21oi_2 _38537_ (.B1(_12617_),
    .Y(_12620_),
    .A2(_12619_),
    .A1(net5402));
 sg13g2_nand2_1 _38538_ (.Y(_12621_),
    .A(net4658),
    .B(_12620_));
 sg13g2_nor2_1 _38539_ (.A(net4546),
    .B(_12620_),
    .Y(_12622_));
 sg13g2_xnor2_1 _38540_ (.Y(_12623_),
    .A(net4594),
    .B(_12620_));
 sg13g2_nand4_1 _38541_ (.B(_12591_),
    .C(_12593_),
    .A(_12590_),
    .Y(_12624_),
    .D(_12608_));
 sg13g2_and3_1 _38542_ (.X(_12625_),
    .A(_12590_),
    .B(_12607_),
    .C(_12624_));
 sg13g2_nand3_1 _38543_ (.B(_12607_),
    .C(_12624_),
    .A(_12590_),
    .Y(_12626_));
 sg13g2_nor2b_1 _38544_ (.A(_12551_),
    .B_N(_12579_),
    .Y(_12627_));
 sg13g2_nand4_1 _38545_ (.B(_12591_),
    .C(_12608_),
    .A(_12590_),
    .Y(_12628_),
    .D(_12627_));
 sg13g2_o21ai_1 _38546_ (.B1(_12625_),
    .Y(_12629_),
    .A1(_12562_),
    .A2(_12628_));
 sg13g2_xor2_1 _38547_ (.B(_12629_),
    .A(_12623_),
    .X(_12630_));
 sg13g2_o21ai_1 _38548_ (.B1(_12621_),
    .Y(_12631_),
    .A1(net4658),
    .A2(_12630_));
 sg13g2_a21oi_1 _38549_ (.A1(net4408),
    .A2(_12631_),
    .Y(_12632_),
    .B1(net5548));
 sg13g2_o21ai_1 _38550_ (.B1(_12632_),
    .Y(_12633_),
    .A1(net4404),
    .A2(_12605_));
 sg13g2_nand2_1 _38551_ (.Y(_00969_),
    .A(_12616_),
    .B(_12633_));
 sg13g2_nand2_1 _38552_ (.Y(_12634_),
    .A(net2238),
    .B(net4171));
 sg13g2_nor2_1 _38553_ (.A(net5402),
    .B(_07125_),
    .Y(_12635_));
 sg13g2_a22oi_1 _38554_ (.Y(_12636_),
    .B1(_07158_),
    .B2(_12603_),
    .A2(_07156_),
    .A1(net4804));
 sg13g2_xnor2_1 _38555_ (.Y(_12637_),
    .A(_07128_),
    .B(_12636_));
 sg13g2_a21oi_2 _38556_ (.B1(_12635_),
    .Y(_12638_),
    .A2(_12637_),
    .A1(net5406));
 sg13g2_xnor2_1 _38557_ (.Y(_12639_),
    .A(net4594),
    .B(_12638_));
 sg13g2_a21oi_1 _38558_ (.A1(_12623_),
    .A2(_12629_),
    .Y(_12640_),
    .B1(_12622_));
 sg13g2_xnor2_1 _38559_ (.Y(_12641_),
    .A(_12639_),
    .B(_12640_));
 sg13g2_nand2_1 _38560_ (.Y(_12642_),
    .A(net4658),
    .B(_12638_));
 sg13g2_o21ai_1 _38561_ (.B1(_12642_),
    .Y(_12643_),
    .A1(net4658),
    .A2(_12641_));
 sg13g2_mux2_1 _38562_ (.A0(_12620_),
    .A1(_12643_),
    .S(net4404),
    .X(_12644_));
 sg13g2_o21ai_1 _38563_ (.B1(_12634_),
    .Y(_00970_),
    .A1(net5548),
    .A2(_12644_));
 sg13g2_nand2_1 _38564_ (.Y(_12645_),
    .A(net5356),
    .B(_07137_));
 sg13g2_a21oi_1 _38565_ (.A1(_07127_),
    .A2(_12636_),
    .Y(_12646_),
    .B1(_07126_));
 sg13g2_xnor2_1 _38566_ (.Y(_12647_),
    .A(_07138_),
    .B(_12646_));
 sg13g2_o21ai_1 _38567_ (.B1(_12645_),
    .Y(_12648_),
    .A1(net5356),
    .A2(_12647_));
 sg13g2_nor2_1 _38568_ (.A(net4546),
    .B(_12648_),
    .Y(_12649_));
 sg13g2_xnor2_1 _38569_ (.Y(_12650_),
    .A(net4594),
    .B(_12648_));
 sg13g2_a21oi_1 _38570_ (.A1(_12620_),
    .A2(_12638_),
    .Y(_12651_),
    .B1(net4546));
 sg13g2_a21oi_1 _38571_ (.A1(_12623_),
    .A2(_12629_),
    .Y(_12652_),
    .B1(_12651_));
 sg13g2_a21oi_1 _38572_ (.A1(net4546),
    .A2(_12638_),
    .Y(_12653_),
    .B1(_12652_));
 sg13g2_and2_1 _38573_ (.A(_12650_),
    .B(_12653_),
    .X(_12654_));
 sg13g2_o21ai_1 _38574_ (.B1(net4700),
    .Y(_12655_),
    .A1(_12650_),
    .A2(_12653_));
 sg13g2_nor2_1 _38575_ (.A(net4702),
    .B(_12648_),
    .Y(_12656_));
 sg13g2_nor2_1 _38576_ (.A(net4358),
    .B(_12656_),
    .Y(_12657_));
 sg13g2_o21ai_1 _38577_ (.B1(_12657_),
    .Y(_12658_),
    .A1(_12654_),
    .A2(_12655_));
 sg13g2_a21oi_1 _38578_ (.A1(net4359),
    .A2(_12638_),
    .Y(_12659_),
    .B1(net5547));
 sg13g2_a22oi_1 _38579_ (.Y(_12660_),
    .B1(_12658_),
    .B2(_12659_),
    .A2(net4170),
    .A1(net2257));
 sg13g2_inv_1 _38580_ (.Y(_00971_),
    .A(_12660_));
 sg13g2_nand2_1 _38581_ (.Y(_12661_),
    .A(net2278),
    .B(net4155));
 sg13g2_nand2_1 _38582_ (.Y(_12662_),
    .A(net5358),
    .B(_07109_));
 sg13g2_o21ai_1 _38583_ (.B1(_07209_),
    .Y(_12663_),
    .A1(_07278_),
    .A2(_09659_));
 sg13g2_nand2b_1 _38584_ (.Y(_12664_),
    .B(_12663_),
    .A_N(_07111_));
 sg13g2_xor2_1 _38585_ (.B(_12663_),
    .A(_07111_),
    .X(_12665_));
 sg13g2_o21ai_1 _38586_ (.B1(_12662_),
    .Y(_12666_),
    .A1(net5358),
    .A2(_12665_));
 sg13g2_xnor2_1 _38587_ (.Y(_12667_),
    .A(net4546),
    .B(_12666_));
 sg13g2_nor2_1 _38588_ (.A(_12649_),
    .B(_12654_),
    .Y(_12668_));
 sg13g2_nor3_1 _38589_ (.A(_12649_),
    .B(_12654_),
    .C(_12667_),
    .Y(_12669_));
 sg13g2_nor2b_1 _38590_ (.A(_12668_),
    .B_N(_12667_),
    .Y(_12670_));
 sg13g2_nor3_1 _38591_ (.A(net4658),
    .B(_12669_),
    .C(_12670_),
    .Y(_12671_));
 sg13g2_and2_1 _38592_ (.A(net4658),
    .B(_12666_),
    .X(_12672_));
 sg13g2_nor3_1 _38593_ (.A(net4357),
    .B(_12671_),
    .C(_12672_),
    .Y(_12673_));
 sg13g2_a21o_1 _38594_ (.A2(_12648_),
    .A1(net4357),
    .B1(net5548),
    .X(_12674_));
 sg13g2_o21ai_1 _38595_ (.B1(_12661_),
    .Y(_00972_),
    .A1(_12673_),
    .A2(_12674_));
 sg13g2_nand2_1 _38596_ (.Y(_12675_),
    .A(net2938),
    .B(net4154));
 sg13g2_nor2_1 _38597_ (.A(net5398),
    .B(_07102_),
    .Y(_12676_));
 sg13g2_nand2_1 _38598_ (.Y(_12677_),
    .A(_07110_),
    .B(_12664_));
 sg13g2_xor2_1 _38599_ (.B(_12677_),
    .A(_07104_),
    .X(_12678_));
 sg13g2_a21oi_2 _38600_ (.B1(_12676_),
    .Y(_12679_),
    .A2(_12678_),
    .A1(net5399));
 sg13g2_xnor2_1 _38601_ (.Y(_12680_),
    .A(net4591),
    .B(_12679_));
 sg13g2_and2_1 _38602_ (.A(_12623_),
    .B(_12639_),
    .X(_12681_));
 sg13g2_nand3_1 _38603_ (.B(_12667_),
    .C(_12681_),
    .A(_12650_),
    .Y(_12682_));
 sg13g2_nand4_1 _38604_ (.B(_12650_),
    .C(_12667_),
    .A(_12626_),
    .Y(_12683_),
    .D(_12681_));
 sg13g2_nand3_1 _38605_ (.B(_12651_),
    .C(_12667_),
    .A(_12650_),
    .Y(_12684_));
 sg13g2_a21oi_1 _38606_ (.A1(net4594),
    .A2(_12666_),
    .Y(_12685_),
    .B1(_12649_));
 sg13g2_nand3_1 _38607_ (.B(_12684_),
    .C(_12685_),
    .A(_12683_),
    .Y(_12686_));
 sg13g2_nor2_1 _38608_ (.A(_12628_),
    .B(_12682_),
    .Y(_12687_));
 sg13g2_a21oi_1 _38609_ (.A1(_12563_),
    .A2(_12687_),
    .Y(_12688_),
    .B1(_12686_));
 sg13g2_nor2_1 _38610_ (.A(_12680_),
    .B(_12688_),
    .Y(_12689_));
 sg13g2_inv_1 _38611_ (.Y(_12690_),
    .A(_12689_));
 sg13g2_nand2_1 _38612_ (.Y(_12691_),
    .A(_12680_),
    .B(_12688_));
 sg13g2_a21o_1 _38613_ (.A2(_12691_),
    .A1(_12690_),
    .B1(net4656),
    .X(_12692_));
 sg13g2_o21ai_1 _38614_ (.B1(_12692_),
    .Y(_12693_),
    .A1(net4698),
    .A2(_12679_));
 sg13g2_a21oi_1 _38615_ (.A1(net4402),
    .A2(_12693_),
    .Y(_12694_),
    .B1(net5538));
 sg13g2_o21ai_1 _38616_ (.B1(_12694_),
    .Y(_12695_),
    .A1(net4402),
    .A2(_12666_));
 sg13g2_nand2_1 _38617_ (.Y(_00973_),
    .A(_12675_),
    .B(_12695_));
 sg13g2_nand2_1 _38618_ (.Y(_12696_),
    .A(net2396),
    .B(net4154));
 sg13g2_nand2_1 _38619_ (.Y(_12697_),
    .A(net5356),
    .B(_07081_));
 sg13g2_a22oi_1 _38620_ (.Y(_12698_),
    .B1(_07215_),
    .B2(_12664_),
    .A2(_07103_),
    .A1(net4802));
 sg13g2_xnor2_1 _38621_ (.Y(_12699_),
    .A(_07083_),
    .B(_12698_));
 sg13g2_o21ai_1 _38622_ (.B1(_12697_),
    .Y(_12700_),
    .A1(net5356),
    .A2(_12699_));
 sg13g2_nor2_1 _38623_ (.A(net4591),
    .B(_12700_),
    .Y(_12701_));
 sg13g2_xnor2_1 _38624_ (.Y(_12702_),
    .A(net4544),
    .B(_12700_));
 sg13g2_a21o_1 _38625_ (.A2(_12679_),
    .A1(net4591),
    .B1(_12689_),
    .X(_12703_));
 sg13g2_xor2_1 _38626_ (.B(_12703_),
    .A(_12702_),
    .X(_12704_));
 sg13g2_nor2_1 _38627_ (.A(net4656),
    .B(_12704_),
    .Y(_12705_));
 sg13g2_nor2_1 _38628_ (.A(net4698),
    .B(_12700_),
    .Y(_12706_));
 sg13g2_o21ai_1 _38629_ (.B1(net4402),
    .Y(_12707_),
    .A1(_12705_),
    .A2(_12706_));
 sg13g2_o21ai_1 _38630_ (.B1(_12707_),
    .Y(_12708_),
    .A1(net4400),
    .A2(_12679_));
 sg13g2_o21ai_1 _38631_ (.B1(_12696_),
    .Y(_00974_),
    .A1(net5538),
    .A2(_12708_));
 sg13g2_nor2_1 _38632_ (.A(net5399),
    .B(_07091_),
    .Y(_12709_));
 sg13g2_a21oi_1 _38633_ (.A1(_07083_),
    .A2(_12698_),
    .Y(_12710_),
    .B1(_07082_));
 sg13g2_xor2_1 _38634_ (.B(_12710_),
    .A(_07092_),
    .X(_12711_));
 sg13g2_a21oi_2 _38635_ (.B1(_12709_),
    .Y(_12712_),
    .A2(_12711_),
    .A1(net5399));
 sg13g2_nand2_1 _38636_ (.Y(_12713_),
    .A(net4591),
    .B(_12712_));
 sg13g2_xnor2_1 _38637_ (.Y(_12714_),
    .A(net4543),
    .B(_12712_));
 sg13g2_o21ai_1 _38638_ (.B1(net4593),
    .Y(_12715_),
    .A1(_12679_),
    .A2(_12700_));
 sg13g2_a21oi_1 _38639_ (.A1(_12690_),
    .A2(_12715_),
    .Y(_12716_),
    .B1(_12701_));
 sg13g2_nand2_1 _38640_ (.Y(_12717_),
    .A(_12714_),
    .B(_12716_));
 sg13g2_xnor2_1 _38641_ (.Y(_12718_),
    .A(_12714_),
    .B(_12716_));
 sg13g2_nand2_1 _38642_ (.Y(_12719_),
    .A(net4698),
    .B(_12718_));
 sg13g2_o21ai_1 _38643_ (.B1(_12719_),
    .Y(_12720_),
    .A1(net4698),
    .A2(_12712_));
 sg13g2_o21ai_1 _38644_ (.B1(net5596),
    .Y(_12721_),
    .A1(net4400),
    .A2(_12700_));
 sg13g2_a21oi_1 _38645_ (.A1(net4400),
    .A2(_12720_),
    .Y(_12722_),
    .B1(_12721_));
 sg13g2_a21o_1 _38646_ (.A2(net4155),
    .A1(net1711),
    .B1(_12722_),
    .X(_00975_));
 sg13g2_nand2_1 _38647_ (.Y(_12723_),
    .A(net2148),
    .B(net4155));
 sg13g2_nor2_1 _38648_ (.A(net5399),
    .B(_07062_),
    .Y(_12724_));
 sg13g2_a21oi_1 _38649_ (.A1(_07112_),
    .A2(_12663_),
    .Y(_12725_),
    .B1(_07217_));
 sg13g2_or2_1 _38650_ (.X(_12726_),
    .B(_12725_),
    .A(_07064_));
 sg13g2_a21oi_1 _38651_ (.A1(_07064_),
    .A2(_12725_),
    .Y(_12727_),
    .B1(net5356));
 sg13g2_a21oi_2 _38652_ (.B1(_12724_),
    .Y(_12728_),
    .A2(_12727_),
    .A1(_12726_));
 sg13g2_xnor2_1 _38653_ (.Y(_12729_),
    .A(net4591),
    .B(_12728_));
 sg13g2_nand2_1 _38654_ (.Y(_12730_),
    .A(_12713_),
    .B(_12717_));
 sg13g2_xor2_1 _38655_ (.B(_12730_),
    .A(_12729_),
    .X(_12731_));
 sg13g2_o21ai_1 _38656_ (.B1(net4400),
    .Y(_12732_),
    .A1(net4699),
    .A2(_12728_));
 sg13g2_a21oi_1 _38657_ (.A1(net4699),
    .A2(_12731_),
    .Y(_12733_),
    .B1(_12732_));
 sg13g2_o21ai_1 _38658_ (.B1(net5596),
    .Y(_12734_),
    .A1(net4400),
    .A2(_12712_));
 sg13g2_o21ai_1 _38659_ (.B1(_12723_),
    .Y(_00976_),
    .A1(_12733_),
    .A2(_12734_));
 sg13g2_a21oi_1 _38660_ (.A1(_07063_),
    .A2(_12726_),
    .Y(_12735_),
    .B1(_07073_));
 sg13g2_and3_1 _38661_ (.X(_12736_),
    .A(_07063_),
    .B(_07073_),
    .C(_12726_));
 sg13g2_nor3_1 _38662_ (.A(net5356),
    .B(_12735_),
    .C(_12736_),
    .Y(_12737_));
 sg13g2_a21oi_2 _38663_ (.B1(_12737_),
    .Y(_12738_),
    .A2(_07072_),
    .A1(net5356));
 sg13g2_nand2_1 _38664_ (.Y(_12739_),
    .A(net4656),
    .B(_12738_));
 sg13g2_nand2_1 _38665_ (.Y(_12740_),
    .A(net4591),
    .B(_12738_));
 sg13g2_xnor2_1 _38666_ (.Y(_12741_),
    .A(net4543),
    .B(_12738_));
 sg13g2_nand2_1 _38667_ (.Y(_12742_),
    .A(_12714_),
    .B(_12729_));
 sg13g2_nor2_1 _38668_ (.A(_12715_),
    .B(_12742_),
    .Y(_12743_));
 sg13g2_o21ai_1 _38669_ (.B1(_12713_),
    .Y(_12744_),
    .A1(net4544),
    .A2(_12728_));
 sg13g2_nor2_1 _38670_ (.A(_12743_),
    .B(_12744_),
    .Y(_12745_));
 sg13g2_nor2b_1 _38671_ (.A(_12680_),
    .B_N(_12702_),
    .Y(_12746_));
 sg13g2_nand3_1 _38672_ (.B(_12729_),
    .C(_12746_),
    .A(_12714_),
    .Y(_12747_));
 sg13g2_o21ai_1 _38673_ (.B1(_12745_),
    .Y(_12748_),
    .A1(_12688_),
    .A2(_12747_));
 sg13g2_nand2_1 _38674_ (.Y(_12749_),
    .A(_12741_),
    .B(_12748_));
 sg13g2_o21ai_1 _38675_ (.B1(net4699),
    .Y(_12750_),
    .A1(_12741_),
    .A2(_12748_));
 sg13g2_nand2b_1 _38676_ (.Y(_12751_),
    .B(_12749_),
    .A_N(_12750_));
 sg13g2_nand3_1 _38677_ (.B(_12739_),
    .C(_12751_),
    .A(net4400),
    .Y(_12752_));
 sg13g2_a21oi_1 _38678_ (.A1(net4357),
    .A2(_12728_),
    .Y(_12753_),
    .B1(net5539));
 sg13g2_a22oi_1 _38679_ (.Y(_12754_),
    .B1(_12752_),
    .B2(_12753_),
    .A2(net4155),
    .A1(net2457));
 sg13g2_inv_1 _38680_ (.Y(_00977_),
    .A(_12754_));
 sg13g2_nand2b_1 _38681_ (.Y(_12755_),
    .B(net5356),
    .A_N(_07045_));
 sg13g2_a22oi_1 _38682_ (.Y(_12756_),
    .B1(_07212_),
    .B2(_12726_),
    .A2(_07072_),
    .A1(net4800));
 sg13g2_xor2_1 _38683_ (.B(_12756_),
    .A(_07048_),
    .X(_12757_));
 sg13g2_o21ai_1 _38684_ (.B1(_12755_),
    .Y(_12758_),
    .A1(net5354),
    .A2(_12757_));
 sg13g2_nand2_1 _38685_ (.Y(_12759_),
    .A(net4591),
    .B(_12758_));
 sg13g2_nor2_1 _38686_ (.A(net4589),
    .B(_12758_),
    .Y(_12760_));
 sg13g2_xnor2_1 _38687_ (.Y(_12761_),
    .A(net4544),
    .B(_12758_));
 sg13g2_nand2_1 _38688_ (.Y(_12762_),
    .A(_12740_),
    .B(_12749_));
 sg13g2_o21ai_1 _38689_ (.B1(net4699),
    .Y(_12763_),
    .A1(_12761_),
    .A2(_12762_));
 sg13g2_a21oi_1 _38690_ (.A1(_12761_),
    .A2(_12762_),
    .Y(_12764_),
    .B1(_12763_));
 sg13g2_a21oi_1 _38691_ (.A1(net4656),
    .A2(_12758_),
    .Y(_12765_),
    .B1(_12764_));
 sg13g2_o21ai_1 _38692_ (.B1(net5596),
    .Y(_12766_),
    .A1(net4400),
    .A2(_12738_));
 sg13g2_a21oi_1 _38693_ (.A1(net4400),
    .A2(_12765_),
    .Y(_12767_),
    .B1(_12766_));
 sg13g2_a21o_1 _38694_ (.A2(net4153),
    .A1(net2110),
    .B1(_12767_),
    .X(_00978_));
 sg13g2_nor2_1 _38695_ (.A(net5397),
    .B(_07056_),
    .Y(_12768_));
 sg13g2_a21oi_1 _38696_ (.A1(_07047_),
    .A2(_12756_),
    .Y(_12769_),
    .B1(_07046_));
 sg13g2_xnor2_1 _38697_ (.Y(_12770_),
    .A(_07057_),
    .B(_12769_));
 sg13g2_a21oi_2 _38698_ (.B1(_12768_),
    .Y(_12771_),
    .A2(_12770_),
    .A1(net5397));
 sg13g2_xnor2_1 _38699_ (.Y(_12772_),
    .A(net4589),
    .B(_12771_));
 sg13g2_nand2_1 _38700_ (.Y(_12773_),
    .A(_12740_),
    .B(_12759_));
 sg13g2_a21oi_1 _38701_ (.A1(_12741_),
    .A2(_12748_),
    .Y(_12774_),
    .B1(_12773_));
 sg13g2_nor3_1 _38702_ (.A(_12760_),
    .B(_12772_),
    .C(_12774_),
    .Y(_12775_));
 sg13g2_o21ai_1 _38703_ (.B1(_12772_),
    .Y(_12776_),
    .A1(_12760_),
    .A2(_12774_));
 sg13g2_nand3b_1 _38704_ (.B(_12776_),
    .C(net4697),
    .Y(_12777_),
    .A_N(_12775_));
 sg13g2_a21oi_1 _38705_ (.A1(net4652),
    .A2(_12771_),
    .Y(_12778_),
    .B1(net4356));
 sg13g2_o21ai_1 _38706_ (.B1(net5595),
    .Y(_12779_),
    .A1(net4398),
    .A2(_12758_));
 sg13g2_a21oi_1 _38707_ (.A1(_12777_),
    .A2(_12778_),
    .Y(_12780_),
    .B1(_12779_));
 sg13g2_a21o_1 _38708_ (.A2(net4153),
    .A1(net1145),
    .B1(_12780_),
    .X(_00979_));
 sg13g2_nand2_1 _38709_ (.Y(_12781_),
    .A(net2216),
    .B(net4153));
 sg13g2_nand2_1 _38710_ (.Y(_12782_),
    .A(net5355),
    .B(_07025_));
 sg13g2_a21oi_2 _38711_ (.B1(_07220_),
    .Y(_12783_),
    .A2(_09660_),
    .A1(_07279_));
 sg13g2_a21o_1 _38712_ (.A2(_09660_),
    .A1(_07279_),
    .B1(_07220_),
    .X(_12784_));
 sg13g2_xnor2_1 _38713_ (.Y(_12785_),
    .A(_07027_),
    .B(_12783_));
 sg13g2_o21ai_1 _38714_ (.B1(_12782_),
    .Y(_12786_),
    .A1(net5355),
    .A2(_12785_));
 sg13g2_xnor2_1 _38715_ (.Y(_12787_),
    .A(net4541),
    .B(_12786_));
 sg13g2_inv_1 _38716_ (.Y(_12788_),
    .A(_12787_));
 sg13g2_a21oi_1 _38717_ (.A1(net4589),
    .A2(_12771_),
    .Y(_12789_),
    .B1(_12775_));
 sg13g2_nand2b_1 _38718_ (.Y(_12790_),
    .B(_12787_),
    .A_N(_12789_));
 sg13g2_a21oi_1 _38719_ (.A1(_12788_),
    .A2(_12789_),
    .Y(_12791_),
    .B1(net4652));
 sg13g2_a221oi_1 _38720_ (.B2(_12791_),
    .C1(net4356),
    .B1(_12790_),
    .A1(net4652),
    .Y(_12792_),
    .A2(_12786_));
 sg13g2_o21ai_1 _38721_ (.B1(net5595),
    .Y(_12793_),
    .A1(net4398),
    .A2(_12771_));
 sg13g2_o21ai_1 _38722_ (.B1(_12781_),
    .Y(_00980_),
    .A1(_12792_),
    .A2(_12793_));
 sg13g2_nand2_1 _38723_ (.Y(_12794_),
    .A(net2691),
    .B(net4152));
 sg13g2_o21ai_1 _38724_ (.B1(_07026_),
    .Y(_12795_),
    .A1(_07027_),
    .A2(_12783_));
 sg13g2_xor2_1 _38725_ (.B(_12795_),
    .A(_07020_),
    .X(_12796_));
 sg13g2_nor2_1 _38726_ (.A(net5397),
    .B(_07017_),
    .Y(_12797_));
 sg13g2_a21oi_2 _38727_ (.B1(_12797_),
    .Y(_12798_),
    .A2(_12796_),
    .A1(net5397));
 sg13g2_nand2_1 _38728_ (.Y(_12799_),
    .A(net4653),
    .B(_12798_));
 sg13g2_nor2_1 _38729_ (.A(net4541),
    .B(_12798_),
    .Y(_12800_));
 sg13g2_xnor2_1 _38730_ (.Y(_12801_),
    .A(net4588),
    .B(_12798_));
 sg13g2_nand2_1 _38731_ (.Y(_12802_),
    .A(_12741_),
    .B(_12761_));
 sg13g2_nor3_1 _38732_ (.A(_12772_),
    .B(_12788_),
    .C(_12802_),
    .Y(_12803_));
 sg13g2_nor2b_1 _38733_ (.A(_12747_),
    .B_N(_12803_),
    .Y(_12804_));
 sg13g2_nand3b_1 _38734_ (.B(_12803_),
    .C(_12686_),
    .Y(_12805_),
    .A_N(_12747_));
 sg13g2_o21ai_1 _38735_ (.B1(_12803_),
    .Y(_12806_),
    .A1(_12743_),
    .A2(_12744_));
 sg13g2_nand3b_1 _38736_ (.B(_12773_),
    .C(_12787_),
    .Y(_12807_),
    .A_N(_12772_));
 sg13g2_o21ai_1 _38737_ (.B1(net4591),
    .Y(_12808_),
    .A1(_12771_),
    .A2(_12786_));
 sg13g2_nand4_1 _38738_ (.B(_12806_),
    .C(_12807_),
    .A(_12805_),
    .Y(_12809_),
    .D(_12808_));
 sg13g2_and2_1 _38739_ (.A(_12687_),
    .B(_12804_),
    .X(_12810_));
 sg13g2_a21oi_2 _38740_ (.B1(_12809_),
    .Y(_12811_),
    .A2(_12810_),
    .A1(_12563_));
 sg13g2_nor2b_1 _38741_ (.A(_12811_),
    .B_N(_12801_),
    .Y(_12812_));
 sg13g2_xnor2_1 _38742_ (.Y(_12813_),
    .A(_12801_),
    .B(_12811_));
 sg13g2_o21ai_1 _38743_ (.B1(_12799_),
    .Y(_12814_),
    .A1(net4653),
    .A2(_12813_));
 sg13g2_a21oi_1 _38744_ (.A1(net4399),
    .A2(_12814_),
    .Y(_12815_),
    .B1(net5538));
 sg13g2_o21ai_1 _38745_ (.B1(_12815_),
    .Y(_12816_),
    .A1(net4399),
    .A2(_12786_));
 sg13g2_nand2_1 _38746_ (.Y(_00981_),
    .A(_12794_),
    .B(_12816_));
 sg13g2_nand2_1 _38747_ (.Y(_12817_),
    .A(net4357),
    .B(_12798_));
 sg13g2_o21ai_1 _38748_ (.B1(_07230_),
    .Y(_12818_),
    .A1(_07027_),
    .A2(_12783_));
 sg13g2_nand3_1 _38749_ (.B(_07019_),
    .C(_12818_),
    .A(_07009_),
    .Y(_12819_));
 sg13g2_a21o_1 _38750_ (.A2(_12818_),
    .A1(_07019_),
    .B1(_07009_),
    .X(_12820_));
 sg13g2_nand2_1 _38751_ (.Y(_12821_),
    .A(_12819_),
    .B(_12820_));
 sg13g2_nor2_1 _38752_ (.A(net5397),
    .B(_07007_),
    .Y(_12822_));
 sg13g2_a21oi_2 _38753_ (.B1(_12822_),
    .Y(_12823_),
    .A2(_12821_),
    .A1(net5400));
 sg13g2_nand2b_1 _38754_ (.Y(_12824_),
    .B(net4541),
    .A_N(_12823_));
 sg13g2_xnor2_1 _38755_ (.Y(_12825_),
    .A(net4542),
    .B(_12823_));
 sg13g2_nor2_1 _38756_ (.A(_12800_),
    .B(_12812_),
    .Y(_12826_));
 sg13g2_a21oi_1 _38757_ (.A1(_12825_),
    .A2(_12826_),
    .Y(_12827_),
    .B1(net4652));
 sg13g2_o21ai_1 _38758_ (.B1(_12827_),
    .Y(_12828_),
    .A1(_12825_),
    .A2(_12826_));
 sg13g2_o21ai_1 _38759_ (.B1(_12828_),
    .Y(_12829_),
    .A1(net4696),
    .A2(_12823_));
 sg13g2_a21oi_1 _38760_ (.A1(net4398),
    .A2(_12829_),
    .Y(_12830_),
    .B1(net5538));
 sg13g2_a22oi_1 _38761_ (.Y(_12831_),
    .B1(_12817_),
    .B2(_12830_),
    .A2(net4153),
    .A1(net2921));
 sg13g2_inv_1 _38762_ (.Y(_00982_),
    .A(_12831_));
 sg13g2_nand2_1 _38763_ (.Y(_12832_),
    .A(net5355),
    .B(_07001_));
 sg13g2_nand2b_1 _38764_ (.Y(_12833_),
    .B(_12819_),
    .A_N(_07008_));
 sg13g2_xnor2_1 _38765_ (.Y(_12834_),
    .A(_07002_),
    .B(_12833_));
 sg13g2_o21ai_1 _38766_ (.B1(_12832_),
    .Y(_12835_),
    .A1(net5355),
    .A2(_12834_));
 sg13g2_nand2_1 _38767_ (.Y(_12836_),
    .A(net4588),
    .B(_12835_));
 sg13g2_xnor2_1 _38768_ (.Y(_12837_),
    .A(net4587),
    .B(_12835_));
 sg13g2_a21o_1 _38769_ (.A2(_12823_),
    .A1(net4588),
    .B1(_12800_),
    .X(_12838_));
 sg13g2_o21ai_1 _38770_ (.B1(_12824_),
    .Y(_12839_),
    .A1(_12812_),
    .A2(_12838_));
 sg13g2_xnor2_1 _38771_ (.Y(_12840_),
    .A(_12837_),
    .B(_12839_));
 sg13g2_nand2_1 _38772_ (.Y(_12841_),
    .A(net4696),
    .B(_12840_));
 sg13g2_o21ai_1 _38773_ (.B1(_12841_),
    .Y(_12842_),
    .A1(net4696),
    .A2(_12835_));
 sg13g2_o21ai_1 _38774_ (.B1(net5595),
    .Y(_12843_),
    .A1(net4398),
    .A2(_12823_));
 sg13g2_a21oi_1 _38775_ (.A1(net4398),
    .A2(_12842_),
    .Y(_12844_),
    .B1(_12843_));
 sg13g2_a21o_1 _38776_ (.A2(net4153),
    .A1(net2737),
    .B1(_12844_),
    .X(_00983_));
 sg13g2_nand2_1 _38777_ (.Y(_12845_),
    .A(net2099),
    .B(net4153));
 sg13g2_a21oi_1 _38778_ (.A1(_07030_),
    .A2(_12784_),
    .Y(_12846_),
    .B1(_07232_));
 sg13g2_xnor2_1 _38779_ (.Y(_12847_),
    .A(_06992_),
    .B(_12846_));
 sg13g2_nor2_1 _38780_ (.A(net5355),
    .B(_12847_),
    .Y(_12848_));
 sg13g2_a21oi_2 _38781_ (.B1(_12848_),
    .Y(_12849_),
    .A2(_06990_),
    .A1(net5355));
 sg13g2_xnor2_1 _38782_ (.Y(_12850_),
    .A(net4587),
    .B(_12849_));
 sg13g2_o21ai_1 _38783_ (.B1(_12836_),
    .Y(_12851_),
    .A1(_12837_),
    .A2(_12839_));
 sg13g2_xor2_1 _38784_ (.B(_12851_),
    .A(_12850_),
    .X(_12852_));
 sg13g2_o21ai_1 _38785_ (.B1(net4398),
    .Y(_12853_),
    .A1(net4696),
    .A2(_12849_));
 sg13g2_a21oi_1 _38786_ (.A1(net4696),
    .A2(_12852_),
    .Y(_12854_),
    .B1(_12853_));
 sg13g2_o21ai_1 _38787_ (.B1(net5595),
    .Y(_12855_),
    .A1(net4398),
    .A2(_12835_));
 sg13g2_o21ai_1 _38788_ (.B1(_12845_),
    .Y(_00984_),
    .A1(_12854_),
    .A2(_12855_));
 sg13g2_o21ai_1 _38789_ (.B1(_06991_),
    .Y(_12856_),
    .A1(_06992_),
    .A2(_12846_));
 sg13g2_xnor2_1 _38790_ (.Y(_12857_),
    .A(_06985_),
    .B(_12856_));
 sg13g2_mux2_1 _38791_ (.A0(_06983_),
    .A1(_12857_),
    .S(net5400),
    .X(_12858_));
 sg13g2_nand2_1 _38792_ (.Y(_12859_),
    .A(net4587),
    .B(_12858_));
 sg13g2_xnor2_1 _38793_ (.Y(_12860_),
    .A(net4542),
    .B(_12858_));
 sg13g2_nor2b_1 _38794_ (.A(_12837_),
    .B_N(_12850_),
    .Y(_12861_));
 sg13g2_o21ai_1 _38795_ (.B1(_12836_),
    .Y(_12862_),
    .A1(net4542),
    .A2(_12849_));
 sg13g2_a21oi_1 _38796_ (.A1(_12838_),
    .A2(_12861_),
    .Y(_12863_),
    .B1(_12862_));
 sg13g2_nand3_1 _38797_ (.B(_12825_),
    .C(_12861_),
    .A(_12801_),
    .Y(_12864_));
 sg13g2_o21ai_1 _38798_ (.B1(_12863_),
    .Y(_12865_),
    .A1(_12811_),
    .A2(_12864_));
 sg13g2_nand2_1 _38799_ (.Y(_12866_),
    .A(_12860_),
    .B(_12865_));
 sg13g2_or2_1 _38800_ (.X(_12867_),
    .B(_12865_),
    .A(_12860_));
 sg13g2_a21o_1 _38801_ (.A2(_12867_),
    .A1(_12866_),
    .B1(net4652),
    .X(_12868_));
 sg13g2_o21ai_1 _38802_ (.B1(_12868_),
    .Y(_12869_),
    .A1(net4696),
    .A2(_12858_));
 sg13g2_nand2_1 _38803_ (.Y(_12870_),
    .A(net4357),
    .B(_12849_));
 sg13g2_a21oi_1 _38804_ (.A1(net4398),
    .A2(_12869_),
    .Y(_12871_),
    .B1(net5538));
 sg13g2_a22oi_1 _38805_ (.Y(_12872_),
    .B1(_12870_),
    .B2(_12871_),
    .A2(net4152),
    .A1(net2496));
 sg13g2_inv_1 _38806_ (.Y(_00985_),
    .A(_12872_));
 sg13g2_nand2_1 _38807_ (.Y(_12873_),
    .A(net1674),
    .B(net4153));
 sg13g2_o21ai_1 _38808_ (.B1(_07233_),
    .Y(_12874_),
    .A1(_06992_),
    .A2(_12846_));
 sg13g2_nand3_1 _38809_ (.B(_06984_),
    .C(_12874_),
    .A(_06964_),
    .Y(_12875_));
 sg13g2_a21oi_1 _38810_ (.A1(_06984_),
    .A2(_12874_),
    .Y(_12876_),
    .B1(_06964_));
 sg13g2_nor2_1 _38811_ (.A(net5351),
    .B(_12876_),
    .Y(_12877_));
 sg13g2_a22oi_1 _38812_ (.Y(_12878_),
    .B1(_12875_),
    .B2(_12877_),
    .A2(_06962_),
    .A1(net5351));
 sg13g2_nor2_1 _38813_ (.A(net4542),
    .B(_12878_),
    .Y(_12879_));
 sg13g2_xnor2_1 _38814_ (.Y(_12880_),
    .A(net4587),
    .B(_12878_));
 sg13g2_nand2_1 _38815_ (.Y(_12881_),
    .A(_12859_),
    .B(_12866_));
 sg13g2_xnor2_1 _38816_ (.Y(_12882_),
    .A(_12880_),
    .B(_12881_));
 sg13g2_nand2_1 _38817_ (.Y(_12883_),
    .A(net4652),
    .B(_12878_));
 sg13g2_a21oi_1 _38818_ (.A1(net4696),
    .A2(_12882_),
    .Y(_12884_),
    .B1(net4356));
 sg13g2_a22oi_1 _38819_ (.Y(_12885_),
    .B1(_12883_),
    .B2(_12884_),
    .A2(_12858_),
    .A1(net4356));
 sg13g2_o21ai_1 _38820_ (.B1(_12873_),
    .Y(_00986_),
    .A1(net5538),
    .A2(_12885_));
 sg13g2_nor2_1 _38821_ (.A(net5394),
    .B(_06972_),
    .Y(_12886_));
 sg13g2_nand2_1 _38822_ (.Y(_12887_),
    .A(_06963_),
    .B(_12875_));
 sg13g2_xnor2_1 _38823_ (.Y(_12888_),
    .A(_06973_),
    .B(_12887_));
 sg13g2_a21oi_2 _38824_ (.B1(_12886_),
    .Y(_12889_),
    .A2(_12888_),
    .A1(net5396));
 sg13g2_xnor2_1 _38825_ (.Y(_12890_),
    .A(net4587),
    .B(_12889_));
 sg13g2_a21oi_1 _38826_ (.A1(net4587),
    .A2(_12858_),
    .Y(_12891_),
    .B1(_12879_));
 sg13g2_a22oi_1 _38827_ (.Y(_12892_),
    .B1(_12891_),
    .B2(_12866_),
    .A2(_12878_),
    .A1(net4542));
 sg13g2_nor2b_1 _38828_ (.A(_12890_),
    .B_N(_12892_),
    .Y(_12893_));
 sg13g2_xnor2_1 _38829_ (.Y(_12894_),
    .A(_12890_),
    .B(_12892_));
 sg13g2_nand2_1 _38830_ (.Y(_12895_),
    .A(net4652),
    .B(_12889_));
 sg13g2_nand2_1 _38831_ (.Y(_12896_),
    .A(net4394),
    .B(_12895_));
 sg13g2_a21oi_1 _38832_ (.A1(net4696),
    .A2(_12894_),
    .Y(_12897_),
    .B1(_12896_));
 sg13g2_a21oi_1 _38833_ (.A1(net4355),
    .A2(_12878_),
    .Y(_12898_),
    .B1(_12897_));
 sg13g2_a22oi_1 _38834_ (.Y(_12899_),
    .B1(_12898_),
    .B2(net5593),
    .A2(net4138),
    .A1(net3177));
 sg13g2_inv_1 _38835_ (.Y(_00987_),
    .A(_12899_));
 sg13g2_nand2_1 _38836_ (.Y(_12900_),
    .A(net3106),
    .B(net4137));
 sg13g2_nand2_1 _38837_ (.Y(_12901_),
    .A(net5351),
    .B(_06945_));
 sg13g2_o21ai_1 _38838_ (.B1(_07235_),
    .Y(_12902_),
    .A1(_07032_),
    .A2(_12783_));
 sg13g2_nand2_1 _38839_ (.Y(_12903_),
    .A(_06948_),
    .B(_12902_));
 sg13g2_xnor2_1 _38840_ (.Y(_12904_),
    .A(_06948_),
    .B(_12902_));
 sg13g2_o21ai_1 _38841_ (.B1(_12901_),
    .Y(_12905_),
    .A1(net5351),
    .A2(_12904_));
 sg13g2_xnor2_1 _38842_ (.Y(_12906_),
    .A(net4585),
    .B(_12905_));
 sg13g2_a21oi_1 _38843_ (.A1(net4587),
    .A2(_12889_),
    .Y(_12907_),
    .B1(_12893_));
 sg13g2_or2_1 _38844_ (.X(_12908_),
    .B(_12907_),
    .A(_12906_));
 sg13g2_a21oi_1 _38845_ (.A1(_12906_),
    .A2(_12907_),
    .Y(_12909_),
    .B1(net4652));
 sg13g2_a221oi_1 _38846_ (.B2(_12909_),
    .C1(net4355),
    .B1(_12908_),
    .A1(net4650),
    .Y(_12910_),
    .A2(_12905_));
 sg13g2_o21ai_1 _38847_ (.B1(net5593),
    .Y(_12911_),
    .A1(net4394),
    .A2(_12889_));
 sg13g2_o21ai_1 _38848_ (.B1(_12900_),
    .Y(_00988_),
    .A1(_12910_),
    .A2(_12911_));
 sg13g2_nand2_1 _38849_ (.Y(_12912_),
    .A(net5352),
    .B(_06937_));
 sg13g2_nand2_1 _38850_ (.Y(_12913_),
    .A(_06946_),
    .B(_12903_));
 sg13g2_xnor2_1 _38851_ (.Y(_12914_),
    .A(_06940_),
    .B(_12913_));
 sg13g2_o21ai_1 _38852_ (.B1(_12912_),
    .Y(_12915_),
    .A1(net5351),
    .A2(_12914_));
 sg13g2_nand2_1 _38853_ (.Y(_12916_),
    .A(net4585),
    .B(_12915_));
 sg13g2_xnor2_1 _38854_ (.Y(_12917_),
    .A(net4538),
    .B(_12915_));
 sg13g2_nor2_1 _38855_ (.A(_12890_),
    .B(_12906_),
    .Y(_12918_));
 sg13g2_and2_1 _38856_ (.A(_12860_),
    .B(_12880_),
    .X(_12919_));
 sg13g2_nand3b_1 _38857_ (.B(_12918_),
    .C(_12919_),
    .Y(_12920_),
    .A_N(_12863_));
 sg13g2_nand2b_1 _38858_ (.Y(_12921_),
    .B(_12918_),
    .A_N(_12891_));
 sg13g2_o21ai_1 _38859_ (.B1(net4587),
    .Y(_12922_),
    .A1(_12889_),
    .A2(_12905_));
 sg13g2_and3_1 _38860_ (.X(_12923_),
    .A(_12920_),
    .B(_12921_),
    .C(_12922_));
 sg13g2_nand3b_1 _38861_ (.B(_12918_),
    .C(_12919_),
    .Y(_12924_),
    .A_N(_12864_));
 sg13g2_o21ai_1 _38862_ (.B1(_12923_),
    .Y(_12925_),
    .A1(_12811_),
    .A2(_12924_));
 sg13g2_nand2_2 _38863_ (.Y(_12926_),
    .A(_12917_),
    .B(_12925_));
 sg13g2_or2_1 _38864_ (.X(_12927_),
    .B(_12925_),
    .A(_12917_));
 sg13g2_a21o_1 _38865_ (.A2(_12927_),
    .A1(_12926_),
    .B1(net4648),
    .X(_12928_));
 sg13g2_o21ai_1 _38866_ (.B1(_12928_),
    .Y(_12929_),
    .A1(net4692),
    .A2(_12915_));
 sg13g2_o21ai_1 _38867_ (.B1(net5594),
    .Y(_12930_),
    .A1(net4395),
    .A2(_12905_));
 sg13g2_a21oi_1 _38868_ (.A1(net4394),
    .A2(_12929_),
    .Y(_12931_),
    .B1(_12930_));
 sg13g2_a21o_1 _38869_ (.A2(net4138),
    .A1(net3095),
    .B1(_12931_),
    .X(_00989_));
 sg13g2_nand2_1 _38870_ (.Y(_12932_),
    .A(net2575),
    .B(net4138));
 sg13g2_nand2_1 _38871_ (.Y(_12933_),
    .A(net5351),
    .B(_06918_));
 sg13g2_a21oi_1 _38872_ (.A1(_06948_),
    .A2(_12902_),
    .Y(_12934_),
    .B1(_07222_));
 sg13g2_nor3_1 _38873_ (.A(_06920_),
    .B(_06939_),
    .C(_12934_),
    .Y(_12935_));
 sg13g2_o21ai_1 _38874_ (.B1(_06920_),
    .Y(_12936_),
    .A1(_06939_),
    .A2(_12934_));
 sg13g2_nand3b_1 _38875_ (.B(_12936_),
    .C(net5394),
    .Y(_12937_),
    .A_N(_12935_));
 sg13g2_and2_1 _38876_ (.A(_12933_),
    .B(_12937_),
    .X(_12938_));
 sg13g2_nor2_1 _38877_ (.A(net4537),
    .B(_12938_),
    .Y(_12939_));
 sg13g2_xnor2_1 _38878_ (.Y(_12940_),
    .A(net4586),
    .B(_12938_));
 sg13g2_nand2_1 _38879_ (.Y(_12941_),
    .A(_12916_),
    .B(_12926_));
 sg13g2_xor2_1 _38880_ (.B(_12941_),
    .A(_12940_),
    .X(_12942_));
 sg13g2_o21ai_1 _38881_ (.B1(net4395),
    .Y(_12943_),
    .A1(net4692),
    .A2(_12938_));
 sg13g2_a21oi_1 _38882_ (.A1(net4693),
    .A2(_12942_),
    .Y(_12944_),
    .B1(_12943_));
 sg13g2_o21ai_1 _38883_ (.B1(net5593),
    .Y(_12945_),
    .A1(net4395),
    .A2(_12915_));
 sg13g2_o21ai_1 _38884_ (.B1(_12932_),
    .Y(_00990_),
    .A1(_12944_),
    .A2(_12945_));
 sg13g2_nand2_1 _38885_ (.Y(_12946_),
    .A(net5351),
    .B(_06928_));
 sg13g2_a21oi_1 _38886_ (.A1(net4739),
    .A2(_06918_),
    .Y(_12947_),
    .B1(_12935_));
 sg13g2_xor2_1 _38887_ (.B(_12947_),
    .A(_06929_),
    .X(_12948_));
 sg13g2_o21ai_1 _38888_ (.B1(_12946_),
    .Y(_12949_),
    .A1(net5351),
    .A2(_12948_));
 sg13g2_and2_1 _38889_ (.A(net4585),
    .B(_12949_),
    .X(_12950_));
 sg13g2_xnor2_1 _38890_ (.Y(_12951_),
    .A(net4537),
    .B(_12949_));
 sg13g2_inv_1 _38891_ (.Y(_12952_),
    .A(_12951_));
 sg13g2_a21oi_1 _38892_ (.A1(net4586),
    .A2(_12915_),
    .Y(_12953_),
    .B1(_12939_));
 sg13g2_a22oi_1 _38893_ (.Y(_12954_),
    .B1(_12953_),
    .B2(_12926_),
    .A2(_12938_),
    .A1(net4537));
 sg13g2_a221oi_1 _38894_ (.B2(_12926_),
    .C1(_12952_),
    .B1(_12953_),
    .A1(net4538),
    .Y(_12955_),
    .A2(_12938_));
 sg13g2_nor2_1 _38895_ (.A(net4648),
    .B(_12955_),
    .Y(_12956_));
 sg13g2_o21ai_1 _38896_ (.B1(_12956_),
    .Y(_12957_),
    .A1(_12951_),
    .A2(_12954_));
 sg13g2_nand2_1 _38897_ (.Y(_12958_),
    .A(net4648),
    .B(_12949_));
 sg13g2_nand3_1 _38898_ (.B(_12957_),
    .C(_12958_),
    .A(net4395),
    .Y(_12959_));
 sg13g2_a21oi_1 _38899_ (.A1(net4355),
    .A2(_12938_),
    .Y(_12960_),
    .B1(net5529));
 sg13g2_a22oi_1 _38900_ (.Y(_12961_),
    .B1(_12959_),
    .B2(_12960_),
    .A2(net4138),
    .A1(net2060));
 sg13g2_inv_1 _38901_ (.Y(_00991_),
    .A(_12961_));
 sg13g2_nor2_1 _38902_ (.A(net5394),
    .B(_06907_),
    .Y(_12962_));
 sg13g2_a21oi_2 _38903_ (.B1(_07225_),
    .Y(_12963_),
    .A2(_12902_),
    .A1(_06949_));
 sg13g2_xnor2_1 _38904_ (.Y(_12964_),
    .A(_06909_),
    .B(_12963_));
 sg13g2_a21oi_2 _38905_ (.B1(_12962_),
    .Y(_12965_),
    .A2(_12964_),
    .A1(net5394));
 sg13g2_nor2_1 _38906_ (.A(net4537),
    .B(_12965_),
    .Y(_12966_));
 sg13g2_xnor2_1 _38907_ (.Y(_12967_),
    .A(net4585),
    .B(_12965_));
 sg13g2_o21ai_1 _38908_ (.B1(_12967_),
    .Y(_12968_),
    .A1(_12950_),
    .A2(_12955_));
 sg13g2_nor3_1 _38909_ (.A(_12950_),
    .B(_12955_),
    .C(_12967_),
    .Y(_12969_));
 sg13g2_nor2_1 _38910_ (.A(net4648),
    .B(_12969_),
    .Y(_12970_));
 sg13g2_nor2_1 _38911_ (.A(net4693),
    .B(_12965_),
    .Y(_12971_));
 sg13g2_a21oi_1 _38912_ (.A1(_12968_),
    .A2(_12970_),
    .Y(_12972_),
    .B1(_12971_));
 sg13g2_o21ai_1 _38913_ (.B1(net5594),
    .Y(_12973_),
    .A1(net4394),
    .A2(_12949_));
 sg13g2_a21oi_1 _38914_ (.A1(net4394),
    .A2(_12972_),
    .Y(_12974_),
    .B1(_12973_));
 sg13g2_a21o_1 _38915_ (.A2(net4138),
    .A1(net2530),
    .B1(_12974_),
    .X(_00992_));
 sg13g2_o21ai_1 _38916_ (.B1(_06908_),
    .Y(_12975_),
    .A1(_06910_),
    .A2(_12963_));
 sg13g2_xnor2_1 _38917_ (.Y(_12976_),
    .A(_06902_),
    .B(_12975_));
 sg13g2_mux2_1 _38918_ (.A0(_06900_),
    .A1(_12976_),
    .S(net5394),
    .X(_12977_));
 sg13g2_nor2_1 _38919_ (.A(net4537),
    .B(_12977_),
    .Y(_12978_));
 sg13g2_xnor2_1 _38920_ (.Y(_12979_),
    .A(net4537),
    .B(_12977_));
 sg13g2_nand2_1 _38921_ (.Y(_12980_),
    .A(_12951_),
    .B(_12967_));
 sg13g2_nor2_1 _38922_ (.A(_12953_),
    .B(_12980_),
    .Y(_12981_));
 sg13g2_nor3_1 _38923_ (.A(_12950_),
    .B(_12966_),
    .C(_12981_),
    .Y(_12982_));
 sg13g2_and4_1 _38924_ (.A(_12917_),
    .B(_12940_),
    .C(_12951_),
    .D(_12967_),
    .X(_12983_));
 sg13g2_nand2_1 _38925_ (.Y(_12984_),
    .A(_12925_),
    .B(_12983_));
 sg13g2_a21o_2 _38926_ (.A2(_12984_),
    .A1(_12982_),
    .B1(_12979_),
    .X(_12985_));
 sg13g2_nand3_1 _38927_ (.B(_12982_),
    .C(_12984_),
    .A(_12979_),
    .Y(_12986_));
 sg13g2_nand3_1 _38928_ (.B(_12985_),
    .C(_12986_),
    .A(net4693),
    .Y(_12987_));
 sg13g2_o21ai_1 _38929_ (.B1(net4394),
    .Y(_12988_),
    .A1(net4693),
    .A2(_12977_));
 sg13g2_nand2b_1 _38930_ (.Y(_12989_),
    .B(_12987_),
    .A_N(_12988_));
 sg13g2_a21oi_1 _38931_ (.A1(net4355),
    .A2(_12965_),
    .Y(_12990_),
    .B1(net5530));
 sg13g2_a22oi_1 _38932_ (.Y(_12991_),
    .B1(_12989_),
    .B2(_12990_),
    .A2(net4137),
    .A1(net3091));
 sg13g2_inv_1 _38933_ (.Y(_00993_),
    .A(_12991_));
 sg13g2_nor2b_1 _38934_ (.A(_12978_),
    .B_N(_12985_),
    .Y(_12992_));
 sg13g2_o21ai_1 _38935_ (.B1(_07227_),
    .Y(_12993_),
    .A1(_06910_),
    .A2(_12963_));
 sg13g2_nand3_1 _38936_ (.B(_06901_),
    .C(_12993_),
    .A(_06881_),
    .Y(_12994_));
 sg13g2_a21o_1 _38937_ (.A2(_12993_),
    .A1(_06901_),
    .B1(_06881_),
    .X(_12995_));
 sg13g2_nand3_1 _38938_ (.B(_12994_),
    .C(_12995_),
    .A(net5394),
    .Y(_12996_));
 sg13g2_o21ai_1 _38939_ (.B1(_12996_),
    .Y(_12997_),
    .A1(net5394),
    .A2(_06879_));
 sg13g2_inv_1 _38940_ (.Y(_12998_),
    .A(_12997_));
 sg13g2_xnor2_1 _38941_ (.Y(_12999_),
    .A(net4585),
    .B(_12997_));
 sg13g2_xnor2_1 _38942_ (.Y(_13000_),
    .A(_12992_),
    .B(_12999_));
 sg13g2_a21oi_1 _38943_ (.A1(net4648),
    .A2(_12997_),
    .Y(_13001_),
    .B1(net4355));
 sg13g2_o21ai_1 _38944_ (.B1(_13001_),
    .Y(_13002_),
    .A1(net4648),
    .A2(_13000_));
 sg13g2_a21oi_1 _38945_ (.A1(net4355),
    .A2(_12977_),
    .Y(_13003_),
    .B1(net5530));
 sg13g2_a22oi_1 _38946_ (.Y(_13004_),
    .B1(_13002_),
    .B2(_13003_),
    .A2(net4138),
    .A1(net2988));
 sg13g2_inv_1 _38947_ (.Y(_00994_),
    .A(_13004_));
 sg13g2_nand2_1 _38948_ (.Y(_13005_),
    .A(_06880_),
    .B(_12994_));
 sg13g2_xor2_1 _38949_ (.B(_13005_),
    .A(_06892_),
    .X(_13006_));
 sg13g2_mux2_1 _38950_ (.A0(_06890_),
    .A1(_13006_),
    .S(net5394),
    .X(_13007_));
 sg13g2_and2_1 _38951_ (.A(net4583),
    .B(_13007_),
    .X(_13008_));
 sg13g2_xnor2_1 _38952_ (.Y(_13009_),
    .A(net4585),
    .B(_13007_));
 sg13g2_a21oi_1 _38953_ (.A1(net4585),
    .A2(_12997_),
    .Y(_13010_),
    .B1(_12978_));
 sg13g2_inv_1 _38954_ (.Y(_13011_),
    .A(_13010_));
 sg13g2_a22oi_1 _38955_ (.Y(_13012_),
    .B1(_13010_),
    .B2(_12985_),
    .A2(_12998_),
    .A1(net4537));
 sg13g2_a221oi_1 _38956_ (.B2(_12985_),
    .C1(_13009_),
    .B1(_13010_),
    .A1(net4537),
    .Y(_13013_),
    .A2(_12998_));
 sg13g2_xnor2_1 _38957_ (.Y(_13014_),
    .A(_13009_),
    .B(_13012_));
 sg13g2_or2_1 _38958_ (.X(_13015_),
    .B(_13007_),
    .A(net4693));
 sg13g2_o21ai_1 _38959_ (.B1(_13015_),
    .Y(_13016_),
    .A1(net4648),
    .A2(_13014_));
 sg13g2_o21ai_1 _38960_ (.B1(net5594),
    .Y(_13017_),
    .A1(net4394),
    .A2(_12997_));
 sg13g2_a21oi_1 _38961_ (.A1(net4394),
    .A2(_13016_),
    .Y(_13018_),
    .B1(_13017_));
 sg13g2_a21o_1 _38962_ (.A2(net4139),
    .A1(net3187),
    .B1(_13018_),
    .X(_00995_));
 sg13g2_nand2_1 _38963_ (.Y(_13019_),
    .A(net2528),
    .B(net4136));
 sg13g2_nand2_1 _38964_ (.Y(_13020_),
    .A(net5350),
    .B(_06838_));
 sg13g2_o21ai_1 _38965_ (.B1(_07237_),
    .Y(_13021_),
    .A1(_07280_),
    .A2(_09659_));
 sg13g2_xnor2_1 _38966_ (.Y(_13022_),
    .A(_06841_),
    .B(_13021_));
 sg13g2_o21ai_1 _38967_ (.B1(_13020_),
    .Y(_13023_),
    .A1(net5353),
    .A2(_13022_));
 sg13g2_xnor2_1 _38968_ (.Y(_13024_),
    .A(net4539),
    .B(_13023_));
 sg13g2_nor3_1 _38969_ (.A(_13008_),
    .B(_13013_),
    .C(_13024_),
    .Y(_13025_));
 sg13g2_o21ai_1 _38970_ (.B1(_13024_),
    .Y(_13026_),
    .A1(_13008_),
    .A2(_13013_));
 sg13g2_nor2_1 _38971_ (.A(net4648),
    .B(_13025_),
    .Y(_13027_));
 sg13g2_a221oi_1 _38972_ (.B2(_13027_),
    .C1(net4354),
    .B1(_13026_),
    .A1(net4650),
    .Y(_13028_),
    .A2(_13023_));
 sg13g2_o21ai_1 _38973_ (.B1(net5594),
    .Y(_13029_),
    .A1(net4391),
    .A2(_13007_));
 sg13g2_o21ai_1 _38974_ (.B1(_13019_),
    .Y(_00996_),
    .A1(_13028_),
    .A2(_13029_));
 sg13g2_nand2_1 _38975_ (.Y(_13030_),
    .A(net2887),
    .B(net4136));
 sg13g2_nand2_1 _38976_ (.Y(_13031_),
    .A(net5348),
    .B(_06850_));
 sg13g2_a21oi_1 _38977_ (.A1(_06841_),
    .A2(_13021_),
    .Y(_13032_),
    .B1(_06840_));
 sg13g2_xnor2_1 _38978_ (.Y(_13033_),
    .A(_06852_),
    .B(_13032_));
 sg13g2_o21ai_1 _38979_ (.B1(_13031_),
    .Y(_13034_),
    .A1(net5348),
    .A2(_13033_));
 sg13g2_nand2_1 _38980_ (.Y(_13035_),
    .A(net4650),
    .B(_13034_));
 sg13g2_nor2_1 _38981_ (.A(net4535),
    .B(_13034_),
    .Y(_13036_));
 sg13g2_xnor2_1 _38982_ (.Y(_13037_),
    .A(net4579),
    .B(_13034_));
 sg13g2_nor2b_1 _38983_ (.A(_13009_),
    .B_N(_13024_),
    .Y(_13038_));
 sg13g2_nor2_1 _38984_ (.A(_12979_),
    .B(_12999_),
    .Y(_13039_));
 sg13g2_and3_2 _38985_ (.X(_13040_),
    .A(_12983_),
    .B(_13038_),
    .C(_13039_));
 sg13g2_nor2b_1 _38986_ (.A(_12924_),
    .B_N(_13040_),
    .Y(_13041_));
 sg13g2_and2_1 _38987_ (.A(_12810_),
    .B(_13041_),
    .X(_13042_));
 sg13g2_nand3b_1 _38988_ (.B(_13040_),
    .C(_12809_),
    .Y(_13043_),
    .A_N(_12924_));
 sg13g2_nand2b_1 _38989_ (.Y(_13044_),
    .B(_13040_),
    .A_N(_12923_));
 sg13g2_nand3b_1 _38990_ (.B(_13038_),
    .C(_13039_),
    .Y(_13045_),
    .A_N(_12982_));
 sg13g2_a221oi_1 _38991_ (.B2(_13011_),
    .C1(_13008_),
    .B1(_13038_),
    .A1(net4585),
    .Y(_13046_),
    .A2(_13023_));
 sg13g2_nand4_1 _38992_ (.B(_13044_),
    .C(_13045_),
    .A(_13043_),
    .Y(_13047_),
    .D(_13046_));
 sg13g2_a21o_2 _38993_ (.A2(_13042_),
    .A1(_12563_),
    .B1(_13047_),
    .X(_13048_));
 sg13g2_nand2_1 _38994_ (.Y(_13049_),
    .A(_13037_),
    .B(_13048_));
 sg13g2_xor2_1 _38995_ (.B(_13048_),
    .A(_13037_),
    .X(_13050_));
 sg13g2_o21ai_1 _38996_ (.B1(_13035_),
    .Y(_13051_),
    .A1(net4650),
    .A2(_13050_));
 sg13g2_a21oi_1 _38997_ (.A1(net4391),
    .A2(_13051_),
    .Y(_13052_),
    .B1(net5529));
 sg13g2_o21ai_1 _38998_ (.B1(_13052_),
    .Y(_13053_),
    .A1(net4391),
    .A2(_13023_));
 sg13g2_nand2_1 _38999_ (.Y(_00997_),
    .A(_13030_),
    .B(_13053_));
 sg13g2_nand2_1 _39000_ (.Y(_13054_),
    .A(net5348),
    .B(_06829_));
 sg13g2_a21oi_1 _39001_ (.A1(_06841_),
    .A2(_13021_),
    .Y(_13055_),
    .B1(_07238_));
 sg13g2_nor3_1 _39002_ (.A(_06833_),
    .B(_06851_),
    .C(_13055_),
    .Y(_13056_));
 sg13g2_o21ai_1 _39003_ (.B1(_06833_),
    .Y(_13057_),
    .A1(_06851_),
    .A2(_13055_));
 sg13g2_nand2_1 _39004_ (.Y(_13058_),
    .A(net5392),
    .B(_13057_));
 sg13g2_o21ai_1 _39005_ (.B1(_13054_),
    .Y(_13059_),
    .A1(_13056_),
    .A2(_13058_));
 sg13g2_nor2_1 _39006_ (.A(net4579),
    .B(_13059_),
    .Y(_13060_));
 sg13g2_xnor2_1 _39007_ (.Y(_13061_),
    .A(net4535),
    .B(_13059_));
 sg13g2_a21oi_1 _39008_ (.A1(_13037_),
    .A2(_13048_),
    .Y(_13062_),
    .B1(_13036_));
 sg13g2_xor2_1 _39009_ (.B(_13062_),
    .A(_13061_),
    .X(_13063_));
 sg13g2_nor2_1 _39010_ (.A(net4688),
    .B(_13059_),
    .Y(_13064_));
 sg13g2_a21oi_1 _39011_ (.A1(net4690),
    .A2(_13063_),
    .Y(_13065_),
    .B1(_13064_));
 sg13g2_nor2_1 _39012_ (.A(net4352),
    .B(_13065_),
    .Y(_13066_));
 sg13g2_a21oi_1 _39013_ (.A1(net4354),
    .A2(_13034_),
    .Y(_13067_),
    .B1(_13066_));
 sg13g2_a22oi_1 _39014_ (.Y(_13068_),
    .B1(_13067_),
    .B2(net5594),
    .A2(net4136),
    .A1(net2949));
 sg13g2_inv_1 _39015_ (.Y(_00998_),
    .A(_13068_));
 sg13g2_or3_1 _39016_ (.A(_06823_),
    .B(_06830_),
    .C(_13056_),
    .X(_13069_));
 sg13g2_o21ai_1 _39017_ (.B1(_06823_),
    .Y(_13070_),
    .A1(_06830_),
    .A2(_13056_));
 sg13g2_a21o_2 _39018_ (.A2(_13070_),
    .A1(_13069_),
    .B1(net5348),
    .X(_13071_));
 sg13g2_nand3_1 _39019_ (.B(_06815_),
    .C(_06820_),
    .A(net5349),
    .Y(_13072_));
 sg13g2_nand2_1 _39020_ (.Y(_13073_),
    .A(_13071_),
    .B(_13072_));
 sg13g2_a21oi_2 _39021_ (.B1(net4535),
    .Y(_13074_),
    .A2(_13072_),
    .A1(_13071_));
 sg13g2_and3_1 _39022_ (.X(_13075_),
    .A(net4540),
    .B(_13071_),
    .C(_13072_));
 sg13g2_or2_1 _39023_ (.X(_13076_),
    .B(_13075_),
    .A(_13074_));
 sg13g2_a21oi_1 _39024_ (.A1(net4579),
    .A2(_13059_),
    .Y(_13077_),
    .B1(_13036_));
 sg13g2_a21oi_1 _39025_ (.A1(_13049_),
    .A2(_13077_),
    .Y(_13078_),
    .B1(_13060_));
 sg13g2_nor2b_1 _39026_ (.A(_13076_),
    .B_N(_13078_),
    .Y(_13079_));
 sg13g2_xor2_1 _39027_ (.B(_13078_),
    .A(_13076_),
    .X(_13080_));
 sg13g2_nand2_1 _39028_ (.Y(_13081_),
    .A(net4690),
    .B(_13080_));
 sg13g2_o21ai_1 _39029_ (.B1(_13081_),
    .Y(_13082_),
    .A1(net4688),
    .A2(_13073_));
 sg13g2_o21ai_1 _39030_ (.B1(net5590),
    .Y(_13083_),
    .A1(net4386),
    .A2(_13059_));
 sg13g2_a21oi_1 _39031_ (.A1(net4386),
    .A2(_13082_),
    .Y(_13084_),
    .B1(_13083_));
 sg13g2_a21o_1 _39032_ (.A2(net4136),
    .A1(net5875),
    .B1(_13084_),
    .X(_00999_));
 sg13g2_nand2_1 _39033_ (.Y(_13085_),
    .A(net2189),
    .B(net4126));
 sg13g2_nand2_1 _39034_ (.Y(_13086_),
    .A(net5348),
    .B(_06796_));
 sg13g2_a21oi_1 _39035_ (.A1(_06854_),
    .A2(_13021_),
    .Y(_13087_),
    .B1(_07240_));
 sg13g2_xnor2_1 _39036_ (.Y(_13088_),
    .A(_06799_),
    .B(_13087_));
 sg13g2_o21ai_1 _39037_ (.B1(_13086_),
    .Y(_13089_),
    .A1(net5348),
    .A2(_13088_));
 sg13g2_xnor2_1 _39038_ (.Y(_13090_),
    .A(net4579),
    .B(_13089_));
 sg13g2_nor2_1 _39039_ (.A(_13074_),
    .B(_13079_),
    .Y(_13091_));
 sg13g2_or2_1 _39040_ (.X(_13092_),
    .B(_13091_),
    .A(_13090_));
 sg13g2_a21oi_1 _39041_ (.A1(_13090_),
    .A2(_13091_),
    .Y(_13093_),
    .B1(net4646));
 sg13g2_a221oi_1 _39042_ (.B2(_13093_),
    .C1(net4352),
    .B1(_13092_),
    .A1(net4646),
    .Y(_13094_),
    .A2(_13089_));
 sg13g2_o21ai_1 _39043_ (.B1(net5591),
    .Y(_13095_),
    .A1(net4387),
    .A2(_13073_));
 sg13g2_o21ai_1 _39044_ (.B1(_13085_),
    .Y(_01000_),
    .A1(_13094_),
    .A2(_13095_));
 sg13g2_o21ai_1 _39045_ (.B1(_06797_),
    .Y(_13096_),
    .A1(_06799_),
    .A2(_13087_));
 sg13g2_a21oi_1 _39046_ (.A1(_06803_),
    .A2(_06806_),
    .Y(_13097_),
    .B1(net5392));
 sg13g2_xnor2_1 _39047_ (.Y(_13098_),
    .A(_06809_),
    .B(_13096_));
 sg13g2_a21oi_2 _39048_ (.B1(_13097_),
    .Y(_13099_),
    .A2(_13098_),
    .A1(net5392));
 sg13g2_and2_1 _39049_ (.A(net4579),
    .B(_13099_),
    .X(_13100_));
 sg13g2_xnor2_1 _39050_ (.Y(_13101_),
    .A(net4535),
    .B(_13099_));
 sg13g2_nor4_1 _39051_ (.A(_13074_),
    .B(_13075_),
    .C(_13077_),
    .D(_13090_),
    .Y(_13102_));
 sg13g2_a21oi_1 _39052_ (.A1(net4580),
    .A2(_13089_),
    .Y(_13103_),
    .B1(_13074_));
 sg13g2_nor2b_1 _39053_ (.A(_13102_),
    .B_N(_13103_),
    .Y(_13104_));
 sg13g2_nand2b_1 _39054_ (.Y(_13105_),
    .B(_13103_),
    .A_N(_13102_));
 sg13g2_nand2_1 _39055_ (.Y(_13106_),
    .A(_13037_),
    .B(_13061_));
 sg13g2_nor3_1 _39056_ (.A(_13076_),
    .B(_13090_),
    .C(_13106_),
    .Y(_13107_));
 sg13g2_a21oi_1 _39057_ (.A1(_13048_),
    .A2(_13107_),
    .Y(_13108_),
    .B1(_13105_));
 sg13g2_nor2b_1 _39058_ (.A(_13108_),
    .B_N(_13101_),
    .Y(_13109_));
 sg13g2_xor2_1 _39059_ (.B(_13108_),
    .A(_13101_),
    .X(_13110_));
 sg13g2_nand2_1 _39060_ (.Y(_13111_),
    .A(net4688),
    .B(_13110_));
 sg13g2_o21ai_1 _39061_ (.B1(_13111_),
    .Y(_13112_),
    .A1(net4688),
    .A2(_13099_));
 sg13g2_o21ai_1 _39062_ (.B1(net5591),
    .Y(_13113_),
    .A1(net4387),
    .A2(_13089_));
 sg13g2_a21oi_1 _39063_ (.A1(net4386),
    .A2(_13112_),
    .Y(_13114_),
    .B1(_13113_));
 sg13g2_a21o_1 _39064_ (.A2(net4126),
    .A1(net3226),
    .B1(_13114_),
    .X(_01001_));
 sg13g2_o21ai_1 _39065_ (.B1(_07242_),
    .Y(_13115_),
    .A1(_06799_),
    .A2(_13087_));
 sg13g2_nand2_1 _39066_ (.Y(_13116_),
    .A(_06808_),
    .B(_13115_));
 sg13g2_or2_1 _39067_ (.X(_13117_),
    .B(_13116_),
    .A(_06789_));
 sg13g2_a21oi_1 _39068_ (.A1(_06789_),
    .A2(_13116_),
    .Y(_13118_),
    .B1(net5348));
 sg13g2_a22oi_1 _39069_ (.Y(_13119_),
    .B1(_13117_),
    .B2(_13118_),
    .A2(_06787_),
    .A1(net5348));
 sg13g2_nor2_1 _39070_ (.A(net4535),
    .B(_13119_),
    .Y(_13120_));
 sg13g2_nand2_1 _39071_ (.Y(_13121_),
    .A(net4535),
    .B(_13119_));
 sg13g2_xnor2_1 _39072_ (.Y(_13122_),
    .A(net4579),
    .B(_13119_));
 sg13g2_nor2_1 _39073_ (.A(_13100_),
    .B(_13109_),
    .Y(_13123_));
 sg13g2_xnor2_1 _39074_ (.Y(_13124_),
    .A(_13122_),
    .B(_13123_));
 sg13g2_nor2_1 _39075_ (.A(net4688),
    .B(_13119_),
    .Y(_13125_));
 sg13g2_a21oi_1 _39076_ (.A1(net4688),
    .A2(_13124_),
    .Y(_13126_),
    .B1(_13125_));
 sg13g2_o21ai_1 _39077_ (.B1(net5591),
    .Y(_13127_),
    .A1(net4386),
    .A2(_13099_));
 sg13g2_a21oi_1 _39078_ (.A1(net4386),
    .A2(_13126_),
    .Y(_13128_),
    .B1(_13127_));
 sg13g2_a21o_1 _39079_ (.A2(net4126),
    .A1(net2649),
    .B1(_13128_),
    .X(_01002_));
 sg13g2_a21oi_1 _39080_ (.A1(_06770_),
    .A2(_06778_),
    .Y(_13129_),
    .B1(net5392));
 sg13g2_o21ai_1 _39081_ (.B1(_06788_),
    .Y(_13130_),
    .A1(_06789_),
    .A2(_13116_));
 sg13g2_xnor2_1 _39082_ (.Y(_13131_),
    .A(_06781_),
    .B(_13130_));
 sg13g2_a21oi_2 _39083_ (.B1(_13129_),
    .Y(_13132_),
    .A2(_13131_),
    .A1(net5392));
 sg13g2_xnor2_1 _39084_ (.Y(_13133_),
    .A(net4535),
    .B(_13132_));
 sg13g2_nor2_1 _39085_ (.A(_13100_),
    .B(_13120_),
    .Y(_13134_));
 sg13g2_nand2b_1 _39086_ (.Y(_13135_),
    .B(_13134_),
    .A_N(_13109_));
 sg13g2_and3_1 _39087_ (.X(_13136_),
    .A(_13121_),
    .B(_13133_),
    .C(_13135_));
 sg13g2_a21oi_1 _39088_ (.A1(_13121_),
    .A2(_13135_),
    .Y(_13137_),
    .B1(_13133_));
 sg13g2_nand2b_1 _39089_ (.Y(_13138_),
    .B(net4688),
    .A_N(_13137_));
 sg13g2_a21oi_1 _39090_ (.A1(net4646),
    .A2(_13132_),
    .Y(_13139_),
    .B1(net4352));
 sg13g2_o21ai_1 _39091_ (.B1(_13139_),
    .Y(_13140_),
    .A1(_13136_),
    .A2(_13138_));
 sg13g2_a21oi_1 _39092_ (.A1(net4352),
    .A2(_13119_),
    .Y(_13141_),
    .B1(net5528));
 sg13g2_a22oi_1 _39093_ (.Y(_13142_),
    .B1(_13140_),
    .B2(_13141_),
    .A2(net4126),
    .A1(net2628));
 sg13g2_inv_1 _39094_ (.Y(_01003_),
    .A(_13142_));
 sg13g2_nand2_1 _39095_ (.Y(_13143_),
    .A(net2901),
    .B(net4126));
 sg13g2_nand2_1 _39096_ (.Y(_13144_),
    .A(net5346),
    .B(_06756_));
 sg13g2_nand2_1 _39097_ (.Y(_13145_),
    .A(_06855_),
    .B(_13021_));
 sg13g2_and2_1 _39098_ (.A(_07244_),
    .B(_13145_),
    .X(_13146_));
 sg13g2_nor2_1 _39099_ (.A(_06758_),
    .B(_13146_),
    .Y(_13147_));
 sg13g2_xnor2_1 _39100_ (.Y(_13148_),
    .A(_06758_),
    .B(_13146_));
 sg13g2_o21ai_1 _39101_ (.B1(_13144_),
    .Y(_13149_),
    .A1(net5346),
    .A2(_13148_));
 sg13g2_xnor2_1 _39102_ (.Y(_13150_),
    .A(net4535),
    .B(_13149_));
 sg13g2_a21oi_1 _39103_ (.A1(net4579),
    .A2(_13132_),
    .Y(_13151_),
    .B1(_13136_));
 sg13g2_xnor2_1 _39104_ (.Y(_13152_),
    .A(_13150_),
    .B(_13151_));
 sg13g2_a21o_1 _39105_ (.A2(_13149_),
    .A1(net4651),
    .B1(net4353),
    .X(_13153_));
 sg13g2_a21oi_1 _39106_ (.A1(net4688),
    .A2(_13152_),
    .Y(_13154_),
    .B1(_13153_));
 sg13g2_o21ai_1 _39107_ (.B1(net5591),
    .Y(_13155_),
    .A1(net4386),
    .A2(_13132_));
 sg13g2_o21ai_1 _39108_ (.B1(_13143_),
    .Y(_01004_),
    .A1(_13154_),
    .A2(_13155_));
 sg13g2_nand2_1 _39109_ (.Y(_13156_),
    .A(net5346),
    .B(_06749_));
 sg13g2_a21oi_1 _39110_ (.A1(net4733),
    .A2(_06756_),
    .Y(_13157_),
    .B1(_13147_));
 sg13g2_xnor2_1 _39111_ (.Y(_13158_),
    .A(_06751_),
    .B(_13157_));
 sg13g2_o21ai_1 _39112_ (.B1(_13156_),
    .Y(_13159_),
    .A1(net5346),
    .A2(_13158_));
 sg13g2_nand2_1 _39113_ (.Y(_13160_),
    .A(net4644),
    .B(_13159_));
 sg13g2_xnor2_1 _39114_ (.Y(_13161_),
    .A(net4533),
    .B(_13159_));
 sg13g2_nand2_1 _39115_ (.Y(_13162_),
    .A(_13101_),
    .B(_13122_));
 sg13g2_o21ai_1 _39116_ (.B1(_13134_),
    .Y(_13163_),
    .A1(_13104_),
    .A2(_13162_));
 sg13g2_nand3_1 _39117_ (.B(_13150_),
    .C(_13163_),
    .A(_13133_),
    .Y(_13164_));
 sg13g2_o21ai_1 _39118_ (.B1(net4579),
    .Y(_13165_),
    .A1(_13132_),
    .A2(_13149_));
 sg13g2_nand2_2 _39119_ (.Y(_13166_),
    .A(_13164_),
    .B(_13165_));
 sg13g2_nand3_1 _39120_ (.B(_13133_),
    .C(_13150_),
    .A(_13107_),
    .Y(_13167_));
 sg13g2_nor2_2 _39121_ (.A(_13162_),
    .B(_13167_),
    .Y(_13168_));
 sg13g2_a21oi_2 _39122_ (.B1(_13166_),
    .Y(_13169_),
    .A2(_13168_),
    .A1(_13048_));
 sg13g2_or2_1 _39123_ (.X(_13170_),
    .B(_13169_),
    .A(_13161_));
 sg13g2_xor2_1 _39124_ (.B(_13169_),
    .A(_13161_),
    .X(_13171_));
 sg13g2_o21ai_1 _39125_ (.B1(_13160_),
    .Y(_13172_),
    .A1(net4644),
    .A2(_13171_));
 sg13g2_o21ai_1 _39126_ (.B1(net5591),
    .Y(_13173_),
    .A1(net4386),
    .A2(_13149_));
 sg13g2_a21oi_1 _39127_ (.A1(net4386),
    .A2(_13172_),
    .Y(_13174_),
    .B1(_13173_));
 sg13g2_a21o_1 _39128_ (.A2(net4126),
    .A1(net2573),
    .B1(_13174_),
    .X(_01005_));
 sg13g2_nand2_1 _39129_ (.Y(_13175_),
    .A(net2791),
    .B(net4126));
 sg13g2_o21ai_1 _39130_ (.B1(_06750_),
    .Y(_13176_),
    .A1(_07246_),
    .A2(_13147_));
 sg13g2_xnor2_1 _39131_ (.Y(_13177_),
    .A(_06739_),
    .B(_13176_));
 sg13g2_mux2_1 _39132_ (.A0(_06737_),
    .A1(_13177_),
    .S(net5388),
    .X(_13178_));
 sg13g2_xnor2_1 _39133_ (.Y(_13179_),
    .A(net4533),
    .B(_13178_));
 sg13g2_o21ai_1 _39134_ (.B1(_13170_),
    .Y(_13180_),
    .A1(net4533),
    .A2(_13159_));
 sg13g2_xor2_1 _39135_ (.B(_13180_),
    .A(_13179_),
    .X(_13181_));
 sg13g2_nor2_1 _39136_ (.A(net4644),
    .B(_13181_),
    .Y(_13182_));
 sg13g2_o21ai_1 _39137_ (.B1(net4383),
    .Y(_13183_),
    .A1(net4687),
    .A2(_13178_));
 sg13g2_a21oi_1 _39138_ (.A1(net4352),
    .A2(_13159_),
    .Y(_13184_),
    .B1(net5527));
 sg13g2_o21ai_1 _39139_ (.B1(_13184_),
    .Y(_13185_),
    .A1(_13182_),
    .A2(_13183_));
 sg13g2_nand2_1 _39140_ (.Y(_01006_),
    .A(_13175_),
    .B(_13185_));
 sg13g2_a21oi_1 _39141_ (.A1(_06725_),
    .A2(_06729_),
    .Y(_13186_),
    .B1(net5389));
 sg13g2_o21ai_1 _39142_ (.B1(_06738_),
    .Y(_13187_),
    .A1(_06739_),
    .A2(_13176_));
 sg13g2_xnor2_1 _39143_ (.Y(_13188_),
    .A(_06732_),
    .B(_13187_));
 sg13g2_a21oi_2 _39144_ (.B1(_13186_),
    .Y(_13189_),
    .A2(_13188_),
    .A1(net5389));
 sg13g2_nand2_1 _39145_ (.Y(_13190_),
    .A(net4578),
    .B(_13189_));
 sg13g2_inv_1 _39146_ (.Y(_13191_),
    .A(_13190_));
 sg13g2_xnor2_1 _39147_ (.Y(_13192_),
    .A(net4578),
    .B(_13189_));
 sg13g2_a21oi_1 _39148_ (.A1(_13159_),
    .A2(_13178_),
    .Y(_13193_),
    .B1(net4533));
 sg13g2_inv_1 _39149_ (.Y(_13194_),
    .A(_13193_));
 sg13g2_a22oi_1 _39150_ (.Y(_13195_),
    .B1(_13194_),
    .B2(_13170_),
    .A2(_13178_),
    .A1(net4533));
 sg13g2_nor2b_1 _39151_ (.A(_13192_),
    .B_N(_13195_),
    .Y(_13196_));
 sg13g2_xnor2_1 _39152_ (.Y(_13197_),
    .A(_13192_),
    .B(_13195_));
 sg13g2_nand2_1 _39153_ (.Y(_13198_),
    .A(net4687),
    .B(_13197_));
 sg13g2_nand2_1 _39154_ (.Y(_13199_),
    .A(net4644),
    .B(_13189_));
 sg13g2_nand3_1 _39155_ (.B(_13198_),
    .C(_13199_),
    .A(net4383),
    .Y(_13200_));
 sg13g2_a21oi_1 _39156_ (.A1(net4350),
    .A2(_13178_),
    .Y(_13201_),
    .B1(net5527));
 sg13g2_a22oi_1 _39157_ (.Y(_13202_),
    .B1(_13200_),
    .B2(_13201_),
    .A2(net4124),
    .A1(net2571));
 sg13g2_inv_1 _39158_ (.Y(_01007_),
    .A(_13202_));
 sg13g2_nand2_1 _39159_ (.Y(_13203_),
    .A(net2378),
    .B(net4124));
 sg13g2_nand2_1 _39160_ (.Y(_13204_),
    .A(net5345),
    .B(_06716_));
 sg13g2_o21ai_1 _39161_ (.B1(_07248_),
    .Y(_13205_),
    .A1(_06760_),
    .A2(_13146_));
 sg13g2_nand2b_1 _39162_ (.Y(_13206_),
    .B(_13205_),
    .A_N(_06718_));
 sg13g2_xor2_1 _39163_ (.B(_13205_),
    .A(_06718_),
    .X(_13207_));
 sg13g2_o21ai_1 _39164_ (.B1(_13204_),
    .Y(_13208_),
    .A1(net5345),
    .A2(_13207_));
 sg13g2_nand2_1 _39165_ (.Y(_13209_),
    .A(net4577),
    .B(_13208_));
 sg13g2_xnor2_1 _39166_ (.Y(_13210_),
    .A(net4532),
    .B(_13208_));
 sg13g2_inv_1 _39167_ (.Y(_13211_),
    .A(_13210_));
 sg13g2_o21ai_1 _39168_ (.B1(_13210_),
    .Y(_13212_),
    .A1(_13191_),
    .A2(_13196_));
 sg13g2_nor3_1 _39169_ (.A(_13191_),
    .B(_13196_),
    .C(_13210_),
    .Y(_13213_));
 sg13g2_nor2_1 _39170_ (.A(net4645),
    .B(_13213_),
    .Y(_13214_));
 sg13g2_a221oi_1 _39171_ (.B2(_13214_),
    .C1(net4350),
    .B1(_13212_),
    .A1(net4643),
    .Y(_13215_),
    .A2(_13208_));
 sg13g2_o21ai_1 _39172_ (.B1(net5589),
    .Y(_13216_),
    .A1(net4383),
    .A2(_13189_));
 sg13g2_o21ai_1 _39173_ (.B1(_13203_),
    .Y(_01008_),
    .A1(_13215_),
    .A2(_13216_));
 sg13g2_a21oi_1 _39174_ (.A1(_06704_),
    .A2(_06708_),
    .Y(_13217_),
    .B1(net5388));
 sg13g2_nor2b_1 _39175_ (.A(_06717_),
    .B_N(_13206_),
    .Y(_13218_));
 sg13g2_xnor2_1 _39176_ (.Y(_13219_),
    .A(_06711_),
    .B(_13218_));
 sg13g2_a21oi_2 _39177_ (.B1(_13217_),
    .Y(_13220_),
    .A2(_13219_),
    .A1(net5388));
 sg13g2_nand2_1 _39178_ (.Y(_13221_),
    .A(net4577),
    .B(_13220_));
 sg13g2_xnor2_1 _39179_ (.Y(_13222_),
    .A(net4532),
    .B(_13220_));
 sg13g2_nand3b_1 _39180_ (.B(_13193_),
    .C(_13210_),
    .Y(_13223_),
    .A_N(_13192_));
 sg13g2_nand3_1 _39181_ (.B(_13209_),
    .C(_13223_),
    .A(_13190_),
    .Y(_13224_));
 sg13g2_nor4_1 _39182_ (.A(_13161_),
    .B(_13179_),
    .C(_13192_),
    .D(_13211_),
    .Y(_13225_));
 sg13g2_nor2b_1 _39183_ (.A(_13169_),
    .B_N(_13225_),
    .Y(_13226_));
 sg13g2_o21ai_1 _39184_ (.B1(_13222_),
    .Y(_13227_),
    .A1(_13224_),
    .A2(_13226_));
 sg13g2_or3_1 _39185_ (.A(_13222_),
    .B(_13224_),
    .C(_13226_),
    .X(_13228_));
 sg13g2_nand3_1 _39186_ (.B(_13227_),
    .C(_13228_),
    .A(net4687),
    .Y(_13229_));
 sg13g2_a21oi_1 _39187_ (.A1(net4644),
    .A2(_13220_),
    .Y(_13230_),
    .B1(net4350));
 sg13g2_o21ai_1 _39188_ (.B1(net5589),
    .Y(_13231_),
    .A1(net4382),
    .A2(_13208_));
 sg13g2_a21oi_1 _39189_ (.A1(_13229_),
    .A2(_13230_),
    .Y(_13232_),
    .B1(_13231_));
 sg13g2_a21o_1 _39190_ (.A2(net4123),
    .A1(net2485),
    .B1(_13232_),
    .X(_01009_));
 sg13g2_nand2_1 _39191_ (.Y(_13233_),
    .A(net3210),
    .B(net4123));
 sg13g2_nand2_1 _39192_ (.Y(_13234_),
    .A(net5345),
    .B(_06683_));
 sg13g2_a21oi_1 _39193_ (.A1(_07250_),
    .A2(_13206_),
    .Y(_13235_),
    .B1(_06710_));
 sg13g2_xnor2_1 _39194_ (.Y(_13236_),
    .A(_06685_),
    .B(_13235_));
 sg13g2_o21ai_1 _39195_ (.B1(_13234_),
    .Y(_13237_),
    .A1(net5345),
    .A2(_13236_));
 sg13g2_inv_1 _39196_ (.Y(_13238_),
    .A(_13237_));
 sg13g2_xnor2_1 _39197_ (.Y(_13239_),
    .A(net4531),
    .B(_13237_));
 sg13g2_nand2_1 _39198_ (.Y(_13240_),
    .A(_13221_),
    .B(_13227_));
 sg13g2_xnor2_1 _39199_ (.Y(_13241_),
    .A(_13239_),
    .B(_13240_));
 sg13g2_a21oi_1 _39200_ (.A1(net4643),
    .A2(_13237_),
    .Y(_13242_),
    .B1(net4350));
 sg13g2_o21ai_1 _39201_ (.B1(_13242_),
    .Y(_13243_),
    .A1(net4643),
    .A2(_13241_));
 sg13g2_o21ai_1 _39202_ (.B1(_13243_),
    .Y(_13244_),
    .A1(net4383),
    .A2(_13220_));
 sg13g2_o21ai_1 _39203_ (.B1(_13233_),
    .Y(_01010_),
    .A1(net5527),
    .A2(_13244_));
 sg13g2_nand2_1 _39204_ (.Y(_13245_),
    .A(net2603),
    .B(net4123));
 sg13g2_a21oi_1 _39205_ (.A1(_06685_),
    .A2(_13235_),
    .Y(_13246_),
    .B1(_06684_));
 sg13g2_xor2_1 _39206_ (.B(_13246_),
    .A(_06698_),
    .X(_13247_));
 sg13g2_mux2_1 _39207_ (.A0(_06695_),
    .A1(_13247_),
    .S(net5388),
    .X(_13248_));
 sg13g2_and2_1 _39208_ (.A(net4577),
    .B(_13248_),
    .X(_13249_));
 sg13g2_xnor2_1 _39209_ (.Y(_13250_),
    .A(net4577),
    .B(_13248_));
 sg13g2_o21ai_1 _39210_ (.B1(net4577),
    .Y(_13251_),
    .A1(_13220_),
    .A2(_13237_));
 sg13g2_a22oi_1 _39211_ (.Y(_13252_),
    .B1(_13251_),
    .B2(_13227_),
    .A2(_13238_),
    .A1(net4531));
 sg13g2_a221oi_1 _39212_ (.B2(_13227_),
    .C1(_13250_),
    .B1(_13251_),
    .A1(net4532),
    .Y(_13253_),
    .A2(_13238_));
 sg13g2_xnor2_1 _39213_ (.Y(_13254_),
    .A(_13250_),
    .B(_13252_));
 sg13g2_a21o_1 _39214_ (.A2(_13248_),
    .A1(net4643),
    .B1(net4350),
    .X(_13255_));
 sg13g2_a21oi_1 _39215_ (.A1(net4687),
    .A2(_13254_),
    .Y(_13256_),
    .B1(_13255_));
 sg13g2_o21ai_1 _39216_ (.B1(net5589),
    .Y(_13257_),
    .A1(net4382),
    .A2(_13237_));
 sg13g2_o21ai_1 _39217_ (.B1(_13245_),
    .Y(_01011_),
    .A1(_13256_),
    .A2(_13257_));
 sg13g2_nand2_1 _39218_ (.Y(_13258_),
    .A(net2294),
    .B(net4123));
 sg13g2_nand2_1 _39219_ (.Y(_13259_),
    .A(net5345),
    .B(_06649_));
 sg13g2_a21oi_1 _39220_ (.A1(_06856_),
    .A2(_13021_),
    .Y(_13260_),
    .B1(_07253_));
 sg13g2_a21o_2 _39221_ (.A2(_13021_),
    .A1(_06856_),
    .B1(_07253_),
    .X(_13261_));
 sg13g2_nand2_1 _39222_ (.Y(_13262_),
    .A(_06651_),
    .B(_13261_));
 sg13g2_xnor2_1 _39223_ (.Y(_13263_),
    .A(_06651_),
    .B(_13261_));
 sg13g2_o21ai_1 _39224_ (.B1(_13259_),
    .Y(_13264_),
    .A1(net5345),
    .A2(_13263_));
 sg13g2_xnor2_1 _39225_ (.Y(_13265_),
    .A(net4532),
    .B(_13264_));
 sg13g2_nor3_1 _39226_ (.A(_13249_),
    .B(_13253_),
    .C(_13265_),
    .Y(_13266_));
 sg13g2_o21ai_1 _39227_ (.B1(_13265_),
    .Y(_13267_),
    .A1(_13249_),
    .A2(_13253_));
 sg13g2_nor2_1 _39228_ (.A(net4644),
    .B(_13266_),
    .Y(_13268_));
 sg13g2_a221oi_1 _39229_ (.B2(_13268_),
    .C1(net4350),
    .B1(_13267_),
    .A1(net4644),
    .Y(_13269_),
    .A2(_13264_));
 sg13g2_o21ai_1 _39230_ (.B1(net5589),
    .Y(_13270_),
    .A1(net4383),
    .A2(_13248_));
 sg13g2_o21ai_1 _39231_ (.B1(_13258_),
    .Y(_01012_),
    .A1(_13269_),
    .A2(_13270_));
 sg13g2_nand2_1 _39232_ (.Y(_13271_),
    .A(net5345),
    .B(_06660_));
 sg13g2_o21ai_1 _39233_ (.B1(_13262_),
    .Y(_13272_),
    .A1(net4789),
    .A2(_06650_));
 sg13g2_xor2_1 _39234_ (.B(_13272_),
    .A(_06662_),
    .X(_13273_));
 sg13g2_o21ai_1 _39235_ (.B1(_13271_),
    .Y(_13274_),
    .A1(net5345),
    .A2(_13273_));
 sg13g2_nand2_1 _39236_ (.Y(_13275_),
    .A(net4643),
    .B(_13274_));
 sg13g2_or2_1 _39237_ (.X(_13276_),
    .B(_13274_),
    .A(net4531));
 sg13g2_xnor2_1 _39238_ (.Y(_13277_),
    .A(net4531),
    .B(_13274_));
 sg13g2_inv_1 _39239_ (.Y(_13278_),
    .A(_13277_));
 sg13g2_nor2b_1 _39240_ (.A(_13250_),
    .B_N(_13265_),
    .Y(_13279_));
 sg13g2_and2_1 _39241_ (.A(_13222_),
    .B(_13239_),
    .X(_13280_));
 sg13g2_nand2_1 _39242_ (.Y(_13281_),
    .A(_13224_),
    .B(_13280_));
 sg13g2_nand3_1 _39243_ (.B(_13225_),
    .C(_13280_),
    .A(_13166_),
    .Y(_13282_));
 sg13g2_nand3_1 _39244_ (.B(_13281_),
    .C(_13282_),
    .A(_13251_),
    .Y(_13283_));
 sg13g2_a21o_1 _39245_ (.A2(_13264_),
    .A1(net4578),
    .B1(_13249_),
    .X(_13284_));
 sg13g2_a21o_1 _39246_ (.A2(_13283_),
    .A1(_13279_),
    .B1(_13284_),
    .X(_13285_));
 sg13g2_and4_1 _39247_ (.A(_13168_),
    .B(_13225_),
    .C(_13279_),
    .D(_13280_),
    .X(_13286_));
 sg13g2_a21oi_2 _39248_ (.B1(_13285_),
    .Y(_13287_),
    .A2(_13286_),
    .A1(_13048_));
 sg13g2_xnor2_1 _39249_ (.Y(_13288_),
    .A(_13278_),
    .B(_13287_));
 sg13g2_o21ai_1 _39250_ (.B1(_13275_),
    .Y(_13289_),
    .A1(net4643),
    .A2(_13288_));
 sg13g2_o21ai_1 _39251_ (.B1(net5589),
    .Y(_13290_),
    .A1(net4382),
    .A2(_13264_));
 sg13g2_a21oi_1 _39252_ (.A1(net4382),
    .A2(_13289_),
    .Y(_13291_),
    .B1(_13290_));
 sg13g2_a21o_1 _39253_ (.A2(net4123),
    .A1(net3022),
    .B1(_13291_),
    .X(_01013_));
 sg13g2_nand2_1 _39254_ (.Y(_13292_),
    .A(net2669),
    .B(net4123));
 sg13g2_nor2_1 _39255_ (.A(net5388),
    .B(_06627_),
    .Y(_13293_));
 sg13g2_a21o_1 _39256_ (.A2(_13262_),
    .A1(_07255_),
    .B1(_06661_),
    .X(_13294_));
 sg13g2_xor2_1 _39257_ (.B(_13294_),
    .A(_06630_),
    .X(_13295_));
 sg13g2_a21oi_2 _39258_ (.B1(_13293_),
    .Y(_13296_),
    .A2(_13295_),
    .A1(net5388));
 sg13g2_nand2_1 _39259_ (.Y(_13297_),
    .A(net4531),
    .B(_13296_));
 sg13g2_xnor2_1 _39260_ (.Y(_13298_),
    .A(net4577),
    .B(_13296_));
 sg13g2_o21ai_1 _39261_ (.B1(_13276_),
    .Y(_13299_),
    .A1(_13277_),
    .A2(_13287_));
 sg13g2_xnor2_1 _39262_ (.Y(_13300_),
    .A(_13298_),
    .B(_13299_));
 sg13g2_and2_1 _39263_ (.A(net4643),
    .B(_13296_),
    .X(_13301_));
 sg13g2_a21oi_1 _39264_ (.A1(net4687),
    .A2(_13300_),
    .Y(_13302_),
    .B1(_13301_));
 sg13g2_nor2_1 _39265_ (.A(net4382),
    .B(_13274_),
    .Y(_13303_));
 sg13g2_a21oi_1 _39266_ (.A1(net4382),
    .A2(_13302_),
    .Y(_13304_),
    .B1(_13303_));
 sg13g2_o21ai_1 _39267_ (.B1(_13292_),
    .Y(_01014_),
    .A1(net5527),
    .A2(_13304_));
 sg13g2_a21oi_1 _39268_ (.A1(_06633_),
    .A2(_06638_),
    .Y(_13305_),
    .B1(net5388));
 sg13g2_o21ai_1 _39269_ (.B1(_06628_),
    .Y(_13306_),
    .A1(_06630_),
    .A2(_13294_));
 sg13g2_xnor2_1 _39270_ (.Y(_13307_),
    .A(_06641_),
    .B(_13306_));
 sg13g2_a21oi_2 _39271_ (.B1(_13305_),
    .Y(_13308_),
    .A2(_13307_),
    .A1(net5388));
 sg13g2_nand2_1 _39272_ (.Y(_13309_),
    .A(net4577),
    .B(_13308_));
 sg13g2_xnor2_1 _39273_ (.Y(_13310_),
    .A(net4531),
    .B(_13308_));
 sg13g2_a21o_1 _39274_ (.A2(_13296_),
    .A1(_13274_),
    .B1(net4531),
    .X(_13311_));
 sg13g2_o21ai_1 _39275_ (.B1(_13311_),
    .Y(_13312_),
    .A1(_13277_),
    .A2(_13287_));
 sg13g2_nand3_1 _39276_ (.B(_13310_),
    .C(_13312_),
    .A(_13297_),
    .Y(_13313_));
 sg13g2_a21o_1 _39277_ (.A2(_13312_),
    .A1(_13297_),
    .B1(_13310_),
    .X(_13314_));
 sg13g2_nand3_1 _39278_ (.B(_13313_),
    .C(_13314_),
    .A(net4687),
    .Y(_13315_));
 sg13g2_a21oi_1 _39279_ (.A1(net4643),
    .A2(_13308_),
    .Y(_13316_),
    .B1(net4350));
 sg13g2_a221oi_1 _39280_ (.B2(_13316_),
    .C1(net5527),
    .B1(_13315_),
    .A1(net4350),
    .Y(_13317_),
    .A2(_13296_));
 sg13g2_a21oi_1 _39281_ (.A1(net2236),
    .A2(net4123),
    .Y(_13318_),
    .B1(_13317_));
 sg13g2_inv_1 _39282_ (.Y(_01015_),
    .A(_13318_));
 sg13g2_nor2_1 _39283_ (.A(net5387),
    .B(_06603_),
    .Y(_13319_));
 sg13g2_nor2_1 _39284_ (.A(_06663_),
    .B(_13260_),
    .Y(_13320_));
 sg13g2_nor2b_1 _39285_ (.A(_13320_),
    .B_N(_07257_),
    .Y(_13321_));
 sg13g2_xor2_1 _39286_ (.B(_13321_),
    .A(_06606_),
    .X(_13322_));
 sg13g2_a21oi_2 _39287_ (.B1(_13319_),
    .Y(_13323_),
    .A2(_13322_),
    .A1(net5387));
 sg13g2_xnor2_1 _39288_ (.Y(_13324_),
    .A(net4577),
    .B(_13323_));
 sg13g2_nand2_1 _39289_ (.Y(_13325_),
    .A(_13309_),
    .B(_13313_));
 sg13g2_xor2_1 _39290_ (.B(_13325_),
    .A(_13324_),
    .X(_13326_));
 sg13g2_nor2_1 _39291_ (.A(net4687),
    .B(_13323_),
    .Y(_13327_));
 sg13g2_a21oi_1 _39292_ (.A1(net4687),
    .A2(_13326_),
    .Y(_13328_),
    .B1(_13327_));
 sg13g2_o21ai_1 _39293_ (.B1(net5588),
    .Y(_13329_),
    .A1(net4382),
    .A2(_13308_));
 sg13g2_a21oi_1 _39294_ (.A1(net4382),
    .A2(_13328_),
    .Y(_13330_),
    .B1(_13329_));
 sg13g2_a21o_1 _39295_ (.A2(net4123),
    .A1(net2476),
    .B1(_13330_),
    .X(_01016_));
 sg13g2_nor2_1 _39296_ (.A(net5387),
    .B(_06615_),
    .Y(_13331_));
 sg13g2_o21ai_1 _39297_ (.B1(_06605_),
    .Y(_13332_),
    .A1(_06606_),
    .A2(_13321_));
 sg13g2_xor2_1 _39298_ (.B(_13332_),
    .A(_06618_),
    .X(_13333_));
 sg13g2_a21oi_2 _39299_ (.B1(_13331_),
    .Y(_13334_),
    .A2(_13333_),
    .A1(net5387));
 sg13g2_nand2_1 _39300_ (.Y(_13335_),
    .A(net4575),
    .B(_13334_));
 sg13g2_xnor2_1 _39301_ (.Y(_13336_),
    .A(net4575),
    .B(_13334_));
 sg13g2_nand3b_1 _39302_ (.B(_13324_),
    .C(_13310_),
    .Y(_13337_),
    .A_N(_13311_));
 sg13g2_o21ai_1 _39303_ (.B1(_13309_),
    .Y(_13338_),
    .A1(net4531),
    .A2(_13323_));
 sg13g2_nor2b_2 _39304_ (.A(_13338_),
    .B_N(_13337_),
    .Y(_13339_));
 sg13g2_nand4_1 _39305_ (.B(_13298_),
    .C(_13310_),
    .A(_13278_),
    .Y(_13340_),
    .D(_13324_));
 sg13g2_o21ai_1 _39306_ (.B1(_13339_),
    .Y(_13341_),
    .A1(_13287_),
    .A2(_13340_));
 sg13g2_nand2b_2 _39307_ (.Y(_13342_),
    .B(_13341_),
    .A_N(_13336_));
 sg13g2_nand2b_1 _39308_ (.Y(_13343_),
    .B(_13336_),
    .A_N(_13341_));
 sg13g2_nand3_1 _39309_ (.B(_13342_),
    .C(_13343_),
    .A(net4686),
    .Y(_13344_));
 sg13g2_nand2_1 _39310_ (.Y(_13345_),
    .A(net4642),
    .B(_13334_));
 sg13g2_nand3_1 _39311_ (.B(_13344_),
    .C(_13345_),
    .A(net4380),
    .Y(_13346_));
 sg13g2_a21oi_1 _39312_ (.A1(net4351),
    .A2(_13323_),
    .Y(_13347_),
    .B1(net5527));
 sg13g2_a22oi_1 _39313_ (.Y(_13348_),
    .B1(_13346_),
    .B2(_13347_),
    .A2(net4122),
    .A1(net2917));
 sg13g2_inv_1 _39314_ (.Y(_01017_),
    .A(_13348_));
 sg13g2_a21oi_1 _39315_ (.A1(_06617_),
    .A2(_13332_),
    .Y(_13349_),
    .B1(_06616_));
 sg13g2_nor2_1 _39316_ (.A(_06597_),
    .B(_13349_),
    .Y(_13350_));
 sg13g2_a21oi_1 _39317_ (.A1(_06597_),
    .A2(_13349_),
    .Y(_13351_),
    .B1(net5344));
 sg13g2_nor2b_1 _39318_ (.A(_13350_),
    .B_N(_13351_),
    .Y(_13352_));
 sg13g2_a21oi_2 _39319_ (.B1(_13352_),
    .Y(_13353_),
    .A2(_06595_),
    .A1(net5344));
 sg13g2_nor2_1 _39320_ (.A(net4530),
    .B(_13353_),
    .Y(_13354_));
 sg13g2_xnor2_1 _39321_ (.Y(_13355_),
    .A(net4530),
    .B(_13353_));
 sg13g2_nand3_1 _39322_ (.B(_13342_),
    .C(_13355_),
    .A(_13335_),
    .Y(_13356_));
 sg13g2_a21oi_1 _39323_ (.A1(_13335_),
    .A2(_13342_),
    .Y(_13357_),
    .B1(_13355_));
 sg13g2_nor2_1 _39324_ (.A(net4642),
    .B(_13357_),
    .Y(_13358_));
 sg13g2_nor2_1 _39325_ (.A(net4686),
    .B(_13353_),
    .Y(_13359_));
 sg13g2_a21oi_1 _39326_ (.A1(_13356_),
    .A2(_13358_),
    .Y(_13360_),
    .B1(_13359_));
 sg13g2_o21ai_1 _39327_ (.B1(net5588),
    .Y(_13361_),
    .A1(net4380),
    .A2(_13334_));
 sg13g2_a21oi_1 _39328_ (.A1(net4380),
    .A2(_13360_),
    .Y(_13362_),
    .B1(_13361_));
 sg13g2_a21o_1 _39329_ (.A2(net4122),
    .A1(net1956),
    .B1(_13362_),
    .X(_01018_));
 sg13g2_nor2_1 _39330_ (.A(net5387),
    .B(_06587_),
    .Y(_13363_));
 sg13g2_nor2_1 _39331_ (.A(_06596_),
    .B(_13350_),
    .Y(_13364_));
 sg13g2_xnor2_1 _39332_ (.Y(_13365_),
    .A(_06589_),
    .B(_13364_));
 sg13g2_a21oi_2 _39333_ (.B1(_13363_),
    .Y(_13366_),
    .A2(_13365_),
    .A1(net5387));
 sg13g2_and2_1 _39334_ (.A(net4575),
    .B(_13366_),
    .X(_13367_));
 sg13g2_xnor2_1 _39335_ (.Y(_13368_),
    .A(net4576),
    .B(_13366_));
 sg13g2_a21oi_1 _39336_ (.A1(net4576),
    .A2(_13334_),
    .Y(_13369_),
    .B1(_13354_));
 sg13g2_a22oi_1 _39337_ (.Y(_13370_),
    .B1(_13369_),
    .B2(_13342_),
    .A2(_13353_),
    .A1(net4530));
 sg13g2_a221oi_1 _39338_ (.B2(_13342_),
    .C1(_13368_),
    .B1(_13369_),
    .A1(net4530),
    .Y(_13371_),
    .A2(_13353_));
 sg13g2_xor2_1 _39339_ (.B(_13370_),
    .A(_13368_),
    .X(_13372_));
 sg13g2_a21oi_1 _39340_ (.A1(net4642),
    .A2(_13366_),
    .Y(_13373_),
    .B1(net4351));
 sg13g2_o21ai_1 _39341_ (.B1(_13373_),
    .Y(_13374_),
    .A1(net4642),
    .A2(_13372_));
 sg13g2_a21oi_1 _39342_ (.A1(net4351),
    .A2(_13353_),
    .Y(_13375_),
    .B1(net5527));
 sg13g2_a22oi_1 _39343_ (.Y(_13376_),
    .B1(_13374_),
    .B2(_13375_),
    .A2(net4122),
    .A1(net2150));
 sg13g2_inv_1 _39344_ (.Y(_01019_),
    .A(_13376_));
 sg13g2_nand2_1 _39345_ (.Y(_13377_),
    .A(net2478),
    .B(net4122));
 sg13g2_nand2_1 _39346_ (.Y(_13378_),
    .A(net5343),
    .B(_06553_));
 sg13g2_a21oi_2 _39347_ (.B1(_07261_),
    .Y(_13379_),
    .A2(_13261_),
    .A1(_06664_));
 sg13g2_nor2_1 _39348_ (.A(_06555_),
    .B(_13379_),
    .Y(_13380_));
 sg13g2_xnor2_1 _39349_ (.Y(_13381_),
    .A(_06555_),
    .B(_13379_));
 sg13g2_o21ai_1 _39350_ (.B1(_13378_),
    .Y(_13382_),
    .A1(net5344),
    .A2(_13381_));
 sg13g2_xnor2_1 _39351_ (.Y(_13383_),
    .A(net4530),
    .B(_13382_));
 sg13g2_nor3_1 _39352_ (.A(_13367_),
    .B(_13371_),
    .C(_13383_),
    .Y(_13384_));
 sg13g2_o21ai_1 _39353_ (.B1(_13383_),
    .Y(_13385_),
    .A1(_13367_),
    .A2(_13371_));
 sg13g2_nor2_1 _39354_ (.A(net4642),
    .B(_13384_),
    .Y(_13386_));
 sg13g2_a221oi_1 _39355_ (.B2(_13386_),
    .C1(net4351),
    .B1(_13385_),
    .A1(net4642),
    .Y(_13387_),
    .A2(_13382_));
 sg13g2_o21ai_1 _39356_ (.B1(net5588),
    .Y(_13388_),
    .A1(net4380),
    .A2(_13366_));
 sg13g2_o21ai_1 _39357_ (.B1(_13377_),
    .Y(_01020_),
    .A1(_13387_),
    .A2(_13388_));
 sg13g2_o21ai_1 _39358_ (.B1(_06554_),
    .Y(_13389_),
    .A1(_06555_),
    .A2(_13379_));
 sg13g2_xnor2_1 _39359_ (.Y(_13390_),
    .A(_06565_),
    .B(_13389_));
 sg13g2_nor2_1 _39360_ (.A(net5343),
    .B(_13390_),
    .Y(_13391_));
 sg13g2_a21oi_2 _39361_ (.B1(_13391_),
    .Y(_13392_),
    .A2(_06563_),
    .A1(net5343));
 sg13g2_nand2_1 _39362_ (.Y(_13393_),
    .A(net4575),
    .B(_13392_));
 sg13g2_xnor2_1 _39363_ (.Y(_13394_),
    .A(net4575),
    .B(_13392_));
 sg13g2_nand2b_1 _39364_ (.Y(_13395_),
    .B(_13383_),
    .A_N(_13368_));
 sg13g2_or4_1 _39365_ (.A(_13336_),
    .B(_13340_),
    .C(_13355_),
    .D(_13395_),
    .X(_13396_));
 sg13g2_or3_1 _39366_ (.A(_13336_),
    .B(_13339_),
    .C(_13355_),
    .X(_13397_));
 sg13g2_a21oi_1 _39367_ (.A1(_13369_),
    .A2(_13397_),
    .Y(_13398_),
    .B1(_13395_));
 sg13g2_o21ai_1 _39368_ (.B1(net4576),
    .Y(_13399_),
    .A1(_13366_),
    .A2(_13382_));
 sg13g2_nor2b_1 _39369_ (.A(_13398_),
    .B_N(_13399_),
    .Y(_13400_));
 sg13g2_o21ai_1 _39370_ (.B1(_13400_),
    .Y(_13401_),
    .A1(_13287_),
    .A2(_13396_));
 sg13g2_nand2b_2 _39371_ (.Y(_13402_),
    .B(_13401_),
    .A_N(_13394_));
 sg13g2_nand2b_1 _39372_ (.Y(_13403_),
    .B(_13394_),
    .A_N(_13401_));
 sg13g2_a21o_1 _39373_ (.A2(_13403_),
    .A1(_13402_),
    .B1(net4642),
    .X(_13404_));
 sg13g2_o21ai_1 _39374_ (.B1(_13404_),
    .Y(_13405_),
    .A1(net4686),
    .A2(_13392_));
 sg13g2_o21ai_1 _39375_ (.B1(net5588),
    .Y(_13406_),
    .A1(net4380),
    .A2(_13382_));
 sg13g2_a21oi_1 _39376_ (.A1(net4380),
    .A2(_13405_),
    .Y(_13407_),
    .B1(_13406_));
 sg13g2_a21o_1 _39377_ (.A2(net4122),
    .A1(net3012),
    .B1(_13407_),
    .X(_01021_));
 sg13g2_nand2_1 _39378_ (.Y(_13408_),
    .A(net2902),
    .B(net4122));
 sg13g2_o21ai_1 _39379_ (.B1(_06564_),
    .Y(_13409_),
    .A1(_07263_),
    .A2(_13380_));
 sg13g2_xnor2_1 _39380_ (.Y(_13410_),
    .A(_06545_),
    .B(_13409_));
 sg13g2_nor2_1 _39381_ (.A(net5343),
    .B(_13410_),
    .Y(_13411_));
 sg13g2_a21oi_2 _39382_ (.B1(_13411_),
    .Y(_13412_),
    .A2(_06543_),
    .A1(net5343));
 sg13g2_nor2_1 _39383_ (.A(net4530),
    .B(_13412_),
    .Y(_13413_));
 sg13g2_xnor2_1 _39384_ (.Y(_13414_),
    .A(net4575),
    .B(_13412_));
 sg13g2_nand2_1 _39385_ (.Y(_13415_),
    .A(_13393_),
    .B(_13402_));
 sg13g2_xor2_1 _39386_ (.B(_13415_),
    .A(_13414_),
    .X(_13416_));
 sg13g2_o21ai_1 _39387_ (.B1(net4380),
    .Y(_13417_),
    .A1(net4686),
    .A2(_13412_));
 sg13g2_a21oi_1 _39388_ (.A1(net4686),
    .A2(_13416_),
    .Y(_13418_),
    .B1(_13417_));
 sg13g2_o21ai_1 _39389_ (.B1(net5588),
    .Y(_13419_),
    .A1(net4380),
    .A2(_13392_));
 sg13g2_o21ai_1 _39390_ (.B1(_13408_),
    .Y(_01022_),
    .A1(_13418_),
    .A2(_13419_));
 sg13g2_o21ai_1 _39391_ (.B1(_06544_),
    .Y(_13420_),
    .A1(_06545_),
    .A2(_13409_));
 sg13g2_xnor2_1 _39392_ (.Y(_13421_),
    .A(_06537_),
    .B(_13420_));
 sg13g2_nor2_1 _39393_ (.A(net5343),
    .B(_13421_),
    .Y(_13422_));
 sg13g2_a21o_1 _39394_ (.A2(_06536_),
    .A1(net5343),
    .B1(_13422_),
    .X(_13423_));
 sg13g2_a21oi_1 _39395_ (.A1(net5343),
    .A2(_06536_),
    .Y(_13424_),
    .B1(_13422_));
 sg13g2_nor2_1 _39396_ (.A(net4534),
    .B(_13423_),
    .Y(_13425_));
 sg13g2_xnor2_1 _39397_ (.Y(_13426_),
    .A(net4575),
    .B(_13423_));
 sg13g2_inv_1 _39398_ (.Y(_13427_),
    .A(_13426_));
 sg13g2_a21oi_1 _39399_ (.A1(net4575),
    .A2(_13392_),
    .Y(_13428_),
    .B1(_13413_));
 sg13g2_a22oi_1 _39400_ (.Y(_13429_),
    .B1(_13428_),
    .B2(_13402_),
    .A2(_13412_),
    .A1(net4530));
 sg13g2_a221oi_1 _39401_ (.B2(_13402_),
    .C1(_13427_),
    .B1(_13428_),
    .A1(net4530),
    .Y(_13430_),
    .A2(_13412_));
 sg13g2_o21ai_1 _39402_ (.B1(net4686),
    .Y(_13431_),
    .A1(_13426_),
    .A2(_13429_));
 sg13g2_a21oi_1 _39403_ (.A1(net4642),
    .A2(_13424_),
    .Y(_13432_),
    .B1(net4351));
 sg13g2_o21ai_1 _39404_ (.B1(_13432_),
    .Y(_13433_),
    .A1(_13430_),
    .A2(_13431_));
 sg13g2_a21oi_1 _39405_ (.A1(net4351),
    .A2(_13412_),
    .Y(_13434_),
    .B1(net5527));
 sg13g2_a22oi_1 _39406_ (.Y(_13435_),
    .B1(_13433_),
    .B2(_13434_),
    .A2(net4122),
    .A1(net2265));
 sg13g2_inv_1 _39407_ (.Y(_01023_),
    .A(_13435_));
 sg13g2_nand2_1 _39408_ (.Y(_13436_),
    .A(net2446),
    .B(net4122));
 sg13g2_nand2_1 _39409_ (.Y(_13437_),
    .A(net5347),
    .B(_06522_));
 sg13g2_o21ai_1 _39410_ (.B1(_07265_),
    .Y(_13438_),
    .A1(_06567_),
    .A2(_13379_));
 sg13g2_nand2_1 _39411_ (.Y(_13439_),
    .A(_06524_),
    .B(_13438_));
 sg13g2_xnor2_1 _39412_ (.Y(_13440_),
    .A(_06524_),
    .B(_13438_));
 sg13g2_o21ai_1 _39413_ (.B1(_13437_),
    .Y(_13441_),
    .A1(net5347),
    .A2(_13440_));
 sg13g2_xnor2_1 _39414_ (.Y(_13442_),
    .A(net4534),
    .B(_13441_));
 sg13g2_nor3_1 _39415_ (.A(_13425_),
    .B(_13430_),
    .C(_13442_),
    .Y(_13443_));
 sg13g2_o21ai_1 _39416_ (.B1(_13442_),
    .Y(_13444_),
    .A1(_13425_),
    .A2(_13430_));
 sg13g2_nor2_1 _39417_ (.A(net4645),
    .B(_13443_),
    .Y(_13445_));
 sg13g2_a221oi_1 _39418_ (.B2(_13445_),
    .C1(net4351),
    .B1(_13444_),
    .A1(net4645),
    .Y(_13446_),
    .A2(_13441_));
 sg13g2_o21ai_1 _39419_ (.B1(net5588),
    .Y(_13447_),
    .A1(net4381),
    .A2(_13424_));
 sg13g2_o21ai_1 _39420_ (.B1(_13436_),
    .Y(_01024_),
    .A1(_13446_),
    .A2(_13447_));
 sg13g2_nor2_1 _39421_ (.A(net5387),
    .B(_06515_),
    .Y(_13448_));
 sg13g2_nand2_1 _39422_ (.Y(_13449_),
    .A(_06523_),
    .B(_13439_));
 sg13g2_xnor2_1 _39423_ (.Y(_13450_),
    .A(_06517_),
    .B(_13449_));
 sg13g2_a21oi_2 _39424_ (.B1(_13448_),
    .Y(_13451_),
    .A2(_13450_),
    .A1(net5387));
 sg13g2_nand2_1 _39425_ (.Y(_13452_),
    .A(net4581),
    .B(_13451_));
 sg13g2_xnor2_1 _39426_ (.Y(_13453_),
    .A(net4576),
    .B(_13451_));
 sg13g2_nand2_1 _39427_ (.Y(_13454_),
    .A(_13426_),
    .B(_13442_));
 sg13g2_nand3_1 _39428_ (.B(_13426_),
    .C(_13442_),
    .A(_13414_),
    .Y(_13455_));
 sg13g2_nor2_1 _39429_ (.A(_13394_),
    .B(_13455_),
    .Y(_13456_));
 sg13g2_o21ai_1 _39430_ (.B1(net4576),
    .Y(_13457_),
    .A1(_13424_),
    .A2(_13441_));
 sg13g2_o21ai_1 _39431_ (.B1(_13457_),
    .Y(_13458_),
    .A1(_13428_),
    .A2(_13454_));
 sg13g2_a21oi_2 _39432_ (.B1(_13458_),
    .Y(_13459_),
    .A2(_13456_),
    .A1(_13401_));
 sg13g2_o21ai_1 _39433_ (.B1(net4686),
    .Y(_13460_),
    .A1(_13453_),
    .A2(_13459_));
 sg13g2_a21oi_1 _39434_ (.A1(_13453_),
    .A2(_13459_),
    .Y(_13461_),
    .B1(_13460_));
 sg13g2_a21oi_1 _39435_ (.A1(net4645),
    .A2(_13451_),
    .Y(_13462_),
    .B1(_13461_));
 sg13g2_o21ai_1 _39436_ (.B1(net5588),
    .Y(_13463_),
    .A1(net4381),
    .A2(_13441_));
 sg13g2_a21oi_1 _39437_ (.A1(net4381),
    .A2(_13462_),
    .Y(_13464_),
    .B1(_13463_));
 sg13g2_a21o_1 _39438_ (.A2(net4124),
    .A1(net2658),
    .B1(_13464_),
    .X(_01025_));
 sg13g2_nand2_1 _39439_ (.Y(_13465_),
    .A(net2506),
    .B(net4125));
 sg13g2_a21oi_1 _39440_ (.A1(_07267_),
    .A2(_13439_),
    .Y(_13466_),
    .B1(_06516_));
 sg13g2_xnor2_1 _39441_ (.Y(_13467_),
    .A(_06494_),
    .B(_13466_));
 sg13g2_nand2_1 _39442_ (.Y(_13468_),
    .A(net5389),
    .B(_13467_));
 sg13g2_o21ai_1 _39443_ (.B1(_13468_),
    .Y(_13469_),
    .A1(net5389),
    .A2(_06492_));
 sg13g2_xnor2_1 _39444_ (.Y(_13470_),
    .A(net4576),
    .B(_13469_));
 sg13g2_o21ai_1 _39445_ (.B1(_13452_),
    .Y(_13471_),
    .A1(_13453_),
    .A2(_13459_));
 sg13g2_xnor2_1 _39446_ (.Y(_13472_),
    .A(_13470_),
    .B(_13471_));
 sg13g2_a21o_1 _39447_ (.A2(_13469_),
    .A1(net4646),
    .B1(net4352),
    .X(_13473_));
 sg13g2_a21oi_1 _39448_ (.A1(net4686),
    .A2(_13472_),
    .Y(_13474_),
    .B1(_13473_));
 sg13g2_o21ai_1 _39449_ (.B1(net5588),
    .Y(_13475_),
    .A1(net4381),
    .A2(_13451_));
 sg13g2_o21ai_1 _39450_ (.B1(_13465_),
    .Y(_01026_),
    .A1(_13474_),
    .A2(_13475_));
 sg13g2_nand2_1 _39451_ (.Y(_13476_),
    .A(net1419),
    .B(net4125));
 sg13g2_or2_1 _39452_ (.X(_13477_),
    .B(_13470_),
    .A(_13453_));
 sg13g2_o21ai_1 _39453_ (.B1(net4576),
    .Y(_13478_),
    .A1(_13451_),
    .A2(_13469_));
 sg13g2_o21ai_1 _39454_ (.B1(_13478_),
    .Y(_13479_),
    .A1(_13459_),
    .A2(_13477_));
 sg13g2_nor2_1 _39455_ (.A(net5391),
    .B(_06503_),
    .Y(_13480_));
 sg13g2_a21oi_1 _39456_ (.A1(_06495_),
    .A2(_13466_),
    .Y(_13481_),
    .B1(_06493_));
 sg13g2_xor2_1 _39457_ (.B(_13481_),
    .A(_06504_),
    .X(_13482_));
 sg13g2_a21oi_2 _39458_ (.B1(_13480_),
    .Y(_13483_),
    .A2(_13482_),
    .A1(net5391));
 sg13g2_and2_1 _39459_ (.A(net4580),
    .B(_13483_),
    .X(_13484_));
 sg13g2_xnor2_1 _39460_ (.Y(_13485_),
    .A(net4536),
    .B(_13483_));
 sg13g2_xor2_1 _39461_ (.B(_13485_),
    .A(_13479_),
    .X(_13486_));
 sg13g2_a21o_1 _39462_ (.A2(_13483_),
    .A1(net4646),
    .B1(net4352),
    .X(_13487_));
 sg13g2_a21oi_1 _39463_ (.A1(net4689),
    .A2(_13486_),
    .Y(_13488_),
    .B1(_13487_));
 sg13g2_o21ai_1 _39464_ (.B1(net5590),
    .Y(_13489_),
    .A1(net4384),
    .A2(_13469_));
 sg13g2_o21ai_1 _39465_ (.B1(_13476_),
    .Y(_01027_),
    .A1(_13488_),
    .A2(_13489_));
 sg13g2_nor2_1 _39466_ (.A(net5390),
    .B(_09666_),
    .Y(_13490_));
 sg13g2_xnor2_1 _39467_ (.Y(_13491_),
    .A(_09661_),
    .B(_09668_));
 sg13g2_a21oi_2 _39468_ (.B1(_13490_),
    .Y(_13492_),
    .A2(_13491_),
    .A1(net5390));
 sg13g2_inv_1 _39469_ (.Y(_13493_),
    .A(_13492_));
 sg13g2_xnor2_1 _39470_ (.Y(_13494_),
    .A(net4536),
    .B(_13492_));
 sg13g2_a21oi_1 _39471_ (.A1(_13479_),
    .A2(_13485_),
    .Y(_13495_),
    .B1(_13484_));
 sg13g2_xnor2_1 _39472_ (.Y(_13496_),
    .A(_13494_),
    .B(_13495_));
 sg13g2_o21ai_1 _39473_ (.B1(net4384),
    .Y(_13497_),
    .A1(net4689),
    .A2(_13493_));
 sg13g2_a21oi_1 _39474_ (.A1(net4689),
    .A2(_13496_),
    .Y(_13498_),
    .B1(_13497_));
 sg13g2_o21ai_1 _39475_ (.B1(net5590),
    .Y(_13499_),
    .A1(net4384),
    .A2(_13483_));
 sg13g2_nand2_1 _39476_ (.Y(_13500_),
    .A(net2962),
    .B(net4125));
 sg13g2_o21ai_1 _39477_ (.B1(_13500_),
    .Y(_01028_),
    .A1(_13498_),
    .A2(_13499_));
 sg13g2_nand2_1 _39478_ (.Y(_13501_),
    .A(net2018),
    .B(net4125));
 sg13g2_nand3_1 _39479_ (.B(_13485_),
    .C(_13494_),
    .A(_13479_),
    .Y(_13502_));
 sg13g2_o21ai_1 _39480_ (.B1(net4580),
    .Y(_13503_),
    .A1(_13483_),
    .A2(_13492_));
 sg13g2_and2_1 _39481_ (.A(net4689),
    .B(_13503_),
    .X(_13504_));
 sg13g2_a22oi_1 _39482_ (.Y(_13505_),
    .B1(_13502_),
    .B2(_13504_),
    .A2(net4580),
    .A1(net4646));
 sg13g2_mux2_1 _39483_ (.A0(_13493_),
    .A1(_13505_),
    .S(net4384),
    .X(_13506_));
 sg13g2_o21ai_1 _39484_ (.B1(_13501_),
    .Y(_01029_),
    .A1(net5528),
    .A2(_13506_));
 sg13g2_nand2_1 _39485_ (.Y(_13507_),
    .A(net2349),
    .B(net4125));
 sg13g2_mux2_1 _39486_ (.A0(net4536),
    .A1(_13505_),
    .S(net4384),
    .X(_13508_));
 sg13g2_o21ai_1 _39487_ (.B1(_13507_),
    .Y(_01030_),
    .A1(net5528),
    .A2(_13508_));
 sg13g2_a21oi_2 _39488_ (.B1(net4130),
    .Y(_13509_),
    .A2(net5025),
    .A1(net5634));
 sg13g2_a21o_2 _39489_ (.A2(net5025),
    .A1(net5634),
    .B1(net4130),
    .X(_13510_));
 sg13g2_nor2_1 _39490_ (.A(net5057),
    .B(net5555),
    .Y(_13511_));
 sg13g2_nand2_1 _39491_ (.Y(_13512_),
    .A(net1384),
    .B(net4833));
 sg13g2_o21ai_1 _39492_ (.B1(_13512_),
    .Y(_01031_),
    .A1(_14552_),
    .A2(net4077));
 sg13g2_nand2_1 _39493_ (.Y(_13513_),
    .A(net2398),
    .B(net4833));
 sg13g2_o21ai_1 _39494_ (.B1(_13513_),
    .Y(_01032_),
    .A1(_14808_),
    .A2(net4077));
 sg13g2_nand2_1 _39495_ (.Y(_13514_),
    .A(net2430),
    .B(net4833));
 sg13g2_o21ai_1 _39496_ (.B1(_13514_),
    .Y(_01033_),
    .A1(_14807_),
    .A2(net4077));
 sg13g2_nand2_1 _39497_ (.Y(_13515_),
    .A(net2563),
    .B(net4835));
 sg13g2_o21ai_1 _39498_ (.B1(_13515_),
    .Y(_01034_),
    .A1(_14806_),
    .A2(net4077));
 sg13g2_nand2_1 _39499_ (.Y(_13516_),
    .A(net2781),
    .B(net4840));
 sg13g2_o21ai_1 _39500_ (.B1(_13516_),
    .Y(_01035_),
    .A1(_14805_),
    .A2(net4082));
 sg13g2_nand2_1 _39501_ (.Y(_13517_),
    .A(net2862),
    .B(net4840));
 sg13g2_o21ai_1 _39502_ (.B1(_13517_),
    .Y(_01036_),
    .A1(_14804_),
    .A2(net4082));
 sg13g2_nand2_1 _39503_ (.Y(_13518_),
    .A(net2543),
    .B(net4840));
 sg13g2_o21ai_1 _39504_ (.B1(_13518_),
    .Y(_01037_),
    .A1(_14803_),
    .A2(net4082));
 sg13g2_nand2_1 _39505_ (.Y(_13519_),
    .A(net2426),
    .B(net4840));
 sg13g2_o21ai_1 _39506_ (.B1(_13519_),
    .Y(_01038_),
    .A1(_14802_),
    .A2(net4082));
 sg13g2_nand2_1 _39507_ (.Y(_13520_),
    .A(net2604),
    .B(net4840));
 sg13g2_o21ai_1 _39508_ (.B1(_13520_),
    .Y(_01039_),
    .A1(_14801_),
    .A2(net4082));
 sg13g2_nand2_1 _39509_ (.Y(_13521_),
    .A(net2503),
    .B(net4840));
 sg13g2_o21ai_1 _39510_ (.B1(_13521_),
    .Y(_01040_),
    .A1(_14800_),
    .A2(net4082));
 sg13g2_nand2_1 _39511_ (.Y(_13522_),
    .A(net3093),
    .B(net4840));
 sg13g2_o21ai_1 _39512_ (.B1(_13522_),
    .Y(_01041_),
    .A1(_14799_),
    .A2(net4082));
 sg13g2_nand2_1 _39513_ (.Y(_13523_),
    .A(net3215),
    .B(net4840));
 sg13g2_o21ai_1 _39514_ (.B1(_13523_),
    .Y(_01042_),
    .A1(_14798_),
    .A2(net4082));
 sg13g2_nand2_1 _39515_ (.Y(_13524_),
    .A(net2523),
    .B(net4843));
 sg13g2_o21ai_1 _39516_ (.B1(_13524_),
    .Y(_01043_),
    .A1(_14797_),
    .A2(net4083));
 sg13g2_nand2_1 _39517_ (.Y(_13525_),
    .A(net2508),
    .B(net4843));
 sg13g2_o21ai_1 _39518_ (.B1(_13525_),
    .Y(_01044_),
    .A1(_14796_),
    .A2(net4083));
 sg13g2_nand2_1 _39519_ (.Y(_13526_),
    .A(net2441),
    .B(net4843));
 sg13g2_o21ai_1 _39520_ (.B1(_13526_),
    .Y(_01045_),
    .A1(_14795_),
    .A2(net4083));
 sg13g2_nand2_1 _39521_ (.Y(_13527_),
    .A(net2619),
    .B(net4843));
 sg13g2_o21ai_1 _39522_ (.B1(_13527_),
    .Y(_01046_),
    .A1(_14794_),
    .A2(net4083));
 sg13g2_nand2_1 _39523_ (.Y(_13528_),
    .A(net2934),
    .B(net4843));
 sg13g2_o21ai_1 _39524_ (.B1(_13528_),
    .Y(_01047_),
    .A1(_14793_),
    .A2(net4083));
 sg13g2_nand2_1 _39525_ (.Y(_13529_),
    .A(net2787),
    .B(net4843));
 sg13g2_o21ai_1 _39526_ (.B1(_13529_),
    .Y(_01048_),
    .A1(_14792_),
    .A2(net4083));
 sg13g2_nand2_1 _39527_ (.Y(_13530_),
    .A(net2704),
    .B(net4843));
 sg13g2_o21ai_1 _39528_ (.B1(_13530_),
    .Y(_01049_),
    .A1(_14791_),
    .A2(net4083));
 sg13g2_nand2_1 _39529_ (.Y(_13531_),
    .A(net2904),
    .B(net4852));
 sg13g2_o21ai_1 _39530_ (.B1(_13531_),
    .Y(_01050_),
    .A1(_14790_),
    .A2(net4088));
 sg13g2_nand2_1 _39531_ (.Y(_13532_),
    .A(net2596),
    .B(net4852));
 sg13g2_o21ai_1 _39532_ (.B1(_13532_),
    .Y(_01051_),
    .A1(_14789_),
    .A2(net4088));
 sg13g2_nand2_1 _39533_ (.Y(_13533_),
    .A(net2299),
    .B(net4852));
 sg13g2_o21ai_1 _39534_ (.B1(_13533_),
    .Y(_01052_),
    .A1(_14788_),
    .A2(net4088));
 sg13g2_nand2_1 _39535_ (.Y(_13534_),
    .A(net2308),
    .B(net4852));
 sg13g2_o21ai_1 _39536_ (.B1(_13534_),
    .Y(_01053_),
    .A1(_14787_),
    .A2(net4088));
 sg13g2_nand2_1 _39537_ (.Y(_13535_),
    .A(net3055),
    .B(net4852));
 sg13g2_o21ai_1 _39538_ (.B1(_13535_),
    .Y(_01054_),
    .A1(_14786_),
    .A2(net4088));
 sg13g2_nand2_1 _39539_ (.Y(_13536_),
    .A(net2473),
    .B(net4852));
 sg13g2_o21ai_1 _39540_ (.B1(_13536_),
    .Y(_01055_),
    .A1(_14785_),
    .A2(net4088));
 sg13g2_nand2_1 _39541_ (.Y(_13537_),
    .A(net1612),
    .B(net4852));
 sg13g2_o21ai_1 _39542_ (.B1(_13537_),
    .Y(_01056_),
    .A1(_14784_),
    .A2(net4088));
 sg13g2_nand2_1 _39543_ (.Y(_13538_),
    .A(net2840),
    .B(net4855));
 sg13g2_o21ai_1 _39544_ (.B1(_13538_),
    .Y(_01057_),
    .A1(_14783_),
    .A2(net4087));
 sg13g2_nand2_1 _39545_ (.Y(_13539_),
    .A(net2970),
    .B(net4855));
 sg13g2_o21ai_1 _39546_ (.B1(_13539_),
    .Y(_01058_),
    .A1(_14782_),
    .A2(net4087));
 sg13g2_nand2_1 _39547_ (.Y(_13540_),
    .A(net1597),
    .B(net4855));
 sg13g2_o21ai_1 _39548_ (.B1(_13540_),
    .Y(_01059_),
    .A1(_14781_),
    .A2(net4087));
 sg13g2_nand2_1 _39549_ (.Y(_13541_),
    .A(net2273),
    .B(net4855));
 sg13g2_o21ai_1 _39550_ (.B1(_13541_),
    .Y(_01060_),
    .A1(_14780_),
    .A2(net4087));
 sg13g2_nand2_1 _39551_ (.Y(_13542_),
    .A(net2055),
    .B(net4855));
 sg13g2_o21ai_1 _39552_ (.B1(_13542_),
    .Y(_01061_),
    .A1(_14779_),
    .A2(net4087));
 sg13g2_nand2_1 _39553_ (.Y(_13543_),
    .A(net2130),
    .B(net4855));
 sg13g2_o21ai_1 _39554_ (.B1(_13543_),
    .Y(_01062_),
    .A1(_14778_),
    .A2(net4087));
 sg13g2_nand2_1 _39555_ (.Y(_13544_),
    .A(net2689),
    .B(net4863));
 sg13g2_o21ai_1 _39556_ (.B1(_13544_),
    .Y(_01063_),
    .A1(_14777_),
    .A2(net4092));
 sg13g2_nand2_1 _39557_ (.Y(_13545_),
    .A(net2984),
    .B(net4863));
 sg13g2_o21ai_1 _39558_ (.B1(_13545_),
    .Y(_01064_),
    .A1(_14776_),
    .A2(net4092));
 sg13g2_nand2_1 _39559_ (.Y(_13546_),
    .A(net2588),
    .B(net4863));
 sg13g2_o21ai_1 _39560_ (.B1(_13546_),
    .Y(_01065_),
    .A1(_14775_),
    .A2(net4092));
 sg13g2_nand2_1 _39561_ (.Y(_13547_),
    .A(net2581),
    .B(net4863));
 sg13g2_o21ai_1 _39562_ (.B1(_13547_),
    .Y(_01066_),
    .A1(_14774_),
    .A2(net4092));
 sg13g2_nand2_1 _39563_ (.Y(_13548_),
    .A(net3217),
    .B(net4863));
 sg13g2_o21ai_1 _39564_ (.B1(_13548_),
    .Y(_01067_),
    .A1(_14773_),
    .A2(net4092));
 sg13g2_nand2_1 _39565_ (.Y(_13549_),
    .A(net2864),
    .B(net4863));
 sg13g2_o21ai_1 _39566_ (.B1(_13549_),
    .Y(_01068_),
    .A1(_14772_),
    .A2(net4092));
 sg13g2_nand2_1 _39567_ (.Y(_13550_),
    .A(net2268),
    .B(net4863));
 sg13g2_o21ai_1 _39568_ (.B1(_13550_),
    .Y(_01069_),
    .A1(_14771_),
    .A2(net4092));
 sg13g2_nand2_1 _39569_ (.Y(_13551_),
    .A(net2261),
    .B(net4863));
 sg13g2_o21ai_1 _39570_ (.B1(_13551_),
    .Y(_01070_),
    .A1(_14770_),
    .A2(net4092));
 sg13g2_nand2_1 _39571_ (.Y(_13552_),
    .A(net2885),
    .B(net4865));
 sg13g2_o21ai_1 _39572_ (.B1(_13552_),
    .Y(_01071_),
    .A1(_14769_),
    .A2(net4093));
 sg13g2_nand2_1 _39573_ (.Y(_13553_),
    .A(net2415),
    .B(net4865));
 sg13g2_o21ai_1 _39574_ (.B1(_13553_),
    .Y(_01072_),
    .A1(_14768_),
    .A2(net4093));
 sg13g2_nand2_1 _39575_ (.Y(_13554_),
    .A(net2343),
    .B(net4865));
 sg13g2_o21ai_1 _39576_ (.B1(_13554_),
    .Y(_01073_),
    .A1(_14767_),
    .A2(net4093));
 sg13g2_nand2_1 _39577_ (.Y(_13555_),
    .A(net2213),
    .B(net4865));
 sg13g2_o21ai_1 _39578_ (.B1(_13555_),
    .Y(_01074_),
    .A1(_14766_),
    .A2(net4093));
 sg13g2_nand2_1 _39579_ (.Y(_13556_),
    .A(net2407),
    .B(net4865));
 sg13g2_o21ai_1 _39580_ (.B1(_13556_),
    .Y(_01075_),
    .A1(_14765_),
    .A2(net4093));
 sg13g2_nand2_1 _39581_ (.Y(_13557_),
    .A(net2104),
    .B(net4865));
 sg13g2_o21ai_1 _39582_ (.B1(_13557_),
    .Y(_01076_),
    .A1(_14764_),
    .A2(net4093));
 sg13g2_nand2_1 _39583_ (.Y(_13558_),
    .A(net2325),
    .B(net4875));
 sg13g2_o21ai_1 _39584_ (.B1(_13558_),
    .Y(_01077_),
    .A1(_14763_),
    .A2(net4099));
 sg13g2_nand2_1 _39585_ (.Y(_13559_),
    .A(net2479),
    .B(net4875));
 sg13g2_o21ai_1 _39586_ (.B1(_13559_),
    .Y(_01078_),
    .A1(_14762_),
    .A2(net4099));
 sg13g2_nand2_1 _39587_ (.Y(_13560_),
    .A(net2881),
    .B(net4888));
 sg13g2_o21ai_1 _39588_ (.B1(_13560_),
    .Y(_01079_),
    .A1(_14761_),
    .A2(net4103));
 sg13g2_nand2_1 _39589_ (.Y(_13561_),
    .A(net2926),
    .B(net4888));
 sg13g2_o21ai_1 _39590_ (.B1(_13561_),
    .Y(_01080_),
    .A1(_14760_),
    .A2(net4103));
 sg13g2_nand2_1 _39591_ (.Y(_13562_),
    .A(net3304),
    .B(net4888));
 sg13g2_o21ai_1 _39592_ (.B1(_13562_),
    .Y(_01081_),
    .A1(_14759_),
    .A2(net4103));
 sg13g2_nand2_1 _39593_ (.Y(_13563_),
    .A(net2645),
    .B(net4888));
 sg13g2_o21ai_1 _39594_ (.B1(_13563_),
    .Y(_01082_),
    .A1(_14758_),
    .A2(net4103));
 sg13g2_nand2_1 _39595_ (.Y(_13564_),
    .A(net2740),
    .B(net4888));
 sg13g2_o21ai_1 _39596_ (.B1(_13564_),
    .Y(_01083_),
    .A1(_14757_),
    .A2(net4103));
 sg13g2_nand2_1 _39597_ (.Y(_13565_),
    .A(net2438),
    .B(net4888));
 sg13g2_o21ai_1 _39598_ (.B1(_13565_),
    .Y(_01084_),
    .A1(_14756_),
    .A2(net4103));
 sg13g2_nand2_1 _39599_ (.Y(_13566_),
    .A(net1726),
    .B(net4888));
 sg13g2_o21ai_1 _39600_ (.B1(_13566_),
    .Y(_01085_),
    .A1(_14755_),
    .A2(net4103));
 sg13g2_nand2_1 _39601_ (.Y(_13567_),
    .A(net2590),
    .B(net4890));
 sg13g2_o21ai_1 _39602_ (.B1(_13567_),
    .Y(_01086_),
    .A1(_14754_),
    .A2(net4104));
 sg13g2_nand2_1 _39603_ (.Y(_13568_),
    .A(net2177),
    .B(net4890));
 sg13g2_o21ai_1 _39604_ (.B1(_13568_),
    .Y(_01087_),
    .A1(_14753_),
    .A2(net4103));
 sg13g2_nand2_1 _39605_ (.Y(_13569_),
    .A(net2624),
    .B(net4890));
 sg13g2_o21ai_1 _39606_ (.B1(_13569_),
    .Y(_01088_),
    .A1(_14752_),
    .A2(net4104));
 sg13g2_nand2_1 _39607_ (.Y(_13570_),
    .A(net2606),
    .B(net4890));
 sg13g2_o21ai_1 _39608_ (.B1(_13570_),
    .Y(_01089_),
    .A1(_14751_),
    .A2(net4104));
 sg13g2_nand2_1 _39609_ (.Y(_13571_),
    .A(net2117),
    .B(net4890));
 sg13g2_o21ai_1 _39610_ (.B1(_13571_),
    .Y(_01090_),
    .A1(_14750_),
    .A2(net4104));
 sg13g2_nand2_1 _39611_ (.Y(_13572_),
    .A(net2347),
    .B(net4890));
 sg13g2_o21ai_1 _39612_ (.B1(_13572_),
    .Y(_01091_),
    .A1(_14749_),
    .A2(net4109));
 sg13g2_nand2_1 _39613_ (.Y(_13573_),
    .A(net2600),
    .B(net4890));
 sg13g2_o21ai_1 _39614_ (.B1(_13573_),
    .Y(_01092_),
    .A1(_14748_),
    .A2(net4109));
 sg13g2_nand2_1 _39615_ (.Y(_13574_),
    .A(net1582),
    .B(net4899));
 sg13g2_o21ai_1 _39616_ (.B1(_13574_),
    .Y(_01093_),
    .A1(_14747_),
    .A2(net4109));
 sg13g2_nand2_1 _39617_ (.Y(_13575_),
    .A(net2678),
    .B(net4899));
 sg13g2_o21ai_1 _39618_ (.B1(_13575_),
    .Y(_01094_),
    .A1(_14746_),
    .A2(net4109));
 sg13g2_nand2_1 _39619_ (.Y(_13576_),
    .A(net2641),
    .B(net4899));
 sg13g2_o21ai_1 _39620_ (.B1(_13576_),
    .Y(_01095_),
    .A1(_14745_),
    .A2(net4109));
 sg13g2_nand2_1 _39621_ (.Y(_13577_),
    .A(net2334),
    .B(net4899));
 sg13g2_o21ai_1 _39622_ (.B1(_13577_),
    .Y(_01096_),
    .A1(_14744_),
    .A2(net4109));
 sg13g2_nand2_1 _39623_ (.Y(_13578_),
    .A(net1260),
    .B(net4899));
 sg13g2_o21ai_1 _39624_ (.B1(_13578_),
    .Y(_01097_),
    .A1(_14743_),
    .A2(net4109));
 sg13g2_nand2_1 _39625_ (.Y(_13579_),
    .A(net2879),
    .B(net4899));
 sg13g2_o21ai_1 _39626_ (.B1(_13579_),
    .Y(_01098_),
    .A1(_14742_),
    .A2(net4109));
 sg13g2_nand2_1 _39627_ (.Y(_13580_),
    .A(net2871),
    .B(net4900));
 sg13g2_o21ai_1 _39628_ (.B1(_13580_),
    .Y(_01099_),
    .A1(_14741_),
    .A2(net4110));
 sg13g2_nand2_1 _39629_ (.Y(_13581_),
    .A(net2952),
    .B(net4900));
 sg13g2_o21ai_1 _39630_ (.B1(_13581_),
    .Y(_01100_),
    .A1(_14740_),
    .A2(net4110));
 sg13g2_nand2_1 _39631_ (.Y(_13582_),
    .A(net1406),
    .B(net4900));
 sg13g2_o21ai_1 _39632_ (.B1(_13582_),
    .Y(_01101_),
    .A1(_14739_),
    .A2(net4110));
 sg13g2_nand2_1 _39633_ (.Y(_13583_),
    .A(net2536),
    .B(net4900));
 sg13g2_o21ai_1 _39634_ (.B1(_13583_),
    .Y(_01102_),
    .A1(_14738_),
    .A2(net4115));
 sg13g2_nand2_1 _39635_ (.Y(_13584_),
    .A(net5878),
    .B(net4900));
 sg13g2_o21ai_1 _39636_ (.B1(_13584_),
    .Y(_01103_),
    .A1(_14737_),
    .A2(net4110));
 sg13g2_nand2_1 _39637_ (.Y(_13585_),
    .A(net2963),
    .B(net4900));
 sg13g2_o21ai_1 _39638_ (.B1(_13585_),
    .Y(_01104_),
    .A1(_14736_),
    .A2(net4110));
 sg13g2_nand2_1 _39639_ (.Y(_13586_),
    .A(net1359),
    .B(net4900));
 sg13g2_o21ai_1 _39640_ (.B1(_13586_),
    .Y(_01105_),
    .A1(_14735_),
    .A2(net4110));
 sg13g2_nand2_1 _39641_ (.Y(_13587_),
    .A(net1954),
    .B(net4908));
 sg13g2_o21ai_1 _39642_ (.B1(_13587_),
    .Y(_01106_),
    .A1(_14734_),
    .A2(net4118));
 sg13g2_nand2_1 _39643_ (.Y(_13588_),
    .A(net2974),
    .B(net4908));
 sg13g2_o21ai_1 _39644_ (.B1(_13588_),
    .Y(_01107_),
    .A1(_14733_),
    .A2(net4118));
 sg13g2_nand2_1 _39645_ (.Y(_13589_),
    .A(net3087),
    .B(net4908));
 sg13g2_o21ai_1 _39646_ (.B1(_13589_),
    .Y(_01108_),
    .A1(_14732_),
    .A2(net4118));
 sg13g2_nand2_1 _39647_ (.Y(_13590_),
    .A(net2306),
    .B(net4908));
 sg13g2_o21ai_1 _39648_ (.B1(_13590_),
    .Y(_01109_),
    .A1(_14731_),
    .A2(net4118));
 sg13g2_nand2_1 _39649_ (.Y(_13591_),
    .A(net3027),
    .B(net4908));
 sg13g2_o21ai_1 _39650_ (.B1(_13591_),
    .Y(_01110_),
    .A1(_14730_),
    .A2(net4118));
 sg13g2_nand2_1 _39651_ (.Y(_13592_),
    .A(net2849),
    .B(net4909));
 sg13g2_o21ai_1 _39652_ (.B1(_13592_),
    .Y(_01111_),
    .A1(_14729_),
    .A2(net4117));
 sg13g2_nand2_1 _39653_ (.Y(_13593_),
    .A(net2928),
    .B(net4908));
 sg13g2_o21ai_1 _39654_ (.B1(_13593_),
    .Y(_01112_),
    .A1(_14728_),
    .A2(net4117));
 sg13g2_nand2_1 _39655_ (.Y(_13594_),
    .A(net2448),
    .B(net4909));
 sg13g2_o21ai_1 _39656_ (.B1(_13594_),
    .Y(_01113_),
    .A1(_14727_),
    .A2(net4117));
 sg13g2_nand2_1 _39657_ (.Y(_13595_),
    .A(net2636),
    .B(net4909));
 sg13g2_o21ai_1 _39658_ (.B1(_13595_),
    .Y(_01114_),
    .A1(_14726_),
    .A2(net4117));
 sg13g2_nand2_1 _39659_ (.Y(_13596_),
    .A(net2810),
    .B(net4909));
 sg13g2_o21ai_1 _39660_ (.B1(_13596_),
    .Y(_01115_),
    .A1(_14725_),
    .A2(net4117));
 sg13g2_nand2_1 _39661_ (.Y(_13597_),
    .A(net2468),
    .B(net4909));
 sg13g2_o21ai_1 _39662_ (.B1(_13597_),
    .Y(_01116_),
    .A1(_14724_),
    .A2(net4117));
 sg13g2_nand2_1 _39663_ (.Y(_13598_),
    .A(net2276),
    .B(net4909));
 sg13g2_o21ai_1 _39664_ (.B1(_13598_),
    .Y(_01117_),
    .A1(_14723_),
    .A2(net4117));
 sg13g2_nand2_1 _39665_ (.Y(_13599_),
    .A(net1524),
    .B(net4909));
 sg13g2_o21ai_1 _39666_ (.B1(_13599_),
    .Y(_01118_),
    .A1(_14722_),
    .A2(net4117));
 sg13g2_nand2_1 _39667_ (.Y(_13600_),
    .A(net3270),
    .B(net4909));
 sg13g2_o21ai_1 _39668_ (.B1(_13600_),
    .Y(_01119_),
    .A1(_14721_),
    .A2(net4116));
 sg13g2_nand2_1 _39669_ (.Y(_13601_),
    .A(net3047),
    .B(net4910));
 sg13g2_o21ai_1 _39670_ (.B1(_13601_),
    .Y(_01120_),
    .A1(_14720_),
    .A2(net4118));
 sg13g2_nand2_1 _39671_ (.Y(_13602_),
    .A(net2853),
    .B(net4910));
 sg13g2_o21ai_1 _39672_ (.B1(_13602_),
    .Y(_01121_),
    .A1(_14719_),
    .A2(net4116));
 sg13g2_nand2_1 _39673_ (.Y(_13603_),
    .A(net2667),
    .B(net4910));
 sg13g2_o21ai_1 _39674_ (.B1(_13603_),
    .Y(_01122_),
    .A1(_14718_),
    .A2(net4116));
 sg13g2_nand2_1 _39675_ (.Y(_13604_),
    .A(net2388),
    .B(net4910));
 sg13g2_o21ai_1 _39676_ (.B1(_13604_),
    .Y(_01123_),
    .A1(_14717_),
    .A2(net4116));
 sg13g2_nand2_1 _39677_ (.Y(_13605_),
    .A(net3315),
    .B(net4910));
 sg13g2_o21ai_1 _39678_ (.B1(_13605_),
    .Y(_01124_),
    .A1(_14716_),
    .A2(net4116));
 sg13g2_nand2_1 _39679_ (.Y(_13606_),
    .A(net2626),
    .B(net4910));
 sg13g2_o21ai_1 _39680_ (.B1(_13606_),
    .Y(_01125_),
    .A1(_14715_),
    .A2(net4120));
 sg13g2_nand2_1 _39681_ (.Y(_13607_),
    .A(net2944),
    .B(net4910));
 sg13g2_o21ai_1 _39682_ (.B1(_13607_),
    .Y(_01126_),
    .A1(_14714_),
    .A2(net4116));
 sg13g2_nand2_1 _39683_ (.Y(_13608_),
    .A(net3044),
    .B(net4907));
 sg13g2_o21ai_1 _39684_ (.B1(_13608_),
    .Y(_01127_),
    .A1(_14713_),
    .A2(net4116));
 sg13g2_nand2_1 _39685_ (.Y(_13609_),
    .A(net3104),
    .B(net4911));
 sg13g2_o21ai_1 _39686_ (.B1(_13609_),
    .Y(_01128_),
    .A1(_14712_),
    .A2(net4116));
 sg13g2_nand2_1 _39687_ (.Y(_13610_),
    .A(\u_inv.d_next[98] ),
    .B(net4911));
 sg13g2_o21ai_1 _39688_ (.B1(_13610_),
    .Y(_01129_),
    .A1(_14711_),
    .A2(net4120));
 sg13g2_nand2_1 _39689_ (.Y(_13611_),
    .A(net2420),
    .B(net4908));
 sg13g2_o21ai_1 _39690_ (.B1(_13611_),
    .Y(_01130_),
    .A1(_14710_),
    .A2(net4119));
 sg13g2_nand2_1 _39691_ (.Y(_13612_),
    .A(net2337),
    .B(net4907));
 sg13g2_o21ai_1 _39692_ (.B1(_13612_),
    .Y(_01131_),
    .A1(_14709_),
    .A2(net4119));
 sg13g2_nand2_1 _39693_ (.Y(_13613_),
    .A(net2612),
    .B(net4907));
 sg13g2_o21ai_1 _39694_ (.B1(_13613_),
    .Y(_01132_),
    .A1(_14708_),
    .A2(net4119));
 sg13g2_nand2_1 _39695_ (.Y(_13614_),
    .A(net2327),
    .B(net4907));
 sg13g2_o21ai_1 _39696_ (.B1(_13614_),
    .Y(_01133_),
    .A1(_14707_),
    .A2(net4119));
 sg13g2_nand2_1 _39697_ (.Y(_13615_),
    .A(net1640),
    .B(net4907));
 sg13g2_o21ai_1 _39698_ (.B1(_13615_),
    .Y(_01134_),
    .A1(_14706_),
    .A2(net4119));
 sg13g2_nand2_1 _39699_ (.Y(_13616_),
    .A(net2321),
    .B(net4907));
 sg13g2_o21ai_1 _39700_ (.B1(_13616_),
    .Y(_01135_),
    .A1(_14705_),
    .A2(net4119));
 sg13g2_nand2_1 _39701_ (.Y(_13617_),
    .A(net2514),
    .B(net4907));
 sg13g2_o21ai_1 _39702_ (.B1(_13617_),
    .Y(_01136_),
    .A1(_14704_),
    .A2(net4119));
 sg13g2_nand2_1 _39703_ (.Y(_13618_),
    .A(net3097),
    .B(net4913));
 sg13g2_o21ai_1 _39704_ (.B1(_13618_),
    .Y(_01137_),
    .A1(_14703_),
    .A2(net4120));
 sg13g2_nand2_1 _39705_ (.Y(_13619_),
    .A(net3231),
    .B(net4907));
 sg13g2_o21ai_1 _39706_ (.B1(_13619_),
    .Y(_01138_),
    .A1(_14702_),
    .A2(net4119));
 sg13g2_nand2_1 _39707_ (.Y(_13620_),
    .A(net2516),
    .B(net4906));
 sg13g2_o21ai_1 _39708_ (.B1(_13620_),
    .Y(_01139_),
    .A1(_14701_),
    .A2(net4113));
 sg13g2_nand2_1 _39709_ (.Y(_13621_),
    .A(net1421),
    .B(net4904));
 sg13g2_o21ai_1 _39710_ (.B1(_13621_),
    .Y(_01140_),
    .A1(_14700_),
    .A2(net4114));
 sg13g2_nand2_1 _39711_ (.Y(_13622_),
    .A(net1534),
    .B(net4900));
 sg13g2_o21ai_1 _39712_ (.B1(_13622_),
    .Y(_01141_),
    .A1(_14699_),
    .A2(net4113));
 sg13g2_nand2_1 _39713_ (.Y(_13623_),
    .A(net2919),
    .B(net4901));
 sg13g2_o21ai_1 _39714_ (.B1(_13623_),
    .Y(_01142_),
    .A1(_14698_),
    .A2(net4113));
 sg13g2_nand2_1 _39715_ (.Y(_13624_),
    .A(net2437),
    .B(net4904));
 sg13g2_o21ai_1 _39716_ (.B1(_13624_),
    .Y(_01143_),
    .A1(_14697_),
    .A2(net4113));
 sg13g2_nand2_1 _39717_ (.Y(_13625_),
    .A(net2569),
    .B(net4906));
 sg13g2_o21ai_1 _39718_ (.B1(_13625_),
    .Y(_01144_),
    .A1(_14696_),
    .A2(net4114));
 sg13g2_nand2_1 _39719_ (.Y(_13626_),
    .A(net2372),
    .B(net4901));
 sg13g2_o21ai_1 _39720_ (.B1(_13626_),
    .Y(_01145_),
    .A1(_14695_),
    .A2(net4114));
 sg13g2_nand2_1 _39721_ (.Y(_13627_),
    .A(net2370),
    .B(net4901));
 sg13g2_o21ai_1 _39722_ (.B1(_13627_),
    .Y(_01146_),
    .A1(_14694_),
    .A2(net4113));
 sg13g2_nand2_1 _39723_ (.Y(_13628_),
    .A(net2906),
    .B(net4904));
 sg13g2_o21ai_1 _39724_ (.B1(_13628_),
    .Y(_01147_),
    .A1(_14693_),
    .A2(net4113));
 sg13g2_nand2_1 _39725_ (.Y(_13629_),
    .A(net3066),
    .B(net4904));
 sg13g2_o21ai_1 _39726_ (.B1(_13629_),
    .Y(_01148_),
    .A1(_14692_),
    .A2(net4113));
 sg13g2_nand2_1 _39727_ (.Y(_13630_),
    .A(net2638),
    .B(net4897));
 sg13g2_o21ai_1 _39728_ (.B1(_13630_),
    .Y(_01149_),
    .A1(_14691_),
    .A2(net4111));
 sg13g2_nand2_1 _39729_ (.Y(_13631_),
    .A(net2883),
    .B(net4897));
 sg13g2_o21ai_1 _39730_ (.B1(_13631_),
    .Y(_01150_),
    .A1(_14690_),
    .A2(net4113));
 sg13g2_nand2_1 _39731_ (.Y(_13632_),
    .A(net3068),
    .B(net4898));
 sg13g2_o21ai_1 _39732_ (.B1(_13632_),
    .Y(_01151_),
    .A1(_14689_),
    .A2(net4112));
 sg13g2_nand2_1 _39733_ (.Y(_13633_),
    .A(net3287),
    .B(net4898));
 sg13g2_o21ai_1 _39734_ (.B1(_13633_),
    .Y(_01152_),
    .A1(_14688_),
    .A2(net4112));
 sg13g2_nand2_1 _39735_ (.Y(_13634_),
    .A(net2137),
    .B(net4898));
 sg13g2_o21ai_1 _39736_ (.B1(_13634_),
    .Y(_01153_),
    .A1(_14687_),
    .A2(net4112));
 sg13g2_nand2_1 _39737_ (.Y(_13635_),
    .A(net2621),
    .B(net4898));
 sg13g2_o21ai_1 _39738_ (.B1(_13635_),
    .Y(_01154_),
    .A1(_14686_),
    .A2(net4111));
 sg13g2_nand2_1 _39739_ (.Y(_13636_),
    .A(net2697),
    .B(net4897));
 sg13g2_o21ai_1 _39740_ (.B1(_13636_),
    .Y(_01155_),
    .A1(_14685_),
    .A2(net4111));
 sg13g2_nand2_1 _39741_ (.Y(_13637_),
    .A(net3222),
    .B(net4898));
 sg13g2_o21ai_1 _39742_ (.B1(_13637_),
    .Y(_01156_),
    .A1(_14684_),
    .A2(net4112));
 sg13g2_nand2_1 _39743_ (.Y(_13638_),
    .A(net2443),
    .B(net4897));
 sg13g2_o21ai_1 _39744_ (.B1(_13638_),
    .Y(_01157_),
    .A1(_14683_),
    .A2(net4111));
 sg13g2_nand2_1 _39745_ (.Y(_13639_),
    .A(net2092),
    .B(net4897));
 sg13g2_o21ai_1 _39746_ (.B1(_13639_),
    .Y(_01158_),
    .A1(_14682_),
    .A2(net4111));
 sg13g2_nand2_1 _39747_ (.Y(_13640_),
    .A(net2976),
    .B(net4897));
 sg13g2_o21ai_1 _39748_ (.B1(_13640_),
    .Y(_01159_),
    .A1(_14681_),
    .A2(net4111));
 sg13g2_nand2_1 _39749_ (.Y(_13641_),
    .A(net2610),
    .B(net4897));
 sg13g2_o21ai_1 _39750_ (.B1(_13641_),
    .Y(_01160_),
    .A1(_14680_),
    .A2(net4111));
 sg13g2_nand2_1 _39751_ (.Y(_13642_),
    .A(net2317),
    .B(net4897));
 sg13g2_o21ai_1 _39752_ (.B1(_13642_),
    .Y(_01161_),
    .A1(_14679_),
    .A2(net4110));
 sg13g2_nand2_1 _39753_ (.Y(_13643_),
    .A(net2693),
    .B(net4889));
 sg13g2_o21ai_1 _39754_ (.B1(_13643_),
    .Y(_01162_),
    .A1(_14678_),
    .A2(net4111));
 sg13g2_nand2_1 _39755_ (.Y(_13644_),
    .A(net2470),
    .B(net4889));
 sg13g2_o21ai_1 _39756_ (.B1(_13644_),
    .Y(_01163_),
    .A1(_14677_),
    .A2(net4106));
 sg13g2_nand2_1 _39757_ (.Y(_13645_),
    .A(net3074),
    .B(net4889));
 sg13g2_o21ai_1 _39758_ (.B1(_13645_),
    .Y(_01164_),
    .A1(_14676_),
    .A2(net4105));
 sg13g2_nand2_1 _39759_ (.Y(_13646_),
    .A(net2632),
    .B(net4889));
 sg13g2_o21ai_1 _39760_ (.B1(_13646_),
    .Y(_01165_),
    .A1(_14675_),
    .A2(net4106));
 sg13g2_nand2_1 _39761_ (.Y(_13647_),
    .A(net2996),
    .B(net4891));
 sg13g2_o21ai_1 _39762_ (.B1(_13647_),
    .Y(_01166_),
    .A1(_14674_),
    .A2(net4106));
 sg13g2_nand2_1 _39763_ (.Y(_13648_),
    .A(net2145),
    .B(net4889));
 sg13g2_o21ai_1 _39764_ (.B1(_13648_),
    .Y(_01167_),
    .A1(_14673_),
    .A2(net4105));
 sg13g2_nand2_1 _39765_ (.Y(_13649_),
    .A(net3235),
    .B(net4889));
 sg13g2_o21ai_1 _39766_ (.B1(_13649_),
    .Y(_01168_),
    .A1(_14672_),
    .A2(net4105));
 sg13g2_nand2_1 _39767_ (.Y(_13650_),
    .A(net1969),
    .B(net4889));
 sg13g2_o21ai_1 _39768_ (.B1(_13650_),
    .Y(_01169_),
    .A1(_14671_),
    .A2(net4105));
 sg13g2_nand2_1 _39769_ (.Y(_13651_),
    .A(net2814),
    .B(net4889));
 sg13g2_o21ai_1 _39770_ (.B1(_13651_),
    .Y(_01170_),
    .A1(_14670_),
    .A2(net4106));
 sg13g2_nand2_1 _39771_ (.Y(_13652_),
    .A(\u_inv.d_next[140] ),
    .B(net4886));
 sg13g2_o21ai_1 _39772_ (.B1(_13652_),
    .Y(_01171_),
    .A1(_14669_),
    .A2(net4105));
 sg13g2_nand2_1 _39773_ (.Y(_13653_),
    .A(net2519),
    .B(net4887));
 sg13g2_o21ai_1 _39774_ (.B1(_13653_),
    .Y(_01172_),
    .A1(_14668_),
    .A2(net4105));
 sg13g2_nand2_1 _39775_ (.Y(_13654_),
    .A(net2552),
    .B(net4887));
 sg13g2_o21ai_1 _39776_ (.B1(_13654_),
    .Y(_01173_),
    .A1(_14667_),
    .A2(net4105));
 sg13g2_nand2_1 _39777_ (.Y(_13655_),
    .A(net2249),
    .B(net4886));
 sg13g2_o21ai_1 _39778_ (.B1(_13655_),
    .Y(_01174_),
    .A1(_14666_),
    .A2(net4105));
 sg13g2_nand2_1 _39779_ (.Y(_13656_),
    .A(net2682),
    .B(net4887));
 sg13g2_o21ai_1 _39780_ (.B1(_13656_),
    .Y(_01175_),
    .A1(_14665_),
    .A2(net4107));
 sg13g2_nand2_1 _39781_ (.Y(_13657_),
    .A(net1222),
    .B(net4887));
 sg13g2_o21ai_1 _39782_ (.B1(_13657_),
    .Y(_01176_),
    .A1(_14664_),
    .A2(net4107));
 sg13g2_nand2_1 _39783_ (.Y(_13658_),
    .A(net2756),
    .B(net4886));
 sg13g2_o21ai_1 _39784_ (.B1(_13658_),
    .Y(_01177_),
    .A1(_14663_),
    .A2(net4107));
 sg13g2_nand2_1 _39785_ (.Y(_13659_),
    .A(net2973),
    .B(net4886));
 sg13g2_o21ai_1 _39786_ (.B1(_13659_),
    .Y(_01178_),
    .A1(_14662_),
    .A2(net4107));
 sg13g2_nand2_1 _39787_ (.Y(_13660_),
    .A(net2942),
    .B(net4886));
 sg13g2_o21ai_1 _39788_ (.B1(_13660_),
    .Y(_01179_),
    .A1(_14661_),
    .A2(net4101));
 sg13g2_nand2_1 _39789_ (.Y(_13661_),
    .A(net2932),
    .B(net4886));
 sg13g2_o21ai_1 _39790_ (.B1(_13661_),
    .Y(_01180_),
    .A1(_14660_),
    .A2(net4107));
 sg13g2_nand2_1 _39791_ (.Y(_13662_),
    .A(net3003),
    .B(net4886));
 sg13g2_o21ai_1 _39792_ (.B1(_13662_),
    .Y(_01181_),
    .A1(_14659_),
    .A2(net4107));
 sg13g2_nand2_1 _39793_ (.Y(_13663_),
    .A(net3220),
    .B(net4886));
 sg13g2_o21ai_1 _39794_ (.B1(_13663_),
    .Y(_01182_),
    .A1(_14658_),
    .A2(net4107));
 sg13g2_nand2_1 _39795_ (.Y(_13664_),
    .A(net2381),
    .B(net4878));
 sg13g2_o21ai_1 _39796_ (.B1(_13664_),
    .Y(_01183_),
    .A1(_14657_),
    .A2(net4101));
 sg13g2_nand2_1 _39797_ (.Y(_13665_),
    .A(net2433),
    .B(net4878));
 sg13g2_o21ai_1 _39798_ (.B1(_13665_),
    .Y(_01184_),
    .A1(_14656_),
    .A2(net4101));
 sg13g2_nand2_1 _39799_ (.Y(_13666_),
    .A(net2406),
    .B(net4878));
 sg13g2_o21ai_1 _39800_ (.B1(_13666_),
    .Y(_01185_),
    .A1(_14655_),
    .A2(net4101));
 sg13g2_nand2_1 _39801_ (.Y(_13667_),
    .A(net2062),
    .B(net4878));
 sg13g2_o21ai_1 _39802_ (.B1(_13667_),
    .Y(_01186_),
    .A1(_14654_),
    .A2(net4101));
 sg13g2_nand2_1 _39803_ (.Y(_13668_),
    .A(net2383),
    .B(net4878));
 sg13g2_o21ai_1 _39804_ (.B1(_13668_),
    .Y(_01187_),
    .A1(_14653_),
    .A2(net4097));
 sg13g2_nand2_1 _39805_ (.Y(_13669_),
    .A(net3029),
    .B(net4878));
 sg13g2_o21ai_1 _39806_ (.B1(_13669_),
    .Y(_01188_),
    .A1(_14652_),
    .A2(net4097));
 sg13g2_nand2_1 _39807_ (.Y(_13670_),
    .A(net3254),
    .B(net4878));
 sg13g2_o21ai_1 _39808_ (.B1(_13670_),
    .Y(_01189_),
    .A1(_14651_),
    .A2(net4101));
 sg13g2_nand2_1 _39809_ (.Y(_13671_),
    .A(net3400),
    .B(net4878));
 sg13g2_o21ai_1 _39810_ (.B1(_13671_),
    .Y(_01190_),
    .A1(_14650_),
    .A2(net4101));
 sg13g2_nand2_1 _39811_ (.Y(_13672_),
    .A(net2732),
    .B(net4877));
 sg13g2_o21ai_1 _39812_ (.B1(_13672_),
    .Y(_01191_),
    .A1(_14649_),
    .A2(net4098));
 sg13g2_nand2_1 _39813_ (.Y(_13673_),
    .A(net2722),
    .B(net4877));
 sg13g2_o21ai_1 _39814_ (.B1(_13673_),
    .Y(_01192_),
    .A1(_14648_),
    .A2(net4098));
 sg13g2_nand2_1 _39815_ (.Y(_13674_),
    .A(net3082),
    .B(net4877));
 sg13g2_o21ai_1 _39816_ (.B1(_13674_),
    .Y(_01193_),
    .A1(_14647_),
    .A2(net4098));
 sg13g2_nand2_1 _39817_ (.Y(_13675_),
    .A(net2908),
    .B(net4877));
 sg13g2_o21ai_1 _39818_ (.B1(_13675_),
    .Y(_01194_),
    .A1(_14646_),
    .A2(net4097));
 sg13g2_nand2_1 _39819_ (.Y(_13676_),
    .A(\u_inv.d_next[164] ),
    .B(net4877));
 sg13g2_o21ai_1 _39820_ (.B1(_13676_),
    .Y(_01195_),
    .A1(_14645_),
    .A2(net4097));
 sg13g2_nand2_1 _39821_ (.Y(_13677_),
    .A(net3130),
    .B(net4877));
 sg13g2_o21ai_1 _39822_ (.B1(_13677_),
    .Y(_01196_),
    .A1(_14644_),
    .A2(net4097));
 sg13g2_nand2_1 _39823_ (.Y(_13678_),
    .A(net2875),
    .B(net4877));
 sg13g2_o21ai_1 _39824_ (.B1(_13678_),
    .Y(_01197_),
    .A1(_14643_),
    .A2(net4097));
 sg13g2_nand2_1 _39825_ (.Y(_13679_),
    .A(net2936),
    .B(net4877));
 sg13g2_o21ai_1 _39826_ (.B1(_13679_),
    .Y(_01198_),
    .A1(_14642_),
    .A2(net4097));
 sg13g2_nand2_1 _39827_ (.Y(_13680_),
    .A(net2561),
    .B(net4875));
 sg13g2_o21ai_1 _39828_ (.B1(_13680_),
    .Y(_01199_),
    .A1(_14641_),
    .A2(net4098));
 sg13g2_nand2_1 _39829_ (.Y(_13681_),
    .A(net2587),
    .B(net4875));
 sg13g2_o21ai_1 _39830_ (.B1(_13681_),
    .Y(_01200_),
    .A1(_14640_),
    .A2(net4099));
 sg13g2_nand2_1 _39831_ (.Y(_13682_),
    .A(net2284),
    .B(net4875));
 sg13g2_o21ai_1 _39832_ (.B1(_13682_),
    .Y(_01201_),
    .A1(_14639_),
    .A2(net4099));
 sg13g2_nand2_1 _39833_ (.Y(_13683_),
    .A(net1581),
    .B(net4875));
 sg13g2_o21ai_1 _39834_ (.B1(_13683_),
    .Y(_01202_),
    .A1(_14638_),
    .A2(net4099));
 sg13g2_nand2_1 _39835_ (.Y(_13684_),
    .A(net2246),
    .B(net4875));
 sg13g2_o21ai_1 _39836_ (.B1(_13684_),
    .Y(_01203_),
    .A1(_14637_),
    .A2(net4099));
 sg13g2_nand2_1 _39837_ (.Y(_13685_),
    .A(net2538),
    .B(net4875));
 sg13g2_o21ai_1 _39838_ (.B1(_13685_),
    .Y(_01204_),
    .A1(_14636_),
    .A2(net4099));
 sg13g2_nand2_1 _39839_ (.Y(_13686_),
    .A(net2707),
    .B(net4876));
 sg13g2_o21ai_1 _39840_ (.B1(_13686_),
    .Y(_01205_),
    .A1(_14635_),
    .A2(net4099));
 sg13g2_nand2_1 _39841_ (.Y(_13687_),
    .A(net1423),
    .B(net4876));
 sg13g2_o21ai_1 _39842_ (.B1(_13687_),
    .Y(_01206_),
    .A1(_14634_),
    .A2(net4097));
 sg13g2_nand2_1 _39843_ (.Y(_13688_),
    .A(net2140),
    .B(net4876));
 sg13g2_o21ai_1 _39844_ (.B1(_13688_),
    .Y(_01207_),
    .A1(_14633_),
    .A2(net4100));
 sg13g2_nand2_1 _39845_ (.Y(_13689_),
    .A(net1982),
    .B(net4876));
 sg13g2_o21ai_1 _39846_ (.B1(_13689_),
    .Y(_01208_),
    .A1(_14632_),
    .A2(net4100));
 sg13g2_nand2_1 _39847_ (.Y(_13690_),
    .A(net2418),
    .B(net4876));
 sg13g2_o21ai_1 _39848_ (.B1(_13690_),
    .Y(_01209_),
    .A1(_14631_),
    .A2(net4100));
 sg13g2_nand2_1 _39849_ (.Y(_13691_),
    .A(net1661),
    .B(net4876));
 sg13g2_o21ai_1 _39850_ (.B1(_13691_),
    .Y(_01210_),
    .A1(_14630_),
    .A2(net4100));
 sg13g2_nand2_1 _39851_ (.Y(_13692_),
    .A(net2836),
    .B(net4879));
 sg13g2_o21ai_1 _39852_ (.B1(_13692_),
    .Y(_01211_),
    .A1(_14629_),
    .A2(net4100));
 sg13g2_nand2_1 _39853_ (.Y(_13693_),
    .A(net2663),
    .B(net4876));
 sg13g2_o21ai_1 _39854_ (.B1(_13693_),
    .Y(_01212_),
    .A1(_14628_),
    .A2(net4100));
 sg13g2_nand2_1 _39855_ (.Y(_13694_),
    .A(net2385),
    .B(net4865));
 sg13g2_o21ai_1 _39856_ (.B1(_13694_),
    .Y(_01213_),
    .A1(_14627_),
    .A2(net4100));
 sg13g2_nand2_1 _39857_ (.Y(_13695_),
    .A(net2802),
    .B(net4879));
 sg13g2_o21ai_1 _39858_ (.B1(_13695_),
    .Y(_01214_),
    .A1(_14626_),
    .A2(net4100));
 sg13g2_nand2_1 _39859_ (.Y(_13696_),
    .A(net2909),
    .B(net4866));
 sg13g2_o21ai_1 _39860_ (.B1(_13696_),
    .Y(_01215_),
    .A1(_14625_),
    .A2(net4095));
 sg13g2_nand2_1 _39861_ (.Y(_13697_),
    .A(net1999),
    .B(net4865));
 sg13g2_o21ai_1 _39862_ (.B1(_13697_),
    .Y(_01216_),
    .A1(_14624_),
    .A2(net4095));
 sg13g2_nand2_1 _39863_ (.Y(_13698_),
    .A(net2205),
    .B(net4866));
 sg13g2_o21ai_1 _39864_ (.B1(_13698_),
    .Y(_01217_),
    .A1(_14623_),
    .A2(net4095));
 sg13g2_nand2_1 _39865_ (.Y(_13699_),
    .A(net3076),
    .B(net4866));
 sg13g2_o21ai_1 _39866_ (.B1(_13699_),
    .Y(_01218_),
    .A1(_14622_),
    .A2(net4095));
 sg13g2_nand2_1 _39867_ (.Y(_13700_),
    .A(net2341),
    .B(net4866));
 sg13g2_o21ai_1 _39868_ (.B1(_13700_),
    .Y(_01219_),
    .A1(_14621_),
    .A2(net4095));
 sg13g2_nand2_1 _39869_ (.Y(_13701_),
    .A(net2021),
    .B(net4866));
 sg13g2_o21ai_1 _39870_ (.B1(_13701_),
    .Y(_01220_),
    .A1(_14620_),
    .A2(net4093));
 sg13g2_nand2_1 _39871_ (.Y(_13702_),
    .A(net2292),
    .B(net4866));
 sg13g2_o21ai_1 _39872_ (.B1(_13702_),
    .Y(_01221_),
    .A1(_14619_),
    .A2(net4093));
 sg13g2_nand2_1 _39873_ (.Y(_13703_),
    .A(net1343),
    .B(net4864));
 sg13g2_o21ai_1 _39874_ (.B1(_13703_),
    .Y(_01222_),
    .A1(_14618_),
    .A2(net4094));
 sg13g2_nand2_1 _39875_ (.Y(_13704_),
    .A(net1725),
    .B(net4864));
 sg13g2_o21ai_1 _39876_ (.B1(_13704_),
    .Y(_01223_),
    .A1(_14617_),
    .A2(net4095));
 sg13g2_nand2_1 _39877_ (.Y(_13705_),
    .A(net2462),
    .B(net4864));
 sg13g2_o21ai_1 _39878_ (.B1(_13705_),
    .Y(_01224_),
    .A1(_14616_),
    .A2(net4095));
 sg13g2_nand2_1 _39879_ (.Y(_13706_),
    .A(net2279),
    .B(net4864));
 sg13g2_o21ai_1 _39880_ (.B1(_13706_),
    .Y(_01225_),
    .A1(_14615_),
    .A2(net4096));
 sg13g2_nand2_1 _39881_ (.Y(_13707_),
    .A(net2305),
    .B(net4864));
 sg13g2_o21ai_1 _39882_ (.B1(_13707_),
    .Y(_01226_),
    .A1(_14614_),
    .A2(net4094));
 sg13g2_nand2_1 _39883_ (.Y(_13708_),
    .A(net2238),
    .B(net4854));
 sg13g2_o21ai_1 _39884_ (.B1(_13708_),
    .Y(_01227_),
    .A1(_14613_),
    .A2(net4089));
 sg13g2_nand2_1 _39885_ (.Y(_13709_),
    .A(net2257),
    .B(net4854));
 sg13g2_o21ai_1 _39886_ (.B1(_13709_),
    .Y(_01228_),
    .A1(_14612_),
    .A2(net4090));
 sg13g2_nand2_1 _39887_ (.Y(_13710_),
    .A(net2278),
    .B(net4854));
 sg13g2_o21ai_1 _39888_ (.B1(_13710_),
    .Y(_01229_),
    .A1(_14611_),
    .A2(net4087));
 sg13g2_nand2_1 _39889_ (.Y(_13711_),
    .A(net2938),
    .B(net4855));
 sg13g2_o21ai_1 _39890_ (.B1(_13711_),
    .Y(_01230_),
    .A1(_14610_),
    .A2(net4091));
 sg13g2_nand2_1 _39891_ (.Y(_13712_),
    .A(net2396),
    .B(net4854));
 sg13g2_o21ai_1 _39892_ (.B1(_13712_),
    .Y(_01231_),
    .A1(_14609_),
    .A2(net4090));
 sg13g2_nand2_1 _39893_ (.Y(_13713_),
    .A(net1711),
    .B(net4854));
 sg13g2_o21ai_1 _39894_ (.B1(_13713_),
    .Y(_01232_),
    .A1(_14608_),
    .A2(net4090));
 sg13g2_nand2_1 _39895_ (.Y(_13714_),
    .A(net2148),
    .B(net4854));
 sg13g2_o21ai_1 _39896_ (.B1(_13714_),
    .Y(_01233_),
    .A1(_14607_),
    .A2(net4090));
 sg13g2_nand2_1 _39897_ (.Y(_13715_),
    .A(net2457),
    .B(net4854));
 sg13g2_o21ai_1 _39898_ (.B1(_13715_),
    .Y(_01234_),
    .A1(_14606_),
    .A2(net4087));
 sg13g2_nand2_1 _39899_ (.Y(_13716_),
    .A(net2110),
    .B(net4854));
 sg13g2_o21ai_1 _39900_ (.B1(_13716_),
    .Y(_01235_),
    .A1(_14605_),
    .A2(net4090));
 sg13g2_nand2_1 _39901_ (.Y(_13717_),
    .A(net1145),
    .B(net4852));
 sg13g2_o21ai_1 _39902_ (.B1(_13717_),
    .Y(_01236_),
    .A1(_14604_),
    .A2(net4091));
 sg13g2_nand2_1 _39903_ (.Y(_13718_),
    .A(net2216),
    .B(net4853));
 sg13g2_o21ai_1 _39904_ (.B1(_13718_),
    .Y(_01237_),
    .A1(_14603_),
    .A2(net4089));
 sg13g2_nand2_1 _39905_ (.Y(_13719_),
    .A(net2691),
    .B(net4853));
 sg13g2_o21ai_1 _39906_ (.B1(_13719_),
    .Y(_01238_),
    .A1(_14602_),
    .A2(net4088));
 sg13g2_nand2_1 _39907_ (.Y(_13720_),
    .A(net2921),
    .B(net4853));
 sg13g2_o21ai_1 _39908_ (.B1(_13720_),
    .Y(_01239_),
    .A1(_14601_),
    .A2(net4089));
 sg13g2_nand2_1 _39909_ (.Y(_13721_),
    .A(net2737),
    .B(net4853));
 sg13g2_o21ai_1 _39910_ (.B1(_13721_),
    .Y(_01240_),
    .A1(_14600_),
    .A2(net4089));
 sg13g2_nand2_1 _39911_ (.Y(_13722_),
    .A(net2099),
    .B(net4853));
 sg13g2_o21ai_1 _39912_ (.B1(_13722_),
    .Y(_01241_),
    .A1(_14599_),
    .A2(net4089));
 sg13g2_nand2_1 _39913_ (.Y(_13723_),
    .A(net2496),
    .B(net4853));
 sg13g2_o21ai_1 _39914_ (.B1(_13723_),
    .Y(_01242_),
    .A1(_14598_),
    .A2(net4089));
 sg13g2_nand2_1 _39915_ (.Y(_13724_),
    .A(net1674),
    .B(net4853));
 sg13g2_o21ai_1 _39916_ (.B1(_13724_),
    .Y(_01243_),
    .A1(_14597_),
    .A2(net4089));
 sg13g2_nand2_1 _39917_ (.Y(_13725_),
    .A(net3177),
    .B(net4842));
 sg13g2_o21ai_1 _39918_ (.B1(_13725_),
    .Y(_01244_),
    .A1(_14596_),
    .A2(net4085));
 sg13g2_nand2_1 _39919_ (.Y(_13726_),
    .A(net3106),
    .B(net4842));
 sg13g2_o21ai_1 _39920_ (.B1(_13726_),
    .Y(_01245_),
    .A1(_14595_),
    .A2(net4085));
 sg13g2_nand2_1 _39921_ (.Y(_13727_),
    .A(net3095),
    .B(net4842));
 sg13g2_o21ai_1 _39922_ (.B1(_13727_),
    .Y(_01246_),
    .A1(_14594_),
    .A2(net4083));
 sg13g2_nand2_1 _39923_ (.Y(_13728_),
    .A(net2575),
    .B(net4842));
 sg13g2_o21ai_1 _39924_ (.B1(_13728_),
    .Y(_01247_),
    .A1(_14593_),
    .A2(net4085));
 sg13g2_nand2_1 _39925_ (.Y(_13729_),
    .A(net2060),
    .B(net4844));
 sg13g2_o21ai_1 _39926_ (.B1(_13729_),
    .Y(_01248_),
    .A1(_14592_),
    .A2(net4085));
 sg13g2_nand2_1 _39927_ (.Y(_13730_),
    .A(net2530),
    .B(net4842));
 sg13g2_o21ai_1 _39928_ (.B1(_13730_),
    .Y(_01249_),
    .A1(_14591_),
    .A2(net4085));
 sg13g2_nand2_1 _39929_ (.Y(_13731_),
    .A(net3091),
    .B(net4842));
 sg13g2_o21ai_1 _39930_ (.B1(_13731_),
    .Y(_01250_),
    .A1(_14590_),
    .A2(net4085));
 sg13g2_nand2_1 _39931_ (.Y(_13732_),
    .A(net2988),
    .B(net4842));
 sg13g2_o21ai_1 _39932_ (.B1(_13732_),
    .Y(_01251_),
    .A1(_14589_),
    .A2(net4086));
 sg13g2_nand2_1 _39933_ (.Y(_13733_),
    .A(net3187),
    .B(net4841));
 sg13g2_o21ai_1 _39934_ (.B1(_13733_),
    .Y(_01252_),
    .A1(_14588_),
    .A2(net4084));
 sg13g2_nand2_1 _39935_ (.Y(_13734_),
    .A(net2528),
    .B(net4841));
 sg13g2_o21ai_1 _39936_ (.B1(_13734_),
    .Y(_01253_),
    .A1(_14587_),
    .A2(net4084));
 sg13g2_nand2_1 _39937_ (.Y(_13735_),
    .A(net2887),
    .B(net4842));
 sg13g2_o21ai_1 _39938_ (.B1(_13735_),
    .Y(_01254_),
    .A1(_14586_),
    .A2(net4086));
 sg13g2_nand2_1 _39939_ (.Y(_13736_),
    .A(net2949),
    .B(net4841));
 sg13g2_o21ai_1 _39940_ (.B1(_13736_),
    .Y(_01255_),
    .A1(_14585_),
    .A2(net4084));
 sg13g2_nand2_1 _39941_ (.Y(_13737_),
    .A(net1331),
    .B(net4841));
 sg13g2_o21ai_1 _39942_ (.B1(_13737_),
    .Y(_01256_),
    .A1(_14584_),
    .A2(net4084));
 sg13g2_nand2_1 _39943_ (.Y(_13738_),
    .A(net2189),
    .B(net4834));
 sg13g2_o21ai_1 _39944_ (.B1(_13738_),
    .Y(_01257_),
    .A1(_14583_),
    .A2(net4080));
 sg13g2_nand2_1 _39945_ (.Y(_13739_),
    .A(net3226),
    .B(net4834));
 sg13g2_o21ai_1 _39946_ (.B1(_13739_),
    .Y(_01258_),
    .A1(_14582_),
    .A2(net4085));
 sg13g2_nand2_1 _39947_ (.Y(_13740_),
    .A(net2649),
    .B(net4835));
 sg13g2_o21ai_1 _39948_ (.B1(_13740_),
    .Y(_01259_),
    .A1(_14581_),
    .A2(net4080));
 sg13g2_nand2_1 _39949_ (.Y(_13741_),
    .A(net2628),
    .B(net4835));
 sg13g2_o21ai_1 _39950_ (.B1(_13741_),
    .Y(_01260_),
    .A1(_14580_),
    .A2(net4080));
 sg13g2_nand2_1 _39951_ (.Y(_13742_),
    .A(net2901),
    .B(net4834));
 sg13g2_o21ai_1 _39952_ (.B1(_13742_),
    .Y(_01261_),
    .A1(_14579_),
    .A2(net4080));
 sg13g2_nand2_1 _39953_ (.Y(_13743_),
    .A(net2573),
    .B(net4834));
 sg13g2_o21ai_1 _39954_ (.B1(_13743_),
    .Y(_01262_),
    .A1(_14578_),
    .A2(net4081));
 sg13g2_nand2_1 _39955_ (.Y(_13744_),
    .A(net2791),
    .B(net4834));
 sg13g2_o21ai_1 _39956_ (.B1(_13744_),
    .Y(_01263_),
    .A1(_14577_),
    .A2(net4081));
 sg13g2_nand2_1 _39957_ (.Y(_13745_),
    .A(net2571),
    .B(net4834));
 sg13g2_o21ai_1 _39958_ (.B1(_13745_),
    .Y(_01264_),
    .A1(_14576_),
    .A2(net4081));
 sg13g2_nand2_1 _39959_ (.Y(_13746_),
    .A(net2378),
    .B(net4836));
 sg13g2_o21ai_1 _39960_ (.B1(_13746_),
    .Y(_01265_),
    .A1(_14575_),
    .A2(net4079));
 sg13g2_nand2_1 _39961_ (.Y(_13747_),
    .A(net2485),
    .B(net4836));
 sg13g2_o21ai_1 _39962_ (.B1(_13747_),
    .Y(_01266_),
    .A1(_14574_),
    .A2(net4079));
 sg13g2_nand2_1 _39963_ (.Y(_13748_),
    .A(net3210),
    .B(net4831));
 sg13g2_o21ai_1 _39964_ (.B1(_13748_),
    .Y(_01267_),
    .A1(_14573_),
    .A2(net4079));
 sg13g2_nand2_1 _39965_ (.Y(_13749_),
    .A(net2603),
    .B(net4831));
 sg13g2_o21ai_1 _39966_ (.B1(_13749_),
    .Y(_01268_),
    .A1(_14572_),
    .A2(net4079));
 sg13g2_nand2_1 _39967_ (.Y(_13750_),
    .A(net2294),
    .B(net4831));
 sg13g2_o21ai_1 _39968_ (.B1(_13750_),
    .Y(_01269_),
    .A1(_14571_),
    .A2(net4079));
 sg13g2_nand2_1 _39969_ (.Y(_13751_),
    .A(net3022),
    .B(net4831));
 sg13g2_o21ai_1 _39970_ (.B1(_13751_),
    .Y(_01270_),
    .A1(_14570_),
    .A2(net4079));
 sg13g2_nand2_1 _39971_ (.Y(_13752_),
    .A(net2669),
    .B(net4831));
 sg13g2_o21ai_1 _39972_ (.B1(_13752_),
    .Y(_01271_),
    .A1(_14569_),
    .A2(net4075));
 sg13g2_nand2_1 _39973_ (.Y(_13753_),
    .A(net2236),
    .B(net4831));
 sg13g2_o21ai_1 _39974_ (.B1(_13753_),
    .Y(_01272_),
    .A1(_14568_),
    .A2(net4075));
 sg13g2_nand2_1 _39975_ (.Y(_13754_),
    .A(net2476),
    .B(net4831));
 sg13g2_o21ai_1 _39976_ (.B1(_13754_),
    .Y(_01273_),
    .A1(_14567_),
    .A2(net4075));
 sg13g2_nand2_1 _39977_ (.Y(_13755_),
    .A(net2917),
    .B(net4831));
 sg13g2_o21ai_1 _39978_ (.B1(_13755_),
    .Y(_01274_),
    .A1(_14566_),
    .A2(net4076));
 sg13g2_nand2_1 _39979_ (.Y(_13756_),
    .A(net1956),
    .B(net4832));
 sg13g2_o21ai_1 _39980_ (.B1(_13756_),
    .Y(_01275_),
    .A1(_14565_),
    .A2(net4076));
 sg13g2_nand2_1 _39981_ (.Y(_13757_),
    .A(net2150),
    .B(net4832));
 sg13g2_o21ai_1 _39982_ (.B1(_13757_),
    .Y(_01276_),
    .A1(_14564_),
    .A2(net4076));
 sg13g2_nand2_1 _39983_ (.Y(_13758_),
    .A(net2478),
    .B(net4832));
 sg13g2_o21ai_1 _39984_ (.B1(_13758_),
    .Y(_01277_),
    .A1(_14563_),
    .A2(net4075));
 sg13g2_nand2_1 _39985_ (.Y(_13759_),
    .A(net3012),
    .B(net4832));
 sg13g2_o21ai_1 _39986_ (.B1(_13759_),
    .Y(_01278_),
    .A1(_14562_),
    .A2(net4076));
 sg13g2_nand2_1 _39987_ (.Y(_13760_),
    .A(net2902),
    .B(net4832));
 sg13g2_o21ai_1 _39988_ (.B1(_13760_),
    .Y(_01279_),
    .A1(_14561_),
    .A2(net4075));
 sg13g2_nand2_1 _39989_ (.Y(_13761_),
    .A(net2265),
    .B(net4832));
 sg13g2_o21ai_1 _39990_ (.B1(_13761_),
    .Y(_01280_),
    .A1(_14560_),
    .A2(net4075));
 sg13g2_nand2_1 _39991_ (.Y(_13762_),
    .A(net2446),
    .B(net4832));
 sg13g2_o21ai_1 _39992_ (.B1(_13762_),
    .Y(_01281_),
    .A1(_14559_),
    .A2(net4075));
 sg13g2_nand2_1 _39993_ (.Y(_13763_),
    .A(net2658),
    .B(net4832));
 sg13g2_o21ai_1 _39994_ (.B1(_13763_),
    .Y(_01282_),
    .A1(_14558_),
    .A2(net4075));
 sg13g2_nand2_1 _39995_ (.Y(_13764_),
    .A(net2506),
    .B(net4833));
 sg13g2_o21ai_1 _39996_ (.B1(_13764_),
    .Y(_01283_),
    .A1(_14557_),
    .A2(net4077));
 sg13g2_nand2_1 _39997_ (.Y(_13765_),
    .A(net1419),
    .B(net4833));
 sg13g2_o21ai_1 _39998_ (.B1(_13765_),
    .Y(_01284_),
    .A1(_14556_),
    .A2(net4077));
 sg13g2_nand2_1 _39999_ (.Y(_13766_),
    .A(net2962),
    .B(net4833));
 sg13g2_o21ai_1 _40000_ (.B1(_13766_),
    .Y(_01285_),
    .A1(_14555_),
    .A2(net4077));
 sg13g2_nand2_1 _40001_ (.Y(_13767_),
    .A(net2018),
    .B(net4833));
 sg13g2_o21ai_1 _40002_ (.B1(_13767_),
    .Y(_01286_),
    .A1(_14554_),
    .A2(net4077));
 sg13g2_nand2_1 _40003_ (.Y(_13768_),
    .A(net2349),
    .B(net4833));
 sg13g2_o21ai_1 _40004_ (.B1(_13768_),
    .Y(_01287_),
    .A1(_14553_),
    .A2(net4078));
 sg13g2_nand2b_1 _40005_ (.Y(_01288_),
    .B(net4034),
    .A_N(net1196));
 sg13g2_a22oi_1 _40006_ (.Y(_01289_),
    .B1(net4839),
    .B2(_14170_),
    .A2(net4034),
    .A1(_14255_));
 sg13g2_a22oi_1 _40007_ (.Y(_01290_),
    .B1(net4839),
    .B2(_14169_),
    .A2(net4034),
    .A1(_14256_));
 sg13g2_a22oi_1 _40008_ (.Y(_01291_),
    .B1(net4839),
    .B2(_14168_),
    .A2(net4034),
    .A1(_14257_));
 sg13g2_nand2_1 _40009_ (.Y(_13769_),
    .A(net2355),
    .B(net4837));
 sg13g2_o21ai_1 _40010_ (.B1(_13769_),
    .Y(_01292_),
    .A1(_14258_),
    .A2(net4079));
 sg13g2_a22oi_1 _40011_ (.Y(_01293_),
    .B1(net4837),
    .B2(_14167_),
    .A2(net4034),
    .A1(_14259_));
 sg13g2_nand2_1 _40012_ (.Y(_13770_),
    .A(\u_inv.f_next[6] ),
    .B(net4837));
 sg13g2_o21ai_1 _40013_ (.B1(_13770_),
    .Y(_01294_),
    .A1(_14260_),
    .A2(net4079));
 sg13g2_nand2_1 _40014_ (.Y(_13771_),
    .A(net2608),
    .B(net4837));
 sg13g2_o21ai_1 _40015_ (.B1(_13771_),
    .Y(_01295_),
    .A1(_14261_),
    .A2(net4080));
 sg13g2_nand2_1 _40016_ (.Y(_13772_),
    .A(net1244),
    .B(net4837));
 sg13g2_o21ai_1 _40017_ (.B1(_13772_),
    .Y(_01296_),
    .A1(_14262_),
    .A2(net4080));
 sg13g2_nand2_1 _40018_ (.Y(_13773_),
    .A(net2526),
    .B(net4837));
 sg13g2_o21ai_1 _40019_ (.B1(_13773_),
    .Y(_01297_),
    .A1(_14263_),
    .A2(net4080));
 sg13g2_a22oi_1 _40020_ (.Y(_01298_),
    .B1(net4837),
    .B2(_14164_),
    .A2(net4034),
    .A1(_14264_));
 sg13g2_a22oi_1 _40021_ (.Y(_01299_),
    .B1(net4837),
    .B2(_14163_),
    .A2(net4034),
    .A1(_14265_));
 sg13g2_a22oi_1 _40022_ (.Y(_01300_),
    .B1(net4838),
    .B2(_14162_),
    .A2(net4032),
    .A1(_14266_));
 sg13g2_a22oi_1 _40023_ (.Y(_01301_),
    .B1(net4838),
    .B2(_14161_),
    .A2(net4032),
    .A1(_14267_));
 sg13g2_a22oi_1 _40024_ (.Y(_01302_),
    .B1(net4838),
    .B2(_14160_),
    .A2(net4032),
    .A1(_14268_));
 sg13g2_a22oi_1 _40025_ (.Y(_01303_),
    .B1(net4838),
    .B2(_14159_),
    .A2(net4033),
    .A1(_14269_));
 sg13g2_a22oi_1 _40026_ (.Y(_01304_),
    .B1(net4838),
    .B2(_14158_),
    .A2(net4032),
    .A1(_14270_));
 sg13g2_a22oi_1 _40027_ (.Y(_01305_),
    .B1(net4847),
    .B2(_14157_),
    .A2(net4037),
    .A1(_14271_));
 sg13g2_a22oi_1 _40028_ (.Y(_01306_),
    .B1(net4838),
    .B2(_14156_),
    .A2(net4032),
    .A1(_14272_));
 sg13g2_a22oi_1 _40029_ (.Y(_01307_),
    .B1(net4838),
    .B2(_14155_),
    .A2(net4032),
    .A1(_14273_));
 sg13g2_a22oi_1 _40030_ (.Y(_01308_),
    .B1(net4834),
    .B2(_14154_),
    .A2(net4032),
    .A1(_14274_));
 sg13g2_a22oi_1 _40031_ (.Y(_01309_),
    .B1(net4834),
    .B2(_14153_),
    .A2(net4032),
    .A1(_14275_));
 sg13g2_a22oi_1 _40032_ (.Y(_01310_),
    .B1(net4841),
    .B2(_14152_),
    .A2(net4037),
    .A1(_14276_));
 sg13g2_a22oi_1 _40033_ (.Y(_01311_),
    .B1(net4847),
    .B2(_14151_),
    .A2(net4037),
    .A1(_14277_));
 sg13g2_a22oi_1 _40034_ (.Y(_01312_),
    .B1(net4847),
    .B2(_14150_),
    .A2(net4037),
    .A1(_14278_));
 sg13g2_a22oi_1 _40035_ (.Y(_01313_),
    .B1(net4847),
    .B2(_14149_),
    .A2(net4037),
    .A1(_14279_));
 sg13g2_a22oi_1 _40036_ (.Y(_01314_),
    .B1(net4847),
    .B2(_14148_),
    .A2(net4037),
    .A1(_14280_));
 sg13g2_a22oi_1 _40037_ (.Y(_01315_),
    .B1(net4850),
    .B2(_14147_),
    .A2(net4040),
    .A1(_14281_));
 sg13g2_a22oi_1 _40038_ (.Y(_01316_),
    .B1(net4850),
    .B2(_14146_),
    .A2(net4040),
    .A1(_14282_));
 sg13g2_a22oi_1 _40039_ (.Y(_01317_),
    .B1(net4850),
    .B2(_14145_),
    .A2(net4040),
    .A1(_14283_));
 sg13g2_a22oi_1 _40040_ (.Y(_01318_),
    .B1(net4850),
    .B2(_14144_),
    .A2(net4040),
    .A1(_14284_));
 sg13g2_a22oi_1 _40041_ (.Y(_01319_),
    .B1(net4850),
    .B2(_14143_),
    .A2(net4040),
    .A1(_14285_));
 sg13g2_nand2_1 _40042_ (.Y(_13774_),
    .A(net1743),
    .B(net4850));
 sg13g2_o21ai_1 _40043_ (.B1(_13774_),
    .Y(_01320_),
    .A1(_14286_),
    .A2(net4089));
 sg13g2_a22oi_1 _40044_ (.Y(_01321_),
    .B1(net4857),
    .B2(_14141_),
    .A2(net4043),
    .A1(_14287_));
 sg13g2_a22oi_1 _40045_ (.Y(_01322_),
    .B1(net4857),
    .B2(_14140_),
    .A2(net4043),
    .A1(_14288_));
 sg13g2_a22oi_1 _40046_ (.Y(_01323_),
    .B1(net4857),
    .B2(_14139_),
    .A2(net4043),
    .A1(_14289_));
 sg13g2_a22oi_1 _40047_ (.Y(_01324_),
    .B1(net4857),
    .B2(_14138_),
    .A2(net4043),
    .A1(_14290_));
 sg13g2_a22oi_1 _40048_ (.Y(_01325_),
    .B1(net4857),
    .B2(_14137_),
    .A2(net4043),
    .A1(_14291_));
 sg13g2_a22oi_1 _40049_ (.Y(_01326_),
    .B1(net4857),
    .B2(_14136_),
    .A2(net4043),
    .A1(_14292_));
 sg13g2_a22oi_1 _40050_ (.Y(_01327_),
    .B1(net4857),
    .B2(_14135_),
    .A2(net4043),
    .A1(_14293_));
 sg13g2_a22oi_1 _40051_ (.Y(_01328_),
    .B1(net4860),
    .B2(_14134_),
    .A2(net4046),
    .A1(_14294_));
 sg13g2_a22oi_1 _40052_ (.Y(_01329_),
    .B1(net4860),
    .B2(_14133_),
    .A2(net4046),
    .A1(_14295_));
 sg13g2_a22oi_1 _40053_ (.Y(_01330_),
    .B1(net4860),
    .B2(_14132_),
    .A2(net4046),
    .A1(_14296_));
 sg13g2_a22oi_1 _40054_ (.Y(_01331_),
    .B1(net4860),
    .B2(_14131_),
    .A2(net4046),
    .A1(_14297_));
 sg13g2_a22oi_1 _40055_ (.Y(_01332_),
    .B1(net4860),
    .B2(_14130_),
    .A2(net4046),
    .A1(_14298_));
 sg13g2_a22oi_1 _40056_ (.Y(_01333_),
    .B1(net4860),
    .B2(_14129_),
    .A2(net4046),
    .A1(_14299_));
 sg13g2_a22oi_1 _40057_ (.Y(_01334_),
    .B1(net4870),
    .B2(_14128_),
    .A2(net4049),
    .A1(_14300_));
 sg13g2_a22oi_1 _40058_ (.Y(_01335_),
    .B1(net4870),
    .B2(_14127_),
    .A2(net4049),
    .A1(_14301_));
 sg13g2_a22oi_1 _40059_ (.Y(_01336_),
    .B1(net4870),
    .B2(_14126_),
    .A2(net4049),
    .A1(_14302_));
 sg13g2_a22oi_1 _40060_ (.Y(_01337_),
    .B1(net4870),
    .B2(_14125_),
    .A2(net4049),
    .A1(_14303_));
 sg13g2_a22oi_1 _40061_ (.Y(_01338_),
    .B1(net4873),
    .B2(_14124_),
    .A2(net4052),
    .A1(_14304_));
 sg13g2_a22oi_1 _40062_ (.Y(_01339_),
    .B1(net4873),
    .B2(_14123_),
    .A2(net4052),
    .A1(_14305_));
 sg13g2_a22oi_1 _40063_ (.Y(_01340_),
    .B1(net4873),
    .B2(_14122_),
    .A2(net4052),
    .A1(_14306_));
 sg13g2_a22oi_1 _40064_ (.Y(_01341_),
    .B1(net4873),
    .B2(_14121_),
    .A2(net4052),
    .A1(_14307_));
 sg13g2_a22oi_1 _40065_ (.Y(_01342_),
    .B1(net4873),
    .B2(_14120_),
    .A2(net4052),
    .A1(_14308_));
 sg13g2_a22oi_1 _40066_ (.Y(_01343_),
    .B1(net4873),
    .B2(_14119_),
    .A2(net4052),
    .A1(_14309_));
 sg13g2_a22oi_1 _40067_ (.Y(_01344_),
    .B1(net4881),
    .B2(_14118_),
    .A2(net4056),
    .A1(_14310_));
 sg13g2_a22oi_1 _40068_ (.Y(_01345_),
    .B1(net4881),
    .B2(_14117_),
    .A2(net4056),
    .A1(_14311_));
 sg13g2_a22oi_1 _40069_ (.Y(_01346_),
    .B1(net4881),
    .B2(_14116_),
    .A2(net4056),
    .A1(_14312_));
 sg13g2_a22oi_1 _40070_ (.Y(_01347_),
    .B1(net4881),
    .B2(_14115_),
    .A2(net4056),
    .A1(_14313_));
 sg13g2_a22oi_1 _40071_ (.Y(_01348_),
    .B1(net4881),
    .B2(_14114_),
    .A2(net4056),
    .A1(_14314_));
 sg13g2_a22oi_1 _40072_ (.Y(_01349_),
    .B1(net4881),
    .B2(_14113_),
    .A2(net4056),
    .A1(_14315_));
 sg13g2_a22oi_1 _40073_ (.Y(_01350_),
    .B1(net4883),
    .B2(_14112_),
    .A2(net4058),
    .A1(_14316_));
 sg13g2_a22oi_1 _40074_ (.Y(_01351_),
    .B1(net4881),
    .B2(_14111_),
    .A2(net4056),
    .A1(_14317_));
 sg13g2_a22oi_1 _40075_ (.Y(_01352_),
    .B1(net4883),
    .B2(_14110_),
    .A2(net4058),
    .A1(_14318_));
 sg13g2_a22oi_1 _40076_ (.Y(_01353_),
    .B1(net4883),
    .B2(_14109_),
    .A2(net4058),
    .A1(_14319_));
 sg13g2_a22oi_1 _40077_ (.Y(_01354_),
    .B1(net4883),
    .B2(_14108_),
    .A2(net4058),
    .A1(_14320_));
 sg13g2_a22oi_1 _40078_ (.Y(_01355_),
    .B1(net4883),
    .B2(_14107_),
    .A2(net4058),
    .A1(_14321_));
 sg13g2_a22oi_1 _40079_ (.Y(_01356_),
    .B1(net4883),
    .B2(_14106_),
    .A2(net4058),
    .A1(_14322_));
 sg13g2_a22oi_1 _40080_ (.Y(_01357_),
    .B1(net4883),
    .B2(_14105_),
    .A2(net4058),
    .A1(_14323_));
 sg13g2_a22oi_1 _40081_ (.Y(_01358_),
    .B1(net4893),
    .B2(_14104_),
    .A2(net4062),
    .A1(_14324_));
 sg13g2_a22oi_1 _40082_ (.Y(_01359_),
    .B1(net4883),
    .B2(_14103_),
    .A2(net4058),
    .A1(_14325_));
 sg13g2_a22oi_1 _40083_ (.Y(_01360_),
    .B1(net4893),
    .B2(_14102_),
    .A2(net4062),
    .A1(_14326_));
 sg13g2_a22oi_1 _40084_ (.Y(_01361_),
    .B1(net4893),
    .B2(_14101_),
    .A2(net4062),
    .A1(_14327_));
 sg13g2_a22oi_1 _40085_ (.Y(_01362_),
    .B1(net4893),
    .B2(_14100_),
    .A2(net4062),
    .A1(_14328_));
 sg13g2_a22oi_1 _40086_ (.Y(_01363_),
    .B1(net4895),
    .B2(_14099_),
    .A2(net4064),
    .A1(_14329_));
 sg13g2_a22oi_1 _40087_ (.Y(_01364_),
    .B1(net4895),
    .B2(_14098_),
    .A2(net4064),
    .A1(_14330_));
 sg13g2_a22oi_1 _40088_ (.Y(_01365_),
    .B1(net4895),
    .B2(_14097_),
    .A2(net4064),
    .A1(_14331_));
 sg13g2_a22oi_1 _40089_ (.Y(_01366_),
    .B1(net4895),
    .B2(_14096_),
    .A2(net4064),
    .A1(_14332_));
 sg13g2_a22oi_1 _40090_ (.Y(_01367_),
    .B1(net4895),
    .B2(_14095_),
    .A2(net4064),
    .A1(_14333_));
 sg13g2_a22oi_1 _40091_ (.Y(_01368_),
    .B1(net4903),
    .B2(_14094_),
    .A2(net4066),
    .A1(_14334_));
 sg13g2_a22oi_1 _40092_ (.Y(_01369_),
    .B1(net4903),
    .B2(_14093_),
    .A2(net4066),
    .A1(_14335_));
 sg13g2_a22oi_1 _40093_ (.Y(_01370_),
    .B1(net4903),
    .B2(_14092_),
    .A2(net4066),
    .A1(_14336_));
 sg13g2_a22oi_1 _40094_ (.Y(_01371_),
    .B1(net4903),
    .B2(_14091_),
    .A2(net4066),
    .A1(_14337_));
 sg13g2_a22oi_1 _40095_ (.Y(_01372_),
    .B1(net4904),
    .B2(_14090_),
    .A2(net4068),
    .A1(_14338_));
 sg13g2_a22oi_1 _40096_ (.Y(_01373_),
    .B1(net4904),
    .B2(_14089_),
    .A2(net4068),
    .A1(_14339_));
 sg13g2_a22oi_1 _40097_ (.Y(_01374_),
    .B1(net4904),
    .B2(_14088_),
    .A2(net4068),
    .A1(_14340_));
 sg13g2_a22oi_1 _40098_ (.Y(_01375_),
    .B1(net4904),
    .B2(_14087_),
    .A2(net4068),
    .A1(_14341_));
 sg13g2_a22oi_1 _40099_ (.Y(_01376_),
    .B1(net4915),
    .B2(_14086_),
    .A2(net4072),
    .A1(_14342_));
 sg13g2_a22oi_1 _40100_ (.Y(_01377_),
    .B1(net4915),
    .B2(_14085_),
    .A2(net4072),
    .A1(_14343_));
 sg13g2_a22oi_1 _40101_ (.Y(_01378_),
    .B1(net4915),
    .B2(_14084_),
    .A2(net4072),
    .A1(_14344_));
 sg13g2_a22oi_1 _40102_ (.Y(_01379_),
    .B1(net4915),
    .B2(_14083_),
    .A2(net4072),
    .A1(_14345_));
 sg13g2_a22oi_1 _40103_ (.Y(_01380_),
    .B1(net4915),
    .B2(_14082_),
    .A2(net4072),
    .A1(_14346_));
 sg13g2_a22oi_1 _40104_ (.Y(_01381_),
    .B1(net4915),
    .B2(_14081_),
    .A2(net4072),
    .A1(_14347_));
 sg13g2_a22oi_1 _40105_ (.Y(_01382_),
    .B1(net4915),
    .B2(_14080_),
    .A2(net4072),
    .A1(_14348_));
 sg13g2_a22oi_1 _40106_ (.Y(_01383_),
    .B1(net4914),
    .B2(_14079_),
    .A2(net4071),
    .A1(_14349_));
 sg13g2_a22oi_1 _40107_ (.Y(_01384_),
    .B1(net4914),
    .B2(_14078_),
    .A2(net4071),
    .A1(_14350_));
 sg13g2_a22oi_1 _40108_ (.Y(_01385_),
    .B1(net4914),
    .B2(_14077_),
    .A2(net4071),
    .A1(_14351_));
 sg13g2_a22oi_1 _40109_ (.Y(_01386_),
    .B1(net4914),
    .B2(_14076_),
    .A2(net4071),
    .A1(_14352_));
 sg13g2_a22oi_1 _40110_ (.Y(_01387_),
    .B1(net4914),
    .B2(_14075_),
    .A2(net4071),
    .A1(_14353_));
 sg13g2_a22oi_1 _40111_ (.Y(_01388_),
    .B1(net4916),
    .B2(_14074_),
    .A2(net4073),
    .A1(_14354_));
 sg13g2_a22oi_1 _40112_ (.Y(_01389_),
    .B1(net4916),
    .B2(_14073_),
    .A2(net4073),
    .A1(_14355_));
 sg13g2_a22oi_1 _40113_ (.Y(_01390_),
    .B1(net4914),
    .B2(_14072_),
    .A2(net4071),
    .A1(_14356_));
 sg13g2_a22oi_1 _40114_ (.Y(_01391_),
    .B1(net4914),
    .B2(_14071_),
    .A2(net4071),
    .A1(_14357_));
 sg13g2_a22oi_1 _40115_ (.Y(_01392_),
    .B1(net4912),
    .B2(_14070_),
    .A2(net4069),
    .A1(_14358_));
 sg13g2_a22oi_1 _40116_ (.Y(_01393_),
    .B1(net4912),
    .B2(_14069_),
    .A2(net4069),
    .A1(_14359_));
 sg13g2_a22oi_1 _40117_ (.Y(_01394_),
    .B1(net4914),
    .B2(_14068_),
    .A2(net4071),
    .A1(_14360_));
 sg13g2_a22oi_1 _40118_ (.Y(_01395_),
    .B1(net4913),
    .B2(_14067_),
    .A2(net4070),
    .A1(_14361_));
 sg13g2_a22oi_1 _40119_ (.Y(_01396_),
    .B1(net4912),
    .B2(_14066_),
    .A2(net4069),
    .A1(_14362_));
 sg13g2_a22oi_1 _40120_ (.Y(_01397_),
    .B1(net4913),
    .B2(_14065_),
    .A2(net4070),
    .A1(_14363_));
 sg13g2_a22oi_1 _40121_ (.Y(_01398_),
    .B1(net4912),
    .B2(_14064_),
    .A2(net4069),
    .A1(_14364_));
 sg13g2_a22oi_1 _40122_ (.Y(_01399_),
    .B1(net4913),
    .B2(_14063_),
    .A2(net4070),
    .A1(_14365_));
 sg13g2_a22oi_1 _40123_ (.Y(_01400_),
    .B1(net4912),
    .B2(_14062_),
    .A2(net4069),
    .A1(_14366_));
 sg13g2_a22oi_1 _40124_ (.Y(_01401_),
    .B1(net4912),
    .B2(_14061_),
    .A2(net4069),
    .A1(_14367_));
 sg13g2_a22oi_1 _40125_ (.Y(_01402_),
    .B1(net4912),
    .B2(_14060_),
    .A2(net4069),
    .A1(_14368_));
 sg13g2_a22oi_1 _40126_ (.Y(_01403_),
    .B1(net4912),
    .B2(_14059_),
    .A2(net4069),
    .A1(_14369_));
 sg13g2_a22oi_1 _40127_ (.Y(_01404_),
    .B1(net4905),
    .B2(_14058_),
    .A2(net4067),
    .A1(_14370_));
 sg13g2_a22oi_1 _40128_ (.Y(_01405_),
    .B1(net4906),
    .B2(_14057_),
    .A2(net4068),
    .A1(_14371_));
 sg13g2_a22oi_1 _40129_ (.Y(_01406_),
    .B1(net4906),
    .B2(_14056_),
    .A2(net4068),
    .A1(_14372_));
 sg13g2_a22oi_1 _40130_ (.Y(_01407_),
    .B1(net4906),
    .B2(_14055_),
    .A2(net4068),
    .A1(_14373_));
 sg13g2_a22oi_1 _40131_ (.Y(_01408_),
    .B1(net4905),
    .B2(_14054_),
    .A2(net4067),
    .A1(_14374_));
 sg13g2_a22oi_1 _40132_ (.Y(_01409_),
    .B1(net4905),
    .B2(_14053_),
    .A2(net4067),
    .A1(_14375_));
 sg13g2_a22oi_1 _40133_ (.Y(_01410_),
    .B1(net4905),
    .B2(_14052_),
    .A2(net4067),
    .A1(_14376_));
 sg13g2_a22oi_1 _40134_ (.Y(_01411_),
    .B1(net4905),
    .B2(_14051_),
    .A2(net4067),
    .A1(_14377_));
 sg13g2_a22oi_1 _40135_ (.Y(_01412_),
    .B1(net4905),
    .B2(_14050_),
    .A2(net4067),
    .A1(_14378_));
 sg13g2_a22oi_1 _40136_ (.Y(_01413_),
    .B1(net4905),
    .B2(_14049_),
    .A2(net4067),
    .A1(_14379_));
 sg13g2_a22oi_1 _40137_ (.Y(_01414_),
    .B1(net4905),
    .B2(_14048_),
    .A2(net4067),
    .A1(_14380_));
 sg13g2_a22oi_1 _40138_ (.Y(_01415_),
    .B1(net4903),
    .B2(_14047_),
    .A2(net4066),
    .A1(_14381_));
 sg13g2_a22oi_1 _40139_ (.Y(_01416_),
    .B1(net4902),
    .B2(_14046_),
    .A2(net4065),
    .A1(_14382_));
 sg13g2_a22oi_1 _40140_ (.Y(_01417_),
    .B1(net4902),
    .B2(_14045_),
    .A2(net4065),
    .A1(_14383_));
 sg13g2_a22oi_1 _40141_ (.Y(_01418_),
    .B1(net4902),
    .B2(_14044_),
    .A2(net4065),
    .A1(_14384_));
 sg13g2_a22oi_1 _40142_ (.Y(_01419_),
    .B1(net4902),
    .B2(_14043_),
    .A2(net4065),
    .A1(_14385_));
 sg13g2_a22oi_1 _40143_ (.Y(_01420_),
    .B1(net4902),
    .B2(_14042_),
    .A2(net4065),
    .A1(_14386_));
 sg13g2_a22oi_1 _40144_ (.Y(_01421_),
    .B1(net4902),
    .B2(_14041_),
    .A2(net4065),
    .A1(_14387_));
 sg13g2_a22oi_1 _40145_ (.Y(_01422_),
    .B1(net4902),
    .B2(_14040_),
    .A2(net4065),
    .A1(_14388_));
 sg13g2_a22oi_1 _40146_ (.Y(_01423_),
    .B1(net4902),
    .B2(_14039_),
    .A2(net4065),
    .A1(_14389_));
 sg13g2_a22oi_1 _40147_ (.Y(_01424_),
    .B1(net4894),
    .B2(_14038_),
    .A2(net4063),
    .A1(_14390_));
 sg13g2_a22oi_1 _40148_ (.Y(_01425_),
    .B1(net4894),
    .B2(_14037_),
    .A2(net4063),
    .A1(_14391_));
 sg13g2_a22oi_1 _40149_ (.Y(_01426_),
    .B1(net4894),
    .B2(_14036_),
    .A2(net4063),
    .A1(_14392_));
 sg13g2_a22oi_1 _40150_ (.Y(_01427_),
    .B1(net4894),
    .B2(_14035_),
    .A2(net4063),
    .A1(_14393_));
 sg13g2_a22oi_1 _40151_ (.Y(_01428_),
    .B1(net4894),
    .B2(_14034_),
    .A2(net4064),
    .A1(_14394_));
 sg13g2_a22oi_1 _40152_ (.Y(_01429_),
    .B1(net4895),
    .B2(_14033_),
    .A2(net4063),
    .A1(_14395_));
 sg13g2_a22oi_1 _40153_ (.Y(_01430_),
    .B1(net4894),
    .B2(_14032_),
    .A2(net4063),
    .A1(_14396_));
 sg13g2_a22oi_1 _40154_ (.Y(_01431_),
    .B1(net4894),
    .B2(_14031_),
    .A2(net4063),
    .A1(_14397_));
 sg13g2_a22oi_1 _40155_ (.Y(_01432_),
    .B1(net4894),
    .B2(_14030_),
    .A2(net4063),
    .A1(_14398_));
 sg13g2_a22oi_1 _40156_ (.Y(_01433_),
    .B1(net4892),
    .B2(_14029_),
    .A2(net4061),
    .A1(_14399_));
 sg13g2_a22oi_1 _40157_ (.Y(_01434_),
    .B1(net4893),
    .B2(_14028_),
    .A2(net4062),
    .A1(_14400_));
 sg13g2_a22oi_1 _40158_ (.Y(_01435_),
    .B1(net4893),
    .B2(_14027_),
    .A2(net4062),
    .A1(_14401_));
 sg13g2_a22oi_1 _40159_ (.Y(_01436_),
    .B1(net4892),
    .B2(_14026_),
    .A2(net4062),
    .A1(_14402_));
 sg13g2_a22oi_1 _40160_ (.Y(_01437_),
    .B1(net4892),
    .B2(_14025_),
    .A2(net4061),
    .A1(_14403_));
 sg13g2_a22oi_1 _40161_ (.Y(_01438_),
    .B1(net4892),
    .B2(_14024_),
    .A2(net4061),
    .A1(_14404_));
 sg13g2_a22oi_1 _40162_ (.Y(_01439_),
    .B1(net4892),
    .B2(_14023_),
    .A2(net4061),
    .A1(_14405_));
 sg13g2_a22oi_1 _40163_ (.Y(_01440_),
    .B1(net4893),
    .B2(_14022_),
    .A2(net4061),
    .A1(_14406_));
 sg13g2_a22oi_1 _40164_ (.Y(_01441_),
    .B1(net4892),
    .B2(_14021_),
    .A2(net4061),
    .A1(_14407_));
 sg13g2_a22oi_1 _40165_ (.Y(_01442_),
    .B1(net4884),
    .B2(_14020_),
    .A2(net4059),
    .A1(_14408_));
 sg13g2_a22oi_1 _40166_ (.Y(_01443_),
    .B1(net4892),
    .B2(_14019_),
    .A2(net4061),
    .A1(_14409_));
 sg13g2_a22oi_1 _40167_ (.Y(_01444_),
    .B1(net4882),
    .B2(_14018_),
    .A2(net4057),
    .A1(_14410_));
 sg13g2_a22oi_1 _40168_ (.Y(_01445_),
    .B1(net4884),
    .B2(_14017_),
    .A2(net4059),
    .A1(_14411_));
 sg13g2_a22oi_1 _40169_ (.Y(_01446_),
    .B1(net4884),
    .B2(_14016_),
    .A2(net4059),
    .A1(_14412_));
 sg13g2_a22oi_1 _40170_ (.Y(_01447_),
    .B1(net4892),
    .B2(_14015_),
    .A2(net4061),
    .A1(_14413_));
 sg13g2_a22oi_1 _40171_ (.Y(_01448_),
    .B1(net4882),
    .B2(_14014_),
    .A2(net4057),
    .A1(_14414_));
 sg13g2_a22oi_1 _40172_ (.Y(_01449_),
    .B1(net4882),
    .B2(_14013_),
    .A2(net4057),
    .A1(_14415_));
 sg13g2_a22oi_1 _40173_ (.Y(_01450_),
    .B1(net4882),
    .B2(_14012_),
    .A2(net4057),
    .A1(_14416_));
 sg13g2_a22oi_1 _40174_ (.Y(_01451_),
    .B1(net4882),
    .B2(_14011_),
    .A2(net4057),
    .A1(_14417_));
 sg13g2_a22oi_1 _40175_ (.Y(_01452_),
    .B1(net4882),
    .B2(_14010_),
    .A2(net4057),
    .A1(_14418_));
 sg13g2_a22oi_1 _40176_ (.Y(_01453_),
    .B1(net4880),
    .B2(_14009_),
    .A2(net4055),
    .A1(_14419_));
 sg13g2_a22oi_1 _40177_ (.Y(_01454_),
    .B1(net4882),
    .B2(_14008_),
    .A2(net4057),
    .A1(_14420_));
 sg13g2_a22oi_1 _40178_ (.Y(_01455_),
    .B1(net4882),
    .B2(_14007_),
    .A2(net4057),
    .A1(_14421_));
 sg13g2_a22oi_1 _40179_ (.Y(_01456_),
    .B1(net4880),
    .B2(_14006_),
    .A2(net4055),
    .A1(_14422_));
 sg13g2_a22oi_1 _40180_ (.Y(_01457_),
    .B1(net4880),
    .B2(_14005_),
    .A2(net4055),
    .A1(_14423_));
 sg13g2_a22oi_1 _40181_ (.Y(_01458_),
    .B1(net4885),
    .B2(_14004_),
    .A2(net4060),
    .A1(_14424_));
 sg13g2_a22oi_1 _40182_ (.Y(_01459_),
    .B1(net4885),
    .B2(_14003_),
    .A2(net4060),
    .A1(_14425_));
 sg13g2_a22oi_1 _40183_ (.Y(_01460_),
    .B1(net4880),
    .B2(_14002_),
    .A2(net4055),
    .A1(_14426_));
 sg13g2_a22oi_1 _40184_ (.Y(_01461_),
    .B1(net4880),
    .B2(_14001_),
    .A2(net4055),
    .A1(_14427_));
 sg13g2_a22oi_1 _40185_ (.Y(_01462_),
    .B1(net4880),
    .B2(_14000_),
    .A2(net4055),
    .A1(_14428_));
 sg13g2_a22oi_1 _40186_ (.Y(_01463_),
    .B1(net4880),
    .B2(_13999_),
    .A2(net4055),
    .A1(_14429_));
 sg13g2_a22oi_1 _40187_ (.Y(_01464_),
    .B1(net4871),
    .B2(_13998_),
    .A2(net4050),
    .A1(_14430_));
 sg13g2_a22oi_1 _40188_ (.Y(_01465_),
    .B1(net4872),
    .B2(_13997_),
    .A2(net4050),
    .A1(_14431_));
 sg13g2_a22oi_1 _40189_ (.Y(_01466_),
    .B1(net4880),
    .B2(_13996_),
    .A2(net4055),
    .A1(_14432_));
 sg13g2_a22oi_1 _40190_ (.Y(_01467_),
    .B1(net4872),
    .B2(_13995_),
    .A2(net4051),
    .A1(_14433_));
 sg13g2_a22oi_1 _40191_ (.Y(_01468_),
    .B1(net4872),
    .B2(_13994_),
    .A2(net4051),
    .A1(_14434_));
 sg13g2_a22oi_1 _40192_ (.Y(_01469_),
    .B1(net4872),
    .B2(_13993_),
    .A2(net4051),
    .A1(_14435_));
 sg13g2_a22oi_1 _40193_ (.Y(_01470_),
    .B1(net4872),
    .B2(_13992_),
    .A2(net4051),
    .A1(_14436_));
 sg13g2_a22oi_1 _40194_ (.Y(_01471_),
    .B1(net4872),
    .B2(_13991_),
    .A2(net4051),
    .A1(_14437_));
 sg13g2_a22oi_1 _40195_ (.Y(_01472_),
    .B1(net4871),
    .B2(_13990_),
    .A2(net4050),
    .A1(_14438_));
 sg13g2_a22oi_1 _40196_ (.Y(_01473_),
    .B1(net4871),
    .B2(_13989_),
    .A2(net4050),
    .A1(_14439_));
 sg13g2_a22oi_1 _40197_ (.Y(_01474_),
    .B1(net4871),
    .B2(_13988_),
    .A2(net4050),
    .A1(_14440_));
 sg13g2_a22oi_1 _40198_ (.Y(_01475_),
    .B1(net4871),
    .B2(_13987_),
    .A2(net4050),
    .A1(_14441_));
 sg13g2_a22oi_1 _40199_ (.Y(_01476_),
    .B1(net4871),
    .B2(_13986_),
    .A2(net4048),
    .A1(_14442_));
 sg13g2_a22oi_1 _40200_ (.Y(_01477_),
    .B1(net4869),
    .B2(_13985_),
    .A2(net4048),
    .A1(_14443_));
 sg13g2_a22oi_1 _40201_ (.Y(_01478_),
    .B1(net4871),
    .B2(_13984_),
    .A2(net4050),
    .A1(_14444_));
 sg13g2_a22oi_1 _40202_ (.Y(_01479_),
    .B1(net4871),
    .B2(_13983_),
    .A2(net4050),
    .A1(_14445_));
 sg13g2_a22oi_1 _40203_ (.Y(_01480_),
    .B1(net4868),
    .B2(_13982_),
    .A2(net4047),
    .A1(_14446_));
 sg13g2_a22oi_1 _40204_ (.Y(_01481_),
    .B1(net4869),
    .B2(_13981_),
    .A2(net4048),
    .A1(_14447_));
 sg13g2_a22oi_1 _40205_ (.Y(_01482_),
    .B1(net4869),
    .B2(_13980_),
    .A2(net4048),
    .A1(_14448_));
 sg13g2_a22oi_1 _40206_ (.Y(_01483_),
    .B1(net4869),
    .B2(_13979_),
    .A2(net4048),
    .A1(_14449_));
 sg13g2_a22oi_1 _40207_ (.Y(_01484_),
    .B1(net4868),
    .B2(_13978_),
    .A2(net4047),
    .A1(_14450_));
 sg13g2_a22oi_1 _40208_ (.Y(_01485_),
    .B1(net4868),
    .B2(_13977_),
    .A2(net4047),
    .A1(_14451_));
 sg13g2_a22oi_1 _40209_ (.Y(_01486_),
    .B1(net4868),
    .B2(_13976_),
    .A2(net4047),
    .A1(_14452_));
 sg13g2_a22oi_1 _40210_ (.Y(_01487_),
    .B1(net4868),
    .B2(_13975_),
    .A2(net4047),
    .A1(_14453_));
 sg13g2_a22oi_1 _40211_ (.Y(_01488_),
    .B1(net4868),
    .B2(_13974_),
    .A2(net4047),
    .A1(_14454_));
 sg13g2_a22oi_1 _40212_ (.Y(_01489_),
    .B1(net4868),
    .B2(_13973_),
    .A2(net4047),
    .A1(_14455_));
 sg13g2_a22oi_1 _40213_ (.Y(_01490_),
    .B1(net4859),
    .B2(_13972_),
    .A2(net4045),
    .A1(_14456_));
 sg13g2_a22oi_1 _40214_ (.Y(_01491_),
    .B1(net4859),
    .B2(_13971_),
    .A2(net4045),
    .A1(_14457_));
 sg13g2_a22oi_1 _40215_ (.Y(_01492_),
    .B1(net4868),
    .B2(_13970_),
    .A2(net4047),
    .A1(_14458_));
 sg13g2_a22oi_1 _40216_ (.Y(_01493_),
    .B1(net4859),
    .B2(_13969_),
    .A2(net4045),
    .A1(_14459_));
 sg13g2_a22oi_1 _40217_ (.Y(_01494_),
    .B1(net4858),
    .B2(_13968_),
    .A2(net4044),
    .A1(_14460_));
 sg13g2_a22oi_1 _40218_ (.Y(_01495_),
    .B1(net4859),
    .B2(_13967_),
    .A2(net4045),
    .A1(_14461_));
 sg13g2_a22oi_1 _40219_ (.Y(_01496_),
    .B1(net4858),
    .B2(_13966_),
    .A2(net4044),
    .A1(_14462_));
 sg13g2_a22oi_1 _40220_ (.Y(_01497_),
    .B1(net4858),
    .B2(_13965_),
    .A2(net4044),
    .A1(_14463_));
 sg13g2_a22oi_1 _40221_ (.Y(_01498_),
    .B1(net4859),
    .B2(_13964_),
    .A2(net4044),
    .A1(_14464_));
 sg13g2_a22oi_1 _40222_ (.Y(_01499_),
    .B1(net4858),
    .B2(_13963_),
    .A2(net4044),
    .A1(_14465_));
 sg13g2_a22oi_1 _40223_ (.Y(_01500_),
    .B1(net4858),
    .B2(_13962_),
    .A2(net4044),
    .A1(_14466_));
 sg13g2_a22oi_1 _40224_ (.Y(_01501_),
    .B1(net4858),
    .B2(_13961_),
    .A2(net4044),
    .A1(_14467_));
 sg13g2_a22oi_1 _40225_ (.Y(_01502_),
    .B1(net4856),
    .B2(_13960_),
    .A2(net4041),
    .A1(_14468_));
 sg13g2_a22oi_1 _40226_ (.Y(_01503_),
    .B1(net4858),
    .B2(_13959_),
    .A2(net4041),
    .A1(_14469_));
 sg13g2_a22oi_1 _40227_ (.Y(_01504_),
    .B1(net4858),
    .B2(_13958_),
    .A2(net4044),
    .A1(_14470_));
 sg13g2_a22oi_1 _40228_ (.Y(_01505_),
    .B1(net4861),
    .B2(_13957_),
    .A2(net4042),
    .A1(_14471_));
 sg13g2_a22oi_1 _40229_ (.Y(_01506_),
    .B1(net4861),
    .B2(_13956_),
    .A2(net4042),
    .A1(_14472_));
 sg13g2_a22oi_1 _40230_ (.Y(_01507_),
    .B1(net4861),
    .B2(_13955_),
    .A2(net4042),
    .A1(_14473_));
 sg13g2_a22oi_1 _40231_ (.Y(_01508_),
    .B1(net4856),
    .B2(_13954_),
    .A2(net4041),
    .A1(_14474_));
 sg13g2_a22oi_1 _40232_ (.Y(_01509_),
    .B1(net4856),
    .B2(_13953_),
    .A2(net4042),
    .A1(_14475_));
 sg13g2_a22oi_1 _40233_ (.Y(_01510_),
    .B1(net4856),
    .B2(_13952_),
    .A2(net4041),
    .A1(_14476_));
 sg13g2_a22oi_1 _40234_ (.Y(_01511_),
    .B1(net4856),
    .B2(_13951_),
    .A2(net4041),
    .A1(_14477_));
 sg13g2_a22oi_1 _40235_ (.Y(_01512_),
    .B1(net4856),
    .B2(_13950_),
    .A2(net4041),
    .A1(_14478_));
 sg13g2_a22oi_1 _40236_ (.Y(_01513_),
    .B1(net4856),
    .B2(_13949_),
    .A2(net4041),
    .A1(_14479_));
 sg13g2_a22oi_1 _40237_ (.Y(_01514_),
    .B1(net4849),
    .B2(_13948_),
    .A2(net4039),
    .A1(_14480_));
 sg13g2_a22oi_1 _40238_ (.Y(_01515_),
    .B1(net4849),
    .B2(_13947_),
    .A2(net4039),
    .A1(_14481_));
 sg13g2_a22oi_1 _40239_ (.Y(_01516_),
    .B1(net4856),
    .B2(_13946_),
    .A2(net4041),
    .A1(_14482_));
 sg13g2_a22oi_1 _40240_ (.Y(_01517_),
    .B1(net4849),
    .B2(_13945_),
    .A2(net4039),
    .A1(_14483_));
 sg13g2_a22oi_1 _40241_ (.Y(_01518_),
    .B1(net4849),
    .B2(_13944_),
    .A2(net4039),
    .A1(_14484_));
 sg13g2_a22oi_1 _40242_ (.Y(_01519_),
    .B1(net4849),
    .B2(_13943_),
    .A2(net4039),
    .A1(_14485_));
 sg13g2_a22oi_1 _40243_ (.Y(_01520_),
    .B1(net4848),
    .B2(_13942_),
    .A2(net4038),
    .A1(_14486_));
 sg13g2_a22oi_1 _40244_ (.Y(_01521_),
    .B1(net4848),
    .B2(_13941_),
    .A2(net4038),
    .A1(_14487_));
 sg13g2_a22oi_1 _40245_ (.Y(_01522_),
    .B1(net4848),
    .B2(_13940_),
    .A2(net4038),
    .A1(_14488_));
 sg13g2_a22oi_1 _40246_ (.Y(_01523_),
    .B1(net4848),
    .B2(_13939_),
    .A2(net4038),
    .A1(_14489_));
 sg13g2_a22oi_1 _40247_ (.Y(_01524_),
    .B1(net4848),
    .B2(_13938_),
    .A2(net4038),
    .A1(_14490_));
 sg13g2_a22oi_1 _40248_ (.Y(_01525_),
    .B1(net4848),
    .B2(_13937_),
    .A2(net4038),
    .A1(_14491_));
 sg13g2_a22oi_1 _40249_ (.Y(_01526_),
    .B1(net4848),
    .B2(_13936_),
    .A2(net4038),
    .A1(_14492_));
 sg13g2_a22oi_1 _40250_ (.Y(_01527_),
    .B1(net4848),
    .B2(_13935_),
    .A2(net4038),
    .A1(_14493_));
 sg13g2_a22oi_1 _40251_ (.Y(_01528_),
    .B1(net4845),
    .B2(_13934_),
    .A2(net4035),
    .A1(_14494_));
 sg13g2_a22oi_1 _40252_ (.Y(_01529_),
    .B1(net4846),
    .B2(_13933_),
    .A2(net4035),
    .A1(_14495_));
 sg13g2_a22oi_1 _40253_ (.Y(_01530_),
    .B1(net4846),
    .B2(_13932_),
    .A2(net4036),
    .A1(_14496_));
 sg13g2_a22oi_1 _40254_ (.Y(_01531_),
    .B1(net4846),
    .B2(_13931_),
    .A2(net4036),
    .A1(_14497_));
 sg13g2_a22oi_1 _40255_ (.Y(_01532_),
    .B1(net4846),
    .B2(_13930_),
    .A2(net4036),
    .A1(_14498_));
 sg13g2_a22oi_1 _40256_ (.Y(_01533_),
    .B1(net4846),
    .B2(_13929_),
    .A2(net4036),
    .A1(_14499_));
 sg13g2_a22oi_1 _40257_ (.Y(_01534_),
    .B1(net4845),
    .B2(_13928_),
    .A2(net4035),
    .A1(_14500_));
 sg13g2_a22oi_1 _40258_ (.Y(_01535_),
    .B1(net4845),
    .B2(_13927_),
    .A2(net4035),
    .A1(_14501_));
 sg13g2_a22oi_1 _40259_ (.Y(_01536_),
    .B1(net4845),
    .B2(_13926_),
    .A2(net4033),
    .A1(_14502_));
 sg13g2_a22oi_1 _40260_ (.Y(_01537_),
    .B1(net4838),
    .B2(_13925_),
    .A2(net4033),
    .A1(_14503_));
 sg13g2_a22oi_1 _40261_ (.Y(_01538_),
    .B1(net4839),
    .B2(_13924_),
    .A2(net4033),
    .A1(_14504_));
 sg13g2_a22oi_1 _40262_ (.Y(_01539_),
    .B1(net4839),
    .B2(_13923_),
    .A2(net4033),
    .A1(_14505_));
 sg13g2_a22oi_1 _40263_ (.Y(_01540_),
    .B1(net4845),
    .B2(_13922_),
    .A2(net4035),
    .A1(_14506_));
 sg13g2_a22oi_1 _40264_ (.Y(_01541_),
    .B1(net4845),
    .B2(_13921_),
    .A2(net4035),
    .A1(_14507_));
 sg13g2_a22oi_1 _40265_ (.Y(_01542_),
    .B1(net4845),
    .B2(_13920_),
    .A2(net4035),
    .A1(_14508_));
 sg13g2_a22oi_1 _40266_ (.Y(_01543_),
    .B1(net4845),
    .B2(_13919_),
    .A2(net4035),
    .A1(_14509_));
 sg13g2_nand2_2 _40267_ (.Y(_13775_),
    .A(net2316),
    .B(net4846));
 sg13g2_o21ai_1 _40268_ (.B1(_13775_),
    .Y(_01544_),
    .A1(net5637),
    .A2(net4085));
 sg13g2_nand2b_1 _40269_ (.Y(_01545_),
    .B(_19025_),
    .A_N(_19024_));
 sg13g2_a21oi_1 _40270_ (.A1(net5628),
    .A2(_19017_),
    .Y(_01546_),
    .B1(_19024_));
 sg13g2_nor2_1 _40271_ (.A(net1172),
    .B(net5236),
    .Y(_13776_));
 sg13g2_a21oi_1 _40272_ (.A1(_14248_),
    .A2(net5235),
    .Y(_01547_),
    .B1(_13776_));
 sg13g2_nor2_1 _40273_ (.A(net1273),
    .B(net5235),
    .Y(_13777_));
 sg13g2_a21oi_1 _40274_ (.A1(_14249_),
    .A2(net5235),
    .Y(_01548_),
    .B1(_13777_));
 sg13g2_mux2_1 _40275_ (.A0(net1656),
    .A1(net5881),
    .S(net5235),
    .X(_01549_));
 sg13g2_nor2_1 _40276_ (.A(net1124),
    .B(net5235),
    .Y(_13778_));
 sg13g2_a21oi_1 _40277_ (.A1(_14250_),
    .A2(net5235),
    .Y(_01550_),
    .B1(_13778_));
 sg13g2_mux2_1 _40278_ (.A0(net1411),
    .A1(\u_inv.counter[4] ),
    .S(net5236),
    .X(_01551_));
 sg13g2_nor2_1 _40279_ (.A(net1270),
    .B(net5236),
    .Y(_13779_));
 sg13g2_a21oi_1 _40280_ (.A1(_14253_),
    .A2(net5236),
    .Y(_01552_),
    .B1(_13779_));
 sg13g2_nor2_1 _40281_ (.A(net1364),
    .B(net5237),
    .Y(_13780_));
 sg13g2_a21oi_1 _40282_ (.A1(_14252_),
    .A2(net5237),
    .Y(_01553_),
    .B1(_13780_));
 sg13g2_nor2_1 _40283_ (.A(net1237),
    .B(net5235),
    .Y(_13781_));
 sg13g2_a21oi_1 _40284_ (.A1(_14251_),
    .A2(net5235),
    .Y(_01554_),
    .B1(_13781_));
 sg13g2_nor2_1 _40285_ (.A(net1132),
    .B(net5237),
    .Y(_13782_));
 sg13g2_a21oi_1 _40286_ (.A1(_14254_),
    .A2(net5237),
    .Y(_01555_),
    .B1(_13782_));
 sg13g2_mux2_1 _40287_ (.A0(net1442),
    .A1(\u_inv.counter[9] ),
    .S(net5237),
    .X(_01556_));
 sg13g2_xnor2_1 _40288_ (.Y(_13783_),
    .A(_14244_),
    .B(net4446));
 sg13g2_a22oi_1 _40289_ (.Y(_01557_),
    .B1(_13783_),
    .B2(net5612),
    .A2(net4244),
    .A1(_14244_));
 sg13g2_o21ai_1 _40290_ (.B1(_15967_),
    .Y(_13784_),
    .A1(\u_inv.delta_double[0] ),
    .A2(net4448));
 sg13g2_nand2_1 _40291_ (.Y(_13785_),
    .A(net2083),
    .B(net4244));
 sg13g2_xor2_1 _40292_ (.B(_13784_),
    .A(net2083),
    .X(_13786_));
 sg13g2_o21ai_1 _40293_ (.B1(_13785_),
    .Y(_01558_),
    .A1(net5579),
    .A2(_13786_));
 sg13g2_nor2b_1 _40294_ (.A(\u_inv.delta_double[0] ),
    .B_N(net2083),
    .Y(_13787_));
 sg13g2_o21ai_1 _40295_ (.B1(net2083),
    .Y(_13788_),
    .A1(\u_inv.delta_double[0] ),
    .A2(_15966_));
 sg13g2_xnor2_1 _40296_ (.Y(_13789_),
    .A(net2842),
    .B(_13788_));
 sg13g2_nand2_1 _40297_ (.Y(_13790_),
    .A(_13787_),
    .B(_13789_));
 sg13g2_nor2_1 _40298_ (.A(net4372),
    .B(_13790_),
    .Y(_13791_));
 sg13g2_a21oi_1 _40299_ (.A1(net4446),
    .A2(_13787_),
    .Y(_13792_),
    .B1(_13789_));
 sg13g2_nor3_1 _40300_ (.A(net5579),
    .B(_13791_),
    .C(_13792_),
    .Y(_13793_));
 sg13g2_a21o_1 _40301_ (.A2(net4244),
    .A1(net2842),
    .B1(_13793_),
    .X(_01559_));
 sg13g2_nand2_1 _40302_ (.Y(_13794_),
    .A(net2198),
    .B(net4245));
 sg13g2_and3_1 _40303_ (.X(_13795_),
    .A(\u_inv.delta_double[0] ),
    .B(\u_inv.delta_reg[1] ),
    .C(\u_inv.delta_reg[2] ));
 sg13g2_a21oi_1 _40304_ (.A1(_15960_),
    .A2(net5009),
    .Y(_13796_),
    .B1(_13795_));
 sg13g2_xnor2_1 _40305_ (.Y(_13797_),
    .A(net2198),
    .B(_13796_));
 sg13g2_nor2_1 _40306_ (.A(_13791_),
    .B(_13797_),
    .Y(_13798_));
 sg13g2_nor2b_1 _40307_ (.A(_13790_),
    .B_N(_13797_),
    .Y(_13799_));
 sg13g2_nand2_1 _40308_ (.Y(_13800_),
    .A(net4448),
    .B(_13799_));
 sg13g2_nand2_1 _40309_ (.Y(_13801_),
    .A(net5613),
    .B(_13800_));
 sg13g2_o21ai_1 _40310_ (.B1(_13794_),
    .Y(_01560_),
    .A1(_13798_),
    .A2(_13801_));
 sg13g2_a21oi_1 _40311_ (.A1(\u_inv.delta_reg[3] ),
    .A2(_13795_),
    .Y(_13802_),
    .B1(\u_inv.delta_reg[4] ));
 sg13g2_and3_2 _40312_ (.X(_13803_),
    .A(\u_inv.delta_reg[3] ),
    .B(\u_inv.delta_reg[4] ),
    .C(_13795_));
 sg13g2_nor2_1 _40313_ (.A(_13802_),
    .B(_13803_),
    .Y(_13804_));
 sg13g2_o21ai_1 _40314_ (.B1(\u_inv.delta_reg[4] ),
    .Y(_13805_),
    .A1(\u_inv.delta_reg[3] ),
    .A2(_15960_));
 sg13g2_nor2_1 _40315_ (.A(_15961_),
    .B(net5095),
    .Y(_13806_));
 sg13g2_a22oi_1 _40316_ (.Y(_13807_),
    .B1(_13805_),
    .B2(_13806_),
    .A2(_13804_),
    .A1(net5095));
 sg13g2_or2_1 _40317_ (.X(_13808_),
    .B(_13807_),
    .A(_13800_));
 sg13g2_a21oi_1 _40318_ (.A1(_13800_),
    .A2(_13807_),
    .Y(_13809_),
    .B1(net5582));
 sg13g2_a22oi_1 _40319_ (.Y(_13810_),
    .B1(_13808_),
    .B2(_13809_),
    .A2(net4244),
    .A1(net2866));
 sg13g2_inv_1 _40320_ (.Y(_01561_),
    .A(_13810_));
 sg13g2_nor2_1 _40321_ (.A(_13803_),
    .B(_13806_),
    .Y(_13811_));
 sg13g2_xnor2_1 _40322_ (.Y(_13812_),
    .A(_14245_),
    .B(_13811_));
 sg13g2_nor2_1 _40323_ (.A(_13807_),
    .B(_13812_),
    .Y(_13813_));
 sg13g2_nand3_1 _40324_ (.B(_13799_),
    .C(_13813_),
    .A(net4448),
    .Y(_13814_));
 sg13g2_a21oi_1 _40325_ (.A1(_13808_),
    .A2(_13812_),
    .Y(_13815_),
    .B1(net5582));
 sg13g2_a22oi_1 _40326_ (.Y(_13816_),
    .B1(_13814_),
    .B2(_13815_),
    .A2(net4252),
    .A1(net2888));
 sg13g2_inv_1 _40327_ (.Y(_01562_),
    .A(net2889));
 sg13g2_a22oi_1 _40328_ (.Y(_13817_),
    .B1(_13803_),
    .B2(\u_inv.delta_reg[5] ),
    .A2(_15962_),
    .A1(_15959_));
 sg13g2_xnor2_1 _40329_ (.Y(_13818_),
    .A(net2990),
    .B(_13817_));
 sg13g2_nor2b_1 _40330_ (.A(_13814_),
    .B_N(_13818_),
    .Y(_13819_));
 sg13g2_nor2b_1 _40331_ (.A(_13818_),
    .B_N(_13814_),
    .Y(_13820_));
 sg13g2_nor3_1 _40332_ (.A(net5584),
    .B(_13819_),
    .C(_13820_),
    .Y(_13821_));
 sg13g2_a21o_1 _40333_ (.A2(net4252),
    .A1(net2990),
    .B1(_13821_),
    .X(_01563_));
 sg13g2_nand2_1 _40334_ (.Y(_13822_),
    .A(net1247),
    .B(net4252));
 sg13g2_nand3_1 _40335_ (.B(\u_inv.delta_reg[6] ),
    .C(_13803_),
    .A(\u_inv.delta_reg[5] ),
    .Y(_13823_));
 sg13g2_a21oi_1 _40336_ (.A1(net5095),
    .A2(_13823_),
    .Y(_13824_),
    .B1(_15963_));
 sg13g2_xor2_1 _40337_ (.B(_13824_),
    .A(net1247),
    .X(_13825_));
 sg13g2_nor2_1 _40338_ (.A(_13819_),
    .B(_13825_),
    .Y(_13826_));
 sg13g2_nand4_1 _40339_ (.B(_13813_),
    .C(_13818_),
    .A(_13799_),
    .Y(_13827_),
    .D(_13825_));
 sg13g2_o21ai_1 _40340_ (.B1(net5613),
    .Y(_13828_),
    .A1(net4372),
    .A2(_13827_));
 sg13g2_o21ai_1 _40341_ (.B1(_13822_),
    .Y(_01564_),
    .A1(_13826_),
    .A2(_13828_));
 sg13g2_nand2_1 _40342_ (.Y(_13829_),
    .A(net1864),
    .B(net4245));
 sg13g2_nand2b_1 _40343_ (.Y(_13830_),
    .B(\u_inv.delta_reg[8] ),
    .A_N(_15964_));
 sg13g2_nand4_1 _40344_ (.B(\u_inv.delta_reg[7] ),
    .C(\u_inv.delta_reg[6] ),
    .A(\u_inv.delta_reg[5] ),
    .Y(_13831_),
    .D(_13803_));
 sg13g2_inv_1 _40345_ (.Y(_13832_),
    .A(_13831_));
 sg13g2_xnor2_1 _40346_ (.Y(_13833_),
    .A(\u_inv.delta_reg[8] ),
    .B(_13831_));
 sg13g2_a22oi_1 _40347_ (.Y(_13834_),
    .B1(_13833_),
    .B2(net5095),
    .A2(_13830_),
    .A1(_15966_));
 sg13g2_o21ai_1 _40348_ (.B1(_13834_),
    .Y(_13835_),
    .A1(net4372),
    .A2(_13827_));
 sg13g2_nand2_1 _40349_ (.Y(_13836_),
    .A(net5613),
    .B(_13835_));
 sg13g2_nor3_1 _40350_ (.A(net4372),
    .B(_13827_),
    .C(_13834_),
    .Y(_13837_));
 sg13g2_o21ai_1 _40351_ (.B1(_13829_),
    .Y(_01565_),
    .A1(_13836_),
    .A2(_13837_));
 sg13g2_nand2_1 _40352_ (.Y(_13838_),
    .A(net1224),
    .B(net4244));
 sg13g2_nand3_1 _40353_ (.B(net1224),
    .C(_13832_),
    .A(\u_inv.delta_reg[8] ),
    .Y(_13839_));
 sg13g2_a21oi_1 _40354_ (.A1(\u_inv.delta_reg[8] ),
    .A2(_13832_),
    .Y(_13840_),
    .B1(net1224));
 sg13g2_nor2_1 _40355_ (.A(net5009),
    .B(_13840_),
    .Y(_13841_));
 sg13g2_a21oi_1 _40356_ (.A1(_13839_),
    .A2(_13841_),
    .Y(_13842_),
    .B1(_15966_));
 sg13g2_xor2_1 _40357_ (.B(_13842_),
    .A(_13837_),
    .X(_13843_));
 sg13g2_o21ai_1 _40358_ (.B1(_13838_),
    .Y(_01566_),
    .A1(net5579),
    .A2(_13843_));
 sg13g2_a22oi_1 _40359_ (.Y(_13844_),
    .B1(_02338_),
    .B2(net5633),
    .A2(net4260),
    .A1(net5829));
 sg13g2_nor2_1 _40360_ (.A(_20877_[0]),
    .B(_13844_),
    .Y(_01567_));
 sg13g2_nor3_2 _40361_ (.A(\u_inv.input_valid ),
    .B(_14511_),
    .C(\u_inv.load_input ),
    .Y(_13845_));
 sg13g2_mux2_1 _40362_ (.A0(net1546),
    .A1(net1397),
    .S(net5297),
    .X(_01568_));
 sg13g2_mux2_1 _40363_ (.A0(net2035),
    .A1(\shift_reg[1] ),
    .S(net5297),
    .X(_01569_));
 sg13g2_mux2_1 _40364_ (.A0(net2285),
    .A1(net1312),
    .S(net5298),
    .X(_01570_));
 sg13g2_mux2_1 _40365_ (.A0(net2204),
    .A1(net1287),
    .S(net5298),
    .X(_01571_));
 sg13g2_mux2_1 _40366_ (.A0(net2510),
    .A1(net1326),
    .S(net5298),
    .X(_01572_));
 sg13g2_mux2_1 _40367_ (.A0(net2139),
    .A1(net1629),
    .S(net5297),
    .X(_01573_));
 sg13g2_mux2_1 _40368_ (.A0(net1697),
    .A1(\shift_reg[6] ),
    .S(net5297),
    .X(_01574_));
 sg13g2_mux2_1 _40369_ (.A0(net2522),
    .A1(net1644),
    .S(net5297),
    .X(_01575_));
 sg13g2_mux2_1 _40370_ (.A0(net1438),
    .A1(\shift_reg[8] ),
    .S(net5297),
    .X(_01576_));
 sg13g2_mux2_1 _40371_ (.A0(net1840),
    .A1(\shift_reg[9] ),
    .S(net5297),
    .X(_01577_));
 sg13g2_nor2_1 _40372_ (.A(net1214),
    .B(net5297),
    .Y(_13846_));
 sg13g2_a21oi_1 _40373_ (.A1(_14512_),
    .A2(net5298),
    .Y(_01578_),
    .B1(_13846_));
 sg13g2_nor2_1 _40374_ (.A(net1148),
    .B(net5299),
    .Y(_13847_));
 sg13g2_a21oi_1 _40375_ (.A1(_14513_),
    .A2(net5299),
    .Y(_01579_),
    .B1(_13847_));
 sg13g2_nor2_1 _40376_ (.A(net1158),
    .B(net5300),
    .Y(_13848_));
 sg13g2_a21oi_1 _40377_ (.A1(_14515_),
    .A2(net5300),
    .Y(_01580_),
    .B1(_13848_));
 sg13g2_nor2_1 _40378_ (.A(net1161),
    .B(net5300),
    .Y(_13849_));
 sg13g2_a21oi_1 _40379_ (.A1(_14516_),
    .A2(net5300),
    .Y(_01581_),
    .B1(_13849_));
 sg13g2_nor2_1 _40380_ (.A(net1295),
    .B(net5302),
    .Y(_13850_));
 sg13g2_a21oi_1 _40381_ (.A1(_14517_),
    .A2(net5301),
    .Y(_01582_),
    .B1(_13850_));
 sg13g2_nor2_1 _40382_ (.A(net1291),
    .B(net5302),
    .Y(_13851_));
 sg13g2_a21oi_1 _40383_ (.A1(_14518_),
    .A2(net5302),
    .Y(_01583_),
    .B1(_13851_));
 sg13g2_mux2_1 _40384_ (.A0(net2727),
    .A1(net2460),
    .S(net5302),
    .X(_01584_));
 sg13g2_mux2_1 _40385_ (.A0(net2209),
    .A1(\shift_reg[17] ),
    .S(net5303),
    .X(_01585_));
 sg13g2_mux2_1 _40386_ (.A0(net2488),
    .A1(net2211),
    .S(net5303),
    .X(_01586_));
 sg13g2_mux2_1 _40387_ (.A0(net2345),
    .A1(net1910),
    .S(net5302),
    .X(_01587_));
 sg13g2_mux2_1 _40388_ (.A0(net2447),
    .A1(net1962),
    .S(net5302),
    .X(_01588_));
 sg13g2_mux2_1 _40389_ (.A0(net2071),
    .A1(\shift_reg[21] ),
    .S(net5303),
    .X(_01589_));
 sg13g2_mux2_1 _40390_ (.A0(net2154),
    .A1(net2028),
    .S(net5303),
    .X(_01590_));
 sg13g2_mux2_1 _40391_ (.A0(net2114),
    .A1(net1465),
    .S(net5303),
    .X(_01591_));
 sg13g2_mux2_1 _40392_ (.A0(net1934),
    .A1(net1731),
    .S(net5303),
    .X(_01592_));
 sg13g2_mux2_1 _40393_ (.A0(net1773),
    .A1(\shift_reg[25] ),
    .S(net5303),
    .X(_01593_));
 sg13g2_mux2_1 _40394_ (.A0(net1924),
    .A1(net1500),
    .S(net5303),
    .X(_01594_));
 sg13g2_mux2_1 _40395_ (.A0(net2384),
    .A1(net1900),
    .S(net5305),
    .X(_01595_));
 sg13g2_mux2_1 _40396_ (.A0(net1990),
    .A1(\shift_reg[28] ),
    .S(net5305),
    .X(_01596_));
 sg13g2_mux2_1 _40397_ (.A0(net2119),
    .A1(\shift_reg[29] ),
    .S(net5305),
    .X(_01597_));
 sg13g2_mux2_1 _40398_ (.A0(net1745),
    .A1(\shift_reg[30] ),
    .S(net5307),
    .X(_01598_));
 sg13g2_mux2_1 _40399_ (.A0(net1838),
    .A1(\shift_reg[31] ),
    .S(net5307),
    .X(_01599_));
 sg13g2_mux2_1 _40400_ (.A0(net1792),
    .A1(\shift_reg[32] ),
    .S(net5307),
    .X(_01600_));
 sg13g2_mux2_1 _40401_ (.A0(net2286),
    .A1(net1558),
    .S(net5307),
    .X(_01601_));
 sg13g2_mux2_1 _40402_ (.A0(net1741),
    .A1(net1378),
    .S(net5310),
    .X(_01602_));
 sg13g2_mux2_1 _40403_ (.A0(net1753),
    .A1(\shift_reg[35] ),
    .S(net5310),
    .X(_01603_));
 sg13g2_mux2_1 _40404_ (.A0(net1529),
    .A1(\shift_reg[36] ),
    .S(net5310),
    .X(_01604_));
 sg13g2_mux2_1 _40405_ (.A0(net1755),
    .A1(net1449),
    .S(net5310),
    .X(_01605_));
 sg13g2_mux2_1 _40406_ (.A0(net1677),
    .A1(net1354),
    .S(net5310),
    .X(_01606_));
 sg13g2_mux2_1 _40407_ (.A0(net1928),
    .A1(\shift_reg[39] ),
    .S(net5310),
    .X(_01607_));
 sg13g2_mux2_1 _40408_ (.A0(net1778),
    .A1(\shift_reg[40] ),
    .S(net5310),
    .X(_01608_));
 sg13g2_mux2_1 _40409_ (.A0(net2048),
    .A1(\shift_reg[41] ),
    .S(net5310),
    .X(_01609_));
 sg13g2_mux2_1 _40410_ (.A0(net1742),
    .A1(net1722),
    .S(net5314),
    .X(_01610_));
 sg13g2_mux2_1 _40411_ (.A0(net1690),
    .A1(\shift_reg[43] ),
    .S(net5314),
    .X(_01611_));
 sg13g2_mux2_1 _40412_ (.A0(net1739),
    .A1(\shift_reg[44] ),
    .S(net5314),
    .X(_01612_));
 sg13g2_mux2_1 _40413_ (.A0(net1797),
    .A1(\shift_reg[45] ),
    .S(net5314),
    .X(_01613_));
 sg13g2_mux2_1 _40414_ (.A0(net1813),
    .A1(net1721),
    .S(net5317),
    .X(_01614_));
 sg13g2_mux2_1 _40415_ (.A0(net1672),
    .A1(\shift_reg[47] ),
    .S(net5317),
    .X(_01615_));
 sg13g2_mux2_1 _40416_ (.A0(net1573),
    .A1(\shift_reg[48] ),
    .S(net5317),
    .X(_01616_));
 sg13g2_mux2_1 _40417_ (.A0(net2187),
    .A1(net1310),
    .S(net5317),
    .X(_01617_));
 sg13g2_mux2_1 _40418_ (.A0(net1807),
    .A1(net1516),
    .S(net5317),
    .X(_01618_));
 sg13g2_mux2_1 _40419_ (.A0(net1750),
    .A1(net1416),
    .S(net5319),
    .X(_01619_));
 sg13g2_mux2_1 _40420_ (.A0(net1455),
    .A1(\shift_reg[52] ),
    .S(net5319),
    .X(_01620_));
 sg13g2_mux2_1 _40421_ (.A0(net1663),
    .A1(\shift_reg[53] ),
    .S(net5319),
    .X(_01621_));
 sg13g2_mux2_1 _40422_ (.A0(net1508),
    .A1(\shift_reg[54] ),
    .S(net5319),
    .X(_01622_));
 sg13g2_mux2_1 _40423_ (.A0(net1483),
    .A1(\shift_reg[55] ),
    .S(net5319),
    .X(_01623_));
 sg13g2_mux2_1 _40424_ (.A0(net2331),
    .A1(\shift_reg[56] ),
    .S(net5319),
    .X(_01624_));
 sg13g2_mux2_1 _40425_ (.A0(net1699),
    .A1(\shift_reg[57] ),
    .S(net5323),
    .X(_01625_));
 sg13g2_mux2_1 _40426_ (.A0(net1654),
    .A1(\shift_reg[58] ),
    .S(net5323),
    .X(_01626_));
 sg13g2_mux2_1 _40427_ (.A0(net2240),
    .A1(net1533),
    .S(net5323),
    .X(_01627_));
 sg13g2_mux2_1 _40428_ (.A0(net1436),
    .A1(\shift_reg[60] ),
    .S(net5323),
    .X(_01628_));
 sg13g2_mux2_1 _40429_ (.A0(net1538),
    .A1(\shift_reg[61] ),
    .S(net5323),
    .X(_01629_));
 sg13g2_mux2_1 _40430_ (.A0(net1488),
    .A1(\shift_reg[62] ),
    .S(net5324),
    .X(_01630_));
 sg13g2_mux2_1 _40431_ (.A0(net1457),
    .A1(\shift_reg[63] ),
    .S(net5323),
    .X(_01631_));
 sg13g2_mux2_1 _40432_ (.A0(net1667),
    .A1(net1479),
    .S(net5324),
    .X(_01632_));
 sg13g2_mux2_1 _40433_ (.A0(net1542),
    .A1(net1463),
    .S(net5326),
    .X(_01633_));
 sg13g2_mux2_1 _40434_ (.A0(net1769),
    .A1(\shift_reg[66] ),
    .S(net5326),
    .X(_01634_));
 sg13g2_mux2_1 _40435_ (.A0(net1802),
    .A1(net1329),
    .S(net5326),
    .X(_01635_));
 sg13g2_mux2_1 _40436_ (.A0(net2435),
    .A1(net2073),
    .S(net5324),
    .X(_01636_));
 sg13g2_mux2_1 _40437_ (.A0(net1547),
    .A1(\shift_reg[69] ),
    .S(net5324),
    .X(_01637_));
 sg13g2_mux2_1 _40438_ (.A0(net1958),
    .A1(net1510),
    .S(net5326),
    .X(_01638_));
 sg13g2_mux2_1 _40439_ (.A0(net1514),
    .A1(\shift_reg[71] ),
    .S(net5326),
    .X(_01639_));
 sg13g2_mux2_1 _40440_ (.A0(net1626),
    .A1(\shift_reg[72] ),
    .S(net5326),
    .X(_01640_));
 sg13g2_mux2_1 _40441_ (.A0(net2079),
    .A1(\shift_reg[73] ),
    .S(net5330),
    .X(_01641_));
 sg13g2_mux2_1 _40442_ (.A0(net1650),
    .A1(\shift_reg[74] ),
    .S(net5330),
    .X(_01642_));
 sg13g2_mux2_1 _40443_ (.A0(net1591),
    .A1(\shift_reg[75] ),
    .S(net5330),
    .X(_01643_));
 sg13g2_mux2_1 _40444_ (.A0(net1569),
    .A1(\shift_reg[76] ),
    .S(net5330),
    .X(_01644_));
 sg13g2_mux2_1 _40445_ (.A0(net1562),
    .A1(\shift_reg[77] ),
    .S(net5330),
    .X(_01645_));
 sg13g2_mux2_1 _40446_ (.A0(net1888),
    .A1(\shift_reg[78] ),
    .S(net5333),
    .X(_01646_));
 sg13g2_mux2_1 _40447_ (.A0(net1461),
    .A1(\shift_reg[79] ),
    .S(net5332),
    .X(_01647_));
 sg13g2_mux2_1 _40448_ (.A0(net1589),
    .A1(\shift_reg[80] ),
    .S(net5333),
    .X(_01648_));
 sg13g2_mux2_1 _40449_ (.A0(net1578),
    .A1(\shift_reg[81] ),
    .S(net5333),
    .X(_01649_));
 sg13g2_mux2_1 _40450_ (.A0(net1856),
    .A1(\shift_reg[82] ),
    .S(net5335),
    .X(_01650_));
 sg13g2_mux2_1 _40451_ (.A0(net1522),
    .A1(\shift_reg[83] ),
    .S(net5335),
    .X(_01651_));
 sg13g2_mux2_1 _40452_ (.A0(net2182),
    .A1(net1376),
    .S(net5337),
    .X(_01652_));
 sg13g2_mux2_1 _40453_ (.A0(net1907),
    .A1(\shift_reg[85] ),
    .S(net5337),
    .X(_01653_));
 sg13g2_mux2_1 _40454_ (.A0(net1782),
    .A1(net1492),
    .S(net5335),
    .X(_01654_));
 sg13g2_mux2_1 _40455_ (.A0(net1575),
    .A1(net1395),
    .S(net5336),
    .X(_01655_));
 sg13g2_mux2_1 _40456_ (.A0(net1822),
    .A1(\shift_reg[88] ),
    .S(net5340),
    .X(_01656_));
 sg13g2_mux2_1 _40457_ (.A0(net2077),
    .A1(\shift_reg[89] ),
    .S(net5340),
    .X(_01657_));
 sg13g2_mux2_1 _40458_ (.A0(net1702),
    .A1(\shift_reg[90] ),
    .S(net5340),
    .X(_01658_));
 sg13g2_mux2_1 _40459_ (.A0(net1599),
    .A1(\shift_reg[91] ),
    .S(net5340),
    .X(_01659_));
 sg13g2_mux2_1 _40460_ (.A0(net1576),
    .A1(\shift_reg[92] ),
    .S(net5340),
    .X(_01660_));
 sg13g2_mux2_1 _40461_ (.A0(net2314),
    .A1(\shift_reg[93] ),
    .S(net5340),
    .X(_01661_));
 sg13g2_mux2_1 _40462_ (.A0(net1707),
    .A1(\shift_reg[94] ),
    .S(net5339),
    .X(_01662_));
 sg13g2_mux2_1 _40463_ (.A0(net1494),
    .A1(\shift_reg[95] ),
    .S(net5339),
    .X(_01663_));
 sg13g2_mux2_1 _40464_ (.A0(net1756),
    .A1(\shift_reg[96] ),
    .S(net5339),
    .X(_01664_));
 sg13g2_mux2_1 _40465_ (.A0(net1728),
    .A1(\shift_reg[97] ),
    .S(net5340),
    .X(_01665_));
 sg13g2_mux2_1 _40466_ (.A0(net2436),
    .A1(net1994),
    .S(net5340),
    .X(_01666_));
 sg13g2_mux2_1 _40467_ (.A0(net1512),
    .A1(\shift_reg[99] ),
    .S(net5339),
    .X(_01667_));
 sg13g2_mux2_1 _40468_ (.A0(net2387),
    .A1(net2259),
    .S(net5339),
    .X(_01668_));
 sg13g2_mux2_1 _40469_ (.A0(net1879),
    .A1(\shift_reg[101] ),
    .S(net5338),
    .X(_01669_));
 sg13g2_mux2_1 _40470_ (.A0(net1984),
    .A1(net1374),
    .S(net5338),
    .X(_01670_));
 sg13g2_mux2_1 _40471_ (.A0(net1485),
    .A1(\shift_reg[103] ),
    .S(net5338),
    .X(_01671_));
 sg13g2_mux2_1 _40472_ (.A0(net1930),
    .A1(\shift_reg[104] ),
    .S(net5338),
    .X(_01672_));
 sg13g2_mux2_1 _40473_ (.A0(net2015),
    .A1(\shift_reg[105] ),
    .S(net5338),
    .X(_01673_));
 sg13g2_mux2_1 _40474_ (.A0(net1633),
    .A1(\shift_reg[106] ),
    .S(net5338),
    .X(_01674_));
 sg13g2_mux2_1 _40475_ (.A0(net1447),
    .A1(\shift_reg[107] ),
    .S(net5338),
    .X(_01675_));
 sg13g2_mux2_1 _40476_ (.A0(net1805),
    .A1(\shift_reg[108] ),
    .S(net5338),
    .X(_01676_));
 sg13g2_mux2_1 _40477_ (.A0(net1717),
    .A1(\shift_reg[109] ),
    .S(net5337),
    .X(_01677_));
 sg13g2_mux2_1 _40478_ (.A0(net1917),
    .A1(\shift_reg[110] ),
    .S(net5337),
    .X(_01678_));
 sg13g2_mux2_1 _40479_ (.A0(net1549),
    .A1(\shift_reg[111] ),
    .S(net5336),
    .X(_01679_));
 sg13g2_mux2_1 _40480_ (.A0(net1913),
    .A1(\shift_reg[112] ),
    .S(net5337),
    .X(_01680_));
 sg13g2_mux2_1 _40481_ (.A0(net1892),
    .A1(\shift_reg[113] ),
    .S(net5336),
    .X(_01681_));
 sg13g2_mux2_1 _40482_ (.A0(net1531),
    .A1(\shift_reg[114] ),
    .S(net5336),
    .X(_01682_));
 sg13g2_mux2_1 _40483_ (.A0(net1527),
    .A1(\shift_reg[115] ),
    .S(net5336),
    .X(_01683_));
 sg13g2_mux2_1 _40484_ (.A0(net1632),
    .A1(net1584),
    .S(net5336),
    .X(_01684_));
 sg13g2_mux2_1 _40485_ (.A0(net2157),
    .A1(\shift_reg[117] ),
    .S(net5336),
    .X(_01685_));
 sg13g2_mux2_1 _40486_ (.A0(net2283),
    .A1(net1784),
    .S(net5336),
    .X(_01686_));
 sg13g2_mux2_1 _40487_ (.A0(net1646),
    .A1(\shift_reg[119] ),
    .S(net5334),
    .X(_01687_));
 sg13g2_mux2_1 _40488_ (.A0(net1855),
    .A1(net1800),
    .S(net5334),
    .X(_01688_));
 sg13g2_mux2_1 _40489_ (.A0(net1681),
    .A1(\shift_reg[121] ),
    .S(net5334),
    .X(_01689_));
 sg13g2_mux2_1 _40490_ (.A0(net1974),
    .A1(\shift_reg[122] ),
    .S(net5335),
    .X(_01690_));
 sg13g2_mux2_1 _40491_ (.A0(net1912),
    .A1(net1477),
    .S(net5334),
    .X(_01691_));
 sg13g2_mux2_1 _40492_ (.A0(net2085),
    .A1(net1471),
    .S(net5334),
    .X(_01692_));
 sg13g2_mux2_1 _40493_ (.A0(net2064),
    .A1(net1413),
    .S(net5334),
    .X(_01693_));
 sg13g2_mux2_1 _40494_ (.A0(net2191),
    .A1(net1964),
    .S(net5334),
    .X(_01694_));
 sg13g2_mux2_1 _40495_ (.A0(net1884),
    .A1(net1389),
    .S(net5334),
    .X(_01695_));
 sg13g2_mux2_1 _40496_ (.A0(net1686),
    .A1(\shift_reg[128] ),
    .S(net5332),
    .X(_01696_));
 sg13g2_mux2_1 _40497_ (.A0(net1715),
    .A1(\shift_reg[129] ),
    .S(net5332),
    .X(_01697_));
 sg13g2_mux2_1 _40498_ (.A0(net1622),
    .A1(\shift_reg[130] ),
    .S(net5333),
    .X(_01698_));
 sg13g2_mux2_1 _40499_ (.A0(net2067),
    .A1(\shift_reg[131] ),
    .S(net5333),
    .X(_01699_));
 sg13g2_mux2_1 _40500_ (.A0(net1587),
    .A1(\shift_reg[132] ),
    .S(net5333),
    .X(_01700_));
 sg13g2_mux2_1 _40501_ (.A0(net1693),
    .A1(\shift_reg[133] ),
    .S(net5332),
    .X(_01701_));
 sg13g2_mux2_1 _40502_ (.A0(net1475),
    .A1(net1398),
    .S(net5332),
    .X(_01702_));
 sg13g2_mux2_1 _40503_ (.A0(net1665),
    .A1(\shift_reg[135] ),
    .S(net5332),
    .X(_01703_));
 sg13g2_mux2_1 _40504_ (.A0(net2135),
    .A1(net1938),
    .S(net5328),
    .X(_01704_));
 sg13g2_mux2_1 _40505_ (.A0(net1556),
    .A1(\shift_reg[137] ),
    .S(net5332),
    .X(_01705_));
 sg13g2_mux2_1 _40506_ (.A0(net1803),
    .A1(\shift_reg[138] ),
    .S(net5329),
    .X(_01706_));
 sg13g2_mux2_1 _40507_ (.A0(net1506),
    .A1(\shift_reg[139] ),
    .S(net5329),
    .X(_01707_));
 sg13g2_mux2_1 _40508_ (.A0(net2025),
    .A1(\shift_reg[140] ),
    .S(net5332),
    .X(_01708_));
 sg13g2_mux2_1 _40509_ (.A0(net2090),
    .A1(\shift_reg[141] ),
    .S(net5329),
    .X(_01709_));
 sg13g2_mux2_1 _40510_ (.A0(net2263),
    .A1(\shift_reg[142] ),
    .S(net5328),
    .X(_01710_));
 sg13g2_mux2_1 _40511_ (.A0(net1652),
    .A1(\shift_reg[143] ),
    .S(net5328),
    .X(_01711_));
 sg13g2_mux2_1 _40512_ (.A0(net1883),
    .A1(net1361),
    .S(net5329),
    .X(_01712_));
 sg13g2_mux2_1 _40513_ (.A0(net1861),
    .A1(net1670),
    .S(net5328),
    .X(_01713_));
 sg13g2_mux2_1 _40514_ (.A0(net2014),
    .A1(net1566),
    .S(net5328),
    .X(_01714_));
 sg13g2_mux2_1 _40515_ (.A0(net1776),
    .A1(\shift_reg[147] ),
    .S(net5328),
    .X(_01715_));
 sg13g2_mux2_1 _40516_ (.A0(net1759),
    .A1(\shift_reg[148] ),
    .S(net5328),
    .X(_01716_));
 sg13g2_mux2_1 _40517_ (.A0(net2046),
    .A1(net1871),
    .S(net5328),
    .X(_01717_));
 sg13g2_mux2_1 _40518_ (.A0(net1851),
    .A1(\shift_reg[150] ),
    .S(net5326),
    .X(_01718_));
 sg13g2_mux2_1 _40519_ (.A0(net1932),
    .A1(\shift_reg[151] ),
    .S(net5326),
    .X(_01719_));
 sg13g2_mux2_1 _40520_ (.A0(net2376),
    .A1(\shift_reg[152] ),
    .S(net5327),
    .X(_01720_));
 sg13g2_mux2_1 _40521_ (.A0(net1859),
    .A1(\shift_reg[153] ),
    .S(net5327),
    .X(_01721_));
 sg13g2_mux2_1 _40522_ (.A0(net1886),
    .A1(\shift_reg[154] ),
    .S(net5327),
    .X(_01722_));
 sg13g2_mux2_1 _40523_ (.A0(net1459),
    .A1(\shift_reg[155] ),
    .S(net5327),
    .X(_01723_));
 sg13g2_mux2_1 _40524_ (.A0(net1816),
    .A1(\shift_reg[156] ),
    .S(net5324),
    .X(_01724_));
 sg13g2_mux2_1 _40525_ (.A0(net2166),
    .A1(net1445),
    .S(net5324),
    .X(_01725_));
 sg13g2_mux2_1 _40526_ (.A0(net1940),
    .A1(\shift_reg[158] ),
    .S(net5325),
    .X(_01726_));
 sg13g2_mux2_1 _40527_ (.A0(net1689),
    .A1(net1400),
    .S(net5327),
    .X(_01727_));
 sg13g2_mux2_1 _40528_ (.A0(net1595),
    .A1(\shift_reg[160] ),
    .S(net5324),
    .X(_01728_));
 sg13g2_mux2_1 _40529_ (.A0(net1620),
    .A1(\shift_reg[161] ),
    .S(net5324),
    .X(_01729_));
 sg13g2_mux2_1 _40530_ (.A0(net1935),
    .A1(net1408),
    .S(net5325),
    .X(_01730_));
 sg13g2_mux2_1 _40531_ (.A0(net1897),
    .A1(net1307),
    .S(net5325),
    .X(_01731_));
 sg13g2_mux2_1 _40532_ (.A0(net1607),
    .A1(\shift_reg[164] ),
    .S(net5322),
    .X(_01732_));
 sg13g2_mux2_1 _40533_ (.A0(net2156),
    .A1(net1998),
    .S(net5321),
    .X(_01733_));
 sg13g2_mux2_1 _40534_ (.A0(net1749),
    .A1(net1391),
    .S(net5322),
    .X(_01734_));
 sg13g2_mux2_1 _40535_ (.A0(net1704),
    .A1(\shift_reg[167] ),
    .S(net5322),
    .X(_01735_));
 sg13g2_mux2_1 _40536_ (.A0(net1723),
    .A1(\shift_reg[168] ),
    .S(net5322),
    .X(_01736_));
 sg13g2_mux2_1 _40537_ (.A0(net2109),
    .A1(net2081),
    .S(net5322),
    .X(_01737_));
 sg13g2_mux2_1 _40538_ (.A0(net1735),
    .A1(\shift_reg[170] ),
    .S(net5321),
    .X(_01738_));
 sg13g2_mux2_1 _40539_ (.A0(net2088),
    .A1(net2012),
    .S(net5322),
    .X(_01739_));
 sg13g2_mux2_1 _40540_ (.A0(net2208),
    .A1(net1902),
    .S(net5321),
    .X(_01740_));
 sg13g2_mux2_1 _40541_ (.A0(net2086),
    .A1(\shift_reg[173] ),
    .S(net5321),
    .X(_01741_));
 sg13g2_mux2_1 _40542_ (.A0(net1440),
    .A1(\shift_reg[174] ),
    .S(net5321),
    .X(_01742_));
 sg13g2_mux2_1 _40543_ (.A0(net1695),
    .A1(\shift_reg[175] ),
    .S(net5321),
    .X(_01743_));
 sg13g2_mux2_1 _40544_ (.A0(net1894),
    .A1(net1762),
    .S(net5318),
    .X(_01744_));
 sg13g2_mux2_1 _40545_ (.A0(net1571),
    .A1(\shift_reg[177] ),
    .S(net5319),
    .X(_01745_));
 sg13g2_mux2_1 _40546_ (.A0(net1858),
    .A1(net1370),
    .S(net5321),
    .X(_01746_));
 sg13g2_mux2_1 _40547_ (.A0(net2098),
    .A1(net2008),
    .S(net5321),
    .X(_01747_));
 sg13g2_mux2_1 _40548_ (.A0(net1680),
    .A1(net1614),
    .S(net5318),
    .X(_01748_));
 sg13g2_mux2_1 _40549_ (.A0(net1536),
    .A1(\shift_reg[181] ),
    .S(net5318),
    .X(_01749_));
 sg13g2_mux2_1 _40550_ (.A0(net1895),
    .A1(\shift_reg[182] ),
    .S(net5320),
    .X(_01750_));
 sg13g2_mux2_1 _40551_ (.A0(net1688),
    .A1(net1601),
    .S(net5318),
    .X(_01751_));
 sg13g2_mux2_1 _40552_ (.A0(net1714),
    .A1(net1393),
    .S(net5318),
    .X(_01752_));
 sg13g2_mux2_1 _40553_ (.A0(net1826),
    .A1(\shift_reg[185] ),
    .S(net5318),
    .X(_01753_));
 sg13g2_mux2_1 _40554_ (.A0(net1943),
    .A1(net1796),
    .S(net5318),
    .X(_01754_));
 sg13g2_mux2_1 _40555_ (.A0(net1875),
    .A1(\shift_reg[187] ),
    .S(net5318),
    .X(_01755_));
 sg13g2_mux2_1 _40556_ (.A0(net1970),
    .A1(\shift_reg[188] ),
    .S(net5316),
    .X(_01756_));
 sg13g2_mux2_1 _40557_ (.A0(net1780),
    .A1(\shift_reg[189] ),
    .S(net5316),
    .X(_01757_));
 sg13g2_mux2_1 _40558_ (.A0(net1944),
    .A1(\shift_reg[190] ),
    .S(net5316),
    .X(_01758_));
 sg13g2_mux2_1 _40559_ (.A0(net1683),
    .A1(\shift_reg[191] ),
    .S(net5315),
    .X(_01759_));
 sg13g2_mux2_1 _40560_ (.A0(net1481),
    .A1(\shift_reg[192] ),
    .S(net5316),
    .X(_01760_));
 sg13g2_mux2_1 _40561_ (.A0(net1564),
    .A1(\shift_reg[193] ),
    .S(net5315),
    .X(_01761_));
 sg13g2_mux2_1 _40562_ (.A0(net1758),
    .A1(net1658),
    .S(net5315),
    .X(_01762_));
 sg13g2_mux2_1 _40563_ (.A0(net2006),
    .A1(\shift_reg[195] ),
    .S(net5315),
    .X(_01763_));
 sg13g2_mux2_1 _40564_ (.A0(net1960),
    .A1(\shift_reg[196] ),
    .S(net5315),
    .X(_01764_));
 sg13g2_mux2_1 _40565_ (.A0(net1978),
    .A1(\shift_reg[197] ),
    .S(net5315),
    .X(_01765_));
 sg13g2_mux2_1 _40566_ (.A0(net1789),
    .A1(net1453),
    .S(net5315),
    .X(_01766_));
 sg13g2_mux2_1 _40567_ (.A0(net1764),
    .A1(\shift_reg[199] ),
    .S(net5315),
    .X(_01767_));
 sg13g2_mux2_1 _40568_ (.A0(net1992),
    .A1(\shift_reg[200] ),
    .S(net5313),
    .X(_01768_));
 sg13g2_mux2_1 _40569_ (.A0(net2065),
    .A1(net1835),
    .S(net5313),
    .X(_01769_));
 sg13g2_mux2_1 _40570_ (.A0(net1771),
    .A1(net1692),
    .S(net5312),
    .X(_01770_));
 sg13g2_mux2_1 _40571_ (.A0(net2001),
    .A1(net1719),
    .S(net5313),
    .X(_01771_));
 sg13g2_mux2_1 _40572_ (.A0(net1675),
    .A1(\shift_reg[204] ),
    .S(net5313),
    .X(_01772_));
 sg13g2_mux2_1 _40573_ (.A0(net1927),
    .A1(net1921),
    .S(net5313),
    .X(_01773_));
 sg13g2_mux2_1 _40574_ (.A0(net1873),
    .A1(\shift_reg[206] ),
    .S(net5312),
    .X(_01774_));
 sg13g2_mux2_1 _40575_ (.A0(net2133),
    .A1(\shift_reg[207] ),
    .S(net5312),
    .X(_01775_));
 sg13g2_mux2_1 _40576_ (.A0(net1603),
    .A1(\shift_reg[208] ),
    .S(net5312),
    .X(_01776_));
 sg13g2_mux2_1 _40577_ (.A0(net1747),
    .A1(\shift_reg[209] ),
    .S(net5312),
    .X(_01777_));
 sg13g2_mux2_1 _40578_ (.A0(net1885),
    .A1(net1543),
    .S(net5312),
    .X(_01778_));
 sg13g2_mux2_1 _40579_ (.A0(net1783),
    .A1(net1518),
    .S(net5312),
    .X(_01779_));
 sg13g2_mux2_1 _40580_ (.A0(net2183),
    .A1(net1845),
    .S(net5312),
    .X(_01780_));
 sg13g2_mux2_1 _40581_ (.A0(net2152),
    .A1(net1942),
    .S(net5309),
    .X(_01781_));
 sg13g2_mux2_1 _40582_ (.A0(net1986),
    .A1(\shift_reg[214] ),
    .S(net5309),
    .X(_01782_));
 sg13g2_mux2_1 _40583_ (.A0(net1844),
    .A1(net1425),
    .S(net5311),
    .X(_01783_));
 sg13g2_mux2_1 _40584_ (.A0(net1618),
    .A1(\shift_reg[216] ),
    .S(net5311),
    .X(_01784_));
 sg13g2_mux2_1 _40585_ (.A0(net1560),
    .A1(\shift_reg[217] ),
    .S(net5311),
    .X(_01785_));
 sg13g2_mux2_1 _40586_ (.A0(net1520),
    .A1(\shift_reg[218] ),
    .S(net5309),
    .X(_01786_));
 sg13g2_mux2_1 _40587_ (.A0(net1540),
    .A1(\shift_reg[219] ),
    .S(net5309),
    .X(_01787_));
 sg13g2_mux2_1 _40588_ (.A0(net1824),
    .A1(\shift_reg[220] ),
    .S(net5309),
    .X(_01788_));
 sg13g2_mux2_1 _40589_ (.A0(net1662),
    .A1(net1451),
    .S(net5309),
    .X(_01789_));
 sg13g2_mux2_1 _40590_ (.A0(net1639),
    .A1(net1434),
    .S(net5309),
    .X(_01790_));
 sg13g2_mux2_1 _40591_ (.A0(net1909),
    .A1(net1788),
    .S(net5309),
    .X(_01791_));
 sg13g2_mux2_1 _40592_ (.A0(net1467),
    .A1(\shift_reg[224] ),
    .S(net5306),
    .X(_01792_));
 sg13g2_mux2_1 _40593_ (.A0(net1985),
    .A1(net1973),
    .S(net5307),
    .X(_01793_));
 sg13g2_mux2_1 _40594_ (.A0(net1685),
    .A1(net1431),
    .S(net5307),
    .X(_01794_));
 sg13g2_mux2_1 _40595_ (.A0(net1905),
    .A1(\shift_reg[227] ),
    .S(net5307),
    .X(_01795_));
 sg13g2_mux2_1 _40596_ (.A0(net1469),
    .A1(\shift_reg[228] ),
    .S(net5306),
    .X(_01796_));
 sg13g2_mux2_1 _40597_ (.A0(net1586),
    .A1(net1429),
    .S(net5306),
    .X(_01797_));
 sg13g2_mux2_1 _40598_ (.A0(net2059),
    .A1(net2047),
    .S(net5306),
    .X(_01798_));
 sg13g2_mux2_1 _40599_ (.A0(net1551),
    .A1(\shift_reg[231] ),
    .S(net5306),
    .X(_01799_));
 sg13g2_mux2_1 _40600_ (.A0(net1919),
    .A1(\shift_reg[232] ),
    .S(net5306),
    .X(_01800_));
 sg13g2_mux2_1 _40601_ (.A0(net1814),
    .A1(\shift_reg[233] ),
    .S(net5306),
    .X(_01801_));
 sg13g2_mux2_1 _40602_ (.A0(net1593),
    .A1(\shift_reg[234] ),
    .S(net5304),
    .X(_01802_));
 sg13g2_mux2_1 _40603_ (.A0(net2179),
    .A1(\shift_reg[235] ),
    .S(net5304),
    .X(_01803_));
 sg13g2_mux2_1 _40604_ (.A0(net1637),
    .A1(\shift_reg[236] ),
    .S(net5306),
    .X(_01804_));
 sg13g2_mux2_1 _40605_ (.A0(net2089),
    .A1(net1487),
    .S(net5304),
    .X(_01805_));
 sg13g2_mux2_1 _40606_ (.A0(net2192),
    .A1(net1980),
    .S(net5305),
    .X(_01806_));
 sg13g2_mux2_1 _40607_ (.A0(net1706),
    .A1(net1427),
    .S(net5305),
    .X(_01807_));
 sg13g2_mux2_1 _40608_ (.A0(net1473),
    .A1(\shift_reg[240] ),
    .S(net5305),
    .X(_01808_));
 sg13g2_mux2_1 _40609_ (.A0(net1498),
    .A1(\shift_reg[241] ),
    .S(net5304),
    .X(_01809_));
 sg13g2_mux2_1 _40610_ (.A0(net1568),
    .A1(net1502),
    .S(net5304),
    .X(_01810_));
 sg13g2_mux2_1 _40611_ (.A0(net1553),
    .A1(net1345),
    .S(net5304),
    .X(_01811_));
 sg13g2_mux2_1 _40612_ (.A0(net1580),
    .A1(net1404),
    .S(net5304),
    .X(_01812_));
 sg13g2_mux2_1 _40613_ (.A0(net1833),
    .A1(\shift_reg[245] ),
    .S(net5304),
    .X(_01813_));
 sg13g2_mux2_1 _40614_ (.A0(net1794),
    .A1(\shift_reg[246] ),
    .S(net5301),
    .X(_01814_));
 sg13g2_mux2_1 _40615_ (.A0(net2215),
    .A1(net1611),
    .S(net5301),
    .X(_01815_));
 sg13g2_mux2_1 _40616_ (.A0(net1642),
    .A1(\shift_reg[248] ),
    .S(net5301),
    .X(_01816_));
 sg13g2_mux2_1 _40617_ (.A0(net2780),
    .A1(net1976),
    .S(net5300),
    .X(_01817_));
 sg13g2_mux2_1 _40618_ (.A0(net1648),
    .A1(\shift_reg[250] ),
    .S(net5301),
    .X(_01818_));
 sg13g2_mux2_1 _40619_ (.A0(net1490),
    .A1(\shift_reg[251] ),
    .S(net5300),
    .X(_01819_));
 sg13g2_mux2_1 _40620_ (.A0(net1635),
    .A1(\shift_reg[252] ),
    .S(net5301),
    .X(_01820_));
 sg13g2_mux2_1 _40621_ (.A0(net2288),
    .A1(\shift_reg[253] ),
    .S(net5300),
    .X(_01821_));
 sg13g2_mux2_1 _40622_ (.A0(net1842),
    .A1(net1402),
    .S(net5300),
    .X(_01822_));
 sg13g2_mux2_1 _40623_ (.A0(net1605),
    .A1(\shift_reg[255] ),
    .S(net5301),
    .X(_01823_));
 sg13g2_nand2_1 _40624_ (.Y(_13852_),
    .A(_14815_),
    .B(_14819_));
 sg13g2_a21o_1 _40625_ (.A2(_13852_),
    .A1(net1965),
    .B1(_14820_),
    .X(_01824_));
 sg13g2_nand2_1 _40626_ (.Y(_13853_),
    .A(_18354_),
    .B(net4353));
 sg13g2_a21oi_1 _40627_ (.A1(_18354_),
    .A2(_18360_),
    .Y(_13854_),
    .B1(net5625));
 sg13g2_a221oi_1 _40628_ (.B2(_13854_),
    .C1(net4128),
    .B1(_13853_),
    .A1(net1546),
    .Y(_13855_),
    .A2(net5625));
 sg13g2_a21oi_1 _40629_ (.A1(net5667),
    .A2(net4128),
    .Y(_01825_),
    .B1(_13855_));
 sg13g2_nand2b_1 _40630_ (.Y(_13856_),
    .B(net4304),
    .A_N(_18360_));
 sg13g2_a221oi_1 _40631_ (.B2(net4263),
    .C1(net4128),
    .B1(_18367_),
    .A1(net2035),
    .Y(_13857_),
    .A2(net5625));
 sg13g2_a22oi_1 _40632_ (.Y(_01826_),
    .B1(_13856_),
    .B2(_13857_),
    .A2(net4127),
    .A1(_14170_));
 sg13g2_nand2_1 _40633_ (.Y(_13858_),
    .A(_18367_),
    .B(net4304));
 sg13g2_a221oi_1 _40634_ (.B2(net4263),
    .C1(net4127),
    .B1(_18349_),
    .A1(net2285),
    .Y(_13859_),
    .A2(net5624));
 sg13g2_a22oi_1 _40635_ (.Y(_01827_),
    .B1(_13858_),
    .B2(_13859_),
    .A2(net4127),
    .A1(_14169_));
 sg13g2_nand2_1 _40636_ (.Y(_13860_),
    .A(_18343_),
    .B(net4263));
 sg13g2_a221oi_1 _40637_ (.B2(net4304),
    .C1(net4127),
    .B1(_18349_),
    .A1(net2204),
    .Y(_13861_),
    .A2(net5625));
 sg13g2_a22oi_1 _40638_ (.Y(_01828_),
    .B1(_13860_),
    .B2(_13861_),
    .A2(net4127),
    .A1(_14168_));
 sg13g2_a22oi_1 _40639_ (.Y(_13862_),
    .B1(_18343_),
    .B2(net4304),
    .A2(net5624),
    .A1(net2510));
 sg13g2_o21ai_1 _40640_ (.B1(_13862_),
    .Y(_13863_),
    .A1(_18375_),
    .A2(net4348));
 sg13g2_mux2_1 _40641_ (.A0(_13863_),
    .A1(net2355),
    .S(net4127),
    .X(_01829_));
 sg13g2_nand2b_1 _40642_ (.Y(_13864_),
    .B(net4304),
    .A_N(_18375_));
 sg13g2_a221oi_1 _40643_ (.B2(net4263),
    .C1(net4127),
    .B1(_18336_),
    .A1(net2139),
    .Y(_13865_),
    .A2(net5624));
 sg13g2_a22oi_1 _40644_ (.Y(_01830_),
    .B1(_13864_),
    .B2(_13865_),
    .A2(net4127),
    .A1(_14167_));
 sg13g2_a22oi_1 _40645_ (.Y(_13866_),
    .B1(_18336_),
    .B2(net4304),
    .A2(net5624),
    .A1(net1697));
 sg13g2_o21ai_1 _40646_ (.B1(_13866_),
    .Y(_13867_),
    .A1(_18330_),
    .A2(net4348));
 sg13g2_mux2_1 _40647_ (.A0(_13867_),
    .A1(net3272),
    .S(net4129),
    .X(_01831_));
 sg13g2_a22oi_1 _40648_ (.Y(_13868_),
    .B1(_18382_),
    .B2(net4263),
    .A2(net5624),
    .A1(net2522));
 sg13g2_o21ai_1 _40649_ (.B1(_13868_),
    .Y(_13869_),
    .A1(_18330_),
    .A2(net4260));
 sg13g2_mux2_1 _40650_ (.A0(_13869_),
    .A1(net2608),
    .S(net4129),
    .X(_01832_));
 sg13g2_nand2_1 _40651_ (.Y(_13870_),
    .A(_18324_),
    .B(net4263));
 sg13g2_a221oi_1 _40652_ (.B2(net4305),
    .C1(net4128),
    .B1(_18382_),
    .A1(net1438),
    .Y(_13871_),
    .A2(net5624));
 sg13g2_a22oi_1 _40653_ (.Y(_01833_),
    .B1(_13870_),
    .B2(_13871_),
    .A2(net4129),
    .A1(_14166_));
 sg13g2_nand2_1 _40654_ (.Y(_13872_),
    .A(_18324_),
    .B(net4305));
 sg13g2_a221oi_1 _40655_ (.B2(net4263),
    .C1(net4129),
    .B1(_18317_),
    .A1(net1840),
    .Y(_13873_),
    .A2(net5624));
 sg13g2_a22oi_1 _40656_ (.Y(_01834_),
    .B1(_13872_),
    .B2(_13873_),
    .A2(net4129),
    .A1(_14165_));
 sg13g2_a22oi_1 _40657_ (.Y(_13874_),
    .B1(_18317_),
    .B2(net4304),
    .A2(net5626),
    .A1(net1214));
 sg13g2_o21ai_1 _40658_ (.B1(_13874_),
    .Y(_13875_),
    .A1(_18311_),
    .A2(net4348));
 sg13g2_nor2_1 _40659_ (.A(net4128),
    .B(_13875_),
    .Y(_13876_));
 sg13g2_a21oi_1 _40660_ (.A1(_14164_),
    .A2(net4128),
    .Y(_01835_),
    .B1(_13876_));
 sg13g2_nand2b_1 _40661_ (.Y(_13877_),
    .B(net4304),
    .A_N(_18311_));
 sg13g2_a221oi_1 _40662_ (.B2(net4263),
    .C1(net4133),
    .B1(_18390_),
    .A1(net1148),
    .Y(_13878_),
    .A2(net5627));
 sg13g2_a22oi_1 _40663_ (.Y(_01836_),
    .B1(_13877_),
    .B2(_13878_),
    .A2(net4128),
    .A1(_14163_));
 sg13g2_nand2_1 _40664_ (.Y(_13879_),
    .A(_18390_),
    .B(net4305));
 sg13g2_a221oi_1 _40665_ (.B2(net4262),
    .C1(net4132),
    .B1(_18305_),
    .A1(net1158),
    .Y(_13880_),
    .A2(net5627));
 sg13g2_a22oi_1 _40666_ (.Y(_01837_),
    .B1(_13879_),
    .B2(_13880_),
    .A2(net4133),
    .A1(_14162_));
 sg13g2_nand2_1 _40667_ (.Y(_13881_),
    .A(_18299_),
    .B(net4261));
 sg13g2_a221oi_1 _40668_ (.B2(net4306),
    .C1(net4130),
    .B1(_18305_),
    .A1(net1161),
    .Y(_13882_),
    .A2(net5627));
 sg13g2_a22oi_1 _40669_ (.Y(_01838_),
    .B1(_13881_),
    .B2(_13882_),
    .A2(net4130),
    .A1(_14161_));
 sg13g2_nand2_1 _40670_ (.Y(_13883_),
    .A(_18299_),
    .B(net4306));
 sg13g2_a221oi_1 _40671_ (.B2(net4261),
    .C1(net4130),
    .B1(_18292_),
    .A1(net1295),
    .Y(_13884_),
    .A2(net5629));
 sg13g2_a22oi_1 _40672_ (.Y(_01839_),
    .B1(_13883_),
    .B2(_13884_),
    .A2(net4131),
    .A1(_14160_));
 sg13g2_nand2_1 _40673_ (.Y(_13885_),
    .A(_18292_),
    .B(net4306));
 sg13g2_a221oi_1 _40674_ (.B2(net4261),
    .C1(net4130),
    .B1(_18278_),
    .A1(net1291),
    .Y(_13886_),
    .A2(net5628));
 sg13g2_a22oi_1 _40675_ (.Y(_01840_),
    .B1(_13885_),
    .B2(_13886_),
    .A2(net4131),
    .A1(_14159_));
 sg13g2_nand2_1 _40676_ (.Y(_13887_),
    .A(_18287_),
    .B(net4261));
 sg13g2_a221oi_1 _40677_ (.B2(net4306),
    .C1(net4130),
    .B1(_18278_),
    .A1(net2727),
    .Y(_13888_),
    .A2(net5628));
 sg13g2_a22oi_1 _40678_ (.Y(_01841_),
    .B1(_13887_),
    .B2(_13888_),
    .A2(net4130),
    .A1(_14158_));
 sg13g2_nand2_1 _40679_ (.Y(_13889_),
    .A(_18287_),
    .B(net4306));
 sg13g2_a221oi_1 _40680_ (.B2(net4265),
    .C1(net4140),
    .B1(_18409_),
    .A1(net2209),
    .Y(_13890_),
    .A2(net5629));
 sg13g2_a22oi_1 _40681_ (.Y(_01842_),
    .B1(_13889_),
    .B2(_13890_),
    .A2(net4140),
    .A1(_14157_));
 sg13g2_nand2_1 _40682_ (.Y(_13891_),
    .A(_18270_),
    .B(net4261));
 sg13g2_a221oi_1 _40683_ (.B2(net4309),
    .C1(net4140),
    .B1(_18409_),
    .A1(net2488),
    .Y(_13892_),
    .A2(net5629));
 sg13g2_a22oi_1 _40684_ (.Y(_01843_),
    .B1(_13891_),
    .B2(_13892_),
    .A2(net4140),
    .A1(_14156_));
 sg13g2_a22oi_1 _40685_ (.Y(_13893_),
    .B1(_18270_),
    .B2(net4306),
    .A2(net5629),
    .A1(net2345));
 sg13g2_o21ai_1 _40686_ (.B1(_13893_),
    .Y(_13894_),
    .A1(_18401_),
    .A2(net4348));
 sg13g2_nor2_1 _40687_ (.A(net4131),
    .B(_13894_),
    .Y(_13895_));
 sg13g2_a21oi_1 _40688_ (.A1(_14155_),
    .A2(net4131),
    .Y(_01844_),
    .B1(_13895_));
 sg13g2_nand2b_1 _40689_ (.Y(_13896_),
    .B(net4306),
    .A_N(_18401_));
 sg13g2_a221oi_1 _40690_ (.B2(net4265),
    .C1(net4140),
    .B1(_18264_),
    .A1(net2447),
    .Y(_13897_),
    .A2(net5629));
 sg13g2_a22oi_1 _40691_ (.Y(_01845_),
    .B1(_13896_),
    .B2(_13897_),
    .A2(net4131),
    .A1(_14154_));
 sg13g2_a22oi_1 _40692_ (.Y(_13898_),
    .B1(_18264_),
    .B2(net4309),
    .A2(net5629),
    .A1(net2071));
 sg13g2_o21ai_1 _40693_ (.B1(_13898_),
    .Y(_13899_),
    .A1(_18420_),
    .A2(net4348));
 sg13g2_nor2_1 _40694_ (.A(net4140),
    .B(_13899_),
    .Y(_13900_));
 sg13g2_a21oi_1 _40695_ (.A1(_14153_),
    .A2(net4131),
    .Y(_01846_),
    .B1(_13900_));
 sg13g2_a22oi_1 _40696_ (.Y(_13901_),
    .B1(_18256_),
    .B2(net4265),
    .A2(net5629),
    .A1(net2154));
 sg13g2_o21ai_1 _40697_ (.B1(_13901_),
    .Y(_13902_),
    .A1(_18420_),
    .A2(net4260));
 sg13g2_mux2_1 _40698_ (.A0(_13902_),
    .A1(net3346),
    .S(net4140),
    .X(_01847_));
 sg13g2_nand2_1 _40699_ (.Y(_13903_),
    .A(_18256_),
    .B(net4309));
 sg13g2_a221oi_1 _40700_ (.B2(net4265),
    .C1(net4141),
    .B1(_18251_),
    .A1(net2114),
    .Y(_13904_),
    .A2(net5630));
 sg13g2_a22oi_1 _40701_ (.Y(_01848_),
    .B1(_13903_),
    .B2(_13904_),
    .A2(net4141),
    .A1(_14151_));
 sg13g2_a22oi_1 _40702_ (.Y(_13905_),
    .B1(_18251_),
    .B2(net4309),
    .A2(net5630),
    .A1(net1934));
 sg13g2_o21ai_1 _40703_ (.B1(_13905_),
    .Y(_13906_),
    .A1(_18428_),
    .A2(net4348));
 sg13g2_nor2_1 _40704_ (.A(net4141),
    .B(_13906_),
    .Y(_13907_));
 sg13g2_a21oi_1 _40705_ (.A1(_14150_),
    .A2(net4141),
    .Y(_01849_),
    .B1(_13907_));
 sg13g2_a22oi_1 _40706_ (.Y(_13908_),
    .B1(_18445_),
    .B2(net4265),
    .A2(net5630),
    .A1(net1773));
 sg13g2_o21ai_1 _40707_ (.B1(_13908_),
    .Y(_13909_),
    .A1(_18428_),
    .A2(net4260));
 sg13g2_mux2_1 _40708_ (.A0(_13909_),
    .A1(net2998),
    .S(net4141),
    .X(_01850_));
 sg13g2_nand2_1 _40709_ (.Y(_13910_),
    .A(_18242_),
    .B(net4265));
 sg13g2_a221oi_1 _40710_ (.B2(net4309),
    .C1(net4145),
    .B1(_18445_),
    .A1(net1924),
    .Y(_13911_),
    .A2(net5629));
 sg13g2_a22oi_1 _40711_ (.Y(_01851_),
    .B1(_13910_),
    .B2(_13911_),
    .A2(net4145),
    .A1(_14148_));
 sg13g2_nand2_1 _40712_ (.Y(_13912_),
    .A(_18242_),
    .B(net4312));
 sg13g2_a221oi_1 _40713_ (.B2(net4268),
    .C1(net4145),
    .B1(_18237_),
    .A1(net2384),
    .Y(_13913_),
    .A2(net5630));
 sg13g2_a22oi_1 _40714_ (.Y(_01852_),
    .B1(_13912_),
    .B2(_13913_),
    .A2(net4145),
    .A1(_14147_));
 sg13g2_a22oi_1 _40715_ (.Y(_13914_),
    .B1(_18237_),
    .B2(net4312),
    .A2(net5630),
    .A1(net1990));
 sg13g2_o21ai_1 _40716_ (.B1(_13914_),
    .Y(_13915_),
    .A1(_18468_),
    .A2(net4348));
 sg13g2_nor2_1 _40717_ (.A(net4145),
    .B(_13915_),
    .Y(_13916_));
 sg13g2_a21oi_1 _40718_ (.A1(_14146_),
    .A2(net4145),
    .Y(_01853_),
    .B1(_13916_));
 sg13g2_nand2b_1 _40719_ (.Y(_13917_),
    .B(net4312),
    .A_N(_18468_));
 sg13g2_a221oi_1 _40720_ (.B2(net4268),
    .C1(net4145),
    .B1(_18497_),
    .A1(net2119),
    .Y(_13918_),
    .A2(net5630));
 sg13g2_a22oi_1 _40721_ (.Y(_01854_),
    .B1(_13917_),
    .B2(_13918_),
    .A2(net4145),
    .A1(_14145_));
 sg13g2_dfrbpq_2 _40722_ (.RESET_B(net25),
    .D(_00001_),
    .Q(\u_inv.f_next[30] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _40723_ (.RESET_B(net250),
    .D(_00002_),
    .Q(\u_inv.f_next[31] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _40724_ (.RESET_B(net249),
    .D(_00003_),
    .Q(\u_inv.f_next[32] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _40725_ (.RESET_B(net248),
    .D(_00004_),
    .Q(\u_inv.f_next[33] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _40726_ (.RESET_B(net247),
    .D(_00005_),
    .Q(\u_inv.f_next[34] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _40727_ (.RESET_B(net246),
    .D(_00006_),
    .Q(\u_inv.f_next[35] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _40728_ (.RESET_B(net245),
    .D(_00007_),
    .Q(\u_inv.f_next[36] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _40729_ (.RESET_B(net244),
    .D(_00008_),
    .Q(\u_inv.f_next[37] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _40730_ (.RESET_B(net243),
    .D(_00009_),
    .Q(\u_inv.f_next[38] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _40731_ (.RESET_B(net242),
    .D(_00010_),
    .Q(\u_inv.f_next[39] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _40732_ (.RESET_B(net241),
    .D(_00011_),
    .Q(\u_inv.f_next[40] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _40733_ (.RESET_B(net240),
    .D(_00012_),
    .Q(\u_inv.f_next[41] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _40734_ (.RESET_B(net239),
    .D(_00013_),
    .Q(\u_inv.f_next[42] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _40735_ (.RESET_B(net238),
    .D(_00014_),
    .Q(\u_inv.f_next[43] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _40736_ (.RESET_B(net237),
    .D(_00015_),
    .Q(\u_inv.f_next[44] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _40737_ (.RESET_B(net236),
    .D(_00016_),
    .Q(\u_inv.f_next[45] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _40738_ (.RESET_B(net235),
    .D(_00017_),
    .Q(\u_inv.f_next[46] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _40739_ (.RESET_B(net234),
    .D(_00018_),
    .Q(\u_inv.f_next[47] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _40740_ (.RESET_B(net233),
    .D(_00019_),
    .Q(\u_inv.f_next[48] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _40741_ (.RESET_B(net232),
    .D(_00020_),
    .Q(\u_inv.f_next[49] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _40742_ (.RESET_B(net231),
    .D(_00021_),
    .Q(\u_inv.f_next[50] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _40743_ (.RESET_B(net230),
    .D(_00022_),
    .Q(\u_inv.f_next[51] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _40744_ (.RESET_B(net229),
    .D(_00023_),
    .Q(\u_inv.f_next[52] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _40745_ (.RESET_B(net228),
    .D(_00024_),
    .Q(\u_inv.f_next[53] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _40746_ (.RESET_B(net227),
    .D(_00025_),
    .Q(\u_inv.f_next[54] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _40747_ (.RESET_B(net226),
    .D(_00026_),
    .Q(\u_inv.f_next[55] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _40748_ (.RESET_B(net225),
    .D(_00027_),
    .Q(\u_inv.f_next[56] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _40749_ (.RESET_B(net224),
    .D(_00028_),
    .Q(\u_inv.f_next[57] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _40750_ (.RESET_B(net223),
    .D(_00029_),
    .Q(\u_inv.f_next[58] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _40751_ (.RESET_B(net222),
    .D(_00030_),
    .Q(\u_inv.f_next[59] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _40752_ (.RESET_B(net221),
    .D(_00031_),
    .Q(\u_inv.f_next[60] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _40753_ (.RESET_B(net220),
    .D(_00032_),
    .Q(\u_inv.f_next[61] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _40754_ (.RESET_B(net219),
    .D(_00033_),
    .Q(\u_inv.f_next[62] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _40755_ (.RESET_B(net218),
    .D(_00034_),
    .Q(\u_inv.f_next[63] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _40756_ (.RESET_B(net217),
    .D(_00035_),
    .Q(\u_inv.f_next[64] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _40757_ (.RESET_B(net216),
    .D(_00036_),
    .Q(\u_inv.f_next[65] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_2 _40758_ (.RESET_B(net215),
    .D(_00037_),
    .Q(\u_inv.f_next[66] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _40759_ (.RESET_B(net214),
    .D(_00038_),
    .Q(\u_inv.f_next[67] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _40760_ (.RESET_B(net213),
    .D(_00039_),
    .Q(\u_inv.f_next[68] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _40761_ (.RESET_B(net212),
    .D(_00040_),
    .Q(\u_inv.f_next[69] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _40762_ (.RESET_B(net211),
    .D(_00041_),
    .Q(\u_inv.f_next[70] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _40763_ (.RESET_B(net210),
    .D(_00042_),
    .Q(\u_inv.f_next[71] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _40764_ (.RESET_B(net209),
    .D(_00043_),
    .Q(\u_inv.f_next[72] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _40765_ (.RESET_B(net208),
    .D(_00044_),
    .Q(\u_inv.f_next[73] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _40766_ (.RESET_B(net207),
    .D(_00045_),
    .Q(\u_inv.f_next[74] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _40767_ (.RESET_B(net206),
    .D(_00046_),
    .Q(\u_inv.f_next[75] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _40768_ (.RESET_B(net205),
    .D(_00047_),
    .Q(\u_inv.f_next[76] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _40769_ (.RESET_B(net204),
    .D(_00048_),
    .Q(\u_inv.f_next[77] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _40770_ (.RESET_B(net203),
    .D(_00049_),
    .Q(\u_inv.f_next[78] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_2 _40771_ (.RESET_B(net202),
    .D(_00050_),
    .Q(\u_inv.f_next[79] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _40772_ (.RESET_B(net201),
    .D(_00051_),
    .Q(\u_inv.f_next[80] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _40773_ (.RESET_B(net200),
    .D(_00052_),
    .Q(\u_inv.f_next[81] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _40774_ (.RESET_B(net199),
    .D(_00053_),
    .Q(\u_inv.f_next[82] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _40775_ (.RESET_B(net198),
    .D(_00054_),
    .Q(\u_inv.f_next[83] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _40776_ (.RESET_B(net197),
    .D(_00055_),
    .Q(\u_inv.f_next[84] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _40777_ (.RESET_B(net196),
    .D(_00056_),
    .Q(\u_inv.f_next[85] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _40778_ (.RESET_B(net195),
    .D(_00057_),
    .Q(\u_inv.f_next[86] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _40779_ (.RESET_B(net194),
    .D(_00058_),
    .Q(\u_inv.f_next[87] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _40780_ (.RESET_B(net193),
    .D(_00059_),
    .Q(\u_inv.f_next[88] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_2 _40781_ (.RESET_B(net192),
    .D(_00060_),
    .Q(\u_inv.f_next[89] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _40782_ (.RESET_B(net191),
    .D(_00061_),
    .Q(\u_inv.f_next[90] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_2 _40783_ (.RESET_B(net190),
    .D(_00062_),
    .Q(\u_inv.f_next[91] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _40784_ (.RESET_B(net189),
    .D(_00063_),
    .Q(\u_inv.f_next[92] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _40785_ (.RESET_B(net188),
    .D(_00064_),
    .Q(\u_inv.f_next[93] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _40786_ (.RESET_B(net187),
    .D(_00065_),
    .Q(\u_inv.f_next[94] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _40787_ (.RESET_B(net186),
    .D(_00066_),
    .Q(\u_inv.f_next[95] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _40788_ (.RESET_B(net185),
    .D(_00067_),
    .Q(\u_inv.f_next[96] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _40789_ (.RESET_B(net184),
    .D(_00068_),
    .Q(\u_inv.f_next[97] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _40790_ (.RESET_B(net183),
    .D(_00069_),
    .Q(\u_inv.f_next[98] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _40791_ (.RESET_B(net182),
    .D(_00070_),
    .Q(\u_inv.f_next[99] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _40792_ (.RESET_B(net181),
    .D(_00071_),
    .Q(\u_inv.f_next[100] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _40793_ (.RESET_B(net180),
    .D(_00072_),
    .Q(\u_inv.f_next[101] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _40794_ (.RESET_B(net179),
    .D(_00073_),
    .Q(\u_inv.f_next[102] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _40795_ (.RESET_B(net178),
    .D(_00074_),
    .Q(\u_inv.f_next[103] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _40796_ (.RESET_B(net177),
    .D(_00075_),
    .Q(\u_inv.f_next[104] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _40797_ (.RESET_B(net176),
    .D(_00076_),
    .Q(\u_inv.f_next[105] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _40798_ (.RESET_B(net175),
    .D(_00077_),
    .Q(\u_inv.f_next[106] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _40799_ (.RESET_B(net174),
    .D(_00078_),
    .Q(\u_inv.f_next[107] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _40800_ (.RESET_B(net173),
    .D(_00079_),
    .Q(\u_inv.f_next[108] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _40801_ (.RESET_B(net172),
    .D(_00080_),
    .Q(\u_inv.f_next[109] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _40802_ (.RESET_B(net171),
    .D(_00081_),
    .Q(\u_inv.f_next[110] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _40803_ (.RESET_B(net170),
    .D(_00082_),
    .Q(\u_inv.f_next[111] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _40804_ (.RESET_B(net169),
    .D(_00083_),
    .Q(\u_inv.f_next[112] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _40805_ (.RESET_B(net168),
    .D(_00084_),
    .Q(\u_inv.f_next[113] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _40806_ (.RESET_B(net167),
    .D(_00085_),
    .Q(\u_inv.f_next[114] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _40807_ (.RESET_B(net166),
    .D(_00086_),
    .Q(\u_inv.f_next[115] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _40808_ (.RESET_B(net165),
    .D(_00087_),
    .Q(\u_inv.f_next[116] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _40809_ (.RESET_B(net164),
    .D(_00088_),
    .Q(\u_inv.f_next[117] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _40810_ (.RESET_B(net163),
    .D(_00089_),
    .Q(\u_inv.f_next[118] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _40811_ (.RESET_B(net162),
    .D(_00090_),
    .Q(\u_inv.f_next[119] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _40812_ (.RESET_B(net161),
    .D(_00091_),
    .Q(\u_inv.f_next[120] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _40813_ (.RESET_B(net160),
    .D(_00092_),
    .Q(\u_inv.f_next[121] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _40814_ (.RESET_B(net159),
    .D(_00093_),
    .Q(\u_inv.f_next[122] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _40815_ (.RESET_B(net158),
    .D(_00094_),
    .Q(\u_inv.f_next[123] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _40816_ (.RESET_B(net157),
    .D(_00095_),
    .Q(\u_inv.f_next[124] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _40817_ (.RESET_B(net156),
    .D(_00096_),
    .Q(\u_inv.f_next[125] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _40818_ (.RESET_B(net155),
    .D(_00097_),
    .Q(\u_inv.f_next[126] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _40819_ (.RESET_B(net154),
    .D(_00098_),
    .Q(\u_inv.f_next[127] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _40820_ (.RESET_B(net153),
    .D(_00099_),
    .Q(\u_inv.f_next[128] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _40821_ (.RESET_B(net152),
    .D(_00100_),
    .Q(\u_inv.f_next[129] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _40822_ (.RESET_B(net151),
    .D(_00101_),
    .Q(\u_inv.f_next[130] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _40823_ (.RESET_B(net150),
    .D(_00102_),
    .Q(\u_inv.f_next[131] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _40824_ (.RESET_B(net149),
    .D(_00103_),
    .Q(\u_inv.f_next[132] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _40825_ (.RESET_B(net148),
    .D(_00104_),
    .Q(\u_inv.f_next[133] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_2 _40826_ (.RESET_B(net147),
    .D(_00105_),
    .Q(\u_inv.f_next[134] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _40827_ (.RESET_B(net146),
    .D(_00106_),
    .Q(\u_inv.f_next[135] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _40828_ (.RESET_B(net145),
    .D(_00107_),
    .Q(\u_inv.f_next[136] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _40829_ (.RESET_B(net144),
    .D(_00108_),
    .Q(\u_inv.f_next[137] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _40830_ (.RESET_B(net143),
    .D(_00109_),
    .Q(\u_inv.f_next[138] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _40831_ (.RESET_B(net142),
    .D(_00110_),
    .Q(\u_inv.f_next[139] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _40832_ (.RESET_B(net141),
    .D(_00111_),
    .Q(\u_inv.f_next[140] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _40833_ (.RESET_B(net140),
    .D(_00112_),
    .Q(\u_inv.f_next[141] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _40834_ (.RESET_B(net139),
    .D(_00113_),
    .Q(\u_inv.f_next[142] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _40835_ (.RESET_B(net138),
    .D(_00114_),
    .Q(\u_inv.f_next[143] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _40836_ (.RESET_B(net137),
    .D(_00115_),
    .Q(\u_inv.f_next[144] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _40837_ (.RESET_B(net136),
    .D(_00116_),
    .Q(\u_inv.f_next[145] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _40838_ (.RESET_B(net135),
    .D(_00117_),
    .Q(\u_inv.f_next[146] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _40839_ (.RESET_B(net134),
    .D(_00118_),
    .Q(\u_inv.f_next[147] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _40840_ (.RESET_B(net133),
    .D(_00119_),
    .Q(\u_inv.f_next[148] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _40841_ (.RESET_B(net132),
    .D(_00120_),
    .Q(\u_inv.f_next[149] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _40842_ (.RESET_B(net131),
    .D(_00121_),
    .Q(\u_inv.f_next[150] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _40843_ (.RESET_B(net130),
    .D(_00122_),
    .Q(\u_inv.f_next[151] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _40844_ (.RESET_B(net129),
    .D(_00123_),
    .Q(\u_inv.f_next[152] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _40845_ (.RESET_B(net128),
    .D(_00124_),
    .Q(\u_inv.f_next[153] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _40846_ (.RESET_B(net127),
    .D(_00125_),
    .Q(\u_inv.f_next[154] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _40847_ (.RESET_B(net126),
    .D(_00126_),
    .Q(\u_inv.f_next[155] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _40848_ (.RESET_B(net125),
    .D(_00127_),
    .Q(\u_inv.f_next[156] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _40849_ (.RESET_B(net124),
    .D(_00128_),
    .Q(\u_inv.f_next[157] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _40850_ (.RESET_B(net123),
    .D(_00129_),
    .Q(\u_inv.f_next[158] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _40851_ (.RESET_B(net122),
    .D(_00130_),
    .Q(\u_inv.f_next[159] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _40852_ (.RESET_B(net121),
    .D(_00131_),
    .Q(\u_inv.f_next[160] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _40853_ (.RESET_B(net120),
    .D(_00132_),
    .Q(\u_inv.f_next[161] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _40854_ (.RESET_B(net119),
    .D(_00133_),
    .Q(\u_inv.f_next[162] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _40855_ (.RESET_B(net118),
    .D(_00134_),
    .Q(\u_inv.f_next[163] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _40856_ (.RESET_B(net117),
    .D(_00135_),
    .Q(\u_inv.f_next[164] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _40857_ (.RESET_B(net116),
    .D(_00136_),
    .Q(\u_inv.f_next[165] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _40858_ (.RESET_B(net115),
    .D(_00137_),
    .Q(\u_inv.f_next[166] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _40859_ (.RESET_B(net114),
    .D(_00138_),
    .Q(\u_inv.f_next[167] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _40860_ (.RESET_B(net113),
    .D(_00139_),
    .Q(\u_inv.f_next[168] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _40861_ (.RESET_B(net112),
    .D(_00140_),
    .Q(\u_inv.f_next[169] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _40862_ (.RESET_B(net111),
    .D(_00141_),
    .Q(\u_inv.f_next[170] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _40863_ (.RESET_B(net110),
    .D(_00142_),
    .Q(\u_inv.f_next[171] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _40864_ (.RESET_B(net109),
    .D(_00143_),
    .Q(\u_inv.f_next[172] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _40865_ (.RESET_B(net108),
    .D(_00144_),
    .Q(\u_inv.f_next[173] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _40866_ (.RESET_B(net107),
    .D(_00145_),
    .Q(\u_inv.f_next[174] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _40867_ (.RESET_B(net106),
    .D(_00146_),
    .Q(\u_inv.f_next[175] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _40868_ (.RESET_B(net105),
    .D(_00147_),
    .Q(\u_inv.f_next[176] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _40869_ (.RESET_B(net104),
    .D(_00148_),
    .Q(\u_inv.f_next[177] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _40870_ (.RESET_B(net103),
    .D(_00149_),
    .Q(\u_inv.f_next[178] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _40871_ (.RESET_B(net102),
    .D(_00150_),
    .Q(\u_inv.f_next[179] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _40872_ (.RESET_B(net101),
    .D(_00151_),
    .Q(\u_inv.f_next[180] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _40873_ (.RESET_B(net100),
    .D(_00152_),
    .Q(\u_inv.f_next[181] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _40874_ (.RESET_B(net99),
    .D(_00153_),
    .Q(\u_inv.f_next[182] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _40875_ (.RESET_B(net98),
    .D(_00154_),
    .Q(\u_inv.f_next[183] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_2 _40876_ (.RESET_B(net97),
    .D(_00155_),
    .Q(\u_inv.f_next[184] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _40877_ (.RESET_B(net96),
    .D(_00156_),
    .Q(\u_inv.f_next[185] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _40878_ (.RESET_B(net95),
    .D(_00157_),
    .Q(\u_inv.f_next[186] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _40879_ (.RESET_B(net94),
    .D(_00158_),
    .Q(\u_inv.f_next[187] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _40880_ (.RESET_B(net93),
    .D(_00159_),
    .Q(\u_inv.f_next[188] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _40881_ (.RESET_B(net92),
    .D(_00160_),
    .Q(\u_inv.f_next[189] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _40882_ (.RESET_B(net91),
    .D(_00161_),
    .Q(\u_inv.f_next[190] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _40883_ (.RESET_B(net90),
    .D(_00162_),
    .Q(\u_inv.f_next[191] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _40884_ (.RESET_B(net89),
    .D(_00163_),
    .Q(\u_inv.f_next[192] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _40885_ (.RESET_B(net88),
    .D(_00164_),
    .Q(\u_inv.f_next[193] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _40886_ (.RESET_B(net87),
    .D(_00165_),
    .Q(\u_inv.f_next[194] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _40887_ (.RESET_B(net86),
    .D(_00166_),
    .Q(\u_inv.f_next[195] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _40888_ (.RESET_B(net85),
    .D(_00167_),
    .Q(\u_inv.f_next[196] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _40889_ (.RESET_B(net84),
    .D(_00168_),
    .Q(\u_inv.f_next[197] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _40890_ (.RESET_B(net83),
    .D(_00169_),
    .Q(\u_inv.f_next[198] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _40891_ (.RESET_B(net82),
    .D(_00170_),
    .Q(\u_inv.f_next[199] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _40892_ (.RESET_B(net81),
    .D(_00171_),
    .Q(\u_inv.f_next[200] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _40893_ (.RESET_B(net80),
    .D(_00172_),
    .Q(\u_inv.f_next[201] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _40894_ (.RESET_B(net79),
    .D(net3301),
    .Q(\u_inv.f_next[202] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _40895_ (.RESET_B(net78),
    .D(_00174_),
    .Q(\u_inv.f_next[203] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _40896_ (.RESET_B(net77),
    .D(_00175_),
    .Q(\u_inv.f_next[204] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _40897_ (.RESET_B(net76),
    .D(_00176_),
    .Q(\u_inv.f_next[205] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _40898_ (.RESET_B(net75),
    .D(_00177_),
    .Q(\u_inv.f_next[206] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _40899_ (.RESET_B(net74),
    .D(_00178_),
    .Q(\u_inv.f_next[207] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _40900_ (.RESET_B(net73),
    .D(_00179_),
    .Q(\u_inv.f_next[208] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _40901_ (.RESET_B(net72),
    .D(_00180_),
    .Q(\u_inv.f_next[209] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _40902_ (.RESET_B(net71),
    .D(_00181_),
    .Q(\u_inv.f_next[210] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _40903_ (.RESET_B(net70),
    .D(_00182_),
    .Q(\u_inv.f_next[211] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _40904_ (.RESET_B(net69),
    .D(_00183_),
    .Q(\u_inv.f_next[212] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _40905_ (.RESET_B(net68),
    .D(_00184_),
    .Q(\u_inv.f_next[213] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _40906_ (.RESET_B(net67),
    .D(_00185_),
    .Q(\u_inv.f_next[214] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _40907_ (.RESET_B(net66),
    .D(_00186_),
    .Q(\u_inv.f_next[215] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _40908_ (.RESET_B(net65),
    .D(_00187_),
    .Q(\u_inv.f_next[216] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _40909_ (.RESET_B(net64),
    .D(_00188_),
    .Q(\u_inv.f_next[217] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _40910_ (.RESET_B(net63),
    .D(_00189_),
    .Q(\u_inv.f_next[218] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _40911_ (.RESET_B(net62),
    .D(_00190_),
    .Q(\u_inv.f_next[219] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _40912_ (.RESET_B(net61),
    .D(_00191_),
    .Q(\u_inv.f_next[220] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_2 _40913_ (.RESET_B(net60),
    .D(_00192_),
    .Q(\u_inv.f_next[221] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _40914_ (.RESET_B(net59),
    .D(_00193_),
    .Q(\u_inv.f_next[222] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _40915_ (.RESET_B(net58),
    .D(_00194_),
    .Q(\u_inv.f_next[223] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _40916_ (.RESET_B(net57),
    .D(_00195_),
    .Q(\u_inv.f_next[224] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _40917_ (.RESET_B(net56),
    .D(_00196_),
    .Q(\u_inv.f_next[225] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _40918_ (.RESET_B(net55),
    .D(_00197_),
    .Q(\u_inv.f_next[226] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _40919_ (.RESET_B(net54),
    .D(_00198_),
    .Q(\u_inv.f_next[227] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _40920_ (.RESET_B(net53),
    .D(_00199_),
    .Q(\u_inv.f_next[228] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _40921_ (.RESET_B(net52),
    .D(_00200_),
    .Q(\u_inv.f_next[229] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _40922_ (.RESET_B(net51),
    .D(_00201_),
    .Q(\u_inv.f_next[230] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _40923_ (.RESET_B(net50),
    .D(_00202_),
    .Q(\u_inv.f_next[231] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _40924_ (.RESET_B(net49),
    .D(_00203_),
    .Q(\u_inv.f_next[232] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _40925_ (.RESET_B(net48),
    .D(_00204_),
    .Q(\u_inv.f_next[233] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _40926_ (.RESET_B(net47),
    .D(_00205_),
    .Q(\u_inv.f_next[234] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _40927_ (.RESET_B(net46),
    .D(_00206_),
    .Q(\u_inv.f_next[235] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _40928_ (.RESET_B(net45),
    .D(_00207_),
    .Q(\u_inv.f_next[236] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _40929_ (.RESET_B(net44),
    .D(_00208_),
    .Q(\u_inv.f_next[237] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _40930_ (.RESET_B(net43),
    .D(_00209_),
    .Q(\u_inv.f_next[238] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _40931_ (.RESET_B(net42),
    .D(_00210_),
    .Q(\u_inv.f_next[239] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _40932_ (.RESET_B(net41),
    .D(_00211_),
    .Q(\u_inv.f_next[240] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _40933_ (.RESET_B(net40),
    .D(_00212_),
    .Q(\u_inv.f_next[241] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _40934_ (.RESET_B(net39),
    .D(_00213_),
    .Q(\u_inv.f_next[242] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _40935_ (.RESET_B(net38),
    .D(_00214_),
    .Q(\u_inv.f_next[243] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _40936_ (.RESET_B(net37),
    .D(_00215_),
    .Q(\u_inv.f_next[244] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _40937_ (.RESET_B(net36),
    .D(_00216_),
    .Q(\u_inv.f_next[245] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _40938_ (.RESET_B(net35),
    .D(_00217_),
    .Q(\u_inv.f_next[246] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _40939_ (.RESET_B(net34),
    .D(_00218_),
    .Q(\u_inv.f_next[247] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _40940_ (.RESET_B(net33),
    .D(_00219_),
    .Q(\u_inv.f_next[248] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _40941_ (.RESET_B(net32),
    .D(_00220_),
    .Q(\u_inv.f_next[249] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _40942_ (.RESET_B(net31),
    .D(_00221_),
    .Q(\u_inv.f_next[250] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _40943_ (.RESET_B(net30),
    .D(_00222_),
    .Q(\u_inv.f_next[251] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _40944_ (.RESET_B(net29),
    .D(_00223_),
    .Q(\u_inv.f_next[252] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _40945_ (.RESET_B(net28),
    .D(_00224_),
    .Q(\u_inv.f_next[253] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _40946_ (.RESET_B(net27),
    .D(net1843),
    .Q(\u_inv.f_next[254] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _40947_ (.RESET_B(net26),
    .D(_00226_),
    .Q(\u_inv.f_next[255] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _40948_ (.RESET_B(net5904),
    .D(net1075),
    .Q(\u_inv.input_valid ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _40949_ (.RESET_B(net5904),
    .D(_00228_),
    .Q(\state[0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _40950_ (.RESET_B(net5897),
    .D(_00229_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _40951_ (.RESET_B(net5904),
    .D(net2549),
    .Q(\byte_cnt[0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _40952_ (.RESET_B(net5904),
    .D(net1183),
    .Q(\byte_cnt[1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _40953_ (.RESET_B(net5906),
    .D(_00232_),
    .Q(\byte_cnt[2] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _40954_ (.RESET_B(net5905),
    .D(_00233_),
    .Q(\byte_cnt[3] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _40955_ (.RESET_B(net5905),
    .D(net1154),
    .Q(\byte_cnt[4] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _40956_ (.RESET_B(net5904),
    .D(_20878_[0]),
    .Q(inv_go),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _40957_ (.RESET_B(net5894),
    .D(_00235_),
    .Q(\shift_reg[0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _40958_ (.RESET_B(net5894),
    .D(_00236_),
    .Q(\shift_reg[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _40959_ (.RESET_B(net5895),
    .D(_00237_),
    .Q(\shift_reg[2] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _40960_ (.RESET_B(net5896),
    .D(_00238_),
    .Q(\shift_reg[3] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _40961_ (.RESET_B(net5896),
    .D(_00239_),
    .Q(\shift_reg[4] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _40962_ (.RESET_B(net5896),
    .D(_00240_),
    .Q(\shift_reg[5] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _40963_ (.RESET_B(net5895),
    .D(_00241_),
    .Q(\shift_reg[6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _40964_ (.RESET_B(net5896),
    .D(_00242_),
    .Q(\shift_reg[7] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _40965_ (.RESET_B(net5893),
    .D(_00243_),
    .Q(\shift_reg[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _40966_ (.RESET_B(net5893),
    .D(_00244_),
    .Q(\shift_reg[9] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _40967_ (.RESET_B(net5895),
    .D(net1313),
    .Q(\shift_reg[10] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _40968_ (.RESET_B(net5891),
    .D(net1288),
    .Q(\shift_reg[11] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _40969_ (.RESET_B(net5901),
    .D(net1327),
    .Q(\shift_reg[12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _40970_ (.RESET_B(net5890),
    .D(net1630),
    .Q(\shift_reg[13] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _40971_ (.RESET_B(net5891),
    .D(net2320),
    .Q(\shift_reg[14] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _40972_ (.RESET_B(net5889),
    .D(_00250_),
    .Q(\shift_reg[15] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _40973_ (.RESET_B(net5885),
    .D(net2461),
    .Q(\shift_reg[16] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _40974_ (.RESET_B(net5885),
    .D(net2229),
    .Q(\shift_reg[17] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _40975_ (.RESET_B(net5886),
    .D(net2212),
    .Q(\shift_reg[18] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _40976_ (.RESET_B(net5910),
    .D(net1911),
    .Q(\shift_reg[19] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _40977_ (.RESET_B(net5909),
    .D(net1963),
    .Q(\shift_reg[20] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _40978_ (.RESET_B(net5909),
    .D(net2127),
    .Q(\shift_reg[21] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _40979_ (.RESET_B(net5909),
    .D(net2029),
    .Q(\shift_reg[22] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _40980_ (.RESET_B(net5910),
    .D(net1466),
    .Q(\shift_reg[23] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _40981_ (.RESET_B(net5909),
    .D(net1732),
    .Q(\shift_reg[24] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _40982_ (.RESET_B(net5911),
    .D(net2162),
    .Q(\shift_reg[25] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _40983_ (.RESET_B(net5911),
    .D(net1501),
    .Q(\shift_reg[26] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _40984_ (.RESET_B(net5911),
    .D(net1901),
    .Q(\shift_reg[27] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _40985_ (.RESET_B(net5911),
    .D(_00263_),
    .Q(\shift_reg[28] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _40986_ (.RESET_B(net5911),
    .D(_00264_),
    .Q(\shift_reg[29] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _40987_ (.RESET_B(net5911),
    .D(_00265_),
    .Q(\shift_reg[30] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _40988_ (.RESET_B(net5911),
    .D(_00266_),
    .Q(\shift_reg[31] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _40989_ (.RESET_B(net5913),
    .D(_00267_),
    .Q(\shift_reg[32] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _40990_ (.RESET_B(net5914),
    .D(net1559),
    .Q(\shift_reg[33] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _40991_ (.RESET_B(net5931),
    .D(net1379),
    .Q(\shift_reg[34] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _40992_ (.RESET_B(net5929),
    .D(_00270_),
    .Q(\shift_reg[35] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _40993_ (.RESET_B(net5929),
    .D(net2076),
    .Q(\shift_reg[36] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _40994_ (.RESET_B(net5929),
    .D(net1450),
    .Q(\shift_reg[37] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _40995_ (.RESET_B(net5930),
    .D(net1355),
    .Q(\shift_reg[38] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _40996_ (.RESET_B(net5930),
    .D(_00274_),
    .Q(\shift_reg[39] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _40997_ (.RESET_B(net5930),
    .D(net2405),
    .Q(\shift_reg[40] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _40998_ (.RESET_B(net5933),
    .D(_00276_),
    .Q(\shift_reg[41] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _40999_ (.RESET_B(net5933),
    .D(_00277_),
    .Q(\shift_reg[42] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _41000_ (.RESET_B(net5934),
    .D(_00278_),
    .Q(\shift_reg[43] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _41001_ (.RESET_B(net5948),
    .D(net1866),
    .Q(\shift_reg[44] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _41002_ (.RESET_B(net5933),
    .D(_00280_),
    .Q(\shift_reg[45] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _41003_ (.RESET_B(net5934),
    .D(_00281_),
    .Q(\shift_reg[46] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _41004_ (.RESET_B(net5934),
    .D(net2313),
    .Q(\shift_reg[47] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _41005_ (.RESET_B(net5948),
    .D(net1968),
    .Q(\shift_reg[48] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _41006_ (.RESET_B(net5946),
    .D(net1311),
    .Q(\shift_reg[49] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _41007_ (.RESET_B(net5946),
    .D(net1517),
    .Q(\shift_reg[50] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _41008_ (.RESET_B(net5946),
    .D(net1417),
    .Q(\shift_reg[51] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _41009_ (.RESET_B(net5946),
    .D(_00287_),
    .Q(\shift_reg[52] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _41010_ (.RESET_B(net5950),
    .D(net2219),
    .Q(\shift_reg[53] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _41011_ (.RESET_B(net5951),
    .D(_00289_),
    .Q(\shift_reg[54] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _41012_ (.RESET_B(net5946),
    .D(_00290_),
    .Q(\shift_reg[55] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _41013_ (.RESET_B(net5947),
    .D(_00291_),
    .Q(\shift_reg[56] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _41014_ (.RESET_B(net5950),
    .D(_00292_),
    .Q(\shift_reg[57] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _41015_ (.RESET_B(net5967),
    .D(_00293_),
    .Q(\shift_reg[58] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _41016_ (.RESET_B(net5967),
    .D(_00294_),
    .Q(\shift_reg[59] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _41017_ (.RESET_B(net5967),
    .D(net1738),
    .Q(\shift_reg[60] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _41018_ (.RESET_B(net5981),
    .D(net1916),
    .Q(\shift_reg[61] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _41019_ (.RESET_B(net5981),
    .D(_00297_),
    .Q(\shift_reg[62] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _41020_ (.RESET_B(net5966),
    .D(net1953),
    .Q(\shift_reg[63] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _41021_ (.RESET_B(net5982),
    .D(net1480),
    .Q(\shift_reg[64] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _41022_ (.RESET_B(net5982),
    .D(net1464),
    .Q(\shift_reg[65] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _41023_ (.RESET_B(net5989),
    .D(_00301_),
    .Q(\shift_reg[66] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _41024_ (.RESET_B(net5982),
    .D(net1330),
    .Q(\shift_reg[67] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _41025_ (.RESET_B(net5982),
    .D(net2074),
    .Q(\shift_reg[68] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_2 _41026_ (.RESET_B(net5968),
    .D(net1854),
    .Q(\shift_reg[69] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _41027_ (.RESET_B(net5988),
    .D(net1511),
    .Q(\shift_reg[70] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _41028_ (.RESET_B(net5983),
    .D(net1811),
    .Q(\shift_reg[71] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _41029_ (.RESET_B(net5988),
    .D(_00307_),
    .Q(\shift_reg[72] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_2 _41030_ (.RESET_B(net5988),
    .D(_00308_),
    .Q(\shift_reg[73] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _41031_ (.RESET_B(net5991),
    .D(_00309_),
    .Q(\shift_reg[74] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _41032_ (.RESET_B(net5984),
    .D(_00310_),
    .Q(\shift_reg[75] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _41033_ (.RESET_B(net5984),
    .D(_00311_),
    .Q(\shift_reg[76] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _41034_ (.RESET_B(net5998),
    .D(_00312_),
    .Q(\shift_reg[77] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _41035_ (.RESET_B(net5992),
    .D(_00313_),
    .Q(\shift_reg[78] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _41036_ (.RESET_B(net5998),
    .D(_00314_),
    .Q(\shift_reg[79] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _41037_ (.RESET_B(net6001),
    .D(net1904),
    .Q(\shift_reg[80] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_2 _41038_ (.RESET_B(net5996),
    .D(net2743),
    .Q(\shift_reg[81] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_2 _41039_ (.RESET_B(net5996),
    .D(net2311),
    .Q(\shift_reg[82] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_2 _41040_ (.RESET_B(net5998),
    .D(_00318_),
    .Q(\shift_reg[83] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _41041_ (.RESET_B(net6019),
    .D(net1377),
    .Q(\shift_reg[84] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _41042_ (.RESET_B(net6005),
    .D(_00320_),
    .Q(\shift_reg[85] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _41043_ (.RESET_B(net6007),
    .D(net1493),
    .Q(\shift_reg[86] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _41044_ (.RESET_B(net6019),
    .D(net1396),
    .Q(\shift_reg[87] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _41045_ (.RESET_B(net6019),
    .D(_00323_),
    .Q(\shift_reg[88] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _41046_ (.RESET_B(net6016),
    .D(net2116),
    .Q(\shift_reg[89] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _41047_ (.RESET_B(net6016),
    .D(_00325_),
    .Q(\shift_reg[90] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_2 _41048_ (.RESET_B(net6023),
    .D(net2375),
    .Q(\shift_reg[91] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_2 _41049_ (.RESET_B(net6020),
    .D(_00327_),
    .Q(\shift_reg[92] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _41050_ (.RESET_B(net6020),
    .D(net2401),
    .Q(\shift_reg[93] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _41051_ (.RESET_B(net6018),
    .D(_00329_),
    .Q(\shift_reg[94] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_2 _41052_ (.RESET_B(net6026),
    .D(_00330_),
    .Q(\shift_reg[95] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _41053_ (.RESET_B(net6027),
    .D(net2231),
    .Q(\shift_reg[96] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _41054_ (.RESET_B(net6013),
    .D(_00332_),
    .Q(\shift_reg[97] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _41055_ (.RESET_B(net6013),
    .D(net1995),
    .Q(\shift_reg[98] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _41056_ (.RESET_B(net6026),
    .D(net1710),
    .Q(\shift_reg[99] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _41057_ (.RESET_B(net6027),
    .D(net2260),
    .Q(\shift_reg[100] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _41058_ (.RESET_B(net6028),
    .D(net2225),
    .Q(\shift_reg[101] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _41059_ (.RESET_B(net6028),
    .D(net1375),
    .Q(\shift_reg[102] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _41060_ (.RESET_B(net6023),
    .D(_00338_),
    .Q(\shift_reg[103] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _41061_ (.RESET_B(net6023),
    .D(net1951),
    .Q(\shift_reg[104] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _41062_ (.RESET_B(net6028),
    .D(net2095),
    .Q(\shift_reg[105] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _41063_ (.RESET_B(net6025),
    .D(_00341_),
    .Q(\shift_reg[106] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _41064_ (.RESET_B(net6023),
    .D(_00342_),
    .Q(\shift_reg[107] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _41065_ (.RESET_B(net6025),
    .D(net1989),
    .Q(\shift_reg[108] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _41066_ (.RESET_B(net6024),
    .D(net1937),
    .Q(\shift_reg[109] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _41067_ (.RESET_B(net6025),
    .D(_00345_),
    .Q(\shift_reg[110] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _41068_ (.RESET_B(net6025),
    .D(net2024),
    .Q(\shift_reg[111] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_2 _41069_ (.RESET_B(net6023),
    .D(_00347_),
    .Q(\shift_reg[112] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _41070_ (.RESET_B(net6024),
    .D(net2011),
    .Q(\shift_reg[113] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _41071_ (.RESET_B(net6022),
    .D(net1734),
    .Q(\shift_reg[114] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _41072_ (.RESET_B(net6020),
    .D(net2005),
    .Q(\shift_reg[115] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_2 _41073_ (.RESET_B(net6021),
    .D(net1585),
    .Q(\shift_reg[116] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _41074_ (.RESET_B(net6021),
    .D(_00352_),
    .Q(\shift_reg[117] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _41075_ (.RESET_B(net6022),
    .D(net1785),
    .Q(\shift_reg[118] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_2 _41076_ (.RESET_B(net6022),
    .D(net1891),
    .Q(\shift_reg[119] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _41077_ (.RESET_B(net6018),
    .D(net1801),
    .Q(\shift_reg[120] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _41078_ (.RESET_B(net6017),
    .D(_00356_),
    .Q(\shift_reg[121] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _41079_ (.RESET_B(net6017),
    .D(_00357_),
    .Q(\shift_reg[122] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _41080_ (.RESET_B(net6006),
    .D(net1478),
    .Q(\shift_reg[123] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _41081_ (.RESET_B(net6008),
    .D(net1472),
    .Q(\shift_reg[124] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _41082_ (.RESET_B(net6008),
    .D(net1414),
    .Q(\shift_reg[125] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_2 _41083_ (.RESET_B(net6008),
    .D(_00361_),
    .Q(\shift_reg[126] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _41084_ (.RESET_B(net6001),
    .D(net1390),
    .Q(\shift_reg[127] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _41085_ (.RESET_B(net6008),
    .D(_00363_),
    .Q(\shift_reg[128] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_2 _41086_ (.RESET_B(net6006),
    .D(_00364_),
    .Q(\shift_reg[129] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _41087_ (.RESET_B(net6002),
    .D(net1791),
    .Q(\shift_reg[130] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _41088_ (.RESET_B(net6005),
    .D(_00366_),
    .Q(\shift_reg[131] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _41089_ (.RESET_B(net6001),
    .D(_00367_),
    .Q(\shift_reg[132] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _41090_ (.RESET_B(net6002),
    .D(_00368_),
    .Q(\shift_reg[133] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _41091_ (.RESET_B(net5999),
    .D(net1399),
    .Q(\shift_reg[134] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_2 _41092_ (.RESET_B(net6004),
    .D(_00370_),
    .Q(\shift_reg[135] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _41093_ (.RESET_B(net5999),
    .D(net1939),
    .Q(\shift_reg[136] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _41094_ (.RESET_B(net5999),
    .D(net2045),
    .Q(\shift_reg[137] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _41095_ (.RESET_B(net5999),
    .D(_00373_),
    .Q(\shift_reg[138] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _41096_ (.RESET_B(net5999),
    .D(_00374_),
    .Q(\shift_reg[139] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _41097_ (.RESET_B(net5999),
    .D(_00375_),
    .Q(\shift_reg[140] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _41098_ (.RESET_B(net5999),
    .D(net2129),
    .Q(\shift_reg[141] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_2 _41099_ (.RESET_B(net5999),
    .D(_00377_),
    .Q(\shift_reg[142] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_2 _41100_ (.RESET_B(net6003),
    .D(_00378_),
    .Q(\shift_reg[143] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _41101_ (.RESET_B(net5992),
    .D(net1362),
    .Q(\shift_reg[144] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _41102_ (.RESET_B(net5992),
    .D(net1671),
    .Q(\shift_reg[145] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _41103_ (.RESET_B(net5993),
    .D(net1567),
    .Q(\shift_reg[146] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _41104_ (.RESET_B(net5991),
    .D(net1947),
    .Q(\shift_reg[147] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _41105_ (.RESET_B(net5993),
    .D(net2143),
    .Q(\shift_reg[148] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _41106_ (.RESET_B(net5993),
    .D(net1872),
    .Q(\shift_reg[149] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _41107_ (.RESET_B(net5993),
    .D(net2233),
    .Q(\shift_reg[150] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _41108_ (.RESET_B(net5987),
    .D(_00386_),
    .Q(\shift_reg[151] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _41109_ (.RESET_B(net5987),
    .D(_00387_),
    .Q(\shift_reg[152] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _41110_ (.RESET_B(net5987),
    .D(net1899),
    .Q(\shift_reg[153] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _41111_ (.RESET_B(net5990),
    .D(_00389_),
    .Q(\shift_reg[154] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _41112_ (.RESET_B(net5989),
    .D(net1767),
    .Q(\shift_reg[155] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _41113_ (.RESET_B(net5987),
    .D(_00391_),
    .Q(\shift_reg[156] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _41114_ (.RESET_B(net5977),
    .D(net1446),
    .Q(\shift_reg[157] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _41115_ (.RESET_B(net5989),
    .D(net2054),
    .Q(\shift_reg[158] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _41116_ (.RESET_B(net5977),
    .D(net1401),
    .Q(\shift_reg[159] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _41117_ (.RESET_B(net5995),
    .D(net2195),
    .Q(\shift_reg[160] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _41118_ (.RESET_B(net5989),
    .D(_00396_),
    .Q(\shift_reg[161] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _41119_ (.RESET_B(net5977),
    .D(net1409),
    .Q(\shift_reg[162] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _41120_ (.RESET_B(net5975),
    .D(net1308),
    .Q(\shift_reg[163] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _41121_ (.RESET_B(net5977),
    .D(net1868),
    .Q(\shift_reg[164] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _41122_ (.RESET_B(net5977),
    .D(_00400_),
    .Q(\shift_reg[165] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _41123_ (.RESET_B(net5975),
    .D(net1392),
    .Q(\shift_reg[166] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _41124_ (.RESET_B(net5975),
    .D(_00402_),
    .Q(\shift_reg[167] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _41125_ (.RESET_B(net5975),
    .D(_00403_),
    .Q(\shift_reg[168] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _41126_ (.RESET_B(net5975),
    .D(net2082),
    .Q(\shift_reg[169] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _41127_ (.RESET_B(net5972),
    .D(_00405_),
    .Q(\shift_reg[170] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _41128_ (.RESET_B(net5972),
    .D(net2013),
    .Q(\shift_reg[171] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _41129_ (.RESET_B(net5971),
    .D(_00407_),
    .Q(\shift_reg[172] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _41130_ (.RESET_B(net5971),
    .D(_00408_),
    .Q(\shift_reg[173] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _41131_ (.RESET_B(net5969),
    .D(_00409_),
    .Q(\shift_reg[174] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _41132_ (.RESET_B(net5971),
    .D(_00410_),
    .Q(\shift_reg[175] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _41133_ (.RESET_B(net5974),
    .D(net1763),
    .Q(\shift_reg[176] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _41134_ (.RESET_B(net5969),
    .D(net1752),
    .Q(\shift_reg[177] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _41135_ (.RESET_B(net5969),
    .D(net1371),
    .Q(\shift_reg[178] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _41136_ (.RESET_B(net5974),
    .D(net2009),
    .Q(\shift_reg[179] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _41137_ (.RESET_B(net5963),
    .D(net1615),
    .Q(\shift_reg[180] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _41138_ (.RESET_B(net5970),
    .D(net2324),
    .Q(\shift_reg[181] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _41139_ (.RESET_B(net5962),
    .D(_00417_),
    .Q(\shift_reg[182] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _41140_ (.RESET_B(net5963),
    .D(net1602),
    .Q(\shift_reg[183] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _41141_ (.RESET_B(net5960),
    .D(net1394),
    .Q(\shift_reg[184] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _41142_ (.RESET_B(net5962),
    .D(_00420_),
    .Q(\shift_reg[185] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _41143_ (.RESET_B(net5964),
    .D(_00421_),
    .Q(\shift_reg[186] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _41144_ (.RESET_B(net5961),
    .D(_00422_),
    .Q(\shift_reg[187] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_2 _41145_ (.RESET_B(net5960),
    .D(_00423_),
    .Q(\shift_reg[188] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _41146_ (.RESET_B(net5958),
    .D(net1882),
    .Q(\shift_reg[189] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _41147_ (.RESET_B(net5961),
    .D(_00425_),
    .Q(\shift_reg[190] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _41148_ (.RESET_B(net5961),
    .D(_00426_),
    .Q(\shift_reg[191] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _41149_ (.RESET_B(net5960),
    .D(_00427_),
    .Q(\shift_reg[192] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _41150_ (.RESET_B(net5955),
    .D(net1863),
    .Q(\shift_reg[193] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _41151_ (.RESET_B(net5957),
    .D(net1659),
    .Q(\shift_reg[194] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _41152_ (.RESET_B(net5957),
    .D(net2108),
    .Q(\shift_reg[195] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _41153_ (.RESET_B(net5956),
    .D(net2125),
    .Q(\shift_reg[196] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _41154_ (.RESET_B(net5955),
    .D(_00432_),
    .Q(\shift_reg[197] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _41155_ (.RESET_B(net5955),
    .D(net1454),
    .Q(\shift_reg[198] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _41156_ (.RESET_B(net5956),
    .D(net2359),
    .Q(\shift_reg[199] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _41157_ (.RESET_B(net5956),
    .D(_00435_),
    .Q(\shift_reg[200] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_2 _41158_ (.RESET_B(net5954),
    .D(net1836),
    .Q(\shift_reg[201] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _41159_ (.RESET_B(net5953),
    .D(_00437_),
    .Q(\shift_reg[202] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _41160_ (.RESET_B(net5953),
    .D(net1720),
    .Q(\shift_reg[203] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _41161_ (.RESET_B(net5942),
    .D(net1848),
    .Q(\shift_reg[204] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _41162_ (.RESET_B(net5954),
    .D(net1922),
    .Q(\shift_reg[205] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _41163_ (.RESET_B(net5954),
    .D(_00441_),
    .Q(\shift_reg[206] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _41164_ (.RESET_B(net5959),
    .D(net2412),
    .Q(\shift_reg[207] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _41165_ (.RESET_B(net5943),
    .D(net2122),
    .Q(\shift_reg[208] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _41166_ (.RESET_B(net5942),
    .D(net1787),
    .Q(\shift_reg[209] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _41167_ (.RESET_B(net5943),
    .D(net1544),
    .Q(\shift_reg[210] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _41168_ (.RESET_B(net5941),
    .D(net1519),
    .Q(\shift_reg[211] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_2 _41169_ (.RESET_B(net5942),
    .D(net1846),
    .Q(\shift_reg[212] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_2 _41170_ (.RESET_B(net5940),
    .D(_00448_),
    .Q(\shift_reg[213] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _41171_ (.RESET_B(net5939),
    .D(net2171),
    .Q(\shift_reg[214] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _41172_ (.RESET_B(net5939),
    .D(net1426),
    .Q(\shift_reg[215] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _41173_ (.RESET_B(net5938),
    .D(_00451_),
    .Q(\shift_reg[216] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _41174_ (.RESET_B(net5937),
    .D(net1669),
    .Q(\shift_reg[217] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _41175_ (.RESET_B(net5937),
    .D(_00453_),
    .Q(\shift_reg[218] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _41176_ (.RESET_B(net5938),
    .D(net2102),
    .Q(\shift_reg[219] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_2 _41177_ (.RESET_B(net5938),
    .D(_00455_),
    .Q(\shift_reg[220] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _41178_ (.RESET_B(net5937),
    .D(net1452),
    .Q(\shift_reg[221] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _41179_ (.RESET_B(net5936),
    .D(net1435),
    .Q(\shift_reg[222] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _41180_ (.RESET_B(net5936),
    .D(_00458_),
    .Q(\shift_reg[223] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _41181_ (.RESET_B(net5923),
    .D(net2057),
    .Q(\shift_reg[224] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _41182_ (.RESET_B(net5925),
    .D(_00460_),
    .Q(\shift_reg[225] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _41183_ (.RESET_B(net5923),
    .D(net1432),
    .Q(\shift_reg[226] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _41184_ (.RESET_B(net5924),
    .D(_00462_),
    .Q(\shift_reg[227] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _41185_ (.RESET_B(net5924),
    .D(net1809),
    .Q(\shift_reg[228] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _41186_ (.RESET_B(net5925),
    .D(net1430),
    .Q(\shift_reg[229] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _41187_ (.RESET_B(net5921),
    .D(_00465_),
    .Q(\shift_reg[230] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _41188_ (.RESET_B(net5926),
    .D(_00466_),
    .Q(\shift_reg[231] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _41189_ (.RESET_B(net5921),
    .D(_00467_),
    .Q(\shift_reg[232] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _41190_ (.RESET_B(net5922),
    .D(net1949),
    .Q(\shift_reg[233] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _41191_ (.RESET_B(net5921),
    .D(_00469_),
    .Q(\shift_reg[234] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _41192_ (.RESET_B(net5919),
    .D(net2644),
    .Q(\shift_reg[235] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _41193_ (.RESET_B(net5919),
    .D(_00471_),
    .Q(\shift_reg[236] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _41194_ (.RESET_B(net5919),
    .D(_00472_),
    .Q(\shift_reg[237] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _41195_ (.RESET_B(net5920),
    .D(net1981),
    .Q(\shift_reg[238] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _41196_ (.RESET_B(net5918),
    .D(net1428),
    .Q(\shift_reg[239] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _41197_ (.RESET_B(net5918),
    .D(net1829),
    .Q(\shift_reg[240] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _41198_ (.RESET_B(net5920),
    .D(_00476_),
    .Q(\shift_reg[241] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _41199_ (.RESET_B(net5916),
    .D(net1503),
    .Q(\shift_reg[242] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _41200_ (.RESET_B(net5917),
    .D(net1346),
    .Q(\shift_reg[243] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _41201_ (.RESET_B(net5916),
    .D(net1405),
    .Q(\shift_reg[244] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _41202_ (.RESET_B(net5917),
    .D(_00480_),
    .Q(\shift_reg[245] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _41203_ (.RESET_B(net5902),
    .D(_00481_),
    .Q(\shift_reg[246] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _41204_ (.RESET_B(net5902),
    .D(_00482_),
    .Q(\shift_reg[247] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _41205_ (.RESET_B(net5900),
    .D(_00483_),
    .Q(\shift_reg[248] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _41206_ (.RESET_B(net5900),
    .D(net1977),
    .Q(\shift_reg[249] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _41207_ (.RESET_B(net5900),
    .D(_00485_),
    .Q(\shift_reg[250] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _41208_ (.RESET_B(net5900),
    .D(_00486_),
    .Q(\shift_reg[251] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _41209_ (.RESET_B(net5916),
    .D(_00487_),
    .Q(\shift_reg[252] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _41210_ (.RESET_B(net5891),
    .D(net2304),
    .Q(\shift_reg[253] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _41211_ (.RESET_B(net5900),
    .D(net1403),
    .Q(\shift_reg[254] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _41212_ (.RESET_B(net5890),
    .D(_00490_),
    .Q(\shift_reg[255] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _41213_ (.RESET_B(net5888),
    .D(net1142),
    .Q(\shift_reg[256] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _41214_ (.RESET_B(net5888),
    .D(net1243),
    .Q(\shift_reg[257] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _41215_ (.RESET_B(net5889),
    .D(net1231),
    .Q(\shift_reg[258] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _41216_ (.RESET_B(net5888),
    .D(net1193),
    .Q(\shift_reg[259] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _41217_ (.RESET_B(net5889),
    .D(net1195),
    .Q(\shift_reg[260] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _41218_ (.RESET_B(net5890),
    .D(net1205),
    .Q(\shift_reg[261] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _41219_ (.RESET_B(net5883),
    .D(net1324),
    .Q(\shift_reg[262] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _41220_ (.RESET_B(net5883),
    .D(net1151),
    .Q(\shift_reg[263] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _41221_ (.RESET_B(net5895),
    .D(net1114),
    .Q(\shift_reg[264] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _41222_ (.RESET_B(net5894),
    .D(net1241),
    .Q(\shift_reg[265] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _41223_ (.RESET_B(net5895),
    .D(net1131),
    .Q(\shift_reg[266] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _41224_ (.RESET_B(net5894),
    .D(net1164),
    .Q(\shift_reg[267] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _41225_ (.RESET_B(net5898),
    .D(_00503_),
    .Q(\shift_reg[268] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _41226_ (.RESET_B(net5894),
    .D(net1218),
    .Q(\shift_reg[269] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _41227_ (.RESET_B(net5894),
    .D(net1116),
    .Q(\shift_reg[270] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _41228_ (.RESET_B(net5894),
    .D(net1118),
    .Q(\shift_reg[271] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _41229_ (.RESET_B(net5897),
    .D(_00507_),
    .Q(next_loaded),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _41230_ (.RESET_B(net5898),
    .D(net9),
    .Q(wr_prev),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _41231_ (.RESET_B(net5898),
    .D(net10),
    .Q(rd_prev),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _41232_ (.RESET_B(net24),
    .D(_00508_),
    .Q(\u_inv.f_next[256] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _41233_ (.RESET_B(net5903),
    .D(net3390),
    .Q(\u_inv.counter[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _41234_ (.RESET_B(net5897),
    .D(net3428),
    .Q(\u_inv.counter[2] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _41235_ (.RESET_B(net5896),
    .D(_00511_),
    .Q(\u_inv.counter[3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _41236_ (.RESET_B(net5897),
    .D(_00512_),
    .Q(\u_inv.counter[4] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _41237_ (.RESET_B(net5897),
    .D(net3073),
    .Q(\u_inv.counter[5] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _41238_ (.RESET_B(net5896),
    .D(_00514_),
    .Q(\u_inv.counter[6] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _41239_ (.RESET_B(net5899),
    .D(_00515_),
    .Q(\u_inv.counter[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _41240_ (.RESET_B(net5903),
    .D(_00516_),
    .Q(\u_inv.counter[8] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _41241_ (.RESET_B(net5903),
    .D(net2635),
    .Q(\u_inv.counter[9] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _41242_ (.RESET_B(net5886),
    .D(net1250),
    .Q(\inv_result[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _41243_ (.RESET_B(net5886),
    .D(_00519_),
    .Q(\inv_result[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _41244_ (.RESET_B(net5887),
    .D(_00520_),
    .Q(\inv_result[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _41245_ (.RESET_B(net5887),
    .D(_00521_),
    .Q(\inv_result[3] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _41246_ (.RESET_B(net5887),
    .D(_00522_),
    .Q(\inv_result[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _41247_ (.RESET_B(net5907),
    .D(_00523_),
    .Q(\inv_result[5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _41248_ (.RESET_B(net5907),
    .D(_00524_),
    .Q(\inv_result[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _41249_ (.RESET_B(net5907),
    .D(_00525_),
    .Q(\inv_result[7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _41250_ (.RESET_B(net5907),
    .D(_00526_),
    .Q(\inv_result[8] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _41251_ (.RESET_B(net5907),
    .D(_00527_),
    .Q(\inv_result[9] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _41252_ (.RESET_B(net5907),
    .D(_00528_),
    .Q(\inv_result[10] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _41253_ (.RESET_B(net5907),
    .D(_00529_),
    .Q(\inv_result[11] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _41254_ (.RESET_B(net5907),
    .D(_00530_),
    .Q(\inv_result[12] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _41255_ (.RESET_B(net5908),
    .D(_00531_),
    .Q(\inv_result[13] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _41256_ (.RESET_B(net5908),
    .D(_00532_),
    .Q(\inv_result[14] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _41257_ (.RESET_B(net5908),
    .D(_00533_),
    .Q(\inv_result[15] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _41258_ (.RESET_B(net5908),
    .D(_00534_),
    .Q(\inv_result[16] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _41259_ (.RESET_B(net5914),
    .D(net2176),
    .Q(\inv_result[17] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _41260_ (.RESET_B(net5929),
    .D(_00536_),
    .Q(\inv_result[18] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _41261_ (.RESET_B(net5932),
    .D(_00537_),
    .Q(\inv_result[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _41262_ (.RESET_B(net5914),
    .D(_00538_),
    .Q(\inv_result[20] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _41263_ (.RESET_B(net5929),
    .D(_00539_),
    .Q(\inv_result[21] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _41264_ (.RESET_B(net5932),
    .D(_00540_),
    .Q(\inv_result[22] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _41265_ (.RESET_B(net5929),
    .D(_00541_),
    .Q(\inv_result[23] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _41266_ (.RESET_B(net5930),
    .D(_00542_),
    .Q(\inv_result[24] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _41267_ (.RESET_B(net5930),
    .D(_00543_),
    .Q(\inv_result[25] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _41268_ (.RESET_B(net5930),
    .D(_00544_),
    .Q(\inv_result[26] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _41269_ (.RESET_B(net5932),
    .D(_00545_),
    .Q(\inv_result[27] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _41270_ (.RESET_B(net5932),
    .D(_00546_),
    .Q(\inv_result[28] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _41271_ (.RESET_B(net5932),
    .D(_00547_),
    .Q(\inv_result[29] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _41272_ (.RESET_B(net5935),
    .D(_00548_),
    .Q(\inv_result[30] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _41273_ (.RESET_B(net5935),
    .D(_00549_),
    .Q(\inv_result[31] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _41274_ (.RESET_B(net5948),
    .D(_00550_),
    .Q(\inv_result[32] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _41275_ (.RESET_B(net5949),
    .D(_00551_),
    .Q(\inv_result[33] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _41276_ (.RESET_B(net5946),
    .D(_00552_),
    .Q(\inv_result[34] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _41277_ (.RESET_B(net5949),
    .D(_00553_),
    .Q(\inv_result[35] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _41278_ (.RESET_B(net5949),
    .D(_00554_),
    .Q(\inv_result[36] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _41279_ (.RESET_B(net5947),
    .D(_00555_),
    .Q(\inv_result[37] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _41280_ (.RESET_B(net5949),
    .D(_00556_),
    .Q(\inv_result[38] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _41281_ (.RESET_B(net5949),
    .D(_00557_),
    .Q(\inv_result[39] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _41282_ (.RESET_B(net5946),
    .D(_00558_),
    .Q(\inv_result[40] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _41283_ (.RESET_B(net5952),
    .D(_00559_),
    .Q(\inv_result[41] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _41284_ (.RESET_B(net5952),
    .D(_00560_),
    .Q(\inv_result[42] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _41285_ (.RESET_B(net5950),
    .D(_00561_),
    .Q(\inv_result[43] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _41286_ (.RESET_B(net5966),
    .D(_00562_),
    .Q(\inv_result[44] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _41287_ (.RESET_B(net5968),
    .D(_00563_),
    .Q(\inv_result[45] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _41288_ (.RESET_B(net5966),
    .D(_00564_),
    .Q(\inv_result[46] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _41289_ (.RESET_B(net5966),
    .D(_00565_),
    .Q(\inv_result[47] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_1 _41290_ (.RESET_B(net5982),
    .D(_00566_),
    .Q(\inv_result[48] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _41291_ (.RESET_B(net5986),
    .D(_00567_),
    .Q(\inv_result[49] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_1 _41292_ (.RESET_B(net5983),
    .D(_00568_),
    .Q(\inv_result[50] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _41293_ (.RESET_B(net5983),
    .D(_00569_),
    .Q(\inv_result[51] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_2 _41294_ (.RESET_B(net5986),
    .D(_00570_),
    .Q(\inv_result[52] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _41295_ (.RESET_B(net5983),
    .D(_00571_),
    .Q(\inv_result[53] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _41296_ (.RESET_B(net5983),
    .D(_00572_),
    .Q(\inv_result[54] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _41297_ (.RESET_B(net5982),
    .D(_00573_),
    .Q(\inv_result[55] ),
    .CLK(clknet_leaf_179_clk));
 sg13g2_dfrbpq_1 _41298_ (.RESET_B(net5983),
    .D(_00574_),
    .Q(\inv_result[56] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _41299_ (.RESET_B(net5988),
    .D(_00575_),
    .Q(\inv_result[57] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _41300_ (.RESET_B(net5984),
    .D(_00576_),
    .Q(\inv_result[58] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _41301_ (.RESET_B(net5985),
    .D(_00577_),
    .Q(\inv_result[59] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _41302_ (.RESET_B(net5984),
    .D(_00578_),
    .Q(\inv_result[60] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _41303_ (.RESET_B(net5984),
    .D(_00579_),
    .Q(\inv_result[61] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _41304_ (.RESET_B(net5984),
    .D(_00580_),
    .Q(\inv_result[62] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _41305_ (.RESET_B(net5996),
    .D(_00581_),
    .Q(\inv_result[63] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _41306_ (.RESET_B(net5997),
    .D(_00582_),
    .Q(\inv_result[64] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _41307_ (.RESET_B(net5996),
    .D(_00583_),
    .Q(\inv_result[65] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _41308_ (.RESET_B(net5997),
    .D(_00584_),
    .Q(\inv_result[66] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _41309_ (.RESET_B(net5996),
    .D(_00585_),
    .Q(\inv_result[67] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _41310_ (.RESET_B(net6005),
    .D(_00586_),
    .Q(\inv_result[68] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _41311_ (.RESET_B(net6012),
    .D(_00587_),
    .Q(\inv_result[69] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _41312_ (.RESET_B(net6007),
    .D(_00588_),
    .Q(\inv_result[70] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _41313_ (.RESET_B(net6007),
    .D(_00589_),
    .Q(\inv_result[71] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _41314_ (.RESET_B(net6012),
    .D(_00590_),
    .Q(\inv_result[72] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _41315_ (.RESET_B(net6016),
    .D(_00591_),
    .Q(\inv_result[73] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _41316_ (.RESET_B(net6016),
    .D(_00592_),
    .Q(\inv_result[74] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_1 _41317_ (.RESET_B(net6020),
    .D(_00593_),
    .Q(\inv_result[75] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _41318_ (.RESET_B(net6020),
    .D(_00594_),
    .Q(\inv_result[76] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _41319_ (.RESET_B(net6019),
    .D(_00595_),
    .Q(\inv_result[77] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _41320_ (.RESET_B(net6019),
    .D(_00596_),
    .Q(\inv_result[78] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _41321_ (.RESET_B(net6019),
    .D(_00597_),
    .Q(\inv_result[79] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _41322_ (.RESET_B(net6015),
    .D(_00598_),
    .Q(\inv_result[80] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _41323_ (.RESET_B(net6015),
    .D(_00599_),
    .Q(\inv_result[81] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _41324_ (.RESET_B(net6015),
    .D(_00600_),
    .Q(\inv_result[82] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _41325_ (.RESET_B(net6013),
    .D(_00601_),
    .Q(\inv_result[83] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _41326_ (.RESET_B(net6027),
    .D(_00602_),
    .Q(\inv_result[84] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _41327_ (.RESET_B(net6014),
    .D(_00603_),
    .Q(\inv_result[85] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _41328_ (.RESET_B(net6014),
    .D(_00604_),
    .Q(\inv_result[86] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _41329_ (.RESET_B(net6014),
    .D(_00605_),
    .Q(\inv_result[87] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _41330_ (.RESET_B(net6014),
    .D(_00606_),
    .Q(\inv_result[88] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_1 _41331_ (.RESET_B(net6015),
    .D(_00607_),
    .Q(\inv_result[89] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _41332_ (.RESET_B(net6014),
    .D(_00608_),
    .Q(\inv_result[90] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _41333_ (.RESET_B(net6013),
    .D(_00609_),
    .Q(\inv_result[91] ),
    .CLK(clknet_leaf_158_clk));
 sg13g2_dfrbpq_1 _41334_ (.RESET_B(net6013),
    .D(_00610_),
    .Q(\inv_result[92] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _41335_ (.RESET_B(net6027),
    .D(_00611_),
    .Q(\inv_result[93] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _41336_ (.RESET_B(net6028),
    .D(_00612_),
    .Q(\inv_result[94] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _41337_ (.RESET_B(net6013),
    .D(_00613_),
    .Q(\inv_result[95] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _41338_ (.RESET_B(net6023),
    .D(_00614_),
    .Q(\inv_result[96] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _41339_ (.RESET_B(net6024),
    .D(_00615_),
    .Q(\inv_result[97] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _41340_ (.RESET_B(net6025),
    .D(_00616_),
    .Q(\inv_result[98] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _41341_ (.RESET_B(net6023),
    .D(_00617_),
    .Q(\inv_result[99] ),
    .CLK(clknet_leaf_162_clk));
 sg13g2_dfrbpq_1 _41342_ (.RESET_B(net6023),
    .D(net1140),
    .Q(\inv_result[100] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _41343_ (.RESET_B(net6021),
    .D(net1301),
    .Q(\inv_result[101] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _41344_ (.RESET_B(net6024),
    .D(_00620_),
    .Q(\inv_result[102] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _41345_ (.RESET_B(net6020),
    .D(_00621_),
    .Q(\inv_result[103] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _41346_ (.RESET_B(net6021),
    .D(_00622_),
    .Q(\inv_result[104] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _41347_ (.RESET_B(net6020),
    .D(_00623_),
    .Q(\inv_result[105] ),
    .CLK(clknet_leaf_161_clk));
 sg13g2_dfrbpq_1 _41348_ (.RESET_B(net6020),
    .D(_00624_),
    .Q(\inv_result[106] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _41349_ (.RESET_B(net6018),
    .D(_00625_),
    .Q(\inv_result[107] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _41350_ (.RESET_B(net6019),
    .D(_00626_),
    .Q(\inv_result[108] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _41351_ (.RESET_B(net6017),
    .D(_00627_),
    .Q(\inv_result[109] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _41352_ (.RESET_B(net6017),
    .D(_00628_),
    .Q(\inv_result[110] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _41353_ (.RESET_B(net6008),
    .D(_00629_),
    .Q(\inv_result[111] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_1 _41354_ (.RESET_B(net6007),
    .D(_00630_),
    .Q(\inv_result[112] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _41355_ (.RESET_B(net6006),
    .D(_00631_),
    .Q(\inv_result[113] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _41356_ (.RESET_B(net6006),
    .D(_00632_),
    .Q(\inv_result[114] ),
    .CLK(clknet_leaf_150_clk));
 sg13g2_dfrbpq_1 _41357_ (.RESET_B(net6005),
    .D(_00633_),
    .Q(\inv_result[115] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _41358_ (.RESET_B(net6005),
    .D(_00634_),
    .Q(\inv_result[116] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _41359_ (.RESET_B(net6005),
    .D(_00635_),
    .Q(\inv_result[117] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _41360_ (.RESET_B(net6001),
    .D(_00636_),
    .Q(\inv_result[118] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _41361_ (.RESET_B(net6002),
    .D(_00637_),
    .Q(\inv_result[119] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _41362_ (.RESET_B(net6000),
    .D(_00638_),
    .Q(\inv_result[120] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _41363_ (.RESET_B(net6000),
    .D(_00639_),
    .Q(\inv_result[121] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _41364_ (.RESET_B(net5997),
    .D(_00640_),
    .Q(\inv_result[122] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _41365_ (.RESET_B(net6001),
    .D(net1625),
    .Q(\inv_result[123] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _41366_ (.RESET_B(net5996),
    .D(net1199),
    .Q(\inv_result[124] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _41367_ (.RESET_B(net6000),
    .D(_00643_),
    .Q(\inv_result[125] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_1 _41368_ (.RESET_B(net5996),
    .D(_00644_),
    .Q(\inv_result[126] ),
    .CLK(clknet_leaf_166_clk));
 sg13g2_dfrbpq_1 _41369_ (.RESET_B(net5996),
    .D(_00645_),
    .Q(\inv_result[127] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _41370_ (.RESET_B(net5998),
    .D(_00646_),
    .Q(\inv_result[128] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _41371_ (.RESET_B(net5998),
    .D(net1383),
    .Q(\inv_result[129] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _41372_ (.RESET_B(net5985),
    .D(_00648_),
    .Q(\inv_result[130] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _41373_ (.RESET_B(net5985),
    .D(_00649_),
    .Q(\inv_result[131] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _41374_ (.RESET_B(net5998),
    .D(_00650_),
    .Q(\inv_result[132] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_2 _41375_ (.RESET_B(net5985),
    .D(_00651_),
    .Q(\inv_result[133] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_1 _41376_ (.RESET_B(net5991),
    .D(_00652_),
    .Q(\inv_result[134] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _41377_ (.RESET_B(net5991),
    .D(_00653_),
    .Q(\inv_result[135] ),
    .CLK(clknet_leaf_176_clk));
 sg13g2_dfrbpq_1 _41378_ (.RESET_B(net5984),
    .D(_00654_),
    .Q(\inv_result[136] ),
    .CLK(clknet_leaf_177_clk));
 sg13g2_dfrbpq_1 _41379_ (.RESET_B(net5984),
    .D(_00655_),
    .Q(\inv_result[137] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _41380_ (.RESET_B(net5991),
    .D(_00656_),
    .Q(\inv_result[138] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _41381_ (.RESET_B(net5993),
    .D(_00657_),
    .Q(\inv_result[139] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _41382_ (.RESET_B(net5990),
    .D(_00658_),
    .Q(\inv_result[140] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _41383_ (.RESET_B(net5987),
    .D(_00659_),
    .Q(\inv_result[141] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _41384_ (.RESET_B(net5987),
    .D(_00660_),
    .Q(\inv_result[142] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _41385_ (.RESET_B(net5987),
    .D(_00661_),
    .Q(\inv_result[143] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _41386_ (.RESET_B(net5989),
    .D(_00662_),
    .Q(\inv_result[144] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _41387_ (.RESET_B(net5982),
    .D(_00663_),
    .Q(\inv_result[145] ),
    .CLK(clknet_leaf_178_clk));
 sg13g2_dfrbpq_1 _41388_ (.RESET_B(net5978),
    .D(_00664_),
    .Q(\inv_result[146] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _41389_ (.RESET_B(net5978),
    .D(_00665_),
    .Q(\inv_result[147] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _41390_ (.RESET_B(net5976),
    .D(_00666_),
    .Q(\inv_result[148] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _41391_ (.RESET_B(net5976),
    .D(_00667_),
    .Q(\inv_result[149] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _41392_ (.RESET_B(net5978),
    .D(_00668_),
    .Q(\inv_result[150] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _41393_ (.RESET_B(net5978),
    .D(_00669_),
    .Q(\inv_result[151] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _41394_ (.RESET_B(net5977),
    .D(_00670_),
    .Q(\inv_result[152] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _41395_ (.RESET_B(net5976),
    .D(_00671_),
    .Q(\inv_result[153] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _41396_ (.RESET_B(net5975),
    .D(_00672_),
    .Q(\inv_result[154] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _41397_ (.RESET_B(net5976),
    .D(_00673_),
    .Q(\inv_result[155] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _41398_ (.RESET_B(net5976),
    .D(_00674_),
    .Q(\inv_result[156] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _41399_ (.RESET_B(net5976),
    .D(_00675_),
    .Q(\inv_result[157] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _41400_ (.RESET_B(net5976),
    .D(_00676_),
    .Q(\inv_result[158] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _41401_ (.RESET_B(net5972),
    .D(_00677_),
    .Q(\inv_result[159] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _41402_ (.RESET_B(net5970),
    .D(_00678_),
    .Q(\inv_result[160] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _41403_ (.RESET_B(net5973),
    .D(_00679_),
    .Q(\inv_result[161] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_1 _41404_ (.RESET_B(net5970),
    .D(_00680_),
    .Q(\inv_result[162] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _41405_ (.RESET_B(net5973),
    .D(_00681_),
    .Q(\inv_result[163] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _41406_ (.RESET_B(net5970),
    .D(_00682_),
    .Q(\inv_result[164] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _41407_ (.RESET_B(net5970),
    .D(_00683_),
    .Q(\inv_result[165] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _41408_ (.RESET_B(net5962),
    .D(_00684_),
    .Q(\inv_result[166] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _41409_ (.RESET_B(net5970),
    .D(_00685_),
    .Q(\inv_result[167] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _41410_ (.RESET_B(net5970),
    .D(_00686_),
    .Q(\inv_result[168] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _41411_ (.RESET_B(net5963),
    .D(_00687_),
    .Q(\inv_result[169] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _41412_ (.RESET_B(net5962),
    .D(_00688_),
    .Q(\inv_result[170] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _41413_ (.RESET_B(net5962),
    .D(_00689_),
    .Q(\inv_result[171] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _41414_ (.RESET_B(net5962),
    .D(_00690_),
    .Q(\inv_result[172] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _41415_ (.RESET_B(net5963),
    .D(_00691_),
    .Q(\inv_result[173] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _41416_ (.RESET_B(net5962),
    .D(_00692_),
    .Q(\inv_result[174] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _41417_ (.RESET_B(net5962),
    .D(_00693_),
    .Q(\inv_result[175] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _41418_ (.RESET_B(net5961),
    .D(_00694_),
    .Q(\inv_result[176] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _41419_ (.RESET_B(net5958),
    .D(_00695_),
    .Q(\inv_result[177] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _41420_ (.RESET_B(net5961),
    .D(_00696_),
    .Q(\inv_result[178] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _41421_ (.RESET_B(net5961),
    .D(_00697_),
    .Q(\inv_result[179] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _41422_ (.RESET_B(net5955),
    .D(_00698_),
    .Q(\inv_result[180] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _41423_ (.RESET_B(net5955),
    .D(_00699_),
    .Q(\inv_result[181] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _41424_ (.RESET_B(net5951),
    .D(net2423),
    .Q(\inv_result[182] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _41425_ (.RESET_B(net5955),
    .D(_00701_),
    .Q(\inv_result[183] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _41426_ (.RESET_B(net5955),
    .D(_00702_),
    .Q(\inv_result[184] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _41427_ (.RESET_B(net5954),
    .D(_00703_),
    .Q(\inv_result[185] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _41428_ (.RESET_B(net5955),
    .D(_00704_),
    .Q(\inv_result[186] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _41429_ (.RESET_B(net5954),
    .D(_00705_),
    .Q(\inv_result[187] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _41430_ (.RESET_B(net5954),
    .D(_00706_),
    .Q(\inv_result[188] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _41431_ (.RESET_B(net5948),
    .D(_00707_),
    .Q(\inv_result[189] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _41432_ (.RESET_B(net5954),
    .D(_00708_),
    .Q(\inv_result[190] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _41433_ (.RESET_B(net5948),
    .D(_00709_),
    .Q(\inv_result[191] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _41434_ (.RESET_B(net5942),
    .D(_00710_),
    .Q(\inv_result[192] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _41435_ (.RESET_B(net5942),
    .D(_00711_),
    .Q(\inv_result[193] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _41436_ (.RESET_B(net5954),
    .D(_00712_),
    .Q(\inv_result[194] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _41437_ (.RESET_B(net5942),
    .D(_00713_),
    .Q(\inv_result[195] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _41438_ (.RESET_B(net5942),
    .D(_00714_),
    .Q(\inv_result[196] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _41439_ (.RESET_B(net5942),
    .D(_00715_),
    .Q(\inv_result[197] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _41440_ (.RESET_B(net5933),
    .D(_00716_),
    .Q(\inv_result[198] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _41441_ (.RESET_B(net5940),
    .D(_00717_),
    .Q(\inv_result[199] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _41442_ (.RESET_B(net5933),
    .D(_00718_),
    .Q(\inv_result[200] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _41443_ (.RESET_B(net5940),
    .D(_00719_),
    .Q(\inv_result[201] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _41444_ (.RESET_B(net5940),
    .D(_00720_),
    .Q(\inv_result[202] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _41445_ (.RESET_B(net5940),
    .D(_00721_),
    .Q(\inv_result[203] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _41446_ (.RESET_B(net5940),
    .D(_00722_),
    .Q(\inv_result[204] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _41447_ (.RESET_B(net5933),
    .D(_00723_),
    .Q(\inv_result[205] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _41448_ (.RESET_B(net5939),
    .D(_00724_),
    .Q(\inv_result[206] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _41449_ (.RESET_B(net5939),
    .D(_00725_),
    .Q(\inv_result[207] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _41450_ (.RESET_B(net5925),
    .D(_00726_),
    .Q(\inv_result[208] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _41451_ (.RESET_B(net5913),
    .D(_00727_),
    .Q(\inv_result[209] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _41452_ (.RESET_B(net5925),
    .D(_00728_),
    .Q(\inv_result[210] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _41453_ (.RESET_B(net5936),
    .D(_00729_),
    .Q(\inv_result[211] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _41454_ (.RESET_B(net5924),
    .D(_00730_),
    .Q(\inv_result[212] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _41455_ (.RESET_B(net5925),
    .D(_00731_),
    .Q(\inv_result[213] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _41456_ (.RESET_B(net5925),
    .D(_00732_),
    .Q(\inv_result[214] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _41457_ (.RESET_B(net5924),
    .D(_00733_),
    .Q(\inv_result[215] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _41458_ (.RESET_B(net5925),
    .D(_00734_),
    .Q(\inv_result[216] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _41459_ (.RESET_B(net5922),
    .D(_00735_),
    .Q(\inv_result[217] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _41460_ (.RESET_B(net5922),
    .D(_00736_),
    .Q(\inv_result[218] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _41461_ (.RESET_B(net5922),
    .D(_00737_),
    .Q(\inv_result[219] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _41462_ (.RESET_B(net5922),
    .D(_00738_),
    .Q(\inv_result[220] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _41463_ (.RESET_B(net5922),
    .D(_00739_),
    .Q(\inv_result[221] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _41464_ (.RESET_B(net5920),
    .D(_00740_),
    .Q(\inv_result[222] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _41465_ (.RESET_B(net5922),
    .D(_00741_),
    .Q(\inv_result[223] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _41466_ (.RESET_B(net5920),
    .D(_00742_),
    .Q(\inv_result[224] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _41467_ (.RESET_B(net5920),
    .D(_00743_),
    .Q(\inv_result[225] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _41468_ (.RESET_B(net5916),
    .D(_00744_),
    .Q(\inv_result[226] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _41469_ (.RESET_B(net5917),
    .D(_00745_),
    .Q(\inv_result[227] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _41470_ (.RESET_B(net5916),
    .D(_00746_),
    .Q(\inv_result[228] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _41471_ (.RESET_B(net5916),
    .D(_00747_),
    .Q(\inv_result[229] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _41472_ (.RESET_B(net5916),
    .D(_00748_),
    .Q(\inv_result[230] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _41473_ (.RESET_B(net5916),
    .D(_00749_),
    .Q(\inv_result[231] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _41474_ (.RESET_B(net5885),
    .D(_00750_),
    .Q(\inv_result[232] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _41475_ (.RESET_B(net5885),
    .D(_00751_),
    .Q(\inv_result[233] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _41476_ (.RESET_B(net5885),
    .D(_00752_),
    .Q(\inv_result[234] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _41477_ (.RESET_B(net5900),
    .D(_00753_),
    .Q(\inv_result[235] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _41478_ (.RESET_B(net5900),
    .D(_00754_),
    .Q(\inv_result[236] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _41479_ (.RESET_B(net5890),
    .D(_00755_),
    .Q(\inv_result[237] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _41480_ (.RESET_B(net5884),
    .D(_00756_),
    .Q(\inv_result[238] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _41481_ (.RESET_B(net5884),
    .D(_00757_),
    .Q(\inv_result[239] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _41482_ (.RESET_B(net5883),
    .D(_00758_),
    .Q(\inv_result[240] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _41483_ (.RESET_B(net5884),
    .D(_00759_),
    .Q(\inv_result[241] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _41484_ (.RESET_B(net5889),
    .D(_00760_),
    .Q(\inv_result[242] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _41485_ (.RESET_B(net5888),
    .D(_00761_),
    .Q(\inv_result[243] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _41486_ (.RESET_B(net5889),
    .D(_00762_),
    .Q(\inv_result[244] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _41487_ (.RESET_B(net5884),
    .D(_00763_),
    .Q(\inv_result[245] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _41488_ (.RESET_B(net5883),
    .D(_00764_),
    .Q(\inv_result[246] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _41489_ (.RESET_B(net5883),
    .D(_00765_),
    .Q(\inv_result[247] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _41490_ (.RESET_B(net5884),
    .D(_00766_),
    .Q(\inv_result[248] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _41491_ (.RESET_B(net5883),
    .D(_00767_),
    .Q(\inv_result[249] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _41492_ (.RESET_B(net5889),
    .D(_00768_),
    .Q(\inv_result[250] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _41493_ (.RESET_B(net5888),
    .D(_00769_),
    .Q(\inv_result[251] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _41494_ (.RESET_B(net5889),
    .D(_00770_),
    .Q(\inv_result[252] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _41495_ (.RESET_B(net5889),
    .D(net1610),
    .Q(\inv_result[253] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _41496_ (.RESET_B(net5883),
    .D(_00772_),
    .Q(\inv_result[254] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _41497_ (.RESET_B(net5883),
    .D(_00773_),
    .Q(\inv_result[255] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _41498_ (.RESET_B(net1061),
    .D(_00774_),
    .Q(\u_inv.d_next[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _41499_ (.RESET_B(net1059),
    .D(_00775_),
    .Q(\u_inv.d_next[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _41500_ (.RESET_B(net1058),
    .D(_00776_),
    .Q(\u_inv.d_next[2] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _41501_ (.RESET_B(net1056),
    .D(_00777_),
    .Q(\u_inv.d_next[3] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _41502_ (.RESET_B(net1055),
    .D(_00778_),
    .Q(\u_inv.d_next[4] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _41503_ (.RESET_B(net1053),
    .D(_00779_),
    .Q(\u_inv.d_next[5] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _41504_ (.RESET_B(net1052),
    .D(_00780_),
    .Q(\u_inv.d_next[6] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _41505_ (.RESET_B(net1050),
    .D(_00781_),
    .Q(\u_inv.d_next[7] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _41506_ (.RESET_B(net1049),
    .D(_00782_),
    .Q(\u_inv.d_next[8] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _41507_ (.RESET_B(net1047),
    .D(_00783_),
    .Q(\u_inv.d_next[9] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _41508_ (.RESET_B(net1046),
    .D(_00784_),
    .Q(\u_inv.d_next[10] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _41509_ (.RESET_B(net1044),
    .D(_00785_),
    .Q(\u_inv.d_next[11] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _41510_ (.RESET_B(net1043),
    .D(_00786_),
    .Q(\u_inv.d_next[12] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _41511_ (.RESET_B(net1041),
    .D(_00787_),
    .Q(\u_inv.d_next[13] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _41512_ (.RESET_B(net1040),
    .D(_00788_),
    .Q(\u_inv.d_next[14] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _41513_ (.RESET_B(net1038),
    .D(_00789_),
    .Q(\u_inv.d_next[15] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _41514_ (.RESET_B(net1037),
    .D(_00790_),
    .Q(\u_inv.d_next[16] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _41515_ (.RESET_B(net1035),
    .D(_00791_),
    .Q(\u_inv.d_next[17] ),
    .CLK(clknet_leaf_234_clk));
 sg13g2_dfrbpq_2 _41516_ (.RESET_B(net1034),
    .D(_00792_),
    .Q(\u_inv.d_next[18] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _41517_ (.RESET_B(net1032),
    .D(_00793_),
    .Q(\u_inv.d_next[19] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _41518_ (.RESET_B(net1031),
    .D(_00794_),
    .Q(\u_inv.d_next[20] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _41519_ (.RESET_B(net1029),
    .D(_00795_),
    .Q(\u_inv.d_next[21] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _41520_ (.RESET_B(net1028),
    .D(_00796_),
    .Q(\u_inv.d_next[22] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _41521_ (.RESET_B(net1026),
    .D(_00797_),
    .Q(\u_inv.d_next[23] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _41522_ (.RESET_B(net1025),
    .D(_00798_),
    .Q(\u_inv.d_next[24] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _41523_ (.RESET_B(net1023),
    .D(_00799_),
    .Q(\u_inv.d_next[25] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _41524_ (.RESET_B(net1022),
    .D(_00800_),
    .Q(\u_inv.d_next[26] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _41525_ (.RESET_B(net1020),
    .D(_00801_),
    .Q(\u_inv.d_next[27] ),
    .CLK(clknet_leaf_230_clk));
 sg13g2_dfrbpq_2 _41526_ (.RESET_B(net1019),
    .D(_00802_),
    .Q(\u_inv.d_next[28] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _41527_ (.RESET_B(net1017),
    .D(_00803_),
    .Q(\u_inv.d_next[29] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _41528_ (.RESET_B(net1016),
    .D(_00804_),
    .Q(\u_inv.d_next[30] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _41529_ (.RESET_B(net1014),
    .D(_00805_),
    .Q(\u_inv.d_next[31] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _41530_ (.RESET_B(net1013),
    .D(_00806_),
    .Q(\u_inv.d_next[32] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _41531_ (.RESET_B(net1011),
    .D(_00807_),
    .Q(\u_inv.d_next[33] ),
    .CLK(clknet_leaf_229_clk));
 sg13g2_dfrbpq_2 _41532_ (.RESET_B(net1010),
    .D(_00808_),
    .Q(\u_inv.d_next[34] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _41533_ (.RESET_B(net1008),
    .D(_00809_),
    .Q(\u_inv.d_next[35] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _41534_ (.RESET_B(net1007),
    .D(_00810_),
    .Q(\u_inv.d_next[36] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _41535_ (.RESET_B(net1005),
    .D(_00811_),
    .Q(\u_inv.d_next[37] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _41536_ (.RESET_B(net1004),
    .D(_00812_),
    .Q(\u_inv.d_next[38] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _41537_ (.RESET_B(net1002),
    .D(_00813_),
    .Q(\u_inv.d_next[39] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _41538_ (.RESET_B(net1001),
    .D(_00814_),
    .Q(\u_inv.d_next[40] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _41539_ (.RESET_B(net999),
    .D(_00815_),
    .Q(\u_inv.d_next[41] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _41540_ (.RESET_B(net998),
    .D(_00816_),
    .Q(\u_inv.d_next[42] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _41541_ (.RESET_B(net996),
    .D(_00817_),
    .Q(\u_inv.d_next[43] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _41542_ (.RESET_B(net995),
    .D(_00818_),
    .Q(\u_inv.d_next[44] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _41543_ (.RESET_B(net993),
    .D(_00819_),
    .Q(\u_inv.d_next[45] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _41544_ (.RESET_B(net992),
    .D(_00820_),
    .Q(\u_inv.d_next[46] ),
    .CLK(clknet_leaf_228_clk));
 sg13g2_dfrbpq_2 _41545_ (.RESET_B(net990),
    .D(_00821_),
    .Q(\u_inv.d_next[47] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _41546_ (.RESET_B(net989),
    .D(_00822_),
    .Q(\u_inv.d_next[48] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _41547_ (.RESET_B(net987),
    .D(_00823_),
    .Q(\u_inv.d_next[49] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _41548_ (.RESET_B(net986),
    .D(_00824_),
    .Q(\u_inv.d_next[50] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _41549_ (.RESET_B(net984),
    .D(_00825_),
    .Q(\u_inv.d_next[51] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _41550_ (.RESET_B(net983),
    .D(_00826_),
    .Q(\u_inv.d_next[52] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _41551_ (.RESET_B(net981),
    .D(_00827_),
    .Q(\u_inv.d_next[53] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _41552_ (.RESET_B(net980),
    .D(_00828_),
    .Q(\u_inv.d_next[54] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _41553_ (.RESET_B(net978),
    .D(_00829_),
    .Q(\u_inv.d_next[55] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _41554_ (.RESET_B(net977),
    .D(_00830_),
    .Q(\u_inv.d_next[56] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _41555_ (.RESET_B(net975),
    .D(_00831_),
    .Q(\u_inv.d_next[57] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _41556_ (.RESET_B(net974),
    .D(_00832_),
    .Q(\u_inv.d_next[58] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _41557_ (.RESET_B(net972),
    .D(_00833_),
    .Q(\u_inv.d_next[59] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _41558_ (.RESET_B(net971),
    .D(_00834_),
    .Q(\u_inv.d_next[60] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _41559_ (.RESET_B(net969),
    .D(_00835_),
    .Q(\u_inv.d_next[61] ),
    .CLK(clknet_leaf_209_clk));
 sg13g2_dfrbpq_2 _41560_ (.RESET_B(net968),
    .D(_00836_),
    .Q(\u_inv.d_next[62] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _41561_ (.RESET_B(net966),
    .D(_00837_),
    .Q(\u_inv.d_next[63] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _41562_ (.RESET_B(net965),
    .D(_00838_),
    .Q(\u_inv.d_next[64] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _41563_ (.RESET_B(net963),
    .D(_00839_),
    .Q(\u_inv.d_next[65] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _41564_ (.RESET_B(net962),
    .D(_00840_),
    .Q(\u_inv.d_next[66] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _41565_ (.RESET_B(net960),
    .D(_00841_),
    .Q(\u_inv.d_next[67] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _41566_ (.RESET_B(net959),
    .D(_00842_),
    .Q(\u_inv.d_next[68] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _41567_ (.RESET_B(net957),
    .D(_00843_),
    .Q(\u_inv.d_next[69] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _41568_ (.RESET_B(net956),
    .D(_00844_),
    .Q(\u_inv.d_next[70] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _41569_ (.RESET_B(net954),
    .D(_00845_),
    .Q(\u_inv.d_next[71] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _41570_ (.RESET_B(net953),
    .D(_00846_),
    .Q(\u_inv.d_next[72] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_2 _41571_ (.RESET_B(net951),
    .D(_00847_),
    .Q(\u_inv.d_next[73] ),
    .CLK(clknet_leaf_204_clk));
 sg13g2_dfrbpq_1 _41572_ (.RESET_B(net950),
    .D(_00848_),
    .Q(\u_inv.d_next[74] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _41573_ (.RESET_B(net948),
    .D(_00849_),
    .Q(\u_inv.d_next[75] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _41574_ (.RESET_B(net947),
    .D(_00850_),
    .Q(\u_inv.d_next[76] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _41575_ (.RESET_B(net945),
    .D(_00851_),
    .Q(\u_inv.d_next[77] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _41576_ (.RESET_B(net944),
    .D(_00852_),
    .Q(\u_inv.d_next[78] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _41577_ (.RESET_B(net942),
    .D(_00853_),
    .Q(\u_inv.d_next[79] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _41578_ (.RESET_B(net941),
    .D(_00854_),
    .Q(\u_inv.d_next[80] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _41579_ (.RESET_B(net939),
    .D(_00855_),
    .Q(\u_inv.d_next[81] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _41580_ (.RESET_B(net938),
    .D(_00856_),
    .Q(\u_inv.d_next[82] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _41581_ (.RESET_B(net936),
    .D(_00857_),
    .Q(\u_inv.d_next[83] ),
    .CLK(clknet_leaf_203_clk));
 sg13g2_dfrbpq_2 _41582_ (.RESET_B(net935),
    .D(_00858_),
    .Q(\u_inv.d_next[84] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _41583_ (.RESET_B(net933),
    .D(_00859_),
    .Q(\u_inv.d_next[85] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _41584_ (.RESET_B(net932),
    .D(_00860_),
    .Q(\u_inv.d_next[86] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _41585_ (.RESET_B(net930),
    .D(_00861_),
    .Q(\u_inv.d_next[87] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _41586_ (.RESET_B(net929),
    .D(_00862_),
    .Q(\u_inv.d_next[88] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _41587_ (.RESET_B(net927),
    .D(_00863_),
    .Q(\u_inv.d_next[89] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _41588_ (.RESET_B(net926),
    .D(_00864_),
    .Q(\u_inv.d_next[90] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _41589_ (.RESET_B(net924),
    .D(_00865_),
    .Q(\u_inv.d_next[91] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _41590_ (.RESET_B(net923),
    .D(_00866_),
    .Q(\u_inv.d_next[92] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _41591_ (.RESET_B(net921),
    .D(_00867_),
    .Q(\u_inv.d_next[93] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _41592_ (.RESET_B(net920),
    .D(_00868_),
    .Q(\u_inv.d_next[94] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _41593_ (.RESET_B(net918),
    .D(_00869_),
    .Q(\u_inv.d_next[95] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _41594_ (.RESET_B(net917),
    .D(_00870_),
    .Q(\u_inv.d_next[96] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _41595_ (.RESET_B(net915),
    .D(_00871_),
    .Q(\u_inv.d_next[97] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _41596_ (.RESET_B(net914),
    .D(_00872_),
    .Q(\u_inv.d_next[98] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _41597_ (.RESET_B(net912),
    .D(_00873_),
    .Q(\u_inv.d_next[99] ),
    .CLK(clknet_leaf_196_clk));
 sg13g2_dfrbpq_2 _41598_ (.RESET_B(net911),
    .D(_00874_),
    .Q(\u_inv.d_next[100] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _41599_ (.RESET_B(net909),
    .D(_00875_),
    .Q(\u_inv.d_next[101] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _41600_ (.RESET_B(net908),
    .D(_00876_),
    .Q(\u_inv.d_next[102] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _41601_ (.RESET_B(net906),
    .D(_00877_),
    .Q(\u_inv.d_next[103] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _41602_ (.RESET_B(net905),
    .D(_00878_),
    .Q(\u_inv.d_next[104] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _41603_ (.RESET_B(net903),
    .D(_00879_),
    .Q(\u_inv.d_next[105] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _41604_ (.RESET_B(net902),
    .D(_00880_),
    .Q(\u_inv.d_next[106] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _41605_ (.RESET_B(net900),
    .D(_00881_),
    .Q(\u_inv.d_next[107] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _41606_ (.RESET_B(net899),
    .D(_00882_),
    .Q(\u_inv.d_next[108] ),
    .CLK(clknet_leaf_197_clk));
 sg13g2_dfrbpq_2 _41607_ (.RESET_B(net897),
    .D(_00883_),
    .Q(\u_inv.d_next[109] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _41608_ (.RESET_B(net896),
    .D(_00884_),
    .Q(\u_inv.d_next[110] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _41609_ (.RESET_B(net894),
    .D(_00885_),
    .Q(\u_inv.d_next[111] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _41610_ (.RESET_B(net893),
    .D(_00886_),
    .Q(\u_inv.d_next[112] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _41611_ (.RESET_B(net891),
    .D(_00887_),
    .Q(\u_inv.d_next[113] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _41612_ (.RESET_B(net890),
    .D(_00888_),
    .Q(\u_inv.d_next[114] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _41613_ (.RESET_B(net888),
    .D(_00889_),
    .Q(\u_inv.d_next[115] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _41614_ (.RESET_B(net887),
    .D(_00890_),
    .Q(\u_inv.d_next[116] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _41615_ (.RESET_B(net885),
    .D(_00891_),
    .Q(\u_inv.d_next[117] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _41616_ (.RESET_B(net884),
    .D(_00892_),
    .Q(\u_inv.d_next[118] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _41617_ (.RESET_B(net882),
    .D(_00893_),
    .Q(\u_inv.d_next[119] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _41618_ (.RESET_B(net881),
    .D(_00894_),
    .Q(\u_inv.d_next[120] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _41619_ (.RESET_B(net879),
    .D(_00895_),
    .Q(\u_inv.d_next[121] ),
    .CLK(clknet_leaf_198_clk));
 sg13g2_dfrbpq_2 _41620_ (.RESET_B(net878),
    .D(_00896_),
    .Q(\u_inv.d_next[122] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _41621_ (.RESET_B(net876),
    .D(_00897_),
    .Q(\u_inv.d_next[123] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _41622_ (.RESET_B(net875),
    .D(_00898_),
    .Q(\u_inv.d_next[124] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _41623_ (.RESET_B(net873),
    .D(_00899_),
    .Q(\u_inv.d_next[125] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _41624_ (.RESET_B(net872),
    .D(_00900_),
    .Q(\u_inv.d_next[126] ),
    .CLK(clknet_leaf_199_clk));
 sg13g2_dfrbpq_2 _41625_ (.RESET_B(net870),
    .D(_00901_),
    .Q(\u_inv.d_next[127] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _41626_ (.RESET_B(net869),
    .D(_00902_),
    .Q(\u_inv.d_next[128] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _41627_ (.RESET_B(net867),
    .D(_00903_),
    .Q(\u_inv.d_next[129] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _41628_ (.RESET_B(net866),
    .D(_00904_),
    .Q(\u_inv.d_next[130] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _41629_ (.RESET_B(net864),
    .D(_00905_),
    .Q(\u_inv.d_next[131] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _41630_ (.RESET_B(net863),
    .D(_00906_),
    .Q(\u_inv.d_next[132] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _41631_ (.RESET_B(net861),
    .D(_00907_),
    .Q(\u_inv.d_next[133] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _41632_ (.RESET_B(net860),
    .D(_00908_),
    .Q(\u_inv.d_next[134] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _41633_ (.RESET_B(net858),
    .D(_00909_),
    .Q(\u_inv.d_next[135] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _41634_ (.RESET_B(net857),
    .D(_00910_),
    .Q(\u_inv.d_next[136] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _41635_ (.RESET_B(net855),
    .D(_00911_),
    .Q(\u_inv.d_next[137] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _41636_ (.RESET_B(net854),
    .D(_00912_),
    .Q(\u_inv.d_next[138] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _41637_ (.RESET_B(net852),
    .D(_00913_),
    .Q(\u_inv.d_next[139] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _41638_ (.RESET_B(net851),
    .D(_00914_),
    .Q(\u_inv.d_next[140] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _41639_ (.RESET_B(net849),
    .D(_00915_),
    .Q(\u_inv.d_next[141] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _41640_ (.RESET_B(net848),
    .D(_00916_),
    .Q(\u_inv.d_next[142] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _41641_ (.RESET_B(net846),
    .D(_00917_),
    .Q(\u_inv.d_next[143] ),
    .CLK(clknet_leaf_215_clk));
 sg13g2_dfrbpq_2 _41642_ (.RESET_B(net845),
    .D(_00918_),
    .Q(\u_inv.d_next[144] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_1 _41643_ (.RESET_B(net843),
    .D(_00919_),
    .Q(\u_inv.d_next[145] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _41644_ (.RESET_B(net842),
    .D(_00920_),
    .Q(\u_inv.d_next[146] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _41645_ (.RESET_B(net840),
    .D(_00921_),
    .Q(\u_inv.d_next[147] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _41646_ (.RESET_B(net839),
    .D(_00922_),
    .Q(\u_inv.d_next[148] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _41647_ (.RESET_B(net837),
    .D(_00923_),
    .Q(\u_inv.d_next[149] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _41648_ (.RESET_B(net836),
    .D(_00924_),
    .Q(\u_inv.d_next[150] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _41649_ (.RESET_B(net834),
    .D(_00925_),
    .Q(\u_inv.d_next[151] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _41650_ (.RESET_B(net833),
    .D(_00926_),
    .Q(\u_inv.d_next[152] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _41651_ (.RESET_B(net831),
    .D(_00927_),
    .Q(\u_inv.d_next[153] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _41652_ (.RESET_B(net830),
    .D(_00928_),
    .Q(\u_inv.d_next[154] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _41653_ (.RESET_B(net828),
    .D(_00929_),
    .Q(\u_inv.d_next[155] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _41654_ (.RESET_B(net827),
    .D(_00930_),
    .Q(\u_inv.d_next[156] ),
    .CLK(clknet_leaf_216_clk));
 sg13g2_dfrbpq_2 _41655_ (.RESET_B(net825),
    .D(_00931_),
    .Q(\u_inv.d_next[157] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _41656_ (.RESET_B(net824),
    .D(_00932_),
    .Q(\u_inv.d_next[158] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _41657_ (.RESET_B(net822),
    .D(_00933_),
    .Q(\u_inv.d_next[159] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _41658_ (.RESET_B(net821),
    .D(_00934_),
    .Q(\u_inv.d_next[160] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _41659_ (.RESET_B(net819),
    .D(_00935_),
    .Q(\u_inv.d_next[161] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _41660_ (.RESET_B(net818),
    .D(_00936_),
    .Q(\u_inv.d_next[162] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _41661_ (.RESET_B(net816),
    .D(_00937_),
    .Q(\u_inv.d_next[163] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _41662_ (.RESET_B(net815),
    .D(_00938_),
    .Q(\u_inv.d_next[164] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _41663_ (.RESET_B(net813),
    .D(_00939_),
    .Q(\u_inv.d_next[165] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _41664_ (.RESET_B(net812),
    .D(_00940_),
    .Q(\u_inv.d_next[166] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _41665_ (.RESET_B(net810),
    .D(_00941_),
    .Q(\u_inv.d_next[167] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _41666_ (.RESET_B(net809),
    .D(_00942_),
    .Q(\u_inv.d_next[168] ),
    .CLK(clknet_leaf_210_clk));
 sg13g2_dfrbpq_2 _41667_ (.RESET_B(net807),
    .D(_00943_),
    .Q(\u_inv.d_next[169] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _41668_ (.RESET_B(net806),
    .D(_00944_),
    .Q(\u_inv.d_next[170] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _41669_ (.RESET_B(net804),
    .D(_00945_),
    .Q(\u_inv.d_next[171] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _41670_ (.RESET_B(net803),
    .D(_00946_),
    .Q(\u_inv.d_next[172] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _41671_ (.RESET_B(net801),
    .D(_00947_),
    .Q(\u_inv.d_next[173] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _41672_ (.RESET_B(net800),
    .D(_00948_),
    .Q(\u_inv.d_next[174] ),
    .CLK(clknet_leaf_227_clk));
 sg13g2_dfrbpq_2 _41673_ (.RESET_B(net798),
    .D(_00949_),
    .Q(\u_inv.d_next[175] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _41674_ (.RESET_B(net797),
    .D(_00950_),
    .Q(\u_inv.d_next[176] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _41675_ (.RESET_B(net795),
    .D(_00951_),
    .Q(\u_inv.d_next[177] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _41676_ (.RESET_B(net794),
    .D(_00952_),
    .Q(\u_inv.d_next[178] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _41677_ (.RESET_B(net792),
    .D(_00953_),
    .Q(\u_inv.d_next[179] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _41678_ (.RESET_B(net791),
    .D(_00954_),
    .Q(\u_inv.d_next[180] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _41679_ (.RESET_B(net789),
    .D(_00955_),
    .Q(\u_inv.d_next[181] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _41680_ (.RESET_B(net788),
    .D(_00956_),
    .Q(\u_inv.d_next[182] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _41681_ (.RESET_B(net786),
    .D(_00957_),
    .Q(\u_inv.d_next[183] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _41682_ (.RESET_B(net785),
    .D(_00958_),
    .Q(\u_inv.d_next[184] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _41683_ (.RESET_B(net783),
    .D(_00959_),
    .Q(\u_inv.d_next[185] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _41684_ (.RESET_B(net782),
    .D(_00960_),
    .Q(\u_inv.d_next[186] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _41685_ (.RESET_B(net780),
    .D(_00961_),
    .Q(\u_inv.d_next[187] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _41686_ (.RESET_B(net779),
    .D(_00962_),
    .Q(\u_inv.d_next[188] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _41687_ (.RESET_B(net777),
    .D(_00963_),
    .Q(\u_inv.d_next[189] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _41688_ (.RESET_B(net776),
    .D(_00964_),
    .Q(\u_inv.d_next[190] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _41689_ (.RESET_B(net774),
    .D(_00965_),
    .Q(\u_inv.d_next[191] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _41690_ (.RESET_B(net773),
    .D(_00966_),
    .Q(\u_inv.d_next[192] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _41691_ (.RESET_B(net771),
    .D(_00967_),
    .Q(\u_inv.d_next[193] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _41692_ (.RESET_B(net770),
    .D(_00968_),
    .Q(\u_inv.d_next[194] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _41693_ (.RESET_B(net768),
    .D(_00969_),
    .Q(\u_inv.d_next[195] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _41694_ (.RESET_B(net767),
    .D(_00970_),
    .Q(\u_inv.d_next[196] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _41695_ (.RESET_B(net765),
    .D(_00971_),
    .Q(\u_inv.d_next[197] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _41696_ (.RESET_B(net764),
    .D(_00972_),
    .Q(\u_inv.d_next[198] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _41697_ (.RESET_B(net762),
    .D(_00973_),
    .Q(\u_inv.d_next[199] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _41698_ (.RESET_B(net761),
    .D(_00974_),
    .Q(\u_inv.d_next[200] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _41699_ (.RESET_B(net759),
    .D(_00975_),
    .Q(\u_inv.d_next[201] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _41700_ (.RESET_B(net758),
    .D(_00976_),
    .Q(\u_inv.d_next[202] ),
    .CLK(clknet_leaf_223_clk));
 sg13g2_dfrbpq_2 _41701_ (.RESET_B(net756),
    .D(_00977_),
    .Q(\u_inv.d_next[203] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _41702_ (.RESET_B(net755),
    .D(_00978_),
    .Q(\u_inv.d_next[204] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _41703_ (.RESET_B(net753),
    .D(_00979_),
    .Q(\u_inv.d_next[205] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _41704_ (.RESET_B(net751),
    .D(_00980_),
    .Q(\u_inv.d_next[206] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _41705_ (.RESET_B(net749),
    .D(_00981_),
    .Q(\u_inv.d_next[207] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _41706_ (.RESET_B(net748),
    .D(_00982_),
    .Q(\u_inv.d_next[208] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _41707_ (.RESET_B(net746),
    .D(_00983_),
    .Q(\u_inv.d_next[209] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _41708_ (.RESET_B(net745),
    .D(_00984_),
    .Q(\u_inv.d_next[210] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _41709_ (.RESET_B(net743),
    .D(_00985_),
    .Q(\u_inv.d_next[211] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _41710_ (.RESET_B(net742),
    .D(_00986_),
    .Q(\u_inv.d_next[212] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _41711_ (.RESET_B(net740),
    .D(_00987_),
    .Q(\u_inv.d_next[213] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _41712_ (.RESET_B(net739),
    .D(_00988_),
    .Q(\u_inv.d_next[214] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _41713_ (.RESET_B(net737),
    .D(_00989_),
    .Q(\u_inv.d_next[215] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _41714_ (.RESET_B(net736),
    .D(_00990_),
    .Q(\u_inv.d_next[216] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _41715_ (.RESET_B(net734),
    .D(_00991_),
    .Q(\u_inv.d_next[217] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _41716_ (.RESET_B(net733),
    .D(_00992_),
    .Q(\u_inv.d_next[218] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _41717_ (.RESET_B(net731),
    .D(_00993_),
    .Q(\u_inv.d_next[219] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _41718_ (.RESET_B(net730),
    .D(_00994_),
    .Q(\u_inv.d_next[220] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _41719_ (.RESET_B(net728),
    .D(_00995_),
    .Q(\u_inv.d_next[221] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _41720_ (.RESET_B(net727),
    .D(_00996_),
    .Q(\u_inv.d_next[222] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _41721_ (.RESET_B(net725),
    .D(_00997_),
    .Q(\u_inv.d_next[223] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _41722_ (.RESET_B(net724),
    .D(_00998_),
    .Q(\u_inv.d_next[224] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _41723_ (.RESET_B(net722),
    .D(_00999_),
    .Q(\u_inv.d_next[225] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _41724_ (.RESET_B(net721),
    .D(_01000_),
    .Q(\u_inv.d_next[226] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _41725_ (.RESET_B(net719),
    .D(_01001_),
    .Q(\u_inv.d_next[227] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _41726_ (.RESET_B(net718),
    .D(_01002_),
    .Q(\u_inv.d_next[228] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _41727_ (.RESET_B(net716),
    .D(_01003_),
    .Q(\u_inv.d_next[229] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _41728_ (.RESET_B(net715),
    .D(_01004_),
    .Q(\u_inv.d_next[230] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _41729_ (.RESET_B(net713),
    .D(_01005_),
    .Q(\u_inv.d_next[231] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _41730_ (.RESET_B(net712),
    .D(_01006_),
    .Q(\u_inv.d_next[232] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _41731_ (.RESET_B(net710),
    .D(_01007_),
    .Q(\u_inv.d_next[233] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _41732_ (.RESET_B(net709),
    .D(_01008_),
    .Q(\u_inv.d_next[234] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _41733_ (.RESET_B(net707),
    .D(_01009_),
    .Q(\u_inv.d_next[235] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _41734_ (.RESET_B(net706),
    .D(_01010_),
    .Q(\u_inv.d_next[236] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _41735_ (.RESET_B(net704),
    .D(_01011_),
    .Q(\u_inv.d_next[237] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _41736_ (.RESET_B(net703),
    .D(_01012_),
    .Q(\u_inv.d_next[238] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _41737_ (.RESET_B(net701),
    .D(_01013_),
    .Q(\u_inv.d_next[239] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _41738_ (.RESET_B(net700),
    .D(_01014_),
    .Q(\u_inv.d_next[240] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _41739_ (.RESET_B(net698),
    .D(_01015_),
    .Q(\u_inv.d_next[241] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _41740_ (.RESET_B(net697),
    .D(_01016_),
    .Q(\u_inv.d_next[242] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _41741_ (.RESET_B(net695),
    .D(_01017_),
    .Q(\u_inv.d_next[243] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _41742_ (.RESET_B(net694),
    .D(_01018_),
    .Q(\u_inv.d_next[244] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _41743_ (.RESET_B(net692),
    .D(_01019_),
    .Q(\u_inv.d_next[245] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _41744_ (.RESET_B(net691),
    .D(_01020_),
    .Q(\u_inv.d_next[246] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _41745_ (.RESET_B(net689),
    .D(_01021_),
    .Q(\u_inv.d_next[247] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _41746_ (.RESET_B(net688),
    .D(_01022_),
    .Q(\u_inv.d_next[248] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _41747_ (.RESET_B(net686),
    .D(_01023_),
    .Q(\u_inv.d_next[249] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _41748_ (.RESET_B(net685),
    .D(_01024_),
    .Q(\u_inv.d_next[250] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _41749_ (.RESET_B(net683),
    .D(_01025_),
    .Q(\u_inv.d_next[251] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _41750_ (.RESET_B(net682),
    .D(_01026_),
    .Q(\u_inv.d_next[252] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _41751_ (.RESET_B(net680),
    .D(_01027_),
    .Q(\u_inv.d_next[253] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _41752_ (.RESET_B(net679),
    .D(_01028_),
    .Q(\u_inv.d_next[254] ),
    .CLK(clknet_leaf_235_clk));
 sg13g2_dfrbpq_2 _41753_ (.RESET_B(net677),
    .D(_01029_),
    .Q(\u_inv.d_next[255] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _41754_ (.RESET_B(net752),
    .D(_01030_),
    .Q(\u_inv.d_next[256] ),
    .CLK(clknet_leaf_233_clk));
 sg13g2_dfrbpq_2 _41755_ (.RESET_B(net5904),
    .D(net3333),
    .Q(inv_done),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _41756_ (.RESET_B(net675),
    .D(net1385),
    .Q(\u_inv.d_reg[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _41757_ (.RESET_B(net674),
    .D(net2399),
    .Q(\u_inv.d_reg[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _41758_ (.RESET_B(net672),
    .D(net2431),
    .Q(\u_inv.d_reg[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _41759_ (.RESET_B(net671),
    .D(net2564),
    .Q(\u_inv.d_reg[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _41760_ (.RESET_B(net669),
    .D(_01035_),
    .Q(\u_inv.d_reg[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _41761_ (.RESET_B(net668),
    .D(net2863),
    .Q(\u_inv.d_reg[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _41762_ (.RESET_B(net666),
    .D(net2544),
    .Q(\u_inv.d_reg[6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _41763_ (.RESET_B(net665),
    .D(net2427),
    .Q(\u_inv.d_reg[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _41764_ (.RESET_B(net663),
    .D(net2605),
    .Q(\u_inv.d_reg[8] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _41765_ (.RESET_B(net662),
    .D(net2504),
    .Q(\u_inv.d_reg[9] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _41766_ (.RESET_B(net660),
    .D(net3094),
    .Q(\u_inv.d_reg[10] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _41767_ (.RESET_B(net659),
    .D(net3216),
    .Q(\u_inv.d_reg[11] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _41768_ (.RESET_B(net657),
    .D(net2524),
    .Q(\u_inv.d_reg[12] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _41769_ (.RESET_B(net656),
    .D(net2509),
    .Q(\u_inv.d_reg[13] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _41770_ (.RESET_B(net654),
    .D(net2442),
    .Q(\u_inv.d_reg[14] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _41771_ (.RESET_B(net653),
    .D(net2620),
    .Q(\u_inv.d_reg[15] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_1 _41772_ (.RESET_B(net651),
    .D(net2935),
    .Q(\u_inv.d_reg[16] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _41773_ (.RESET_B(net650),
    .D(net2788),
    .Q(\u_inv.d_reg[17] ),
    .CLK(clknet_leaf_232_clk));
 sg13g2_dfrbpq_2 _41774_ (.RESET_B(net648),
    .D(net2705),
    .Q(\u_inv.d_reg[18] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _41775_ (.RESET_B(net647),
    .D(net2905),
    .Q(\u_inv.d_reg[19] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _41776_ (.RESET_B(net645),
    .D(net2597),
    .Q(\u_inv.d_reg[20] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _41777_ (.RESET_B(net644),
    .D(net2300),
    .Q(\u_inv.d_reg[21] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _41778_ (.RESET_B(net642),
    .D(_01053_),
    .Q(\u_inv.d_reg[22] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _41779_ (.RESET_B(net641),
    .D(net3056),
    .Q(\u_inv.d_reg[23] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _41780_ (.RESET_B(net639),
    .D(net2474),
    .Q(\u_inv.d_reg[24] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _41781_ (.RESET_B(net638),
    .D(net1613),
    .Q(\u_inv.d_reg[25] ),
    .CLK(clknet_leaf_231_clk));
 sg13g2_dfrbpq_2 _41782_ (.RESET_B(net636),
    .D(net2841),
    .Q(\u_inv.d_reg[26] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _41783_ (.RESET_B(net635),
    .D(net2971),
    .Q(\u_inv.d_reg[27] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _41784_ (.RESET_B(net633),
    .D(net1598),
    .Q(\u_inv.d_reg[28] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _41785_ (.RESET_B(net632),
    .D(net2274),
    .Q(\u_inv.d_reg[29] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _41786_ (.RESET_B(net630),
    .D(_01061_),
    .Q(\u_inv.d_reg[30] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _41787_ (.RESET_B(net629),
    .D(net2131),
    .Q(\u_inv.d_reg[31] ),
    .CLK(clknet_leaf_224_clk));
 sg13g2_dfrbpq_2 _41788_ (.RESET_B(net627),
    .D(net2690),
    .Q(\u_inv.d_reg[32] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _41789_ (.RESET_B(net626),
    .D(net2985),
    .Q(\u_inv.d_reg[33] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _41790_ (.RESET_B(net624),
    .D(net2589),
    .Q(\u_inv.d_reg[34] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _41791_ (.RESET_B(net623),
    .D(net2582),
    .Q(\u_inv.d_reg[35] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _41792_ (.RESET_B(net621),
    .D(net3218),
    .Q(\u_inv.d_reg[36] ),
    .CLK(clknet_leaf_222_clk));
 sg13g2_dfrbpq_2 _41793_ (.RESET_B(net620),
    .D(net2865),
    .Q(\u_inv.d_reg[37] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _41794_ (.RESET_B(net618),
    .D(net2269),
    .Q(\u_inv.d_reg[38] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _41795_ (.RESET_B(net617),
    .D(net2262),
    .Q(\u_inv.d_reg[39] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _41796_ (.RESET_B(net615),
    .D(net2886),
    .Q(\u_inv.d_reg[40] ),
    .CLK(clknet_leaf_225_clk));
 sg13g2_dfrbpq_2 _41797_ (.RESET_B(net614),
    .D(net2416),
    .Q(\u_inv.d_reg[41] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _41798_ (.RESET_B(net612),
    .D(net2344),
    .Q(\u_inv.d_reg[42] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _41799_ (.RESET_B(net611),
    .D(net2214),
    .Q(\u_inv.d_reg[43] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _41800_ (.RESET_B(net609),
    .D(net2408),
    .Q(\u_inv.d_reg[44] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _41801_ (.RESET_B(net608),
    .D(net2105),
    .Q(\u_inv.d_reg[45] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _41802_ (.RESET_B(net606),
    .D(net2326),
    .Q(\u_inv.d_reg[46] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _41803_ (.RESET_B(net605),
    .D(net2480),
    .Q(\u_inv.d_reg[47] ),
    .CLK(clknet_leaf_226_clk));
 sg13g2_dfrbpq_2 _41804_ (.RESET_B(net603),
    .D(net2882),
    .Q(\u_inv.d_reg[48] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _41805_ (.RESET_B(net602),
    .D(net2927),
    .Q(\u_inv.d_reg[49] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _41806_ (.RESET_B(net600),
    .D(net3305),
    .Q(\u_inv.d_reg[50] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _41807_ (.RESET_B(net599),
    .D(net2646),
    .Q(\u_inv.d_reg[51] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _41808_ (.RESET_B(net597),
    .D(net2741),
    .Q(\u_inv.d_reg[52] ),
    .CLK(clknet_leaf_214_clk));
 sg13g2_dfrbpq_2 _41809_ (.RESET_B(net596),
    .D(net2439),
    .Q(\u_inv.d_reg[53] ),
    .CLK(clknet_leaf_208_clk));
 sg13g2_dfrbpq_2 _41810_ (.RESET_B(net594),
    .D(net1727),
    .Q(\u_inv.d_reg[54] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _41811_ (.RESET_B(net593),
    .D(net2591),
    .Q(\u_inv.d_reg[55] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _41812_ (.RESET_B(net591),
    .D(net2178),
    .Q(\u_inv.d_reg[56] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _41813_ (.RESET_B(net590),
    .D(net2625),
    .Q(\u_inv.d_reg[57] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _41814_ (.RESET_B(net588),
    .D(net2607),
    .Q(\u_inv.d_reg[58] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _41815_ (.RESET_B(net587),
    .D(net2118),
    .Q(\u_inv.d_reg[59] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _41816_ (.RESET_B(net585),
    .D(net2348),
    .Q(\u_inv.d_reg[60] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _41817_ (.RESET_B(net584),
    .D(net2601),
    .Q(\u_inv.d_reg[61] ),
    .CLK(clknet_leaf_207_clk));
 sg13g2_dfrbpq_2 _41818_ (.RESET_B(net582),
    .D(net1583),
    .Q(\u_inv.d_reg[62] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _41819_ (.RESET_B(net581),
    .D(net2679),
    .Q(\u_inv.d_reg[63] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _41820_ (.RESET_B(net579),
    .D(net2642),
    .Q(\u_inv.d_reg[64] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _41821_ (.RESET_B(net578),
    .D(net2335),
    .Q(\u_inv.d_reg[65] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _41822_ (.RESET_B(net576),
    .D(net1261),
    .Q(\u_inv.d_reg[66] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _41823_ (.RESET_B(net575),
    .D(net2880),
    .Q(\u_inv.d_reg[67] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _41824_ (.RESET_B(net573),
    .D(net2872),
    .Q(\u_inv.d_reg[68] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _41825_ (.RESET_B(net572),
    .D(net2953),
    .Q(\u_inv.d_reg[69] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _41826_ (.RESET_B(net570),
    .D(net1407),
    .Q(\u_inv.d_reg[70] ),
    .CLK(clknet_leaf_206_clk));
 sg13g2_dfrbpq_2 _41827_ (.RESET_B(net569),
    .D(net2537),
    .Q(\u_inv.d_reg[71] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _41828_ (.RESET_B(net567),
    .D(net3419),
    .Q(\u_inv.d_reg[72] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _41829_ (.RESET_B(net566),
    .D(net2964),
    .Q(\u_inv.d_reg[73] ),
    .CLK(clknet_leaf_205_clk));
 sg13g2_dfrbpq_2 _41830_ (.RESET_B(net564),
    .D(net1360),
    .Q(\u_inv.d_reg[74] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _41831_ (.RESET_B(net563),
    .D(net1955),
    .Q(\u_inv.d_reg[75] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _41832_ (.RESET_B(net561),
    .D(net2975),
    .Q(\u_inv.d_reg[76] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_1 _41833_ (.RESET_B(net560),
    .D(net3088),
    .Q(\u_inv.d_reg[77] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _41834_ (.RESET_B(net558),
    .D(net2307),
    .Q(\u_inv.d_reg[78] ),
    .CLK(clknet_leaf_202_clk));
 sg13g2_dfrbpq_2 _41835_ (.RESET_B(net557),
    .D(net3028),
    .Q(\u_inv.d_reg[79] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _41836_ (.RESET_B(net555),
    .D(net2850),
    .Q(\u_inv.d_reg[80] ),
    .CLK(clknet_leaf_200_clk));
 sg13g2_dfrbpq_2 _41837_ (.RESET_B(net554),
    .D(net2929),
    .Q(\u_inv.d_reg[81] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _41838_ (.RESET_B(net552),
    .D(net2449),
    .Q(\u_inv.d_reg[82] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _41839_ (.RESET_B(net551),
    .D(net2637),
    .Q(\u_inv.d_reg[83] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _41840_ (.RESET_B(net549),
    .D(net2811),
    .Q(\u_inv.d_reg[84] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _41841_ (.RESET_B(net548),
    .D(net2469),
    .Q(\u_inv.d_reg[85] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _41842_ (.RESET_B(net546),
    .D(net2277),
    .Q(\u_inv.d_reg[86] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _41843_ (.RESET_B(net545),
    .D(net1525),
    .Q(\u_inv.d_reg[87] ),
    .CLK(clknet_leaf_201_clk));
 sg13g2_dfrbpq_2 _41844_ (.RESET_B(net543),
    .D(net3271),
    .Q(\u_inv.d_reg[88] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _41845_ (.RESET_B(net542),
    .D(net3048),
    .Q(\u_inv.d_reg[89] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _41846_ (.RESET_B(net540),
    .D(_01121_),
    .Q(\u_inv.d_reg[90] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _41847_ (.RESET_B(net539),
    .D(net2668),
    .Q(\u_inv.d_reg[91] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _41848_ (.RESET_B(net537),
    .D(net2389),
    .Q(\u_inv.d_reg[92] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _41849_ (.RESET_B(net536),
    .D(net3316),
    .Q(\u_inv.d_reg[93] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _41850_ (.RESET_B(net534),
    .D(net2627),
    .Q(\u_inv.d_reg[94] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _41851_ (.RESET_B(net533),
    .D(net2945),
    .Q(\u_inv.d_reg[95] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_2 _41852_ (.RESET_B(net531),
    .D(net3045),
    .Q(\u_inv.d_reg[96] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _41853_ (.RESET_B(net530),
    .D(net3105),
    .Q(\u_inv.d_reg[97] ),
    .CLK(clknet_leaf_195_clk));
 sg13g2_dfrbpq_1 _41854_ (.RESET_B(net528),
    .D(net2186),
    .Q(\u_inv.d_reg[98] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _41855_ (.RESET_B(net527),
    .D(net2421),
    .Q(\u_inv.d_reg[99] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _41856_ (.RESET_B(net525),
    .D(net2338),
    .Q(\u_inv.d_reg[100] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _41857_ (.RESET_B(net524),
    .D(net2613),
    .Q(\u_inv.d_reg[101] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _41858_ (.RESET_B(net522),
    .D(net2328),
    .Q(\u_inv.d_reg[102] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _41859_ (.RESET_B(net521),
    .D(net1641),
    .Q(\u_inv.d_reg[103] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _41860_ (.RESET_B(net519),
    .D(net2322),
    .Q(\u_inv.d_reg[104] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _41861_ (.RESET_B(net518),
    .D(net2515),
    .Q(\u_inv.d_reg[105] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _41862_ (.RESET_B(net516),
    .D(net3098),
    .Q(\u_inv.d_reg[106] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _41863_ (.RESET_B(net515),
    .D(net3232),
    .Q(\u_inv.d_reg[107] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _41864_ (.RESET_B(net513),
    .D(net2517),
    .Q(\u_inv.d_reg[108] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _41865_ (.RESET_B(net512),
    .D(net1422),
    .Q(\u_inv.d_reg[109] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _41866_ (.RESET_B(net510),
    .D(net1535),
    .Q(\u_inv.d_reg[110] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _41867_ (.RESET_B(net509),
    .D(net2920),
    .Q(\u_inv.d_reg[111] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _41868_ (.RESET_B(net507),
    .D(_01143_),
    .Q(\u_inv.d_reg[112] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_2 _41869_ (.RESET_B(net506),
    .D(net2570),
    .Q(\u_inv.d_reg[113] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _41870_ (.RESET_B(net504),
    .D(net2373),
    .Q(\u_inv.d_reg[114] ),
    .CLK(clknet_leaf_191_clk));
 sg13g2_dfrbpq_2 _41871_ (.RESET_B(net503),
    .D(net2371),
    .Q(\u_inv.d_reg[115] ),
    .CLK(clknet_leaf_192_clk));
 sg13g2_dfrbpq_2 _41872_ (.RESET_B(net501),
    .D(net2907),
    .Q(\u_inv.d_reg[116] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _41873_ (.RESET_B(net500),
    .D(net3067),
    .Q(\u_inv.d_reg[117] ),
    .CLK(clknet_leaf_165_clk));
 sg13g2_dfrbpq_2 _41874_ (.RESET_B(net498),
    .D(net2639),
    .Q(\u_inv.d_reg[118] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _41875_ (.RESET_B(net497),
    .D(net2884),
    .Q(\u_inv.d_reg[119] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _41876_ (.RESET_B(net495),
    .D(net3069),
    .Q(\u_inv.d_reg[120] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _41877_ (.RESET_B(net494),
    .D(net3288),
    .Q(\u_inv.d_reg[121] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _41878_ (.RESET_B(net492),
    .D(_01153_),
    .Q(\u_inv.d_reg[122] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _41879_ (.RESET_B(net491),
    .D(net2622),
    .Q(\u_inv.d_reg[123] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _41880_ (.RESET_B(net489),
    .D(_01155_),
    .Q(\u_inv.d_reg[124] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _41881_ (.RESET_B(net488),
    .D(net3223),
    .Q(\u_inv.d_reg[125] ),
    .CLK(clknet_leaf_190_clk));
 sg13g2_dfrbpq_2 _41882_ (.RESET_B(net486),
    .D(net2444),
    .Q(\u_inv.d_reg[126] ),
    .CLK(clknet_leaf_189_clk));
 sg13g2_dfrbpq_2 _41883_ (.RESET_B(net485),
    .D(net2093),
    .Q(\u_inv.d_reg[127] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _41884_ (.RESET_B(net483),
    .D(net2977),
    .Q(\u_inv.d_reg[128] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _41885_ (.RESET_B(net482),
    .D(net2611),
    .Q(\u_inv.d_reg[129] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _41886_ (.RESET_B(net480),
    .D(net2318),
    .Q(\u_inv.d_reg[130] ),
    .CLK(clknet_leaf_188_clk));
 sg13g2_dfrbpq_2 _41887_ (.RESET_B(net479),
    .D(net2694),
    .Q(\u_inv.d_reg[131] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _41888_ (.RESET_B(net477),
    .D(_01163_),
    .Q(\u_inv.d_reg[132] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _41889_ (.RESET_B(net476),
    .D(net3075),
    .Q(\u_inv.d_reg[133] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _41890_ (.RESET_B(net474),
    .D(_01165_),
    .Q(\u_inv.d_reg[134] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _41891_ (.RESET_B(net473),
    .D(net2997),
    .Q(\u_inv.d_reg[135] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _41892_ (.RESET_B(net471),
    .D(net2146),
    .Q(\u_inv.d_reg[136] ),
    .CLK(clknet_leaf_187_clk));
 sg13g2_dfrbpq_2 _41893_ (.RESET_B(net470),
    .D(net3236),
    .Q(\u_inv.d_reg[137] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _41894_ (.RESET_B(net468),
    .D(_01169_),
    .Q(\u_inv.d_reg[138] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _41895_ (.RESET_B(net467),
    .D(net2815),
    .Q(\u_inv.d_reg[139] ),
    .CLK(clknet_leaf_186_clk));
 sg13g2_dfrbpq_2 _41896_ (.RESET_B(net465),
    .D(net2558),
    .Q(\u_inv.d_reg[140] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _41897_ (.RESET_B(net464),
    .D(net2520),
    .Q(\u_inv.d_reg[141] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _41898_ (.RESET_B(net462),
    .D(net2553),
    .Q(\u_inv.d_reg[142] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _41899_ (.RESET_B(net461),
    .D(net2250),
    .Q(\u_inv.d_reg[143] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _41900_ (.RESET_B(net459),
    .D(net2683),
    .Q(\u_inv.d_reg[144] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _41901_ (.RESET_B(net458),
    .D(net1223),
    .Q(\u_inv.d_reg[145] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _41902_ (.RESET_B(net456),
    .D(net2757),
    .Q(\u_inv.d_reg[146] ),
    .CLK(clknet_leaf_185_clk));
 sg13g2_dfrbpq_2 _41903_ (.RESET_B(net455),
    .D(_01178_),
    .Q(\u_inv.d_reg[147] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _41904_ (.RESET_B(net453),
    .D(net2943),
    .Q(\u_inv.d_reg[148] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _41905_ (.RESET_B(net452),
    .D(net2933),
    .Q(\u_inv.d_reg[149] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _41906_ (.RESET_B(net450),
    .D(net3004),
    .Q(\u_inv.d_reg[150] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _41907_ (.RESET_B(net449),
    .D(net3221),
    .Q(\u_inv.d_reg[151] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _41908_ (.RESET_B(net447),
    .D(net2382),
    .Q(\u_inv.d_reg[152] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _41909_ (.RESET_B(net446),
    .D(_01184_),
    .Q(\u_inv.d_reg[153] ),
    .CLK(clknet_leaf_184_clk));
 sg13g2_dfrbpq_2 _41910_ (.RESET_B(net444),
    .D(_01185_),
    .Q(\u_inv.d_reg[154] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _41911_ (.RESET_B(net443),
    .D(net2063),
    .Q(\u_inv.d_reg[155] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _41912_ (.RESET_B(net441),
    .D(_01187_),
    .Q(\u_inv.d_reg[156] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _41913_ (.RESET_B(net440),
    .D(_01188_),
    .Q(\u_inv.d_reg[157] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _41914_ (.RESET_B(net438),
    .D(net3255),
    .Q(\u_inv.d_reg[158] ),
    .CLK(clknet_leaf_183_clk));
 sg13g2_dfrbpq_2 _41915_ (.RESET_B(net437),
    .D(_01190_),
    .Q(\u_inv.d_reg[159] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _41916_ (.RESET_B(net435),
    .D(_01191_),
    .Q(\u_inv.d_reg[160] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _41917_ (.RESET_B(net434),
    .D(net2723),
    .Q(\u_inv.d_reg[161] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _41918_ (.RESET_B(net432),
    .D(net3083),
    .Q(\u_inv.d_reg[162] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _41919_ (.RESET_B(net430),
    .D(_01194_),
    .Q(\u_inv.d_reg[163] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_1 _41920_ (.RESET_B(net428),
    .D(net2726),
    .Q(\u_inv.d_reg[164] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _41921_ (.RESET_B(net426),
    .D(net3131),
    .Q(\u_inv.d_reg[165] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _41922_ (.RESET_B(net424),
    .D(net2876),
    .Q(\u_inv.d_reg[166] ),
    .CLK(clknet_leaf_218_clk));
 sg13g2_dfrbpq_2 _41923_ (.RESET_B(net422),
    .D(net2937),
    .Q(\u_inv.d_reg[167] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _41924_ (.RESET_B(net420),
    .D(net2562),
    .Q(\u_inv.d_reg[168] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _41925_ (.RESET_B(net418),
    .D(_01200_),
    .Q(\u_inv.d_reg[169] ),
    .CLK(clknet_leaf_211_clk));
 sg13g2_dfrbpq_2 _41926_ (.RESET_B(net416),
    .D(_01201_),
    .Q(\u_inv.d_reg[170] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _41927_ (.RESET_B(net414),
    .D(_01202_),
    .Q(\u_inv.d_reg[171] ),
    .CLK(clknet_leaf_212_clk));
 sg13g2_dfrbpq_2 _41928_ (.RESET_B(net412),
    .D(net2247),
    .Q(\u_inv.d_reg[172] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _41929_ (.RESET_B(net410),
    .D(_01204_),
    .Q(\u_inv.d_reg[173] ),
    .CLK(clknet_leaf_213_clk));
 sg13g2_dfrbpq_2 _41930_ (.RESET_B(net408),
    .D(net2708),
    .Q(\u_inv.d_reg[174] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _41931_ (.RESET_B(net406),
    .D(net1424),
    .Q(\u_inv.d_reg[175] ),
    .CLK(clknet_leaf_217_clk));
 sg13g2_dfrbpq_2 _41932_ (.RESET_B(net404),
    .D(_01207_),
    .Q(\u_inv.d_reg[176] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _41933_ (.RESET_B(net402),
    .D(net1983),
    .Q(\u_inv.d_reg[177] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _41934_ (.RESET_B(net400),
    .D(net2419),
    .Q(\u_inv.d_reg[178] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _41935_ (.RESET_B(net398),
    .D(_01210_),
    .Q(\u_inv.d_reg[179] ),
    .CLK(clknet_leaf_219_clk));
 sg13g2_dfrbpq_2 _41936_ (.RESET_B(net396),
    .D(net2837),
    .Q(\u_inv.d_reg[180] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _41937_ (.RESET_B(net394),
    .D(net2664),
    .Q(\u_inv.d_reg[181] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _41938_ (.RESET_B(net392),
    .D(_01213_),
    .Q(\u_inv.d_reg[182] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _41939_ (.RESET_B(net390),
    .D(_01214_),
    .Q(\u_inv.d_reg[183] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _41940_ (.RESET_B(net388),
    .D(net2910),
    .Q(\u_inv.d_reg[184] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _41941_ (.RESET_B(net386),
    .D(_01216_),
    .Q(\u_inv.d_reg[185] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _41942_ (.RESET_B(net384),
    .D(net2206),
    .Q(\u_inv.d_reg[186] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _41943_ (.RESET_B(net382),
    .D(net3077),
    .Q(\u_inv.d_reg[187] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _41944_ (.RESET_B(net380),
    .D(net2342),
    .Q(\u_inv.d_reg[188] ),
    .CLK(clknet_leaf_220_clk));
 sg13g2_dfrbpq_2 _41945_ (.RESET_B(net378),
    .D(net2022),
    .Q(\u_inv.d_reg[189] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _41946_ (.RESET_B(net376),
    .D(net2293),
    .Q(\u_inv.d_reg[190] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _41947_ (.RESET_B(net374),
    .D(net1344),
    .Q(\u_inv.d_reg[191] ),
    .CLK(clknet_leaf_221_clk));
 sg13g2_dfrbpq_2 _41948_ (.RESET_B(net372),
    .D(_01223_),
    .Q(\u_inv.d_reg[192] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _41949_ (.RESET_B(net370),
    .D(net2463),
    .Q(\u_inv.d_reg[193] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _41950_ (.RESET_B(net368),
    .D(net2280),
    .Q(\u_inv.d_reg[194] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _41951_ (.RESET_B(net366),
    .D(_01226_),
    .Q(\u_inv.d_reg[195] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _41952_ (.RESET_B(net364),
    .D(net2239),
    .Q(\u_inv.d_reg[196] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _41953_ (.RESET_B(net362),
    .D(net2258),
    .Q(\u_inv.d_reg[197] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _41954_ (.RESET_B(net360),
    .D(_01229_),
    .Q(\u_inv.d_reg[198] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _41955_ (.RESET_B(net358),
    .D(_01230_),
    .Q(\u_inv.d_reg[199] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _41956_ (.RESET_B(net356),
    .D(_01231_),
    .Q(\u_inv.d_reg[200] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _41957_ (.RESET_B(net354),
    .D(net1712),
    .Q(\u_inv.d_reg[201] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _41958_ (.RESET_B(net352),
    .D(_01233_),
    .Q(\u_inv.d_reg[202] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _41959_ (.RESET_B(net350),
    .D(net2458),
    .Q(\u_inv.d_reg[203] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _41960_ (.RESET_B(net349),
    .D(net2111),
    .Q(\u_inv.d_reg[204] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _41961_ (.RESET_B(net348),
    .D(net1146),
    .Q(\u_inv.d_reg[205] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _41962_ (.RESET_B(net347),
    .D(net2217),
    .Q(\u_inv.d_reg[206] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _41963_ (.RESET_B(net346),
    .D(net2692),
    .Q(\u_inv.d_reg[207] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _41964_ (.RESET_B(net345),
    .D(net2922),
    .Q(\u_inv.d_reg[208] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _41965_ (.RESET_B(net344),
    .D(net2738),
    .Q(\u_inv.d_reg[209] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _41966_ (.RESET_B(net343),
    .D(_01241_),
    .Q(\u_inv.d_reg[210] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _41967_ (.RESET_B(net342),
    .D(net2497),
    .Q(\u_inv.d_reg[211] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _41968_ (.RESET_B(net341),
    .D(_01243_),
    .Q(\u_inv.d_reg[212] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _41969_ (.RESET_B(net340),
    .D(net3178),
    .Q(\u_inv.d_reg[213] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _41970_ (.RESET_B(net339),
    .D(_01245_),
    .Q(\u_inv.d_reg[214] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _41971_ (.RESET_B(net338),
    .D(net3096),
    .Q(\u_inv.d_reg[215] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _41972_ (.RESET_B(net336),
    .D(net2576),
    .Q(\u_inv.d_reg[216] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _41973_ (.RESET_B(net334),
    .D(net2061),
    .Q(\u_inv.d_reg[217] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _41974_ (.RESET_B(net332),
    .D(net2531),
    .Q(\u_inv.d_reg[218] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _41975_ (.RESET_B(net330),
    .D(net3092),
    .Q(\u_inv.d_reg[219] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _41976_ (.RESET_B(net328),
    .D(net2989),
    .Q(\u_inv.d_reg[220] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _41977_ (.RESET_B(net326),
    .D(net3188),
    .Q(\u_inv.d_reg[221] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _41978_ (.RESET_B(net324),
    .D(net2529),
    .Q(\u_inv.d_reg[222] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _41979_ (.RESET_B(net322),
    .D(_01254_),
    .Q(\u_inv.d_reg[223] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _41980_ (.RESET_B(net320),
    .D(net2950),
    .Q(\u_inv.d_reg[224] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _41981_ (.RESET_B(net318),
    .D(net1332),
    .Q(\u_inv.d_reg[225] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _41982_ (.RESET_B(net316),
    .D(_01257_),
    .Q(\u_inv.d_reg[226] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _41983_ (.RESET_B(net314),
    .D(net3227),
    .Q(\u_inv.d_reg[227] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _41984_ (.RESET_B(net312),
    .D(net2650),
    .Q(\u_inv.d_reg[228] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _41985_ (.RESET_B(net310),
    .D(net2629),
    .Q(\u_inv.d_reg[229] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _41986_ (.RESET_B(net308),
    .D(_01261_),
    .Q(\u_inv.d_reg[230] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _41987_ (.RESET_B(net306),
    .D(net2574),
    .Q(\u_inv.d_reg[231] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _41988_ (.RESET_B(net304),
    .D(net2792),
    .Q(\u_inv.d_reg[232] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _41989_ (.RESET_B(net302),
    .D(net2572),
    .Q(\u_inv.d_reg[233] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _41990_ (.RESET_B(net300),
    .D(net2379),
    .Q(\u_inv.d_reg[234] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _41991_ (.RESET_B(net298),
    .D(_01266_),
    .Q(\u_inv.d_reg[235] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _41992_ (.RESET_B(net297),
    .D(_01267_),
    .Q(\u_inv.d_reg[236] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _41993_ (.RESET_B(net296),
    .D(_01268_),
    .Q(\u_inv.d_reg[237] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _41994_ (.RESET_B(net295),
    .D(_01269_),
    .Q(\u_inv.d_reg[238] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _41995_ (.RESET_B(net294),
    .D(net3023),
    .Q(\u_inv.d_reg[239] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _41996_ (.RESET_B(net293),
    .D(_01271_),
    .Q(\u_inv.d_reg[240] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _41997_ (.RESET_B(net292),
    .D(net2237),
    .Q(\u_inv.d_reg[241] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _41998_ (.RESET_B(net291),
    .D(net2477),
    .Q(\u_inv.d_reg[242] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _41999_ (.RESET_B(net290),
    .D(net2918),
    .Q(\u_inv.d_reg[243] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _42000_ (.RESET_B(net289),
    .D(net1957),
    .Q(\u_inv.d_reg[244] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _42001_ (.RESET_B(net288),
    .D(net2151),
    .Q(\u_inv.d_reg[245] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _42002_ (.RESET_B(net287),
    .D(_01277_),
    .Q(\u_inv.d_reg[246] ),
    .CLK(clknet_leaf_236_clk));
 sg13g2_dfrbpq_2 _42003_ (.RESET_B(net286),
    .D(net3013),
    .Q(\u_inv.d_reg[247] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _42004_ (.RESET_B(net285),
    .D(net2903),
    .Q(\u_inv.d_reg[248] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _42005_ (.RESET_B(net284),
    .D(net2266),
    .Q(\u_inv.d_reg[249] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _42006_ (.RESET_B(net283),
    .D(_01281_),
    .Q(\u_inv.d_reg[250] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _42007_ (.RESET_B(net282),
    .D(net2659),
    .Q(\u_inv.d_reg[251] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _42008_ (.RESET_B(net281),
    .D(net2507),
    .Q(\u_inv.d_reg[252] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _42009_ (.RESET_B(net280),
    .D(net1420),
    .Q(\u_inv.d_reg[253] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _42010_ (.RESET_B(net279),
    .D(_01285_),
    .Q(\u_inv.d_reg[254] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _42011_ (.RESET_B(net278),
    .D(net2019),
    .Q(\u_inv.d_reg[255] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _42012_ (.RESET_B(net299),
    .D(_01287_),
    .Q(\u_inv.d_reg[256] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _42013_ (.RESET_B(net5904),
    .D(_20877_[0]),
    .Q(\u_inv.load_input ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _42014_ (.RESET_B(net277),
    .D(_01288_),
    .Q(\u_inv.f_reg[0] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _42015_ (.RESET_B(net276),
    .D(net2361),
    .Q(\u_inv.f_reg[1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _42016_ (.RESET_B(net275),
    .D(net2254),
    .Q(\u_inv.f_reg[2] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _42017_ (.RESET_B(net274),
    .D(net2834),
    .Q(\u_inv.f_reg[3] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _42018_ (.RESET_B(net273),
    .D(net2356),
    .Q(\u_inv.f_reg[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _42019_ (.RESET_B(net272),
    .D(net2857),
    .Q(\u_inv.f_reg[5] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _42020_ (.RESET_B(net271),
    .D(net2164),
    .Q(\u_inv.f_reg[6] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _42021_ (.RESET_B(net270),
    .D(net2609),
    .Q(\u_inv.f_reg[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _42022_ (.RESET_B(net269),
    .D(net1245),
    .Q(\u_inv.f_reg[8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _42023_ (.RESET_B(net268),
    .D(net2527),
    .Q(\u_inv.f_reg[9] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _42024_ (.RESET_B(net267),
    .D(net2925),
    .Q(\u_inv.f_reg[10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _42025_ (.RESET_B(net266),
    .D(net2861),
    .Q(\u_inv.f_reg[11] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _42026_ (.RESET_B(net265),
    .D(net3170),
    .Q(\u_inv.f_reg[12] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _42027_ (.RESET_B(net264),
    .D(_01301_),
    .Q(\u_inv.f_reg[13] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _42028_ (.RESET_B(net263),
    .D(net2818),
    .Q(\u_inv.f_reg[14] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _42029_ (.RESET_B(net262),
    .D(net2502),
    .Q(\u_inv.f_reg[15] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _42030_ (.RESET_B(net261),
    .D(net3090),
    .Q(\u_inv.f_reg[16] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _42031_ (.RESET_B(net260),
    .D(net3118),
    .Q(\u_inv.f_reg[17] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _42032_ (.RESET_B(net259),
    .D(net3035),
    .Q(\u_inv.f_reg[18] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _42033_ (.RESET_B(net258),
    .D(net2981),
    .Q(\u_inv.f_reg[19] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _42034_ (.RESET_B(net257),
    .D(net2594),
    .Q(\u_inv.f_reg[20] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _42035_ (.RESET_B(net256),
    .D(net1555),
    .Q(\u_inv.f_reg[21] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _42036_ (.RESET_B(net255),
    .D(net2671),
    .Q(\u_inv.f_reg[22] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _42037_ (.RESET_B(net254),
    .D(_01311_),
    .Q(\u_inv.f_reg[23] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _42038_ (.RESET_B(net253),
    .D(net2852),
    .Q(\u_inv.f_reg[24] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _42039_ (.RESET_B(net252),
    .D(net2999),
    .Q(\u_inv.f_reg[25] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _42040_ (.RESET_B(net251),
    .D(net2465),
    .Q(\u_inv.f_reg[26] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _42041_ (.RESET_B(net1060),
    .D(net2761),
    .Q(\u_inv.f_reg[27] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _42042_ (.RESET_B(net1057),
    .D(net3162),
    .Q(\u_inv.f_reg[28] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _42043_ (.RESET_B(net1054),
    .D(net3148),
    .Q(\u_inv.f_reg[29] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _42044_ (.RESET_B(net1051),
    .D(net3040),
    .Q(\u_inv.f_reg[30] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _42045_ (.RESET_B(net1048),
    .D(net3193),
    .Q(\u_inv.f_reg[31] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _42046_ (.RESET_B(net1045),
    .D(net1744),
    .Q(\u_inv.f_reg[32] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _42047_ (.RESET_B(net1042),
    .D(net3054),
    .Q(\u_inv.f_reg[33] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _42048_ (.RESET_B(net1039),
    .D(net2893),
    .Q(\u_inv.f_reg[34] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _42049_ (.RESET_B(net1036),
    .D(_01323_),
    .Q(\u_inv.f_reg[35] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _42050_ (.RESET_B(net1033),
    .D(net2940),
    .Q(\u_inv.f_reg[36] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_2 _42051_ (.RESET_B(net1030),
    .D(net3285),
    .Q(\u_inv.f_reg[37] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _42052_ (.RESET_B(net1027),
    .D(net2767),
    .Q(\u_inv.f_reg[38] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _42053_ (.RESET_B(net1024),
    .D(net3303),
    .Q(\u_inv.f_reg[39] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _42054_ (.RESET_B(net1021),
    .D(net2891),
    .Q(\u_inv.f_reg[40] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _42055_ (.RESET_B(net1018),
    .D(net3071),
    .Q(\u_inv.f_reg[41] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _42056_ (.RESET_B(net1015),
    .D(net2410),
    .Q(\u_inv.f_reg[42] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _42057_ (.RESET_B(net1012),
    .D(net2699),
    .Q(\u_inv.f_reg[43] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _42058_ (.RESET_B(net1009),
    .D(net2900),
    .Q(\u_inv.f_reg[44] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _42059_ (.RESET_B(net1006),
    .D(net2685),
    .Q(\u_inv.f_reg[45] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _42060_ (.RESET_B(net1003),
    .D(net2243),
    .Q(\u_inv.f_reg[46] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _42061_ (.RESET_B(net1000),
    .D(net2779),
    .Q(\u_inv.f_reg[47] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_2 _42062_ (.RESET_B(net997),
    .D(net3042),
    .Q(\u_inv.f_reg[48] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _42063_ (.RESET_B(net994),
    .D(_01337_),
    .Q(\u_inv.f_reg[49] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _42064_ (.RESET_B(net991),
    .D(net2513),
    .Q(\u_inv.f_reg[50] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _42065_ (.RESET_B(net988),
    .D(net2560),
    .Q(\u_inv.f_reg[51] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _42066_ (.RESET_B(net985),
    .D(net2302),
    .Q(\u_inv.f_reg[52] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _42067_ (.RESET_B(net982),
    .D(net3180),
    .Q(\u_inv.f_reg[53] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _42068_ (.RESET_B(net979),
    .D(net3124),
    .Q(\u_inv.f_reg[54] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _42069_ (.RESET_B(net976),
    .D(net3133),
    .Q(\u_inv.f_reg[55] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _42070_ (.RESET_B(net973),
    .D(net2547),
    .Q(\u_inv.f_reg[56] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _42071_ (.RESET_B(net970),
    .D(_01345_),
    .Q(\u_inv.f_reg[57] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_2 _42072_ (.RESET_B(net967),
    .D(net2878),
    .Q(\u_inv.f_reg[58] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _42073_ (.RESET_B(net964),
    .D(net3110),
    .Q(\u_inv.f_reg[59] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _42074_ (.RESET_B(net961),
    .D(_01348_),
    .Q(\u_inv.f_reg[60] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _42075_ (.RESET_B(net958),
    .D(net2914),
    .Q(\u_inv.f_reg[61] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_2 _42076_ (.RESET_B(net955),
    .D(net1878),
    .Q(\u_inv.f_reg[62] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _42077_ (.RESET_B(net952),
    .D(net2710),
    .Q(\u_inv.f_reg[63] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _42078_ (.RESET_B(net949),
    .D(net2968),
    .Q(\u_inv.f_reg[64] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _42079_ (.RESET_B(net946),
    .D(net2160),
    .Q(\u_inv.f_reg[65] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_2 _42080_ (.RESET_B(net943),
    .D(net2753),
    .Q(\u_inv.f_reg[66] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _42081_ (.RESET_B(net940),
    .D(net3081),
    .Q(\u_inv.f_reg[67] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _42082_ (.RESET_B(net937),
    .D(net2221),
    .Q(\u_inv.f_reg[68] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _42083_ (.RESET_B(net934),
    .D(net2759),
    .Q(\u_inv.f_reg[69] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _42084_ (.RESET_B(net931),
    .D(net2467),
    .Q(\u_inv.f_reg[70] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _42085_ (.RESET_B(net928),
    .D(net3238),
    .Q(\u_inv.f_reg[71] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_2 _42086_ (.RESET_B(net925),
    .D(net3167),
    .Q(\u_inv.f_reg[72] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_2 _42087_ (.RESET_B(net922),
    .D(net3002),
    .Q(\u_inv.f_reg[73] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _42088_ (.RESET_B(net919),
    .D(net3058),
    .Q(\u_inv.f_reg[74] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _42089_ (.RESET_B(net916),
    .D(net3038),
    .Q(\u_inv.f_reg[75] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _42090_ (.RESET_B(net913),
    .D(net2895),
    .Q(\u_inv.f_reg[76] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_1 _42091_ (.RESET_B(net910),
    .D(net3146),
    .Q(\u_inv.f_reg[77] ),
    .CLK(clknet_leaf_172_clk));
 sg13g2_dfrbpq_2 _42092_ (.RESET_B(net907),
    .D(net2696),
    .Q(\u_inv.f_reg[78] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _42093_ (.RESET_B(net904),
    .D(net3103),
    .Q(\u_inv.f_reg[79] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _42094_ (.RESET_B(net901),
    .D(net2772),
    .Q(\u_inv.f_reg[80] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_2 _42095_ (.RESET_B(net898),
    .D(net2826),
    .Q(\u_inv.f_reg[81] ),
    .CLK(clknet_leaf_149_clk));
 sg13g2_dfrbpq_1 _42096_ (.RESET_B(net895),
    .D(net1821),
    .Q(\u_inv.f_reg[82] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _42097_ (.RESET_B(net892),
    .D(net2839),
    .Q(\u_inv.f_reg[83] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _42098_ (.RESET_B(net889),
    .D(net2674),
    .Q(\u_inv.f_reg[84] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_2 _42099_ (.RESET_B(net886),
    .D(net2003),
    .Q(\u_inv.f_reg[85] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_1 _42100_ (.RESET_B(net883),
    .D(net2813),
    .Q(\u_inv.f_reg[86] ),
    .CLK(clknet_leaf_170_clk));
 sg13g2_dfrbpq_2 _42101_ (.RESET_B(net880),
    .D(_01375_),
    .Q(\u_inv.f_reg[87] ),
    .CLK(clknet_leaf_151_clk));
 sg13g2_dfrbpq_2 _42102_ (.RESET_B(net877),
    .D(net2912),
    .Q(\u_inv.f_reg[88] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _42103_ (.RESET_B(net874),
    .D(net2296),
    .Q(\u_inv.f_reg[89] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _42104_ (.RESET_B(net871),
    .D(_01378_),
    .Q(\u_inv.f_reg[90] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_2 _42105_ (.RESET_B(net868),
    .D(net2648),
    .Q(\u_inv.f_reg[91] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _42106_ (.RESET_B(net865),
    .D(net3309),
    .Q(\u_inv.f_reg[92] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_2 _42107_ (.RESET_B(net862),
    .D(net3261),
    .Q(\u_inv.f_reg[93] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _42108_ (.RESET_B(net859),
    .D(net2392),
    .Q(\u_inv.f_reg[94] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _42109_ (.RESET_B(net856),
    .D(net2586),
    .Q(\u_inv.f_reg[95] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _42110_ (.RESET_B(net853),
    .D(_01384_),
    .Q(\u_inv.f_reg[96] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _42111_ (.RESET_B(net850),
    .D(net2615),
    .Q(\u_inv.f_reg[97] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _42112_ (.RESET_B(net847),
    .D(net3209),
    .Q(\u_inv.f_reg[98] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _42113_ (.RESET_B(net844),
    .D(_01387_),
    .Q(\u_inv.f_reg[99] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _42114_ (.RESET_B(net841),
    .D(net2492),
    .Q(\u_inv.f_reg[100] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _42115_ (.RESET_B(net838),
    .D(net2688),
    .Q(\u_inv.f_reg[101] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _42116_ (.RESET_B(net835),
    .D(net3135),
    .Q(\u_inv.f_reg[102] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _42117_ (.RESET_B(net832),
    .D(net3243),
    .Q(\u_inv.f_reg[103] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _42118_ (.RESET_B(net829),
    .D(net2790),
    .Q(\u_inv.f_reg[104] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _42119_ (.RESET_B(net826),
    .D(net3205),
    .Q(\u_inv.f_reg[105] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _42120_ (.RESET_B(net823),
    .D(net2916),
    .Q(\u_inv.f_reg[106] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _42121_ (.RESET_B(net820),
    .D(net3345),
    .Q(\u_inv.f_reg[107] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _42122_ (.RESET_B(net817),
    .D(net1298),
    .Q(\u_inv.f_reg[108] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _42123_ (.RESET_B(net814),
    .D(net3151),
    .Q(\u_inv.f_reg[109] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _42124_ (.RESET_B(net811),
    .D(net2490),
    .Q(\u_inv.f_reg[110] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _42125_ (.RESET_B(net808),
    .D(net3112),
    .Q(\u_inv.f_reg[111] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _42126_ (.RESET_B(net805),
    .D(net3108),
    .Q(\u_inv.f_reg[112] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _42127_ (.RESET_B(net802),
    .D(_01401_),
    .Q(\u_inv.f_reg[113] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _42128_ (.RESET_B(net799),
    .D(net2830),
    .Q(\u_inv.f_reg[114] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _42129_ (.RESET_B(net796),
    .D(net2987),
    .Q(\u_inv.f_reg[115] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _42130_ (.RESET_B(net793),
    .D(net3031),
    .Q(\u_inv.f_reg[116] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _42131_ (.RESET_B(net790),
    .D(net2555),
    .Q(\u_inv.f_reg[117] ),
    .CLK(clknet_leaf_145_clk));
 sg13g2_dfrbpq_2 _42132_ (.RESET_B(net787),
    .D(net2051),
    .Q(\u_inv.f_reg[118] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _42133_ (.RESET_B(net784),
    .D(net3354),
    .Q(\u_inv.f_reg[119] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_2 _42134_ (.RESET_B(net781),
    .D(net2931),
    .Q(\u_inv.f_reg[120] ),
    .CLK(clknet_leaf_138_clk));
 sg13g2_dfrbpq_1 _42135_ (.RESET_B(net778),
    .D(net3203),
    .Q(\u_inv.f_reg[121] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _42136_ (.RESET_B(net775),
    .D(net2039),
    .Q(\u_inv.f_reg[122] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_2 _42137_ (.RESET_B(net772),
    .D(net2235),
    .Q(\u_inv.f_reg[123] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _42138_ (.RESET_B(net769),
    .D(net3114),
    .Q(\u_inv.f_reg[124] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _42139_ (.RESET_B(net766),
    .D(net2847),
    .Q(\u_inv.f_reg[125] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _42140_ (.RESET_B(net763),
    .D(net2747),
    .Q(\u_inv.f_reg[126] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _42141_ (.RESET_B(net760),
    .D(net3176),
    .Q(\u_inv.f_reg[127] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _42142_ (.RESET_B(net757),
    .D(net2784),
    .Q(\u_inv.f_reg[128] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _42143_ (.RESET_B(net754),
    .D(net2666),
    .Q(\u_inv.f_reg[129] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _42144_ (.RESET_B(net750),
    .D(net2472),
    .Q(\u_inv.f_reg[130] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _42145_ (.RESET_B(net747),
    .D(net2500),
    .Q(\u_inv.f_reg[131] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _42146_ (.RESET_B(net744),
    .D(net2662),
    .Q(\u_inv.f_reg[132] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _42147_ (.RESET_B(net741),
    .D(net2456),
    .Q(\u_inv.f_reg[133] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _42148_ (.RESET_B(net738),
    .D(net2959),
    .Q(\u_inv.f_reg[134] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _42149_ (.RESET_B(net735),
    .D(net3164),
    .Q(\u_inv.f_reg[135] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_1 _42150_ (.RESET_B(net732),
    .D(net2566),
    .Q(\u_inv.f_reg[136] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _42151_ (.RESET_B(net729),
    .D(net1369),
    .Q(\u_inv.f_reg[137] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _42152_ (.RESET_B(net726),
    .D(_01426_),
    .Q(\u_inv.f_reg[138] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _42153_ (.RESET_B(net723),
    .D(_01427_),
    .Q(\u_inv.f_reg[139] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _42154_ (.RESET_B(net720),
    .D(net2821),
    .Q(\u_inv.f_reg[140] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _42155_ (.RESET_B(net717),
    .D(net3213),
    .Q(\u_inv.f_reg[141] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _42156_ (.RESET_B(net714),
    .D(net3269),
    .Q(\u_inv.f_reg[142] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _42157_ (.RESET_B(net711),
    .D(net2701),
    .Q(\u_inv.f_reg[143] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _42158_ (.RESET_B(net708),
    .D(net2806),
    .Q(\u_inv.f_reg[144] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _42159_ (.RESET_B(net705),
    .D(net2425),
    .Q(\u_inv.f_reg[145] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _42160_ (.RESET_B(net702),
    .D(net2947),
    .Q(\u_inv.f_reg[146] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _42161_ (.RESET_B(net699),
    .D(net2799),
    .Q(\u_inv.f_reg[147] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _42162_ (.RESET_B(net696),
    .D(net1850),
    .Q(\u_inv.f_reg[148] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _42163_ (.RESET_B(net693),
    .D(_01437_),
    .Q(\u_inv.f_reg[149] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _42164_ (.RESET_B(net690),
    .D(net1926),
    .Q(\u_inv.f_reg[150] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _42165_ (.RESET_B(net687),
    .D(net3182),
    .Q(\u_inv.f_reg[151] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _42166_ (.RESET_B(net684),
    .D(_01440_),
    .Q(\u_inv.f_reg[152] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _42167_ (.RESET_B(net681),
    .D(net3278),
    .Q(\u_inv.f_reg[153] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _42168_ (.RESET_B(net678),
    .D(net3015),
    .Q(\u_inv.f_reg[154] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _42169_ (.RESET_B(net676),
    .D(net3142),
    .Q(\u_inv.f_reg[155] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _42170_ (.RESET_B(net673),
    .D(net2599),
    .Q(\u_inv.f_reg[156] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _42171_ (.RESET_B(net670),
    .D(net3281),
    .Q(\u_inv.f_reg[157] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _42172_ (.RESET_B(net667),
    .D(net2983),
    .Q(\u_inv.f_reg[158] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_1 _42173_ (.RESET_B(net664),
    .D(net3101),
    .Q(\u_inv.f_reg[159] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _42174_ (.RESET_B(net661),
    .D(net3144),
    .Q(\u_inv.f_reg[160] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _42175_ (.RESET_B(net658),
    .D(net2655),
    .Q(\u_inv.f_reg[161] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _42176_ (.RESET_B(net655),
    .D(net2720),
    .Q(\u_inv.f_reg[162] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _42177_ (.RESET_B(net652),
    .D(net2745),
    .Q(\u_inv.f_reg[163] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _42178_ (.RESET_B(net649),
    .D(net2870),
    .Q(\u_inv.f_reg[164] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _42179_ (.RESET_B(net646),
    .D(net2855),
    .Q(\u_inv.f_reg[165] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _42180_ (.RESET_B(net643),
    .D(net1819),
    .Q(\u_inv.f_reg[166] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _42181_ (.RESET_B(net640),
    .D(net3155),
    .Q(\u_inv.f_reg[167] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _42182_ (.RESET_B(net637),
    .D(net3356),
    .Q(\u_inv.f_reg[168] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _42183_ (.RESET_B(net634),
    .D(net3195),
    .Q(\u_inv.f_reg[169] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _42184_ (.RESET_B(net631),
    .D(net2749),
    .Q(\u_inv.f_reg[170] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _42185_ (.RESET_B(net628),
    .D(net3377),
    .Q(\u_inv.f_reg[171] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _42186_ (.RESET_B(net625),
    .D(net3063),
    .Q(\u_inv.f_reg[172] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _42187_ (.RESET_B(net622),
    .D(net3325),
    .Q(\u_inv.f_reg[173] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _42188_ (.RESET_B(net619),
    .D(net2808),
    .Q(\u_inv.f_reg[174] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _42189_ (.RESET_B(net616),
    .D(net3245),
    .Q(\u_inv.f_reg[175] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _42190_ (.RESET_B(net613),
    .D(net3191),
    .Q(\u_inv.f_reg[176] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _42191_ (.RESET_B(net610),
    .D(net3026),
    .Q(\u_inv.f_reg[177] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _42192_ (.RESET_B(net607),
    .D(net3011),
    .Q(\u_inv.f_reg[178] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _42193_ (.RESET_B(net604),
    .D(net2715),
    .Q(\u_inv.f_reg[179] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _42194_ (.RESET_B(net601),
    .D(net3019),
    .Q(\u_inv.f_reg[180] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _42195_ (.RESET_B(net598),
    .D(net2774),
    .Q(\u_inv.f_reg[181] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _42196_ (.RESET_B(net595),
    .D(net2031),
    .Q(\u_inv.f_reg[182] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _42197_ (.RESET_B(net592),
    .D(net2736),
    .Q(\u_inv.f_reg[183] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _42198_ (.RESET_B(net589),
    .D(net3017),
    .Q(\u_inv.f_reg[184] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _42199_ (.RESET_B(net586),
    .D(net2797),
    .Q(\u_inv.f_reg[185] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _42200_ (.RESET_B(net583),
    .D(net2354),
    .Q(\u_inv.f_reg[186] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _42201_ (.RESET_B(net580),
    .D(net2677),
    .Q(\u_inv.f_reg[187] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _42202_ (.RESET_B(net577),
    .D(net2271),
    .Q(\u_inv.f_reg[188] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _42203_ (.RESET_B(net574),
    .D(net3322),
    .Q(\u_inv.f_reg[189] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _42204_ (.RESET_B(net571),
    .D(net2584),
    .Q(\u_inv.f_reg[190] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _42205_ (.RESET_B(net568),
    .D(_01479_),
    .Q(\u_inv.f_reg[191] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_2 _42206_ (.RESET_B(net565),
    .D(net3184),
    .Q(\u_inv.f_reg[192] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _42207_ (.RESET_B(net562),
    .D(net3086),
    .Q(\u_inv.f_reg[193] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _42208_ (.RESET_B(net559),
    .D(net2794),
    .Q(\u_inv.f_reg[194] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _42209_ (.RESET_B(net556),
    .D(net3198),
    .Q(\u_inv.f_reg[195] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _42210_ (.RESET_B(net553),
    .D(net2828),
    .Q(\u_inv.f_reg[196] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _42211_ (.RESET_B(net550),
    .D(net2580),
    .Q(\u_inv.f_reg[197] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_2 _42212_ (.RESET_B(net547),
    .D(net2653),
    .Q(\u_inv.f_reg[198] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _42213_ (.RESET_B(net544),
    .D(net2494),
    .Q(\u_inv.f_reg[199] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_2 _42214_ (.RESET_B(net541),
    .D(net3007),
    .Q(\u_inv.f_reg[200] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _42215_ (.RESET_B(net538),
    .D(_01489_),
    .Q(\u_inv.f_reg[201] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _42216_ (.RESET_B(net535),
    .D(net2804),
    .Q(\u_inv.f_reg[202] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _42217_ (.RESET_B(net532),
    .D(net2256),
    .Q(\u_inv.f_reg[203] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _42218_ (.RESET_B(net529),
    .D(net2282),
    .Q(\u_inv.f_reg[204] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _42219_ (.RESET_B(net526),
    .D(net2352),
    .Q(\u_inv.f_reg[205] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _42220_ (.RESET_B(net523),
    .D(net2765),
    .Q(\u_inv.f_reg[206] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _42221_ (.RESET_B(net520),
    .D(net3229),
    .Q(\u_inv.f_reg[207] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _42222_ (.RESET_B(net517),
    .D(net2414),
    .Q(\u_inv.f_reg[208] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _42223_ (.RESET_B(net514),
    .D(net3240),
    .Q(\u_inv.f_reg[209] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _42224_ (.RESET_B(net511),
    .D(net2482),
    .Q(\u_inv.f_reg[210] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _42225_ (.RESET_B(net508),
    .D(net2533),
    .Q(\u_inv.f_reg[211] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _42226_ (.RESET_B(net505),
    .D(net2298),
    .Q(\u_inv.f_reg[212] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _42227_ (.RESET_B(net502),
    .D(net2541),
    .Q(\u_inv.f_reg[213] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _42228_ (.RESET_B(net499),
    .D(_01502_),
    .Q(\u_inv.f_reg[214] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _42229_ (.RESET_B(net496),
    .D(net2957),
    .Q(\u_inv.f_reg[215] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _42230_ (.RESET_B(net493),
    .D(net3173),
    .Q(\u_inv.f_reg[216] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _42231_ (.RESET_B(net490),
    .D(net3122),
    .Q(\u_inv.f_reg[217] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _42232_ (.RESET_B(net487),
    .D(net3033),
    .Q(\u_inv.f_reg[218] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _42233_ (.RESET_B(net484),
    .D(net3128),
    .Q(\u_inv.f_reg[219] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _42234_ (.RESET_B(net481),
    .D(net1505),
    .Q(\u_inv.f_reg[220] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _42235_ (.RESET_B(net478),
    .D(_01509_),
    .Q(\u_inv.f_reg[221] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _42236_ (.RESET_B(net475),
    .D(net1679),
    .Q(\u_inv.f_reg[222] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _42237_ (.RESET_B(net472),
    .D(net2578),
    .Q(\u_inv.f_reg[223] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _42238_ (.RESET_B(net469),
    .D(net2786),
    .Q(\u_inv.f_reg[224] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _42239_ (.RESET_B(net466),
    .D(net2730),
    .Q(\u_inv.f_reg[225] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _42240_ (.RESET_B(net463),
    .D(net2484),
    .Q(\u_inv.f_reg[226] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _42241_ (.RESET_B(net460),
    .D(net3120),
    .Q(\u_inv.f_reg[227] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _42242_ (.RESET_B(net457),
    .D(net3050),
    .Q(\u_inv.f_reg[228] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _42243_ (.RESET_B(net454),
    .D(net2618),
    .Q(\u_inv.f_reg[229] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _42244_ (.RESET_B(net451),
    .D(net2777),
    .Q(\u_inv.f_reg[230] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _42245_ (.RESET_B(net448),
    .D(net2734),
    .Q(\u_inv.f_reg[231] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _42246_ (.RESET_B(net445),
    .D(net3160),
    .Q(\u_inv.f_reg[232] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _42247_ (.RESET_B(net442),
    .D(net3158),
    .Q(\u_inv.f_reg[233] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _42248_ (.RESET_B(net439),
    .D(net2034),
    .Q(\u_inv.f_reg[234] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _42249_ (.RESET_B(net436),
    .D(net2993),
    .Q(\u_inv.f_reg[235] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _42250_ (.RESET_B(net433),
    .D(net2366),
    .Q(\u_inv.f_reg[236] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _42251_ (.RESET_B(net429),
    .D(net3116),
    .Q(\u_inv.f_reg[237] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _42252_ (.RESET_B(net425),
    .D(net2657),
    .Q(\u_inv.f_reg[238] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _42253_ (.RESET_B(net421),
    .D(net3348),
    .Q(\u_inv.f_reg[239] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _42254_ (.RESET_B(net417),
    .D(net2070),
    .Q(\u_inv.f_reg[240] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _42255_ (.RESET_B(net413),
    .D(net2451),
    .Q(\u_inv.f_reg[241] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _42256_ (.RESET_B(net409),
    .D(net1870),
    .Q(\u_inv.f_reg[242] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _42257_ (.RESET_B(net405),
    .D(net2995),
    .Q(\u_inv.f_reg[243] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _42258_ (.RESET_B(net401),
    .D(net2718),
    .Q(\u_inv.f_reg[244] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _42259_ (.RESET_B(net397),
    .D(net2801),
    .Q(\u_inv.f_reg[245] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _42260_ (.RESET_B(net393),
    .D(net2874),
    .Q(\u_inv.f_reg[246] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _42261_ (.RESET_B(net389),
    .D(net3265),
    .Q(\u_inv.f_reg[247] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _42262_ (.RESET_B(net385),
    .D(net2202),
    .Q(\u_inv.f_reg[248] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _42263_ (.RESET_B(net381),
    .D(net2712),
    .Q(\u_inv.f_reg[249] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _42264_ (.RESET_B(net377),
    .D(net2769),
    .Q(\u_inv.f_reg[250] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _42265_ (.RESET_B(net373),
    .D(net2755),
    .Q(\u_inv.f_reg[251] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _42266_ (.RESET_B(net369),
    .D(net2369),
    .Q(\u_inv.f_reg[252] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _42267_ (.RESET_B(net365),
    .D(net2097),
    .Q(\u_inv.f_reg[253] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _42268_ (.RESET_B(net361),
    .D(net2197),
    .Q(\u_inv.f_reg[254] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _42269_ (.RESET_B(net357),
    .D(net2252),
    .Q(\u_inv.f_reg[255] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _42270_ (.RESET_B(net353),
    .D(_01544_),
    .Q(\u_inv.f_reg[256] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _42271_ (.RESET_B(net5903),
    .D(_01545_),
    .Q(\u_inv.state[0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _42272_ (.RESET_B(net5905),
    .D(_01546_),
    .Q(\u_inv.state[1] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _42273_ (.RESET_B(net5897),
    .D(net1173),
    .Q(\inv_cycles[0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _42274_ (.RESET_B(net5898),
    .D(net1274),
    .Q(\inv_cycles[1] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _42275_ (.RESET_B(net5897),
    .D(net1657),
    .Q(\inv_cycles[2] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _42276_ (.RESET_B(net5896),
    .D(net1125),
    .Q(\inv_cycles[3] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _42277_ (.RESET_B(net5897),
    .D(net1412),
    .Q(\inv_cycles[4] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _42278_ (.RESET_B(net5898),
    .D(net1271),
    .Q(\inv_cycles[5] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _42279_ (.RESET_B(net5898),
    .D(net1365),
    .Q(\inv_cycles[6] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _42280_ (.RESET_B(net5896),
    .D(net1238),
    .Q(\inv_cycles[7] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _42281_ (.RESET_B(net5893),
    .D(net1133),
    .Q(\inv_cycles[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _42282_ (.RESET_B(net5893),
    .D(net1443),
    .Q(\inv_cycles[9] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _42283_ (.RESET_B(net337),
    .D(_01557_),
    .Q(\u_inv.delta_double[0] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _42284_ (.RESET_B(net333),
    .D(net2084),
    .Q(\u_inv.delta_reg[1] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_1 _42285_ (.RESET_B(net329),
    .D(net2843),
    .Q(\u_inv.delta_reg[2] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _42286_ (.RESET_B(net325),
    .D(net2199),
    .Q(\u_inv.delta_reg[3] ),
    .CLK(clknet_leaf_193_clk));
 sg13g2_dfrbpq_2 _42287_ (.RESET_B(net321),
    .D(_01561_),
    .Q(\u_inv.delta_reg[4] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _42288_ (.RESET_B(net317),
    .D(_01562_),
    .Q(\u_inv.delta_reg[5] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _42289_ (.RESET_B(net313),
    .D(_01563_),
    .Q(\u_inv.delta_reg[6] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _42290_ (.RESET_B(net309),
    .D(_01564_),
    .Q(\u_inv.delta_reg[7] ),
    .CLK(clknet_leaf_160_clk));
 sg13g2_dfrbpq_2 _42291_ (.RESET_B(net305),
    .D(_01565_),
    .Q(\u_inv.delta_reg[8] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _42292_ (.RESET_B(net301),
    .D(net1225),
    .Q(\u_inv.delta_reg[9] ),
    .CLK(clknet_leaf_194_clk));
 sg13g2_dfrbpq_2 _42293_ (.RESET_B(net5903),
    .D(_01567_),
    .Q(\u_inv.counter[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _42294_ (.RESET_B(net5894),
    .D(_01568_),
    .Q(\u_inv.input_reg[0] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _42295_ (.RESET_B(net5893),
    .D(net2036),
    .Q(\u_inv.input_reg[1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _42296_ (.RESET_B(net5893),
    .D(_01570_),
    .Q(\u_inv.input_reg[2] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _42297_ (.RESET_B(net5893),
    .D(_01571_),
    .Q(\u_inv.input_reg[3] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _42298_ (.RESET_B(net5893),
    .D(_01572_),
    .Q(\u_inv.input_reg[4] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _42299_ (.RESET_B(net5888),
    .D(_01573_),
    .Q(\u_inv.input_reg[5] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _42300_ (.RESET_B(net5888),
    .D(net1698),
    .Q(\u_inv.input_reg[6] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _42301_ (.RESET_B(net5892),
    .D(_01575_),
    .Q(\u_inv.input_reg[7] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _42302_ (.RESET_B(net5888),
    .D(net1439),
    .Q(\u_inv.input_reg[8] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _42303_ (.RESET_B(net5892),
    .D(net1841),
    .Q(\u_inv.input_reg[9] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _42304_ (.RESET_B(net5892),
    .D(net1215),
    .Q(\u_inv.input_reg[10] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _42305_ (.RESET_B(net5891),
    .D(net1149),
    .Q(\u_inv.input_reg[11] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _42306_ (.RESET_B(net5901),
    .D(net1159),
    .Q(\u_inv.input_reg[12] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _42307_ (.RESET_B(net5901),
    .D(net1162),
    .Q(\u_inv.input_reg[13] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _42308_ (.RESET_B(net5902),
    .D(net1296),
    .Q(\u_inv.input_reg[14] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _42309_ (.RESET_B(net5901),
    .D(net1292),
    .Q(\u_inv.input_reg[15] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _42310_ (.RESET_B(net5886),
    .D(_01584_),
    .Q(\u_inv.input_reg[16] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _42311_ (.RESET_B(net5910),
    .D(net2210),
    .Q(\u_inv.input_reg[17] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _42312_ (.RESET_B(net5910),
    .D(_01586_),
    .Q(\u_inv.input_reg[18] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _42313_ (.RESET_B(net5885),
    .D(_01587_),
    .Q(\u_inv.input_reg[19] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _42314_ (.RESET_B(net5887),
    .D(_01588_),
    .Q(\u_inv.input_reg[20] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _42315_ (.RESET_B(net5909),
    .D(net2072),
    .Q(\u_inv.input_reg[21] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _42316_ (.RESET_B(net5909),
    .D(_01590_),
    .Q(\u_inv.input_reg[22] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _42317_ (.RESET_B(net5909),
    .D(_01591_),
    .Q(\u_inv.input_reg[23] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _42318_ (.RESET_B(net5909),
    .D(_01592_),
    .Q(\u_inv.input_reg[24] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _42319_ (.RESET_B(net5912),
    .D(net1774),
    .Q(\u_inv.input_reg[25] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _42320_ (.RESET_B(net5912),
    .D(_01594_),
    .Q(\u_inv.input_reg[26] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _42321_ (.RESET_B(net5913),
    .D(_01595_),
    .Q(\u_inv.input_reg[27] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _42322_ (.RESET_B(net5911),
    .D(net1991),
    .Q(\u_inv.input_reg[28] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _42323_ (.RESET_B(net5913),
    .D(net2120),
    .Q(\u_inv.input_reg[29] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _42324_ (.RESET_B(net5913),
    .D(net1746),
    .Q(\u_inv.input_reg[30] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _42325_ (.RESET_B(net5913),
    .D(net1839),
    .Q(\u_inv.input_reg[31] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _42326_ (.RESET_B(net5913),
    .D(net1793),
    .Q(\u_inv.input_reg[32] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _42327_ (.RESET_B(net5913),
    .D(_01601_),
    .Q(\u_inv.input_reg[33] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _42328_ (.RESET_B(net5929),
    .D(_01602_),
    .Q(\u_inv.input_reg[34] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _42329_ (.RESET_B(net5929),
    .D(net1754),
    .Q(\u_inv.input_reg[35] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _42330_ (.RESET_B(net5931),
    .D(net1530),
    .Q(\u_inv.input_reg[36] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _42331_ (.RESET_B(net5931),
    .D(_01605_),
    .Q(\u_inv.input_reg[37] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _42332_ (.RESET_B(net5931),
    .D(_01606_),
    .Q(\u_inv.input_reg[38] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _42333_ (.RESET_B(net5931),
    .D(net1929),
    .Q(\u_inv.input_reg[39] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _42334_ (.RESET_B(net5930),
    .D(net1779),
    .Q(\u_inv.input_reg[40] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _42335_ (.RESET_B(net5930),
    .D(net2049),
    .Q(\u_inv.input_reg[41] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _42336_ (.RESET_B(net5933),
    .D(_01610_),
    .Q(\u_inv.input_reg[42] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _42337_ (.RESET_B(net5933),
    .D(net1691),
    .Q(\u_inv.input_reg[43] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _42338_ (.RESET_B(net5934),
    .D(net1740),
    .Q(\u_inv.input_reg[44] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _42339_ (.RESET_B(net5934),
    .D(net1798),
    .Q(\u_inv.input_reg[45] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _42340_ (.RESET_B(net5948),
    .D(_01614_),
    .Q(\u_inv.input_reg[46] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _42341_ (.RESET_B(net5948),
    .D(net1673),
    .Q(\u_inv.input_reg[47] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _42342_ (.RESET_B(net5948),
    .D(net1574),
    .Q(\u_inv.input_reg[48] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _42343_ (.RESET_B(net5947),
    .D(_01617_),
    .Q(\u_inv.input_reg[49] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _42344_ (.RESET_B(net5946),
    .D(_01618_),
    .Q(\u_inv.input_reg[50] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _42345_ (.RESET_B(net5950),
    .D(_01619_),
    .Q(\u_inv.input_reg[51] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _42346_ (.RESET_B(net5950),
    .D(net1456),
    .Q(\u_inv.input_reg[52] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _42347_ (.RESET_B(net5950),
    .D(net1664),
    .Q(\u_inv.input_reg[53] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _42348_ (.RESET_B(net5950),
    .D(net1509),
    .Q(\u_inv.input_reg[54] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _42349_ (.RESET_B(net5950),
    .D(net1484),
    .Q(\u_inv.input_reg[55] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _42350_ (.RESET_B(net5951),
    .D(net2332),
    .Q(\u_inv.input_reg[56] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _42351_ (.RESET_B(net5967),
    .D(net1700),
    .Q(\u_inv.input_reg[57] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _42352_ (.RESET_B(net5967),
    .D(net1655),
    .Q(\u_inv.input_reg[58] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _42353_ (.RESET_B(net5966),
    .D(_01627_),
    .Q(\u_inv.input_reg[59] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_1 _42354_ (.RESET_B(net5966),
    .D(net1437),
    .Q(\u_inv.input_reg[60] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _42355_ (.RESET_B(net5966),
    .D(net1539),
    .Q(\u_inv.input_reg[61] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _42356_ (.RESET_B(net5968),
    .D(net1489),
    .Q(\u_inv.input_reg[62] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _42357_ (.RESET_B(net5966),
    .D(net1458),
    .Q(\u_inv.input_reg[63] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _42358_ (.RESET_B(net5968),
    .D(_01632_),
    .Q(\u_inv.input_reg[64] ),
    .CLK(clknet_leaf_181_clk));
 sg13g2_dfrbpq_1 _42359_ (.RESET_B(net5982),
    .D(_01633_),
    .Q(\u_inv.input_reg[65] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _42360_ (.RESET_B(net5989),
    .D(net1770),
    .Q(\u_inv.input_reg[66] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _42361_ (.RESET_B(net5968),
    .D(_01635_),
    .Q(\u_inv.input_reg[67] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _42362_ (.RESET_B(net5968),
    .D(_01636_),
    .Q(\u_inv.input_reg[68] ),
    .CLK(clknet_leaf_182_clk));
 sg13g2_dfrbpq_1 _42363_ (.RESET_B(net5968),
    .D(net1548),
    .Q(\u_inv.input_reg[69] ),
    .CLK(clknet_leaf_180_clk));
 sg13g2_dfrbpq_1 _42364_ (.RESET_B(net5988),
    .D(_01638_),
    .Q(\u_inv.input_reg[70] ),
    .CLK(clknet_leaf_173_clk));
 sg13g2_dfrbpq_1 _42365_ (.RESET_B(net5989),
    .D(net1515),
    .Q(\u_inv.input_reg[71] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _42366_ (.RESET_B(net5988),
    .D(net1627),
    .Q(\u_inv.input_reg[72] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _42367_ (.RESET_B(net5991),
    .D(net2080),
    .Q(\u_inv.input_reg[73] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _42368_ (.RESET_B(net5988),
    .D(net1651),
    .Q(\u_inv.input_reg[74] ),
    .CLK(clknet_leaf_174_clk));
 sg13g2_dfrbpq_1 _42369_ (.RESET_B(net5992),
    .D(net1592),
    .Q(\u_inv.input_reg[75] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _42370_ (.RESET_B(net5992),
    .D(net1570),
    .Q(\u_inv.input_reg[76] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _42371_ (.RESET_B(net5992),
    .D(net1563),
    .Q(\u_inv.input_reg[77] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _42372_ (.RESET_B(net5998),
    .D(net1889),
    .Q(\u_inv.input_reg[78] ),
    .CLK(clknet_leaf_175_clk));
 sg13g2_dfrbpq_1 _42373_ (.RESET_B(net5998),
    .D(net1462),
    .Q(\u_inv.input_reg[79] ),
    .CLK(clknet_leaf_171_clk));
 sg13g2_dfrbpq_1 _42374_ (.RESET_B(net6001),
    .D(net1590),
    .Q(\u_inv.input_reg[80] ),
    .CLK(clknet_leaf_167_clk));
 sg13g2_dfrbpq_1 _42375_ (.RESET_B(net6001),
    .D(net1579),
    .Q(\u_inv.input_reg[81] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _42376_ (.RESET_B(net6005),
    .D(net1857),
    .Q(\u_inv.input_reg[82] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _42377_ (.RESET_B(net6001),
    .D(net1523),
    .Q(\u_inv.input_reg[83] ),
    .CLK(clknet_leaf_168_clk));
 sg13g2_dfrbpq_1 _42378_ (.RESET_B(net6007),
    .D(_01652_),
    .Q(\u_inv.input_reg[84] ),
    .CLK(clknet_leaf_163_clk));
 sg13g2_dfrbpq_1 _42379_ (.RESET_B(net6007),
    .D(net1908),
    .Q(\u_inv.input_reg[85] ),
    .CLK(clknet_leaf_169_clk));
 sg13g2_dfrbpq_1 _42380_ (.RESET_B(net6007),
    .D(_01654_),
    .Q(\u_inv.input_reg[86] ),
    .CLK(clknet_leaf_164_clk));
 sg13g2_dfrbpq_1 _42381_ (.RESET_B(net6019),
    .D(_01655_),
    .Q(\u_inv.input_reg[87] ),
    .CLK(clknet_leaf_152_clk));
 sg13g2_dfrbpq_1 _42382_ (.RESET_B(net6026),
    .D(net1823),
    .Q(\u_inv.input_reg[88] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _42383_ (.RESET_B(net6015),
    .D(net2078),
    .Q(\u_inv.input_reg[89] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _42384_ (.RESET_B(net6013),
    .D(net1703),
    .Q(\u_inv.input_reg[90] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _42385_ (.RESET_B(net6027),
    .D(net1600),
    .Q(\u_inv.input_reg[91] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _42386_ (.RESET_B(net6027),
    .D(net1577),
    .Q(\u_inv.input_reg[92] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _42387_ (.RESET_B(net6027),
    .D(net2315),
    .Q(\u_inv.input_reg[93] ),
    .CLK(clknet_leaf_156_clk));
 sg13g2_dfrbpq_1 _42388_ (.RESET_B(net6028),
    .D(net1708),
    .Q(\u_inv.input_reg[94] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _42389_ (.RESET_B(net6028),
    .D(net1495),
    .Q(\u_inv.input_reg[95] ),
    .CLK(clknet_leaf_154_clk));
 sg13g2_dfrbpq_1 _42390_ (.RESET_B(net6028),
    .D(net1757),
    .Q(\u_inv.input_reg[96] ),
    .CLK(clknet_leaf_155_clk));
 sg13g2_dfrbpq_1 _42391_ (.RESET_B(net6013),
    .D(net1729),
    .Q(\u_inv.input_reg[97] ),
    .CLK(clknet_leaf_159_clk));
 sg13g2_dfrbpq_1 _42392_ (.RESET_B(net6027),
    .D(_01666_),
    .Q(\u_inv.input_reg[98] ),
    .CLK(clknet_leaf_157_clk));
 sg13g2_dfrbpq_1 _42393_ (.RESET_B(net6029),
    .D(net1513),
    .Q(\u_inv.input_reg[99] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _42394_ (.RESET_B(net6029),
    .D(_01668_),
    .Q(\u_inv.input_reg[100] ),
    .CLK(clknet_leaf_153_clk));
 sg13g2_dfrbpq_1 _42395_ (.RESET_B(net6030),
    .D(net1880),
    .Q(\u_inv.input_reg[101] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _42396_ (.RESET_B(net6029),
    .D(_01670_),
    .Q(\u_inv.input_reg[102] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _42397_ (.RESET_B(net6029),
    .D(net1486),
    .Q(\u_inv.input_reg[103] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _42398_ (.RESET_B(net6024),
    .D(net1931),
    .Q(\u_inv.input_reg[104] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _42399_ (.RESET_B(net6024),
    .D(net2016),
    .Q(\u_inv.input_reg[105] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _42400_ (.RESET_B(net6029),
    .D(net1634),
    .Q(\u_inv.input_reg[106] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _42401_ (.RESET_B(net6024),
    .D(net1448),
    .Q(\u_inv.input_reg[107] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _42402_ (.RESET_B(net6024),
    .D(net1806),
    .Q(\u_inv.input_reg[108] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _42403_ (.RESET_B(net6021),
    .D(net1718),
    .Q(\u_inv.input_reg[109] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _42404_ (.RESET_B(net6030),
    .D(net1918),
    .Q(\u_inv.input_reg[110] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _42405_ (.RESET_B(net6021),
    .D(net1550),
    .Q(\u_inv.input_reg[111] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_1 _42406_ (.RESET_B(net6021),
    .D(net1914),
    .Q(\u_inv.input_reg[112] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_1 _42407_ (.RESET_B(net6017),
    .D(net1893),
    .Q(\u_inv.input_reg[113] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _42408_ (.RESET_B(net6017),
    .D(net1532),
    .Q(\u_inv.input_reg[114] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _42409_ (.RESET_B(net6018),
    .D(net1528),
    .Q(\u_inv.input_reg[115] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _42410_ (.RESET_B(net6017),
    .D(_01684_),
    .Q(\u_inv.input_reg[116] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _42411_ (.RESET_B(net6017),
    .D(net2158),
    .Q(\u_inv.input_reg[117] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _42412_ (.RESET_B(net6018),
    .D(_01686_),
    .Q(\u_inv.input_reg[118] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _42413_ (.RESET_B(net6007),
    .D(net1647),
    .Q(\u_inv.input_reg[119] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _42414_ (.RESET_B(net6010),
    .D(_01688_),
    .Q(\u_inv.input_reg[120] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _42415_ (.RESET_B(net6010),
    .D(net1682),
    .Q(\u_inv.input_reg[121] ),
    .CLK(clknet_leaf_146_clk));
 sg13g2_dfrbpq_1 _42416_ (.RESET_B(net6008),
    .D(net1975),
    .Q(\u_inv.input_reg[122] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _42417_ (.RESET_B(net6010),
    .D(_01691_),
    .Q(\u_inv.input_reg[123] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _42418_ (.RESET_B(net6005),
    .D(_01692_),
    .Q(\u_inv.input_reg[124] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _42419_ (.RESET_B(net6010),
    .D(_01693_),
    .Q(\u_inv.input_reg[125] ),
    .CLK(clknet_leaf_147_clk));
 sg13g2_dfrbpq_1 _42420_ (.RESET_B(net6010),
    .D(_01694_),
    .Q(\u_inv.input_reg[126] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _42421_ (.RESET_B(net6003),
    .D(_01695_),
    .Q(\u_inv.input_reg[127] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _42422_ (.RESET_B(net6003),
    .D(net1687),
    .Q(\u_inv.input_reg[128] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _42423_ (.RESET_B(net6004),
    .D(net1716),
    .Q(\u_inv.input_reg[129] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _42424_ (.RESET_B(net6004),
    .D(net1623),
    .Q(\u_inv.input_reg[130] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _42425_ (.RESET_B(net6004),
    .D(net2068),
    .Q(\u_inv.input_reg[131] ),
    .CLK(clknet_leaf_148_clk));
 sg13g2_dfrbpq_1 _42426_ (.RESET_B(net6003),
    .D(net1588),
    .Q(\u_inv.input_reg[132] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _42427_ (.RESET_B(net6003),
    .D(net1694),
    .Q(\u_inv.input_reg[133] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _42428_ (.RESET_B(net6003),
    .D(_01702_),
    .Q(\u_inv.input_reg[134] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _42429_ (.RESET_B(net6003),
    .D(net1666),
    .Q(\u_inv.input_reg[135] ),
    .CLK(clknet_leaf_133_clk));
 sg13g2_dfrbpq_1 _42430_ (.RESET_B(net5992),
    .D(_01704_),
    .Q(\u_inv.input_reg[136] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _42431_ (.RESET_B(net5994),
    .D(net1557),
    .Q(\u_inv.input_reg[137] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _42432_ (.RESET_B(net5994),
    .D(net1804),
    .Q(\u_inv.input_reg[138] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _42433_ (.RESET_B(net5994),
    .D(net1507),
    .Q(\u_inv.input_reg[139] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _42434_ (.RESET_B(net5994),
    .D(net2026),
    .Q(\u_inv.input_reg[140] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _42435_ (.RESET_B(net5992),
    .D(net2091),
    .Q(\u_inv.input_reg[141] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _42436_ (.RESET_B(net5991),
    .D(net2264),
    .Q(\u_inv.input_reg[142] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _42437_ (.RESET_B(net5994),
    .D(net1653),
    .Q(\u_inv.input_reg[143] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _42438_ (.RESET_B(net6003),
    .D(_01712_),
    .Q(\u_inv.input_reg[144] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _42439_ (.RESET_B(net5994),
    .D(_01713_),
    .Q(\u_inv.input_reg[145] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _42440_ (.RESET_B(net5991),
    .D(_01714_),
    .Q(\u_inv.input_reg[146] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _42441_ (.RESET_B(net5994),
    .D(net1777),
    .Q(\u_inv.input_reg[147] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _42442_ (.RESET_B(net5995),
    .D(net1760),
    .Q(\u_inv.input_reg[148] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _42443_ (.RESET_B(net5990),
    .D(_01717_),
    .Q(\u_inv.input_reg[149] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_dfrbpq_1 _42444_ (.RESET_B(net5987),
    .D(net1852),
    .Q(\u_inv.input_reg[150] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _42445_ (.RESET_B(net5990),
    .D(net1933),
    .Q(\u_inv.input_reg[151] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _42446_ (.RESET_B(net5990),
    .D(net2377),
    .Q(\u_inv.input_reg[152] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _42447_ (.RESET_B(net5990),
    .D(net1860),
    .Q(\u_inv.input_reg[153] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _42448_ (.RESET_B(net5990),
    .D(net1887),
    .Q(\u_inv.input_reg[154] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _42449_ (.RESET_B(net5995),
    .D(net1460),
    .Q(\u_inv.input_reg[155] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _42450_ (.RESET_B(net5979),
    .D(net1817),
    .Q(\u_inv.input_reg[156] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _42451_ (.RESET_B(net5977),
    .D(_01725_),
    .Q(\u_inv.input_reg[157] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _42452_ (.RESET_B(net5979),
    .D(net1941),
    .Q(\u_inv.input_reg[158] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _42453_ (.RESET_B(net5979),
    .D(_01727_),
    .Q(\u_inv.input_reg[159] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _42454_ (.RESET_B(net5979),
    .D(net1596),
    .Q(\u_inv.input_reg[160] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _42455_ (.RESET_B(net5979),
    .D(net1621),
    .Q(\u_inv.input_reg[161] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _42456_ (.RESET_B(net5975),
    .D(_01730_),
    .Q(\u_inv.input_reg[162] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _42457_ (.RESET_B(net5975),
    .D(_01731_),
    .Q(\u_inv.input_reg[163] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _42458_ (.RESET_B(net5971),
    .D(net1608),
    .Q(\u_inv.input_reg[164] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _42459_ (.RESET_B(net5972),
    .D(_01733_),
    .Q(\u_inv.input_reg[165] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _42460_ (.RESET_B(net5971),
    .D(_01734_),
    .Q(\u_inv.input_reg[166] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _42461_ (.RESET_B(net5971),
    .D(net1705),
    .Q(\u_inv.input_reg[167] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_1 _42462_ (.RESET_B(net5971),
    .D(net1724),
    .Q(\u_inv.input_reg[168] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _42463_ (.RESET_B(net5971),
    .D(_01737_),
    .Q(\u_inv.input_reg[169] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _42464_ (.RESET_B(net5980),
    .D(net1736),
    .Q(\u_inv.input_reg[170] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _42465_ (.RESET_B(net5980),
    .D(_01739_),
    .Q(\u_inv.input_reg[171] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _42466_ (.RESET_B(net5974),
    .D(_01740_),
    .Q(\u_inv.input_reg[172] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _42467_ (.RESET_B(net5969),
    .D(net2087),
    .Q(\u_inv.input_reg[173] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _42468_ (.RESET_B(net5969),
    .D(net1441),
    .Q(\u_inv.input_reg[174] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _42469_ (.RESET_B(net5969),
    .D(net1696),
    .Q(\u_inv.input_reg[175] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _42470_ (.RESET_B(net5963),
    .D(_01744_),
    .Q(\u_inv.input_reg[176] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _42471_ (.RESET_B(net5963),
    .D(net1572),
    .Q(\u_inv.input_reg[177] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _42472_ (.RESET_B(net5969),
    .D(_01746_),
    .Q(\u_inv.input_reg[178] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _42473_ (.RESET_B(net5969),
    .D(_01747_),
    .Q(\u_inv.input_reg[179] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _42474_ (.RESET_B(net5963),
    .D(_01748_),
    .Q(\u_inv.input_reg[180] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _42475_ (.RESET_B(net5964),
    .D(net1537),
    .Q(\u_inv.input_reg[181] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _42476_ (.RESET_B(net5960),
    .D(net1896),
    .Q(\u_inv.input_reg[182] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _42477_ (.RESET_B(net5960),
    .D(_01751_),
    .Q(\u_inv.input_reg[183] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _42478_ (.RESET_B(net5960),
    .D(_01752_),
    .Q(\u_inv.input_reg[184] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _42479_ (.RESET_B(net5960),
    .D(net1827),
    .Q(\u_inv.input_reg[185] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _42480_ (.RESET_B(net5960),
    .D(_01754_),
    .Q(\u_inv.input_reg[186] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _42481_ (.RESET_B(net5956),
    .D(net1876),
    .Q(\u_inv.input_reg[187] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _42482_ (.RESET_B(net5956),
    .D(net1971),
    .Q(\u_inv.input_reg[188] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _42483_ (.RESET_B(net5957),
    .D(net1781),
    .Q(\u_inv.input_reg[189] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _42484_ (.RESET_B(net5957),
    .D(net1945),
    .Q(\u_inv.input_reg[190] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _42485_ (.RESET_B(net5956),
    .D(net1684),
    .Q(\u_inv.input_reg[191] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _42486_ (.RESET_B(net5956),
    .D(net1482),
    .Q(\u_inv.input_reg[192] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _42487_ (.RESET_B(net5956),
    .D(net1565),
    .Q(\u_inv.input_reg[193] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _42488_ (.RESET_B(net5953),
    .D(_01762_),
    .Q(\u_inv.input_reg[194] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _42489_ (.RESET_B(net5953),
    .D(net2007),
    .Q(\u_inv.input_reg[195] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _42490_ (.RESET_B(net5953),
    .D(net1961),
    .Q(\u_inv.input_reg[196] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _42491_ (.RESET_B(net5953),
    .D(net1979),
    .Q(\u_inv.input_reg[197] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _42492_ (.RESET_B(net5953),
    .D(_01766_),
    .Q(\u_inv.input_reg[198] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _42493_ (.RESET_B(net5953),
    .D(net1765),
    .Q(\u_inv.input_reg[199] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _42494_ (.RESET_B(net5943),
    .D(net1993),
    .Q(\u_inv.input_reg[200] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _42495_ (.RESET_B(net5943),
    .D(_01769_),
    .Q(\u_inv.input_reg[201] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _42496_ (.RESET_B(net5943),
    .D(_01770_),
    .Q(\u_inv.input_reg[202] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _42497_ (.RESET_B(net5943),
    .D(_01771_),
    .Q(\u_inv.input_reg[203] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _42498_ (.RESET_B(net5943),
    .D(net1676),
    .Q(\u_inv.input_reg[204] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _42499_ (.RESET_B(net5943),
    .D(_01773_),
    .Q(\u_inv.input_reg[205] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _42500_ (.RESET_B(net5940),
    .D(net1874),
    .Q(\u_inv.input_reg[206] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _42501_ (.RESET_B(net5940),
    .D(net2134),
    .Q(\u_inv.input_reg[207] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _42502_ (.RESET_B(net5941),
    .D(net1604),
    .Q(\u_inv.input_reg[208] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _42503_ (.RESET_B(net5941),
    .D(net1748),
    .Q(\u_inv.input_reg[209] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _42504_ (.RESET_B(net5941),
    .D(_01778_),
    .Q(\u_inv.input_reg[210] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _42505_ (.RESET_B(net5941),
    .D(_01779_),
    .Q(\u_inv.input_reg[211] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _42506_ (.RESET_B(net5941),
    .D(_01780_),
    .Q(\u_inv.input_reg[212] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _42507_ (.RESET_B(net5938),
    .D(_01781_),
    .Q(\u_inv.input_reg[213] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _42508_ (.RESET_B(net5938),
    .D(net1987),
    .Q(\u_inv.input_reg[214] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _42509_ (.RESET_B(net5938),
    .D(_01783_),
    .Q(\u_inv.input_reg[215] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _42510_ (.RESET_B(net5938),
    .D(net1619),
    .Q(\u_inv.input_reg[216] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _42511_ (.RESET_B(net5938),
    .D(net1561),
    .Q(\u_inv.input_reg[217] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _42512_ (.RESET_B(net5936),
    .D(net1521),
    .Q(\u_inv.input_reg[218] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _42513_ (.RESET_B(net5936),
    .D(net1541),
    .Q(\u_inv.input_reg[219] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _42514_ (.RESET_B(net5937),
    .D(net1825),
    .Q(\u_inv.input_reg[220] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _42515_ (.RESET_B(net5936),
    .D(_01789_),
    .Q(\u_inv.input_reg[221] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _42516_ (.RESET_B(net5936),
    .D(_01790_),
    .Q(\u_inv.input_reg[222] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _42517_ (.RESET_B(net5936),
    .D(_01791_),
    .Q(\u_inv.input_reg[223] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _42518_ (.RESET_B(net5923),
    .D(net1468),
    .Q(\u_inv.input_reg[224] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _42519_ (.RESET_B(net5923),
    .D(_01793_),
    .Q(\u_inv.input_reg[225] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _42520_ (.RESET_B(net5923),
    .D(_01794_),
    .Q(\u_inv.input_reg[226] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _42521_ (.RESET_B(net5923),
    .D(net1906),
    .Q(\u_inv.input_reg[227] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _42522_ (.RESET_B(net5923),
    .D(net1470),
    .Q(\u_inv.input_reg[228] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _42523_ (.RESET_B(net5923),
    .D(_01797_),
    .Q(\u_inv.input_reg[229] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _42524_ (.RESET_B(net5921),
    .D(_01798_),
    .Q(\u_inv.input_reg[230] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _42525_ (.RESET_B(net5921),
    .D(net1552),
    .Q(\u_inv.input_reg[231] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _42526_ (.RESET_B(net5921),
    .D(net1920),
    .Q(\u_inv.input_reg[232] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _42527_ (.RESET_B(net5921),
    .D(net1815),
    .Q(\u_inv.input_reg[233] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _42528_ (.RESET_B(net5918),
    .D(net1594),
    .Q(\u_inv.input_reg[234] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _42529_ (.RESET_B(net5918),
    .D(net2180),
    .Q(\u_inv.input_reg[235] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _42530_ (.RESET_B(net5921),
    .D(net1638),
    .Q(\u_inv.input_reg[236] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _42531_ (.RESET_B(net5919),
    .D(_01805_),
    .Q(\u_inv.input_reg[237] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _42532_ (.RESET_B(net5918),
    .D(_01806_),
    .Q(\u_inv.input_reg[238] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _42533_ (.RESET_B(net5918),
    .D(_01807_),
    .Q(\u_inv.input_reg[239] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _42534_ (.RESET_B(net5918),
    .D(net1474),
    .Q(\u_inv.input_reg[240] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _42535_ (.RESET_B(net5918),
    .D(net1499),
    .Q(\u_inv.input_reg[241] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _42536_ (.RESET_B(net5917),
    .D(_01810_),
    .Q(\u_inv.input_reg[242] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _42537_ (.RESET_B(net5917),
    .D(_01811_),
    .Q(\u_inv.input_reg[243] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _42538_ (.RESET_B(net5917),
    .D(_01812_),
    .Q(\u_inv.input_reg[244] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _42539_ (.RESET_B(net5917),
    .D(net1834),
    .Q(\u_inv.input_reg[245] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _42540_ (.RESET_B(net5917),
    .D(net1795),
    .Q(\u_inv.input_reg[246] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _42541_ (.RESET_B(net5902),
    .D(_01815_),
    .Q(\u_inv.input_reg[247] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _42542_ (.RESET_B(net5903),
    .D(net1643),
    .Q(\u_inv.input_reg[248] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _42543_ (.RESET_B(net5900),
    .D(_01817_),
    .Q(\u_inv.input_reg[249] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _42544_ (.RESET_B(net5903),
    .D(net1649),
    .Q(\u_inv.input_reg[250] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _42545_ (.RESET_B(net5901),
    .D(net1491),
    .Q(\u_inv.input_reg[251] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _42546_ (.RESET_B(net5902),
    .D(net1636),
    .Q(\u_inv.input_reg[252] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _42547_ (.RESET_B(net5902),
    .D(net2289),
    .Q(\u_inv.input_reg[253] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _42548_ (.RESET_B(net5901),
    .D(_01822_),
    .Q(\u_inv.input_reg[254] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _42549_ (.RESET_B(net5902),
    .D(net1606),
    .Q(\u_inv.input_reg[255] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _42550_ (.RESET_B(net5904),
    .D(net1966),
    .Q(pipe_pending),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _42551_ (.RESET_B(net431),
    .D(_01825_),
    .Q(\u_inv.f_next[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _42552_ (.RESET_B(net427),
    .D(_01826_),
    .Q(\u_inv.f_next[1] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _42553_ (.RESET_B(net423),
    .D(_01827_),
    .Q(\u_inv.f_next[2] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _42554_ (.RESET_B(net419),
    .D(_01828_),
    .Q(\u_inv.f_next[3] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _42555_ (.RESET_B(net415),
    .D(_01829_),
    .Q(\u_inv.f_next[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _42556_ (.RESET_B(net411),
    .D(_01830_),
    .Q(\u_inv.f_next[5] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _42557_ (.RESET_B(net407),
    .D(_01831_),
    .Q(\u_inv.f_next[6] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _42558_ (.RESET_B(net403),
    .D(_01832_),
    .Q(\u_inv.f_next[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _42559_ (.RESET_B(net399),
    .D(_01833_),
    .Q(\u_inv.f_next[8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _42560_ (.RESET_B(net395),
    .D(_01834_),
    .Q(\u_inv.f_next[9] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _42561_ (.RESET_B(net391),
    .D(_01835_),
    .Q(\u_inv.f_next[10] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _42562_ (.RESET_B(net387),
    .D(_01836_),
    .Q(\u_inv.f_next[11] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _42563_ (.RESET_B(net383),
    .D(_01837_),
    .Q(\u_inv.f_next[12] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _42564_ (.RESET_B(net379),
    .D(_01838_),
    .Q(\u_inv.f_next[13] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _42565_ (.RESET_B(net375),
    .D(_01839_),
    .Q(\u_inv.f_next[14] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _42566_ (.RESET_B(net371),
    .D(_01840_),
    .Q(\u_inv.f_next[15] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _42567_ (.RESET_B(net367),
    .D(_01841_),
    .Q(\u_inv.f_next[16] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _42568_ (.RESET_B(net363),
    .D(_01842_),
    .Q(\u_inv.f_next[17] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _42569_ (.RESET_B(net359),
    .D(_01843_),
    .Q(\u_inv.f_next[18] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _42570_ (.RESET_B(net355),
    .D(_01844_),
    .Q(\u_inv.f_next[19] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _42571_ (.RESET_B(net351),
    .D(_01845_),
    .Q(\u_inv.f_next[20] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _42572_ (.RESET_B(net335),
    .D(_01846_),
    .Q(\u_inv.f_next[21] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _42573_ (.RESET_B(net331),
    .D(_01847_),
    .Q(\u_inv.f_next[22] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _42574_ (.RESET_B(net327),
    .D(_01848_),
    .Q(\u_inv.f_next[23] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _42575_ (.RESET_B(net323),
    .D(_01849_),
    .Q(\u_inv.f_next[24] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _42576_ (.RESET_B(net319),
    .D(_01850_),
    .Q(\u_inv.f_next[25] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _42577_ (.RESET_B(net315),
    .D(_01851_),
    .Q(\u_inv.f_next[26] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _42578_ (.RESET_B(net311),
    .D(_01852_),
    .Q(\u_inv.f_next[27] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _42579_ (.RESET_B(net307),
    .D(_01853_),
    .Q(\u_inv.f_next[28] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _42580_ (.RESET_B(net303),
    .D(_01854_),
    .Q(\u_inv.f_next[29] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_tiehi _40722__25 (.L_HI(net25));
 sg13g2_tiehi _40947__26 (.L_HI(net26));
 sg13g2_tiehi _40946__27 (.L_HI(net27));
 sg13g2_tiehi _40945__28 (.L_HI(net28));
 sg13g2_tiehi _40944__29 (.L_HI(net29));
 sg13g2_tiehi _40943__30 (.L_HI(net30));
 sg13g2_tiehi _40942__31 (.L_HI(net31));
 sg13g2_tiehi _40941__32 (.L_HI(net32));
 sg13g2_tiehi _40940__33 (.L_HI(net33));
 sg13g2_tiehi _40939__34 (.L_HI(net34));
 sg13g2_tiehi _40938__35 (.L_HI(net35));
 sg13g2_tiehi _40937__36 (.L_HI(net36));
 sg13g2_tiehi _40936__37 (.L_HI(net37));
 sg13g2_tiehi _40935__38 (.L_HI(net38));
 sg13g2_tiehi _40934__39 (.L_HI(net39));
 sg13g2_tiehi _40933__40 (.L_HI(net40));
 sg13g2_tiehi _40932__41 (.L_HI(net41));
 sg13g2_tiehi _40931__42 (.L_HI(net42));
 sg13g2_tiehi _40930__43 (.L_HI(net43));
 sg13g2_tiehi _40929__44 (.L_HI(net44));
 sg13g2_tiehi _40928__45 (.L_HI(net45));
 sg13g2_tiehi _40927__46 (.L_HI(net46));
 sg13g2_tiehi _40926__47 (.L_HI(net47));
 sg13g2_tiehi _40925__48 (.L_HI(net48));
 sg13g2_tiehi _40924__49 (.L_HI(net49));
 sg13g2_tiehi _40923__50 (.L_HI(net50));
 sg13g2_tiehi _40922__51 (.L_HI(net51));
 sg13g2_tiehi _40921__52 (.L_HI(net52));
 sg13g2_tiehi _40920__53 (.L_HI(net53));
 sg13g2_tiehi _40919__54 (.L_HI(net54));
 sg13g2_tiehi _40918__55 (.L_HI(net55));
 sg13g2_tiehi _40917__56 (.L_HI(net56));
 sg13g2_tiehi _40916__57 (.L_HI(net57));
 sg13g2_tiehi _40915__58 (.L_HI(net58));
 sg13g2_tiehi _40914__59 (.L_HI(net59));
 sg13g2_tiehi _40913__60 (.L_HI(net60));
 sg13g2_tiehi _40912__61 (.L_HI(net61));
 sg13g2_tiehi _40911__62 (.L_HI(net62));
 sg13g2_tiehi _40910__63 (.L_HI(net63));
 sg13g2_tiehi _40909__64 (.L_HI(net64));
 sg13g2_tiehi _40908__65 (.L_HI(net65));
 sg13g2_tiehi _40907__66 (.L_HI(net66));
 sg13g2_tiehi _40906__67 (.L_HI(net67));
 sg13g2_tiehi _40905__68 (.L_HI(net68));
 sg13g2_tiehi _40904__69 (.L_HI(net69));
 sg13g2_tiehi _40903__70 (.L_HI(net70));
 sg13g2_tiehi _40902__71 (.L_HI(net71));
 sg13g2_tiehi _40901__72 (.L_HI(net72));
 sg13g2_tiehi _40900__73 (.L_HI(net73));
 sg13g2_tiehi _40899__74 (.L_HI(net74));
 sg13g2_tiehi _40898__75 (.L_HI(net75));
 sg13g2_tiehi _40897__76 (.L_HI(net76));
 sg13g2_tiehi _40896__77 (.L_HI(net77));
 sg13g2_tiehi _40895__78 (.L_HI(net78));
 sg13g2_tiehi _40894__79 (.L_HI(net79));
 sg13g2_tiehi _40893__80 (.L_HI(net80));
 sg13g2_tiehi _40892__81 (.L_HI(net81));
 sg13g2_tiehi _40891__82 (.L_HI(net82));
 sg13g2_tiehi _40890__83 (.L_HI(net83));
 sg13g2_tiehi _40889__84 (.L_HI(net84));
 sg13g2_tiehi _40888__85 (.L_HI(net85));
 sg13g2_tiehi _40887__86 (.L_HI(net86));
 sg13g2_tiehi _40886__87 (.L_HI(net87));
 sg13g2_tiehi _40885__88 (.L_HI(net88));
 sg13g2_tiehi _40884__89 (.L_HI(net89));
 sg13g2_tiehi _40883__90 (.L_HI(net90));
 sg13g2_tiehi _40882__91 (.L_HI(net91));
 sg13g2_tiehi _40881__92 (.L_HI(net92));
 sg13g2_tiehi _40880__93 (.L_HI(net93));
 sg13g2_tiehi _40879__94 (.L_HI(net94));
 sg13g2_tiehi _40878__95 (.L_HI(net95));
 sg13g2_tiehi _40877__96 (.L_HI(net96));
 sg13g2_tiehi _40876__97 (.L_HI(net97));
 sg13g2_tiehi _40875__98 (.L_HI(net98));
 sg13g2_tiehi _40874__99 (.L_HI(net99));
 sg13g2_tiehi _40873__100 (.L_HI(net100));
 sg13g2_tiehi _40872__101 (.L_HI(net101));
 sg13g2_tiehi _40871__102 (.L_HI(net102));
 sg13g2_tiehi _40870__103 (.L_HI(net103));
 sg13g2_tiehi _40869__104 (.L_HI(net104));
 sg13g2_tiehi _40868__105 (.L_HI(net105));
 sg13g2_tiehi _40867__106 (.L_HI(net106));
 sg13g2_tiehi _40866__107 (.L_HI(net107));
 sg13g2_tiehi _40865__108 (.L_HI(net108));
 sg13g2_tiehi _40864__109 (.L_HI(net109));
 sg13g2_tiehi _40863__110 (.L_HI(net110));
 sg13g2_tiehi _40862__111 (.L_HI(net111));
 sg13g2_tiehi _40861__112 (.L_HI(net112));
 sg13g2_tiehi _40860__113 (.L_HI(net113));
 sg13g2_tiehi _40859__114 (.L_HI(net114));
 sg13g2_tiehi _40858__115 (.L_HI(net115));
 sg13g2_tiehi _40857__116 (.L_HI(net116));
 sg13g2_tiehi _40856__117 (.L_HI(net117));
 sg13g2_tiehi _40855__118 (.L_HI(net118));
 sg13g2_tiehi _40854__119 (.L_HI(net119));
 sg13g2_tiehi _40853__120 (.L_HI(net120));
 sg13g2_tiehi _40852__121 (.L_HI(net121));
 sg13g2_tiehi _40851__122 (.L_HI(net122));
 sg13g2_tiehi _40850__123 (.L_HI(net123));
 sg13g2_tiehi _40849__124 (.L_HI(net124));
 sg13g2_tiehi _40848__125 (.L_HI(net125));
 sg13g2_tiehi _40847__126 (.L_HI(net126));
 sg13g2_tiehi _40846__127 (.L_HI(net127));
 sg13g2_tiehi _40845__128 (.L_HI(net128));
 sg13g2_tiehi _40844__129 (.L_HI(net129));
 sg13g2_tiehi _40843__130 (.L_HI(net130));
 sg13g2_tiehi _40842__131 (.L_HI(net131));
 sg13g2_tiehi _40841__132 (.L_HI(net132));
 sg13g2_tiehi _40840__133 (.L_HI(net133));
 sg13g2_tiehi _40839__134 (.L_HI(net134));
 sg13g2_tiehi _40838__135 (.L_HI(net135));
 sg13g2_tiehi _40837__136 (.L_HI(net136));
 sg13g2_tiehi _40836__137 (.L_HI(net137));
 sg13g2_tiehi _40835__138 (.L_HI(net138));
 sg13g2_tiehi _40834__139 (.L_HI(net139));
 sg13g2_tiehi _40833__140 (.L_HI(net140));
 sg13g2_tiehi _40832__141 (.L_HI(net141));
 sg13g2_tiehi _40831__142 (.L_HI(net142));
 sg13g2_tiehi _40830__143 (.L_HI(net143));
 sg13g2_tiehi _40829__144 (.L_HI(net144));
 sg13g2_tiehi _40828__145 (.L_HI(net145));
 sg13g2_tiehi _40827__146 (.L_HI(net146));
 sg13g2_tiehi _40826__147 (.L_HI(net147));
 sg13g2_tiehi _40825__148 (.L_HI(net148));
 sg13g2_tiehi _40824__149 (.L_HI(net149));
 sg13g2_tiehi _40823__150 (.L_HI(net150));
 sg13g2_tiehi _40822__151 (.L_HI(net151));
 sg13g2_tiehi _40821__152 (.L_HI(net152));
 sg13g2_tiehi _40820__153 (.L_HI(net153));
 sg13g2_tiehi _40819__154 (.L_HI(net154));
 sg13g2_tiehi _40818__155 (.L_HI(net155));
 sg13g2_tiehi _40817__156 (.L_HI(net156));
 sg13g2_tiehi _40816__157 (.L_HI(net157));
 sg13g2_tiehi _40815__158 (.L_HI(net158));
 sg13g2_tiehi _40814__159 (.L_HI(net159));
 sg13g2_tiehi _40813__160 (.L_HI(net160));
 sg13g2_tiehi _40812__161 (.L_HI(net161));
 sg13g2_tiehi _40811__162 (.L_HI(net162));
 sg13g2_tiehi _40810__163 (.L_HI(net163));
 sg13g2_tiehi _40809__164 (.L_HI(net164));
 sg13g2_tiehi _40808__165 (.L_HI(net165));
 sg13g2_tiehi _40807__166 (.L_HI(net166));
 sg13g2_tiehi _40806__167 (.L_HI(net167));
 sg13g2_tiehi _40805__168 (.L_HI(net168));
 sg13g2_tiehi _40804__169 (.L_HI(net169));
 sg13g2_tiehi _40803__170 (.L_HI(net170));
 sg13g2_tiehi _40802__171 (.L_HI(net171));
 sg13g2_tiehi _40801__172 (.L_HI(net172));
 sg13g2_tiehi _40800__173 (.L_HI(net173));
 sg13g2_tiehi _40799__174 (.L_HI(net174));
 sg13g2_tiehi _40798__175 (.L_HI(net175));
 sg13g2_tiehi _40797__176 (.L_HI(net176));
 sg13g2_tiehi _40796__177 (.L_HI(net177));
 sg13g2_tiehi _40795__178 (.L_HI(net178));
 sg13g2_tiehi _40794__179 (.L_HI(net179));
 sg13g2_tiehi _40793__180 (.L_HI(net180));
 sg13g2_tiehi _40792__181 (.L_HI(net181));
 sg13g2_tiehi _40791__182 (.L_HI(net182));
 sg13g2_tiehi _40790__183 (.L_HI(net183));
 sg13g2_tiehi _40789__184 (.L_HI(net184));
 sg13g2_tiehi _40788__185 (.L_HI(net185));
 sg13g2_tiehi _40787__186 (.L_HI(net186));
 sg13g2_tiehi _40786__187 (.L_HI(net187));
 sg13g2_tiehi _40785__188 (.L_HI(net188));
 sg13g2_tiehi _40784__189 (.L_HI(net189));
 sg13g2_tiehi _40783__190 (.L_HI(net190));
 sg13g2_tiehi _40782__191 (.L_HI(net191));
 sg13g2_tiehi _40781__192 (.L_HI(net192));
 sg13g2_tiehi _40780__193 (.L_HI(net193));
 sg13g2_tiehi _40779__194 (.L_HI(net194));
 sg13g2_tiehi _40778__195 (.L_HI(net195));
 sg13g2_tiehi _40777__196 (.L_HI(net196));
 sg13g2_tiehi _40776__197 (.L_HI(net197));
 sg13g2_tiehi _40775__198 (.L_HI(net198));
 sg13g2_tiehi _40774__199 (.L_HI(net199));
 sg13g2_tiehi _40773__200 (.L_HI(net200));
 sg13g2_tiehi _40772__201 (.L_HI(net201));
 sg13g2_tiehi _40771__202 (.L_HI(net202));
 sg13g2_tiehi _40770__203 (.L_HI(net203));
 sg13g2_tiehi _40769__204 (.L_HI(net204));
 sg13g2_tiehi _40768__205 (.L_HI(net205));
 sg13g2_tiehi _40767__206 (.L_HI(net206));
 sg13g2_tiehi _40766__207 (.L_HI(net207));
 sg13g2_tiehi _40765__208 (.L_HI(net208));
 sg13g2_tiehi _40764__209 (.L_HI(net209));
 sg13g2_tiehi _40763__210 (.L_HI(net210));
 sg13g2_tiehi _40762__211 (.L_HI(net211));
 sg13g2_tiehi _40761__212 (.L_HI(net212));
 sg13g2_tiehi _40760__213 (.L_HI(net213));
 sg13g2_tiehi _40759__214 (.L_HI(net214));
 sg13g2_tiehi _40758__215 (.L_HI(net215));
 sg13g2_tiehi _40757__216 (.L_HI(net216));
 sg13g2_tiehi _40756__217 (.L_HI(net217));
 sg13g2_tiehi _40755__218 (.L_HI(net218));
 sg13g2_tiehi _40754__219 (.L_HI(net219));
 sg13g2_tiehi _40753__220 (.L_HI(net220));
 sg13g2_tiehi _40752__221 (.L_HI(net221));
 sg13g2_tiehi _40751__222 (.L_HI(net222));
 sg13g2_tiehi _40750__223 (.L_HI(net223));
 sg13g2_tiehi _40749__224 (.L_HI(net224));
 sg13g2_tiehi _40748__225 (.L_HI(net225));
 sg13g2_tiehi _40747__226 (.L_HI(net226));
 sg13g2_tiehi _40746__227 (.L_HI(net227));
 sg13g2_tiehi _40745__228 (.L_HI(net228));
 sg13g2_tiehi _40744__229 (.L_HI(net229));
 sg13g2_tiehi _40743__230 (.L_HI(net230));
 sg13g2_tiehi _40742__231 (.L_HI(net231));
 sg13g2_tiehi _40741__232 (.L_HI(net232));
 sg13g2_tiehi _40740__233 (.L_HI(net233));
 sg13g2_tiehi _40739__234 (.L_HI(net234));
 sg13g2_tiehi _40738__235 (.L_HI(net235));
 sg13g2_tiehi _40737__236 (.L_HI(net236));
 sg13g2_tiehi _40736__237 (.L_HI(net237));
 sg13g2_tiehi _40735__238 (.L_HI(net238));
 sg13g2_tiehi _40734__239 (.L_HI(net239));
 sg13g2_tiehi _40733__240 (.L_HI(net240));
 sg13g2_tiehi _40732__241 (.L_HI(net241));
 sg13g2_tiehi _40731__242 (.L_HI(net242));
 sg13g2_tiehi _40730__243 (.L_HI(net243));
 sg13g2_tiehi _40729__244 (.L_HI(net244));
 sg13g2_tiehi _40728__245 (.L_HI(net245));
 sg13g2_tiehi _40727__246 (.L_HI(net246));
 sg13g2_tiehi _40726__247 (.L_HI(net247));
 sg13g2_tiehi _40725__248 (.L_HI(net248));
 sg13g2_tiehi _40724__249 (.L_HI(net249));
 sg13g2_tiehi _40723__250 (.L_HI(net250));
 sg13g2_tiehi _42040__251 (.L_HI(net251));
 sg13g2_tiehi _42039__252 (.L_HI(net252));
 sg13g2_tiehi _42038__253 (.L_HI(net253));
 sg13g2_tiehi _42037__254 (.L_HI(net254));
 sg13g2_tiehi _42036__255 (.L_HI(net255));
 sg13g2_tiehi _42035__256 (.L_HI(net256));
 sg13g2_tiehi _42034__257 (.L_HI(net257));
 sg13g2_tiehi _42033__258 (.L_HI(net258));
 sg13g2_tiehi _42032__259 (.L_HI(net259));
 sg13g2_tiehi _42031__260 (.L_HI(net260));
 sg13g2_tiehi _42030__261 (.L_HI(net261));
 sg13g2_tiehi _42029__262 (.L_HI(net262));
 sg13g2_tiehi _42028__263 (.L_HI(net263));
 sg13g2_tiehi _42027__264 (.L_HI(net264));
 sg13g2_tiehi _42026__265 (.L_HI(net265));
 sg13g2_tiehi _42025__266 (.L_HI(net266));
 sg13g2_tiehi _42024__267 (.L_HI(net267));
 sg13g2_tiehi _42023__268 (.L_HI(net268));
 sg13g2_tiehi _42022__269 (.L_HI(net269));
 sg13g2_tiehi _42021__270 (.L_HI(net270));
 sg13g2_tiehi _42020__271 (.L_HI(net271));
 sg13g2_tiehi _42019__272 (.L_HI(net272));
 sg13g2_tiehi _42018__273 (.L_HI(net273));
 sg13g2_tiehi _42017__274 (.L_HI(net274));
 sg13g2_tiehi _42016__275 (.L_HI(net275));
 sg13g2_tiehi _42015__276 (.L_HI(net276));
 sg13g2_tiehi _42014__277 (.L_HI(net277));
 sg13g2_tiehi _42011__278 (.L_HI(net278));
 sg13g2_tiehi _42010__279 (.L_HI(net279));
 sg13g2_tiehi _42009__280 (.L_HI(net280));
 sg13g2_tiehi _42008__281 (.L_HI(net281));
 sg13g2_tiehi _42007__282 (.L_HI(net282));
 sg13g2_tiehi _42006__283 (.L_HI(net283));
 sg13g2_tiehi _42005__284 (.L_HI(net284));
 sg13g2_tiehi _42004__285 (.L_HI(net285));
 sg13g2_tiehi _42003__286 (.L_HI(net286));
 sg13g2_tiehi _42002__287 (.L_HI(net287));
 sg13g2_tiehi _42001__288 (.L_HI(net288));
 sg13g2_tiehi _42000__289 (.L_HI(net289));
 sg13g2_tiehi _41999__290 (.L_HI(net290));
 sg13g2_tiehi _41998__291 (.L_HI(net291));
 sg13g2_tiehi _41997__292 (.L_HI(net292));
 sg13g2_tiehi _41996__293 (.L_HI(net293));
 sg13g2_tiehi _41995__294 (.L_HI(net294));
 sg13g2_tiehi _41994__295 (.L_HI(net295));
 sg13g2_tiehi _41993__296 (.L_HI(net296));
 sg13g2_tiehi _41992__297 (.L_HI(net297));
 sg13g2_tiehi _41991__298 (.L_HI(net298));
 sg13g2_tiehi _42012__299 (.L_HI(net299));
 sg13g2_tiehi _41990__300 (.L_HI(net300));
 sg13g2_tiehi _42292__301 (.L_HI(net301));
 sg13g2_tiehi _41989__302 (.L_HI(net302));
 sg13g2_tiehi _42580__303 (.L_HI(net303));
 sg13g2_tiehi _41988__304 (.L_HI(net304));
 sg13g2_tiehi _42291__305 (.L_HI(net305));
 sg13g2_tiehi _41987__306 (.L_HI(net306));
 sg13g2_tiehi _42579__307 (.L_HI(net307));
 sg13g2_tiehi _41986__308 (.L_HI(net308));
 sg13g2_tiehi _42290__309 (.L_HI(net309));
 sg13g2_tiehi _41985__310 (.L_HI(net310));
 sg13g2_tiehi _42578__311 (.L_HI(net311));
 sg13g2_tiehi _41984__312 (.L_HI(net312));
 sg13g2_tiehi _42289__313 (.L_HI(net313));
 sg13g2_tiehi _41983__314 (.L_HI(net314));
 sg13g2_tiehi _42577__315 (.L_HI(net315));
 sg13g2_tiehi _41982__316 (.L_HI(net316));
 sg13g2_tiehi _42288__317 (.L_HI(net317));
 sg13g2_tiehi _41981__318 (.L_HI(net318));
 sg13g2_tiehi _42576__319 (.L_HI(net319));
 sg13g2_tiehi _41980__320 (.L_HI(net320));
 sg13g2_tiehi _42287__321 (.L_HI(net321));
 sg13g2_tiehi _41979__322 (.L_HI(net322));
 sg13g2_tiehi _42575__323 (.L_HI(net323));
 sg13g2_tiehi _41978__324 (.L_HI(net324));
 sg13g2_tiehi _42286__325 (.L_HI(net325));
 sg13g2_tiehi _41977__326 (.L_HI(net326));
 sg13g2_tiehi _42574__327 (.L_HI(net327));
 sg13g2_tiehi _41976__328 (.L_HI(net328));
 sg13g2_tiehi _42285__329 (.L_HI(net329));
 sg13g2_tiehi _41975__330 (.L_HI(net330));
 sg13g2_tiehi _42573__331 (.L_HI(net331));
 sg13g2_tiehi _41974__332 (.L_HI(net332));
 sg13g2_tiehi _42284__333 (.L_HI(net333));
 sg13g2_tiehi _41973__334 (.L_HI(net334));
 sg13g2_tiehi _42572__335 (.L_HI(net335));
 sg13g2_tiehi _41972__336 (.L_HI(net336));
 sg13g2_tiehi _42283__337 (.L_HI(net337));
 sg13g2_tiehi _41971__338 (.L_HI(net338));
 sg13g2_tiehi _41970__339 (.L_HI(net339));
 sg13g2_tiehi _41969__340 (.L_HI(net340));
 sg13g2_tiehi _41968__341 (.L_HI(net341));
 sg13g2_tiehi _41967__342 (.L_HI(net342));
 sg13g2_tiehi _41966__343 (.L_HI(net343));
 sg13g2_tiehi _41965__344 (.L_HI(net344));
 sg13g2_tiehi _41964__345 (.L_HI(net345));
 sg13g2_tiehi _41963__346 (.L_HI(net346));
 sg13g2_tiehi _41962__347 (.L_HI(net347));
 sg13g2_tiehi _41961__348 (.L_HI(net348));
 sg13g2_tiehi _41960__349 (.L_HI(net349));
 sg13g2_tiehi _41959__350 (.L_HI(net350));
 sg13g2_tiehi _42571__351 (.L_HI(net351));
 sg13g2_tiehi _41958__352 (.L_HI(net352));
 sg13g2_tiehi _42270__353 (.L_HI(net353));
 sg13g2_tiehi _41957__354 (.L_HI(net354));
 sg13g2_tiehi _42570__355 (.L_HI(net355));
 sg13g2_tiehi _41956__356 (.L_HI(net356));
 sg13g2_tiehi _42269__357 (.L_HI(net357));
 sg13g2_tiehi _41955__358 (.L_HI(net358));
 sg13g2_tiehi _42569__359 (.L_HI(net359));
 sg13g2_tiehi _41954__360 (.L_HI(net360));
 sg13g2_tiehi _42268__361 (.L_HI(net361));
 sg13g2_tiehi _41953__362 (.L_HI(net362));
 sg13g2_tiehi _42568__363 (.L_HI(net363));
 sg13g2_tiehi _41952__364 (.L_HI(net364));
 sg13g2_tiehi _42267__365 (.L_HI(net365));
 sg13g2_tiehi _41951__366 (.L_HI(net366));
 sg13g2_tiehi _42567__367 (.L_HI(net367));
 sg13g2_tiehi _41950__368 (.L_HI(net368));
 sg13g2_tiehi _42266__369 (.L_HI(net369));
 sg13g2_tiehi _41949__370 (.L_HI(net370));
 sg13g2_tiehi _42566__371 (.L_HI(net371));
 sg13g2_tiehi _41948__372 (.L_HI(net372));
 sg13g2_tiehi _42265__373 (.L_HI(net373));
 sg13g2_tiehi _41947__374 (.L_HI(net374));
 sg13g2_tiehi _42565__375 (.L_HI(net375));
 sg13g2_tiehi _41946__376 (.L_HI(net376));
 sg13g2_tiehi _42264__377 (.L_HI(net377));
 sg13g2_tiehi _41945__378 (.L_HI(net378));
 sg13g2_tiehi _42564__379 (.L_HI(net379));
 sg13g2_tiehi _41944__380 (.L_HI(net380));
 sg13g2_tiehi _42263__381 (.L_HI(net381));
 sg13g2_tiehi _41943__382 (.L_HI(net382));
 sg13g2_tiehi _42563__383 (.L_HI(net383));
 sg13g2_tiehi _41942__384 (.L_HI(net384));
 sg13g2_tiehi _42262__385 (.L_HI(net385));
 sg13g2_tiehi _41941__386 (.L_HI(net386));
 sg13g2_tiehi _42562__387 (.L_HI(net387));
 sg13g2_tiehi _41940__388 (.L_HI(net388));
 sg13g2_tiehi _42261__389 (.L_HI(net389));
 sg13g2_tiehi _41939__390 (.L_HI(net390));
 sg13g2_tiehi _42561__391 (.L_HI(net391));
 sg13g2_tiehi _41938__392 (.L_HI(net392));
 sg13g2_tiehi _42260__393 (.L_HI(net393));
 sg13g2_tiehi _41937__394 (.L_HI(net394));
 sg13g2_tiehi _42560__395 (.L_HI(net395));
 sg13g2_tiehi _41936__396 (.L_HI(net396));
 sg13g2_tiehi _42259__397 (.L_HI(net397));
 sg13g2_tiehi _41935__398 (.L_HI(net398));
 sg13g2_tiehi _42559__399 (.L_HI(net399));
 sg13g2_tiehi _41934__400 (.L_HI(net400));
 sg13g2_tiehi _42258__401 (.L_HI(net401));
 sg13g2_tiehi _41933__402 (.L_HI(net402));
 sg13g2_tiehi _42558__403 (.L_HI(net403));
 sg13g2_tiehi _41932__404 (.L_HI(net404));
 sg13g2_tiehi _42257__405 (.L_HI(net405));
 sg13g2_tiehi _41931__406 (.L_HI(net406));
 sg13g2_tiehi _42557__407 (.L_HI(net407));
 sg13g2_tiehi _41930__408 (.L_HI(net408));
 sg13g2_tiehi _42256__409 (.L_HI(net409));
 sg13g2_tiehi _41929__410 (.L_HI(net410));
 sg13g2_tiehi _42556__411 (.L_HI(net411));
 sg13g2_tiehi _41928__412 (.L_HI(net412));
 sg13g2_tiehi _42255__413 (.L_HI(net413));
 sg13g2_tiehi _41927__414 (.L_HI(net414));
 sg13g2_tiehi _42555__415 (.L_HI(net415));
 sg13g2_tiehi _41926__416 (.L_HI(net416));
 sg13g2_tiehi _42254__417 (.L_HI(net417));
 sg13g2_tiehi _41925__418 (.L_HI(net418));
 sg13g2_tiehi _42554__419 (.L_HI(net419));
 sg13g2_tiehi _41924__420 (.L_HI(net420));
 sg13g2_tiehi _42253__421 (.L_HI(net421));
 sg13g2_tiehi _41923__422 (.L_HI(net422));
 sg13g2_tiehi _42553__423 (.L_HI(net423));
 sg13g2_tiehi _41922__424 (.L_HI(net424));
 sg13g2_tiehi _42252__425 (.L_HI(net425));
 sg13g2_tiehi _41921__426 (.L_HI(net426));
 sg13g2_tiehi _42552__427 (.L_HI(net427));
 sg13g2_tiehi _41920__428 (.L_HI(net428));
 sg13g2_tiehi _42251__429 (.L_HI(net429));
 sg13g2_tiehi _41919__430 (.L_HI(net430));
 sg13g2_tiehi _42551__431 (.L_HI(net431));
 sg13g2_tiehi _41918__432 (.L_HI(net432));
 sg13g2_tiehi _42250__433 (.L_HI(net433));
 sg13g2_tiehi _41917__434 (.L_HI(net434));
 sg13g2_tiehi _41916__435 (.L_HI(net435));
 sg13g2_tiehi _42249__436 (.L_HI(net436));
 sg13g2_tiehi _41915__437 (.L_HI(net437));
 sg13g2_tiehi _41914__438 (.L_HI(net438));
 sg13g2_tiehi _42248__439 (.L_HI(net439));
 sg13g2_tiehi _41913__440 (.L_HI(net440));
 sg13g2_tiehi _41912__441 (.L_HI(net441));
 sg13g2_tiehi _42247__442 (.L_HI(net442));
 sg13g2_tiehi _41911__443 (.L_HI(net443));
 sg13g2_tiehi _41910__444 (.L_HI(net444));
 sg13g2_tiehi _42246__445 (.L_HI(net445));
 sg13g2_tiehi _41909__446 (.L_HI(net446));
 sg13g2_tiehi _41908__447 (.L_HI(net447));
 sg13g2_tiehi _42245__448 (.L_HI(net448));
 sg13g2_tiehi _41907__449 (.L_HI(net449));
 sg13g2_tiehi _41906__450 (.L_HI(net450));
 sg13g2_tiehi _42244__451 (.L_HI(net451));
 sg13g2_tiehi _41905__452 (.L_HI(net452));
 sg13g2_tiehi _41904__453 (.L_HI(net453));
 sg13g2_tiehi _42243__454 (.L_HI(net454));
 sg13g2_tiehi _41903__455 (.L_HI(net455));
 sg13g2_tiehi _41902__456 (.L_HI(net456));
 sg13g2_tiehi _42242__457 (.L_HI(net457));
 sg13g2_tiehi _41901__458 (.L_HI(net458));
 sg13g2_tiehi _41900__459 (.L_HI(net459));
 sg13g2_tiehi _42241__460 (.L_HI(net460));
 sg13g2_tiehi _41899__461 (.L_HI(net461));
 sg13g2_tiehi _41898__462 (.L_HI(net462));
 sg13g2_tiehi _42240__463 (.L_HI(net463));
 sg13g2_tiehi _41897__464 (.L_HI(net464));
 sg13g2_tiehi _41896__465 (.L_HI(net465));
 sg13g2_tiehi _42239__466 (.L_HI(net466));
 sg13g2_tiehi _41895__467 (.L_HI(net467));
 sg13g2_tiehi _41894__468 (.L_HI(net468));
 sg13g2_tiehi _42238__469 (.L_HI(net469));
 sg13g2_tiehi _41893__470 (.L_HI(net470));
 sg13g2_tiehi _41892__471 (.L_HI(net471));
 sg13g2_tiehi _42237__472 (.L_HI(net472));
 sg13g2_tiehi _41891__473 (.L_HI(net473));
 sg13g2_tiehi _41890__474 (.L_HI(net474));
 sg13g2_tiehi _42236__475 (.L_HI(net475));
 sg13g2_tiehi _41889__476 (.L_HI(net476));
 sg13g2_tiehi _41888__477 (.L_HI(net477));
 sg13g2_tiehi _42235__478 (.L_HI(net478));
 sg13g2_tiehi _41887__479 (.L_HI(net479));
 sg13g2_tiehi _41886__480 (.L_HI(net480));
 sg13g2_tiehi _42234__481 (.L_HI(net481));
 sg13g2_tiehi _41885__482 (.L_HI(net482));
 sg13g2_tiehi _41884__483 (.L_HI(net483));
 sg13g2_tiehi _42233__484 (.L_HI(net484));
 sg13g2_tiehi _41883__485 (.L_HI(net485));
 sg13g2_tiehi _41882__486 (.L_HI(net486));
 sg13g2_tiehi _42232__487 (.L_HI(net487));
 sg13g2_tiehi _41881__488 (.L_HI(net488));
 sg13g2_tiehi _41880__489 (.L_HI(net489));
 sg13g2_tiehi _42231__490 (.L_HI(net490));
 sg13g2_tiehi _41879__491 (.L_HI(net491));
 sg13g2_tiehi _41878__492 (.L_HI(net492));
 sg13g2_tiehi _42230__493 (.L_HI(net493));
 sg13g2_tiehi _41877__494 (.L_HI(net494));
 sg13g2_tiehi _41876__495 (.L_HI(net495));
 sg13g2_tiehi _42229__496 (.L_HI(net496));
 sg13g2_tiehi _41875__497 (.L_HI(net497));
 sg13g2_tiehi _41874__498 (.L_HI(net498));
 sg13g2_tiehi _42228__499 (.L_HI(net499));
 sg13g2_tiehi _41873__500 (.L_HI(net500));
 sg13g2_tiehi _41872__501 (.L_HI(net501));
 sg13g2_tiehi _42227__502 (.L_HI(net502));
 sg13g2_tiehi _41871__503 (.L_HI(net503));
 sg13g2_tiehi _41870__504 (.L_HI(net504));
 sg13g2_tiehi _42226__505 (.L_HI(net505));
 sg13g2_tiehi _41869__506 (.L_HI(net506));
 sg13g2_tiehi _41868__507 (.L_HI(net507));
 sg13g2_tiehi _42225__508 (.L_HI(net508));
 sg13g2_tiehi _41867__509 (.L_HI(net509));
 sg13g2_tiehi _41866__510 (.L_HI(net510));
 sg13g2_tiehi _42224__511 (.L_HI(net511));
 sg13g2_tiehi _41865__512 (.L_HI(net512));
 sg13g2_tiehi _41864__513 (.L_HI(net513));
 sg13g2_tiehi _42223__514 (.L_HI(net514));
 sg13g2_tiehi _41863__515 (.L_HI(net515));
 sg13g2_tiehi _41862__516 (.L_HI(net516));
 sg13g2_tiehi _42222__517 (.L_HI(net517));
 sg13g2_tiehi _41861__518 (.L_HI(net518));
 sg13g2_tiehi _41860__519 (.L_HI(net519));
 sg13g2_tiehi _42221__520 (.L_HI(net520));
 sg13g2_tiehi _41859__521 (.L_HI(net521));
 sg13g2_tiehi _41858__522 (.L_HI(net522));
 sg13g2_tiehi _42220__523 (.L_HI(net523));
 sg13g2_tiehi _41857__524 (.L_HI(net524));
 sg13g2_tiehi _41856__525 (.L_HI(net525));
 sg13g2_tiehi _42219__526 (.L_HI(net526));
 sg13g2_tiehi _41855__527 (.L_HI(net527));
 sg13g2_tiehi _41854__528 (.L_HI(net528));
 sg13g2_tiehi _42218__529 (.L_HI(net529));
 sg13g2_tiehi _41853__530 (.L_HI(net530));
 sg13g2_tiehi _41852__531 (.L_HI(net531));
 sg13g2_tiehi _42217__532 (.L_HI(net532));
 sg13g2_tiehi _41851__533 (.L_HI(net533));
 sg13g2_tiehi _41850__534 (.L_HI(net534));
 sg13g2_tiehi _42216__535 (.L_HI(net535));
 sg13g2_tiehi _41849__536 (.L_HI(net536));
 sg13g2_tiehi _41848__537 (.L_HI(net537));
 sg13g2_tiehi _42215__538 (.L_HI(net538));
 sg13g2_tiehi _41847__539 (.L_HI(net539));
 sg13g2_tiehi _41846__540 (.L_HI(net540));
 sg13g2_tiehi _42214__541 (.L_HI(net541));
 sg13g2_tiehi _41845__542 (.L_HI(net542));
 sg13g2_tiehi _41844__543 (.L_HI(net543));
 sg13g2_tiehi _42213__544 (.L_HI(net544));
 sg13g2_tiehi _41843__545 (.L_HI(net545));
 sg13g2_tiehi _41842__546 (.L_HI(net546));
 sg13g2_tiehi _42212__547 (.L_HI(net547));
 sg13g2_tiehi _41841__548 (.L_HI(net548));
 sg13g2_tiehi _41840__549 (.L_HI(net549));
 sg13g2_tiehi _42211__550 (.L_HI(net550));
 sg13g2_tiehi _41839__551 (.L_HI(net551));
 sg13g2_tiehi _41838__552 (.L_HI(net552));
 sg13g2_tiehi _42210__553 (.L_HI(net553));
 sg13g2_tiehi _41837__554 (.L_HI(net554));
 sg13g2_tiehi _41836__555 (.L_HI(net555));
 sg13g2_tiehi _42209__556 (.L_HI(net556));
 sg13g2_tiehi _41835__557 (.L_HI(net557));
 sg13g2_tiehi _41834__558 (.L_HI(net558));
 sg13g2_tiehi _42208__559 (.L_HI(net559));
 sg13g2_tiehi _41833__560 (.L_HI(net560));
 sg13g2_tiehi _41832__561 (.L_HI(net561));
 sg13g2_tiehi _42207__562 (.L_HI(net562));
 sg13g2_tiehi _41831__563 (.L_HI(net563));
 sg13g2_tiehi _41830__564 (.L_HI(net564));
 sg13g2_tiehi _42206__565 (.L_HI(net565));
 sg13g2_tiehi _41829__566 (.L_HI(net566));
 sg13g2_tiehi _41828__567 (.L_HI(net567));
 sg13g2_tiehi _42205__568 (.L_HI(net568));
 sg13g2_tiehi _41827__569 (.L_HI(net569));
 sg13g2_tiehi _41826__570 (.L_HI(net570));
 sg13g2_tiehi _42204__571 (.L_HI(net571));
 sg13g2_tiehi _41825__572 (.L_HI(net572));
 sg13g2_tiehi _41824__573 (.L_HI(net573));
 sg13g2_tiehi _42203__574 (.L_HI(net574));
 sg13g2_tiehi _41823__575 (.L_HI(net575));
 sg13g2_tiehi _41822__576 (.L_HI(net576));
 sg13g2_tiehi _42202__577 (.L_HI(net577));
 sg13g2_tiehi _41821__578 (.L_HI(net578));
 sg13g2_tiehi _41820__579 (.L_HI(net579));
 sg13g2_tiehi _42201__580 (.L_HI(net580));
 sg13g2_tiehi _41819__581 (.L_HI(net581));
 sg13g2_tiehi _41818__582 (.L_HI(net582));
 sg13g2_tiehi _42200__583 (.L_HI(net583));
 sg13g2_tiehi _41817__584 (.L_HI(net584));
 sg13g2_tiehi _41816__585 (.L_HI(net585));
 sg13g2_tiehi _42199__586 (.L_HI(net586));
 sg13g2_tiehi _41815__587 (.L_HI(net587));
 sg13g2_tiehi _41814__588 (.L_HI(net588));
 sg13g2_tiehi _42198__589 (.L_HI(net589));
 sg13g2_tiehi _41813__590 (.L_HI(net590));
 sg13g2_tiehi _41812__591 (.L_HI(net591));
 sg13g2_tiehi _42197__592 (.L_HI(net592));
 sg13g2_tiehi _41811__593 (.L_HI(net593));
 sg13g2_tiehi _41810__594 (.L_HI(net594));
 sg13g2_tiehi _42196__595 (.L_HI(net595));
 sg13g2_tiehi _41809__596 (.L_HI(net596));
 sg13g2_tiehi _41808__597 (.L_HI(net597));
 sg13g2_tiehi _42195__598 (.L_HI(net598));
 sg13g2_tiehi _41807__599 (.L_HI(net599));
 sg13g2_tiehi _41806__600 (.L_HI(net600));
 sg13g2_tiehi _42194__601 (.L_HI(net601));
 sg13g2_tiehi _41805__602 (.L_HI(net602));
 sg13g2_tiehi _41804__603 (.L_HI(net603));
 sg13g2_tiehi _42193__604 (.L_HI(net604));
 sg13g2_tiehi _41803__605 (.L_HI(net605));
 sg13g2_tiehi _41802__606 (.L_HI(net606));
 sg13g2_tiehi _42192__607 (.L_HI(net607));
 sg13g2_tiehi _41801__608 (.L_HI(net608));
 sg13g2_tiehi _41800__609 (.L_HI(net609));
 sg13g2_tiehi _42191__610 (.L_HI(net610));
 sg13g2_tiehi _41799__611 (.L_HI(net611));
 sg13g2_tiehi _41798__612 (.L_HI(net612));
 sg13g2_tiehi _42190__613 (.L_HI(net613));
 sg13g2_tiehi _41797__614 (.L_HI(net614));
 sg13g2_tiehi _41796__615 (.L_HI(net615));
 sg13g2_tiehi _42189__616 (.L_HI(net616));
 sg13g2_tiehi _41795__617 (.L_HI(net617));
 sg13g2_tiehi _41794__618 (.L_HI(net618));
 sg13g2_tiehi _42188__619 (.L_HI(net619));
 sg13g2_tiehi _41793__620 (.L_HI(net620));
 sg13g2_tiehi _41792__621 (.L_HI(net621));
 sg13g2_tiehi _42187__622 (.L_HI(net622));
 sg13g2_tiehi _41791__623 (.L_HI(net623));
 sg13g2_tiehi _41790__624 (.L_HI(net624));
 sg13g2_tiehi _42186__625 (.L_HI(net625));
 sg13g2_tiehi _41789__626 (.L_HI(net626));
 sg13g2_tiehi _41788__627 (.L_HI(net627));
 sg13g2_tiehi _42185__628 (.L_HI(net628));
 sg13g2_tiehi _41787__629 (.L_HI(net629));
 sg13g2_tiehi _41786__630 (.L_HI(net630));
 sg13g2_tiehi _42184__631 (.L_HI(net631));
 sg13g2_tiehi _41785__632 (.L_HI(net632));
 sg13g2_tiehi _41784__633 (.L_HI(net633));
 sg13g2_tiehi _42183__634 (.L_HI(net634));
 sg13g2_tiehi _41783__635 (.L_HI(net635));
 sg13g2_tiehi _41782__636 (.L_HI(net636));
 sg13g2_tiehi _42182__637 (.L_HI(net637));
 sg13g2_tiehi _41781__638 (.L_HI(net638));
 sg13g2_tiehi _41780__639 (.L_HI(net639));
 sg13g2_tiehi _42181__640 (.L_HI(net640));
 sg13g2_tiehi _41779__641 (.L_HI(net641));
 sg13g2_tiehi _41778__642 (.L_HI(net642));
 sg13g2_tiehi _42180__643 (.L_HI(net643));
 sg13g2_tiehi _41777__644 (.L_HI(net644));
 sg13g2_tiehi _41776__645 (.L_HI(net645));
 sg13g2_tiehi _42179__646 (.L_HI(net646));
 sg13g2_tiehi _41775__647 (.L_HI(net647));
 sg13g2_tiehi _41774__648 (.L_HI(net648));
 sg13g2_tiehi _42178__649 (.L_HI(net649));
 sg13g2_tiehi _41773__650 (.L_HI(net650));
 sg13g2_tiehi _41772__651 (.L_HI(net651));
 sg13g2_tiehi _42177__652 (.L_HI(net652));
 sg13g2_tiehi _41771__653 (.L_HI(net653));
 sg13g2_tiehi _41770__654 (.L_HI(net654));
 sg13g2_tiehi _42176__655 (.L_HI(net655));
 sg13g2_tiehi _41769__656 (.L_HI(net656));
 sg13g2_tiehi _41768__657 (.L_HI(net657));
 sg13g2_tiehi _42175__658 (.L_HI(net658));
 sg13g2_tiehi _41767__659 (.L_HI(net659));
 sg13g2_tiehi _41766__660 (.L_HI(net660));
 sg13g2_tiehi _42174__661 (.L_HI(net661));
 sg13g2_tiehi _41765__662 (.L_HI(net662));
 sg13g2_tiehi _41764__663 (.L_HI(net663));
 sg13g2_tiehi _42173__664 (.L_HI(net664));
 sg13g2_tiehi _41763__665 (.L_HI(net665));
 sg13g2_tiehi _41762__666 (.L_HI(net666));
 sg13g2_tiehi _42172__667 (.L_HI(net667));
 sg13g2_tiehi _41761__668 (.L_HI(net668));
 sg13g2_tiehi _41760__669 (.L_HI(net669));
 sg13g2_tiehi _42171__670 (.L_HI(net670));
 sg13g2_tiehi _41759__671 (.L_HI(net671));
 sg13g2_tiehi _41758__672 (.L_HI(net672));
 sg13g2_tiehi _42170__673 (.L_HI(net673));
 sg13g2_tiehi _41757__674 (.L_HI(net674));
 sg13g2_tiehi _41756__675 (.L_HI(net675));
 sg13g2_tiehi _42169__676 (.L_HI(net676));
 sg13g2_tiehi _41753__677 (.L_HI(net677));
 sg13g2_tiehi _42168__678 (.L_HI(net678));
 sg13g2_tiehi _41752__679 (.L_HI(net679));
 sg13g2_tiehi _41751__680 (.L_HI(net680));
 sg13g2_tiehi _42167__681 (.L_HI(net681));
 sg13g2_tiehi _41750__682 (.L_HI(net682));
 sg13g2_tiehi _41749__683 (.L_HI(net683));
 sg13g2_tiehi _42166__684 (.L_HI(net684));
 sg13g2_tiehi _41748__685 (.L_HI(net685));
 sg13g2_tiehi _41747__686 (.L_HI(net686));
 sg13g2_tiehi _42165__687 (.L_HI(net687));
 sg13g2_tiehi _41746__688 (.L_HI(net688));
 sg13g2_tiehi _41745__689 (.L_HI(net689));
 sg13g2_tiehi _42164__690 (.L_HI(net690));
 sg13g2_tiehi _41744__691 (.L_HI(net691));
 sg13g2_tiehi _41743__692 (.L_HI(net692));
 sg13g2_tiehi _42163__693 (.L_HI(net693));
 sg13g2_tiehi _41742__694 (.L_HI(net694));
 sg13g2_tiehi _41741__695 (.L_HI(net695));
 sg13g2_tiehi _42162__696 (.L_HI(net696));
 sg13g2_tiehi _41740__697 (.L_HI(net697));
 sg13g2_tiehi _41739__698 (.L_HI(net698));
 sg13g2_tiehi _42161__699 (.L_HI(net699));
 sg13g2_tiehi _41738__700 (.L_HI(net700));
 sg13g2_tiehi _41737__701 (.L_HI(net701));
 sg13g2_tiehi _42160__702 (.L_HI(net702));
 sg13g2_tiehi _41736__703 (.L_HI(net703));
 sg13g2_tiehi _41735__704 (.L_HI(net704));
 sg13g2_tiehi _42159__705 (.L_HI(net705));
 sg13g2_tiehi _41734__706 (.L_HI(net706));
 sg13g2_tiehi _41733__707 (.L_HI(net707));
 sg13g2_tiehi _42158__708 (.L_HI(net708));
 sg13g2_tiehi _41732__709 (.L_HI(net709));
 sg13g2_tiehi _41731__710 (.L_HI(net710));
 sg13g2_tiehi _42157__711 (.L_HI(net711));
 sg13g2_tiehi _41730__712 (.L_HI(net712));
 sg13g2_tiehi _41729__713 (.L_HI(net713));
 sg13g2_tiehi _42156__714 (.L_HI(net714));
 sg13g2_tiehi _41728__715 (.L_HI(net715));
 sg13g2_tiehi _41727__716 (.L_HI(net716));
 sg13g2_tiehi _42155__717 (.L_HI(net717));
 sg13g2_tiehi _41726__718 (.L_HI(net718));
 sg13g2_tiehi _41725__719 (.L_HI(net719));
 sg13g2_tiehi _42154__720 (.L_HI(net720));
 sg13g2_tiehi _41724__721 (.L_HI(net721));
 sg13g2_tiehi _41723__722 (.L_HI(net722));
 sg13g2_tiehi _42153__723 (.L_HI(net723));
 sg13g2_tiehi _41722__724 (.L_HI(net724));
 sg13g2_tiehi _41721__725 (.L_HI(net725));
 sg13g2_tiehi _42152__726 (.L_HI(net726));
 sg13g2_tiehi _41720__727 (.L_HI(net727));
 sg13g2_tiehi _41719__728 (.L_HI(net728));
 sg13g2_tiehi _42151__729 (.L_HI(net729));
 sg13g2_tiehi _41718__730 (.L_HI(net730));
 sg13g2_tiehi _41717__731 (.L_HI(net731));
 sg13g2_tiehi _42150__732 (.L_HI(net732));
 sg13g2_tiehi _41716__733 (.L_HI(net733));
 sg13g2_tiehi _41715__734 (.L_HI(net734));
 sg13g2_tiehi _42149__735 (.L_HI(net735));
 sg13g2_tiehi _41714__736 (.L_HI(net736));
 sg13g2_tiehi _41713__737 (.L_HI(net737));
 sg13g2_tiehi _42148__738 (.L_HI(net738));
 sg13g2_tiehi _41712__739 (.L_HI(net739));
 sg13g2_tiehi _41711__740 (.L_HI(net740));
 sg13g2_tiehi _42147__741 (.L_HI(net741));
 sg13g2_tiehi _41710__742 (.L_HI(net742));
 sg13g2_tiehi _41709__743 (.L_HI(net743));
 sg13g2_tiehi _42146__744 (.L_HI(net744));
 sg13g2_tiehi _41708__745 (.L_HI(net745));
 sg13g2_tiehi _41707__746 (.L_HI(net746));
 sg13g2_tiehi _42145__747 (.L_HI(net747));
 sg13g2_tiehi _41706__748 (.L_HI(net748));
 sg13g2_tiehi _41705__749 (.L_HI(net749));
 sg13g2_tiehi _42144__750 (.L_HI(net750));
 sg13g2_tiehi _41704__751 (.L_HI(net751));
 sg13g2_tiehi _41754__752 (.L_HI(net752));
 sg13g2_tiehi _41703__753 (.L_HI(net753));
 sg13g2_tiehi _42143__754 (.L_HI(net754));
 sg13g2_tiehi _41702__755 (.L_HI(net755));
 sg13g2_tiehi _41701__756 (.L_HI(net756));
 sg13g2_tiehi _42142__757 (.L_HI(net757));
 sg13g2_tiehi _41700__758 (.L_HI(net758));
 sg13g2_tiehi _41699__759 (.L_HI(net759));
 sg13g2_tiehi _42141__760 (.L_HI(net760));
 sg13g2_tiehi _41698__761 (.L_HI(net761));
 sg13g2_tiehi _41697__762 (.L_HI(net762));
 sg13g2_tiehi _42140__763 (.L_HI(net763));
 sg13g2_tiehi _41696__764 (.L_HI(net764));
 sg13g2_tiehi _41695__765 (.L_HI(net765));
 sg13g2_tiehi _42139__766 (.L_HI(net766));
 sg13g2_tiehi _41694__767 (.L_HI(net767));
 sg13g2_tiehi _41693__768 (.L_HI(net768));
 sg13g2_tiehi _42138__769 (.L_HI(net769));
 sg13g2_tiehi _41692__770 (.L_HI(net770));
 sg13g2_tiehi _41691__771 (.L_HI(net771));
 sg13g2_tiehi _42137__772 (.L_HI(net772));
 sg13g2_tiehi _41690__773 (.L_HI(net773));
 sg13g2_tiehi _41689__774 (.L_HI(net774));
 sg13g2_tiehi _42136__775 (.L_HI(net775));
 sg13g2_tiehi _41688__776 (.L_HI(net776));
 sg13g2_tiehi _41687__777 (.L_HI(net777));
 sg13g2_tiehi _42135__778 (.L_HI(net778));
 sg13g2_tiehi _41686__779 (.L_HI(net779));
 sg13g2_tiehi _41685__780 (.L_HI(net780));
 sg13g2_tiehi _42134__781 (.L_HI(net781));
 sg13g2_tiehi _41684__782 (.L_HI(net782));
 sg13g2_tiehi _41683__783 (.L_HI(net783));
 sg13g2_tiehi _42133__784 (.L_HI(net784));
 sg13g2_tiehi _41682__785 (.L_HI(net785));
 sg13g2_tiehi _41681__786 (.L_HI(net786));
 sg13g2_tiehi _42132__787 (.L_HI(net787));
 sg13g2_tiehi _41680__788 (.L_HI(net788));
 sg13g2_tiehi _41679__789 (.L_HI(net789));
 sg13g2_tiehi _42131__790 (.L_HI(net790));
 sg13g2_tiehi _41678__791 (.L_HI(net791));
 sg13g2_tiehi _41677__792 (.L_HI(net792));
 sg13g2_tiehi _42130__793 (.L_HI(net793));
 sg13g2_tiehi _41676__794 (.L_HI(net794));
 sg13g2_tiehi _41675__795 (.L_HI(net795));
 sg13g2_tiehi _42129__796 (.L_HI(net796));
 sg13g2_tiehi _41674__797 (.L_HI(net797));
 sg13g2_tiehi _41673__798 (.L_HI(net798));
 sg13g2_tiehi _42128__799 (.L_HI(net799));
 sg13g2_tiehi _41672__800 (.L_HI(net800));
 sg13g2_tiehi _41671__801 (.L_HI(net801));
 sg13g2_tiehi _42127__802 (.L_HI(net802));
 sg13g2_tiehi _41670__803 (.L_HI(net803));
 sg13g2_tiehi _41669__804 (.L_HI(net804));
 sg13g2_tiehi _42126__805 (.L_HI(net805));
 sg13g2_tiehi _41668__806 (.L_HI(net806));
 sg13g2_tiehi _41667__807 (.L_HI(net807));
 sg13g2_tiehi _42125__808 (.L_HI(net808));
 sg13g2_tiehi _41666__809 (.L_HI(net809));
 sg13g2_tiehi _41665__810 (.L_HI(net810));
 sg13g2_tiehi _42124__811 (.L_HI(net811));
 sg13g2_tiehi _41664__812 (.L_HI(net812));
 sg13g2_tiehi _41663__813 (.L_HI(net813));
 sg13g2_tiehi _42123__814 (.L_HI(net814));
 sg13g2_tiehi _41662__815 (.L_HI(net815));
 sg13g2_tiehi _41661__816 (.L_HI(net816));
 sg13g2_tiehi _42122__817 (.L_HI(net817));
 sg13g2_tiehi _41660__818 (.L_HI(net818));
 sg13g2_tiehi _41659__819 (.L_HI(net819));
 sg13g2_tiehi _42121__820 (.L_HI(net820));
 sg13g2_tiehi _41658__821 (.L_HI(net821));
 sg13g2_tiehi _41657__822 (.L_HI(net822));
 sg13g2_tiehi _42120__823 (.L_HI(net823));
 sg13g2_tiehi _41656__824 (.L_HI(net824));
 sg13g2_tiehi _41655__825 (.L_HI(net825));
 sg13g2_tiehi _42119__826 (.L_HI(net826));
 sg13g2_tiehi _41654__827 (.L_HI(net827));
 sg13g2_tiehi _41653__828 (.L_HI(net828));
 sg13g2_tiehi _42118__829 (.L_HI(net829));
 sg13g2_tiehi _41652__830 (.L_HI(net830));
 sg13g2_tiehi _41651__831 (.L_HI(net831));
 sg13g2_tiehi _42117__832 (.L_HI(net832));
 sg13g2_tiehi _41650__833 (.L_HI(net833));
 sg13g2_tiehi _41649__834 (.L_HI(net834));
 sg13g2_tiehi _42116__835 (.L_HI(net835));
 sg13g2_tiehi _41648__836 (.L_HI(net836));
 sg13g2_tiehi _41647__837 (.L_HI(net837));
 sg13g2_tiehi _42115__838 (.L_HI(net838));
 sg13g2_tiehi _41646__839 (.L_HI(net839));
 sg13g2_tiehi _41645__840 (.L_HI(net840));
 sg13g2_tiehi _42114__841 (.L_HI(net841));
 sg13g2_tiehi _41644__842 (.L_HI(net842));
 sg13g2_tiehi _41643__843 (.L_HI(net843));
 sg13g2_tiehi _42113__844 (.L_HI(net844));
 sg13g2_tiehi _41642__845 (.L_HI(net845));
 sg13g2_tiehi _41641__846 (.L_HI(net846));
 sg13g2_tiehi _42112__847 (.L_HI(net847));
 sg13g2_tiehi _41640__848 (.L_HI(net848));
 sg13g2_tiehi _41639__849 (.L_HI(net849));
 sg13g2_tiehi _42111__850 (.L_HI(net850));
 sg13g2_tiehi _41638__851 (.L_HI(net851));
 sg13g2_tiehi _41637__852 (.L_HI(net852));
 sg13g2_tiehi _42110__853 (.L_HI(net853));
 sg13g2_tiehi _41636__854 (.L_HI(net854));
 sg13g2_tiehi _41635__855 (.L_HI(net855));
 sg13g2_tiehi _42109__856 (.L_HI(net856));
 sg13g2_tiehi _41634__857 (.L_HI(net857));
 sg13g2_tiehi _41633__858 (.L_HI(net858));
 sg13g2_tiehi _42108__859 (.L_HI(net859));
 sg13g2_tiehi _41632__860 (.L_HI(net860));
 sg13g2_tiehi _41631__861 (.L_HI(net861));
 sg13g2_tiehi _42107__862 (.L_HI(net862));
 sg13g2_tiehi _41630__863 (.L_HI(net863));
 sg13g2_tiehi _41629__864 (.L_HI(net864));
 sg13g2_tiehi _42106__865 (.L_HI(net865));
 sg13g2_tiehi _41628__866 (.L_HI(net866));
 sg13g2_tiehi _41627__867 (.L_HI(net867));
 sg13g2_tiehi _42105__868 (.L_HI(net868));
 sg13g2_tiehi _41626__869 (.L_HI(net869));
 sg13g2_tiehi _41625__870 (.L_HI(net870));
 sg13g2_tiehi _42104__871 (.L_HI(net871));
 sg13g2_tiehi _41624__872 (.L_HI(net872));
 sg13g2_tiehi _41623__873 (.L_HI(net873));
 sg13g2_tiehi _42103__874 (.L_HI(net874));
 sg13g2_tiehi _41622__875 (.L_HI(net875));
 sg13g2_tiehi _41621__876 (.L_HI(net876));
 sg13g2_tiehi _42102__877 (.L_HI(net877));
 sg13g2_tiehi _41620__878 (.L_HI(net878));
 sg13g2_tiehi _41619__879 (.L_HI(net879));
 sg13g2_tiehi _42101__880 (.L_HI(net880));
 sg13g2_tiehi _41618__881 (.L_HI(net881));
 sg13g2_tiehi _41617__882 (.L_HI(net882));
 sg13g2_tiehi _42100__883 (.L_HI(net883));
 sg13g2_tiehi _41616__884 (.L_HI(net884));
 sg13g2_tiehi _41615__885 (.L_HI(net885));
 sg13g2_tiehi _42099__886 (.L_HI(net886));
 sg13g2_tiehi _41614__887 (.L_HI(net887));
 sg13g2_tiehi _41613__888 (.L_HI(net888));
 sg13g2_tiehi _42098__889 (.L_HI(net889));
 sg13g2_tiehi _41612__890 (.L_HI(net890));
 sg13g2_tiehi _41611__891 (.L_HI(net891));
 sg13g2_tiehi _42097__892 (.L_HI(net892));
 sg13g2_tiehi _41610__893 (.L_HI(net893));
 sg13g2_tiehi _41609__894 (.L_HI(net894));
 sg13g2_tiehi _42096__895 (.L_HI(net895));
 sg13g2_tiehi _41608__896 (.L_HI(net896));
 sg13g2_tiehi _41607__897 (.L_HI(net897));
 sg13g2_tiehi _42095__898 (.L_HI(net898));
 sg13g2_tiehi _41606__899 (.L_HI(net899));
 sg13g2_tiehi _41605__900 (.L_HI(net900));
 sg13g2_tiehi _42094__901 (.L_HI(net901));
 sg13g2_tiehi _41604__902 (.L_HI(net902));
 sg13g2_tiehi _41603__903 (.L_HI(net903));
 sg13g2_tiehi _42093__904 (.L_HI(net904));
 sg13g2_tiehi _41602__905 (.L_HI(net905));
 sg13g2_tiehi _41601__906 (.L_HI(net906));
 sg13g2_tiehi _42092__907 (.L_HI(net907));
 sg13g2_tiehi _41600__908 (.L_HI(net908));
 sg13g2_tiehi _41599__909 (.L_HI(net909));
 sg13g2_tiehi _42091__910 (.L_HI(net910));
 sg13g2_tiehi _41598__911 (.L_HI(net911));
 sg13g2_tiehi _41597__912 (.L_HI(net912));
 sg13g2_tiehi _42090__913 (.L_HI(net913));
 sg13g2_tiehi _41596__914 (.L_HI(net914));
 sg13g2_tiehi _41595__915 (.L_HI(net915));
 sg13g2_tiehi _42089__916 (.L_HI(net916));
 sg13g2_tiehi _41594__917 (.L_HI(net917));
 sg13g2_tiehi _41593__918 (.L_HI(net918));
 sg13g2_tiehi _42088__919 (.L_HI(net919));
 sg13g2_tiehi _41592__920 (.L_HI(net920));
 sg13g2_tiehi _41591__921 (.L_HI(net921));
 sg13g2_tiehi _42087__922 (.L_HI(net922));
 sg13g2_tiehi _41590__923 (.L_HI(net923));
 sg13g2_tiehi _41589__924 (.L_HI(net924));
 sg13g2_tiehi _42086__925 (.L_HI(net925));
 sg13g2_tiehi _41588__926 (.L_HI(net926));
 sg13g2_tiehi _41587__927 (.L_HI(net927));
 sg13g2_tiehi _42085__928 (.L_HI(net928));
 sg13g2_tiehi _41586__929 (.L_HI(net929));
 sg13g2_tiehi _41585__930 (.L_HI(net930));
 sg13g2_tiehi _42084__931 (.L_HI(net931));
 sg13g2_tiehi _41584__932 (.L_HI(net932));
 sg13g2_tiehi _41583__933 (.L_HI(net933));
 sg13g2_tiehi _42083__934 (.L_HI(net934));
 sg13g2_tiehi _41582__935 (.L_HI(net935));
 sg13g2_tiehi _41581__936 (.L_HI(net936));
 sg13g2_tiehi _42082__937 (.L_HI(net937));
 sg13g2_tiehi _41580__938 (.L_HI(net938));
 sg13g2_tiehi _41579__939 (.L_HI(net939));
 sg13g2_tiehi _42081__940 (.L_HI(net940));
 sg13g2_tiehi _41578__941 (.L_HI(net941));
 sg13g2_tiehi _41577__942 (.L_HI(net942));
 sg13g2_tiehi _42080__943 (.L_HI(net943));
 sg13g2_tiehi _41576__944 (.L_HI(net944));
 sg13g2_tiehi _41575__945 (.L_HI(net945));
 sg13g2_tiehi _42079__946 (.L_HI(net946));
 sg13g2_tiehi _41574__947 (.L_HI(net947));
 sg13g2_tiehi _41573__948 (.L_HI(net948));
 sg13g2_tiehi _42078__949 (.L_HI(net949));
 sg13g2_tiehi _41572__950 (.L_HI(net950));
 sg13g2_tiehi _41571__951 (.L_HI(net951));
 sg13g2_tiehi _42077__952 (.L_HI(net952));
 sg13g2_tiehi _41570__953 (.L_HI(net953));
 sg13g2_tiehi _41569__954 (.L_HI(net954));
 sg13g2_tiehi _42076__955 (.L_HI(net955));
 sg13g2_tiehi _41568__956 (.L_HI(net956));
 sg13g2_tiehi _41567__957 (.L_HI(net957));
 sg13g2_tiehi _42075__958 (.L_HI(net958));
 sg13g2_tiehi _41566__959 (.L_HI(net959));
 sg13g2_tiehi _41565__960 (.L_HI(net960));
 sg13g2_tiehi _42074__961 (.L_HI(net961));
 sg13g2_tiehi _41564__962 (.L_HI(net962));
 sg13g2_tiehi _41563__963 (.L_HI(net963));
 sg13g2_tiehi _42073__964 (.L_HI(net964));
 sg13g2_tiehi _41562__965 (.L_HI(net965));
 sg13g2_tiehi _41561__966 (.L_HI(net966));
 sg13g2_tiehi _42072__967 (.L_HI(net967));
 sg13g2_tiehi _41560__968 (.L_HI(net968));
 sg13g2_tiehi _41559__969 (.L_HI(net969));
 sg13g2_tiehi _42071__970 (.L_HI(net970));
 sg13g2_tiehi _41558__971 (.L_HI(net971));
 sg13g2_tiehi _41557__972 (.L_HI(net972));
 sg13g2_tiehi _42070__973 (.L_HI(net973));
 sg13g2_tiehi _41556__974 (.L_HI(net974));
 sg13g2_tiehi _41555__975 (.L_HI(net975));
 sg13g2_tiehi _42069__976 (.L_HI(net976));
 sg13g2_tiehi _41554__977 (.L_HI(net977));
 sg13g2_tiehi _41553__978 (.L_HI(net978));
 sg13g2_tiehi _42068__979 (.L_HI(net979));
 sg13g2_tiehi _41552__980 (.L_HI(net980));
 sg13g2_tiehi _41551__981 (.L_HI(net981));
 sg13g2_tiehi _42067__982 (.L_HI(net982));
 sg13g2_tiehi _41550__983 (.L_HI(net983));
 sg13g2_tiehi _41549__984 (.L_HI(net984));
 sg13g2_tiehi _42066__985 (.L_HI(net985));
 sg13g2_tiehi _41548__986 (.L_HI(net986));
 sg13g2_tiehi _41547__987 (.L_HI(net987));
 sg13g2_tiehi _42065__988 (.L_HI(net988));
 sg13g2_tiehi _41546__989 (.L_HI(net989));
 sg13g2_tiehi _41545__990 (.L_HI(net990));
 sg13g2_tiehi _42064__991 (.L_HI(net991));
 sg13g2_tiehi _41544__992 (.L_HI(net992));
 sg13g2_tiehi _41543__993 (.L_HI(net993));
 sg13g2_tiehi _42063__994 (.L_HI(net994));
 sg13g2_tiehi _41542__995 (.L_HI(net995));
 sg13g2_tiehi _41541__996 (.L_HI(net996));
 sg13g2_tiehi _42062__997 (.L_HI(net997));
 sg13g2_tiehi _41540__998 (.L_HI(net998));
 sg13g2_tiehi _41539__999 (.L_HI(net999));
 sg13g2_tiehi _42061__1000 (.L_HI(net1000));
 sg13g2_tiehi _41538__1001 (.L_HI(net1001));
 sg13g2_tiehi _41537__1002 (.L_HI(net1002));
 sg13g2_tiehi _42060__1003 (.L_HI(net1003));
 sg13g2_tiehi _41536__1004 (.L_HI(net1004));
 sg13g2_tiehi _41535__1005 (.L_HI(net1005));
 sg13g2_tiehi _42059__1006 (.L_HI(net1006));
 sg13g2_tiehi _41534__1007 (.L_HI(net1007));
 sg13g2_tiehi _41533__1008 (.L_HI(net1008));
 sg13g2_tiehi _42058__1009 (.L_HI(net1009));
 sg13g2_tiehi _41532__1010 (.L_HI(net1010));
 sg13g2_tiehi _41531__1011 (.L_HI(net1011));
 sg13g2_tiehi _42057__1012 (.L_HI(net1012));
 sg13g2_tiehi _41530__1013 (.L_HI(net1013));
 sg13g2_tiehi _41529__1014 (.L_HI(net1014));
 sg13g2_tiehi _42056__1015 (.L_HI(net1015));
 sg13g2_tiehi _41528__1016 (.L_HI(net1016));
 sg13g2_tiehi _41527__1017 (.L_HI(net1017));
 sg13g2_tiehi _42055__1018 (.L_HI(net1018));
 sg13g2_tiehi _41526__1019 (.L_HI(net1019));
 sg13g2_tiehi _41525__1020 (.L_HI(net1020));
 sg13g2_tiehi _42054__1021 (.L_HI(net1021));
 sg13g2_tiehi _41524__1022 (.L_HI(net1022));
 sg13g2_tiehi _41523__1023 (.L_HI(net1023));
 sg13g2_tiehi _42053__1024 (.L_HI(net1024));
 sg13g2_tiehi _41522__1025 (.L_HI(net1025));
 sg13g2_tiehi _41521__1026 (.L_HI(net1026));
 sg13g2_tiehi _42052__1027 (.L_HI(net1027));
 sg13g2_tiehi _41520__1028 (.L_HI(net1028));
 sg13g2_tiehi _41519__1029 (.L_HI(net1029));
 sg13g2_tiehi _42051__1030 (.L_HI(net1030));
 sg13g2_tiehi _41518__1031 (.L_HI(net1031));
 sg13g2_tiehi _41517__1032 (.L_HI(net1032));
 sg13g2_tiehi _42050__1033 (.L_HI(net1033));
 sg13g2_tiehi _41516__1034 (.L_HI(net1034));
 sg13g2_tiehi _41515__1035 (.L_HI(net1035));
 sg13g2_tiehi _42049__1036 (.L_HI(net1036));
 sg13g2_tiehi _41514__1037 (.L_HI(net1037));
 sg13g2_tiehi _41513__1038 (.L_HI(net1038));
 sg13g2_tiehi _42048__1039 (.L_HI(net1039));
 sg13g2_tiehi _41512__1040 (.L_HI(net1040));
 sg13g2_tiehi _41511__1041 (.L_HI(net1041));
 sg13g2_tiehi _42047__1042 (.L_HI(net1042));
 sg13g2_tiehi _41510__1043 (.L_HI(net1043));
 sg13g2_tiehi _41509__1044 (.L_HI(net1044));
 sg13g2_tiehi _42046__1045 (.L_HI(net1045));
 sg13g2_tiehi _41508__1046 (.L_HI(net1046));
 sg13g2_tiehi _41507__1047 (.L_HI(net1047));
 sg13g2_tiehi _42045__1048 (.L_HI(net1048));
 sg13g2_tiehi _41506__1049 (.L_HI(net1049));
 sg13g2_tiehi _41505__1050 (.L_HI(net1050));
 sg13g2_tiehi _42044__1051 (.L_HI(net1051));
 sg13g2_tiehi _41504__1052 (.L_HI(net1052));
 sg13g2_tiehi _41503__1053 (.L_HI(net1053));
 sg13g2_tiehi _42043__1054 (.L_HI(net1054));
 sg13g2_tiehi _41502__1055 (.L_HI(net1055));
 sg13g2_tiehi _41501__1056 (.L_HI(net1056));
 sg13g2_tiehi _42042__1057 (.L_HI(net1057));
 sg13g2_tiehi _41500__1058 (.L_HI(net1058));
 sg13g2_tiehi _41499__1059 (.L_HI(net1059));
 sg13g2_tiehi _42041__1060 (.L_HI(net1060));
 sg13g2_tiehi _41498__1061 (.L_HI(net1061));
 sg13g2_tiehi tt_um_corey_1062 (.L_HI(net1062));
 sg13g2_tiehi tt_um_corey_1063 (.L_HI(net1063));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_corey_13 (.L_LO(net13));
 sg13g2_tielo tt_um_corey_14 (.L_LO(net14));
 sg13g2_tielo tt_um_corey_15 (.L_LO(net15));
 sg13g2_tielo tt_um_corey_16 (.L_LO(net16));
 sg13g2_tielo tt_um_corey_17 (.L_LO(net17));
 sg13g2_tielo tt_um_corey_18 (.L_LO(net18));
 sg13g2_tielo tt_um_corey_19 (.L_LO(net19));
 sg13g2_tielo tt_um_corey_20 (.L_LO(net20));
 sg13g2_tielo tt_um_corey_21 (.L_LO(net21));
 sg13g2_tielo tt_um_corey_22 (.L_LO(net22));
 sg13g2_tielo tt_um_corey_23 (.L_LO(net23));
 sg13g2_tiehi _41232__24 (.L_HI(net24));
 sg13g2_buf_1 _43633_ (.A(accepting),
    .X(uio_out[0]));
 sg13g2_buf_1 _43634_ (.A(\shift_reg[264] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _43635_ (.A(\shift_reg[265] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _43636_ (.A(\shift_reg[266] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _43637_ (.A(\shift_reg[267] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _43638_ (.A(\shift_reg[268] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _43639_ (.A(\shift_reg[269] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _43640_ (.A(\shift_reg[270] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _43641_ (.A(\shift_reg[271] ),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout4032 (.A(net4033),
    .X(net4032));
 sg13g2_buf_8 fanout4033 (.A(net4034),
    .X(net4033));
 sg13g2_buf_8 fanout4034 (.A(net4054),
    .X(net4034));
 sg13g2_buf_8 fanout4035 (.A(net4037),
    .X(net4035));
 sg13g2_buf_1 fanout4036 (.A(net4037),
    .X(net4036));
 sg13g2_buf_8 fanout4037 (.A(net4054),
    .X(net4037));
 sg13g2_buf_8 fanout4038 (.A(net4040),
    .X(net4038));
 sg13g2_buf_2 fanout4039 (.A(net4040),
    .X(net4039));
 sg13g2_buf_8 fanout4040 (.A(net4054),
    .X(net4040));
 sg13g2_buf_8 fanout4041 (.A(net4053),
    .X(net4041));
 sg13g2_buf_1 fanout4042 (.A(net4043),
    .X(net4042));
 sg13g2_buf_8 fanout4043 (.A(net4053),
    .X(net4043));
 sg13g2_buf_8 fanout4044 (.A(net4046),
    .X(net4044));
 sg13g2_buf_1 fanout4045 (.A(net4046),
    .X(net4045));
 sg13g2_buf_8 fanout4046 (.A(net4053),
    .X(net4046));
 sg13g2_buf_8 fanout4047 (.A(net4049),
    .X(net4047));
 sg13g2_buf_2 fanout4048 (.A(net4049),
    .X(net4048));
 sg13g2_buf_8 fanout4049 (.A(net4053),
    .X(net4049));
 sg13g2_buf_8 fanout4050 (.A(net4052),
    .X(net4050));
 sg13g2_buf_1 fanout4051 (.A(net4052),
    .X(net4051));
 sg13g2_buf_8 fanout4052 (.A(net4053),
    .X(net4052));
 sg13g2_buf_8 fanout4053 (.A(net4054),
    .X(net4053));
 sg13g2_buf_8 fanout4054 (.A(_13510_),
    .X(net4054));
 sg13g2_buf_8 fanout4055 (.A(net4056),
    .X(net4055));
 sg13g2_buf_8 fanout4056 (.A(net4060),
    .X(net4056));
 sg13g2_buf_8 fanout4057 (.A(net4059),
    .X(net4057));
 sg13g2_buf_8 fanout4058 (.A(net4060),
    .X(net4058));
 sg13g2_buf_2 fanout4059 (.A(net4060),
    .X(net4059));
 sg13g2_buf_8 fanout4060 (.A(net4074),
    .X(net4060));
 sg13g2_buf_8 fanout4061 (.A(net4062),
    .X(net4061));
 sg13g2_buf_8 fanout4062 (.A(net4074),
    .X(net4062));
 sg13g2_buf_8 fanout4063 (.A(net4064),
    .X(net4063));
 sg13g2_buf_8 fanout4064 (.A(net4074),
    .X(net4064));
 sg13g2_buf_8 fanout4065 (.A(net4066),
    .X(net4065));
 sg13g2_buf_8 fanout4066 (.A(net4074),
    .X(net4066));
 sg13g2_buf_8 fanout4067 (.A(net4068),
    .X(net4067));
 sg13g2_buf_8 fanout4068 (.A(net4074),
    .X(net4068));
 sg13g2_buf_8 fanout4069 (.A(net4070),
    .X(net4069));
 sg13g2_buf_1 fanout4070 (.A(net4073),
    .X(net4070));
 sg13g2_buf_8 fanout4071 (.A(net4072),
    .X(net4071));
 sg13g2_buf_8 fanout4072 (.A(net4073),
    .X(net4072));
 sg13g2_buf_8 fanout4073 (.A(net4074),
    .X(net4073));
 sg13g2_buf_8 fanout4074 (.A(_13510_),
    .X(net4074));
 sg13g2_buf_8 fanout4075 (.A(net4078),
    .X(net4075));
 sg13g2_buf_1 fanout4076 (.A(net4078),
    .X(net4076));
 sg13g2_buf_8 fanout4077 (.A(net4078),
    .X(net4077));
 sg13g2_buf_8 fanout4078 (.A(net4081),
    .X(net4078));
 sg13g2_buf_8 fanout4079 (.A(net4080),
    .X(net4079));
 sg13g2_buf_8 fanout4080 (.A(net4081),
    .X(net4080));
 sg13g2_buf_8 fanout4081 (.A(net4096),
    .X(net4081));
 sg13g2_buf_8 fanout4082 (.A(net4084),
    .X(net4082));
 sg13g2_buf_8 fanout4083 (.A(net4084),
    .X(net4083));
 sg13g2_buf_8 fanout4084 (.A(net4086),
    .X(net4084));
 sg13g2_buf_8 fanout4085 (.A(net4086),
    .X(net4085));
 sg13g2_buf_2 fanout4086 (.A(net4096),
    .X(net4086));
 sg13g2_buf_8 fanout4087 (.A(net4091),
    .X(net4087));
 sg13g2_buf_8 fanout4088 (.A(net4091),
    .X(net4088));
 sg13g2_buf_8 fanout4089 (.A(net4091),
    .X(net4089));
 sg13g2_buf_2 fanout4090 (.A(net4091),
    .X(net4090));
 sg13g2_buf_8 fanout4091 (.A(net4096),
    .X(net4091));
 sg13g2_buf_8 fanout4092 (.A(net4094),
    .X(net4092));
 sg13g2_buf_8 fanout4093 (.A(net4094),
    .X(net4093));
 sg13g2_buf_8 fanout4094 (.A(net4095),
    .X(net4094));
 sg13g2_buf_8 fanout4095 (.A(net4096),
    .X(net4095));
 sg13g2_buf_8 fanout4096 (.A(_13509_),
    .X(net4096));
 sg13g2_buf_8 fanout4097 (.A(net4098),
    .X(net4097));
 sg13g2_buf_8 fanout4098 (.A(net4102),
    .X(net4098));
 sg13g2_buf_8 fanout4099 (.A(net4102),
    .X(net4099));
 sg13g2_buf_8 fanout4100 (.A(net4102),
    .X(net4100));
 sg13g2_buf_8 fanout4101 (.A(net4102),
    .X(net4101));
 sg13g2_buf_8 fanout4102 (.A(net4121),
    .X(net4102));
 sg13g2_buf_8 fanout4103 (.A(net4108),
    .X(net4103));
 sg13g2_buf_1 fanout4104 (.A(net4108),
    .X(net4104));
 sg13g2_buf_8 fanout4105 (.A(net4107),
    .X(net4105));
 sg13g2_buf_1 fanout4106 (.A(net4108),
    .X(net4106));
 sg13g2_buf_8 fanout4107 (.A(net4108),
    .X(net4107));
 sg13g2_buf_8 fanout4108 (.A(net4121),
    .X(net4108));
 sg13g2_buf_8 fanout4109 (.A(net4110),
    .X(net4109));
 sg13g2_buf_8 fanout4110 (.A(net4115),
    .X(net4110));
 sg13g2_buf_8 fanout4111 (.A(net4115),
    .X(net4111));
 sg13g2_buf_1 fanout4112 (.A(net4115),
    .X(net4112));
 sg13g2_buf_8 fanout4113 (.A(net4114),
    .X(net4113));
 sg13g2_buf_1 fanout4114 (.A(net4115),
    .X(net4114));
 sg13g2_buf_8 fanout4115 (.A(net4121),
    .X(net4115));
 sg13g2_buf_8 fanout4116 (.A(net4118),
    .X(net4116));
 sg13g2_buf_8 fanout4117 (.A(net4118),
    .X(net4117));
 sg13g2_buf_8 fanout4118 (.A(net4121),
    .X(net4118));
 sg13g2_buf_8 fanout4119 (.A(net4120),
    .X(net4119));
 sg13g2_buf_8 fanout4120 (.A(net4121),
    .X(net4120));
 sg13g2_buf_8 fanout4121 (.A(_13509_),
    .X(net4121));
 sg13g2_buf_8 fanout4122 (.A(net4124),
    .X(net4122));
 sg13g2_buf_8 fanout4123 (.A(net4124),
    .X(net4123));
 sg13g2_buf_8 fanout4124 (.A(net4134),
    .X(net4124));
 sg13g2_buf_8 fanout4125 (.A(net4134),
    .X(net4125));
 sg13g2_buf_8 fanout4126 (.A(net4134),
    .X(net4126));
 sg13g2_buf_8 fanout4127 (.A(net4128),
    .X(net4127));
 sg13g2_buf_8 fanout4128 (.A(net4129),
    .X(net4128));
 sg13g2_buf_8 fanout4129 (.A(net4134),
    .X(net4129));
 sg13g2_buf_8 fanout4130 (.A(net4131),
    .X(net4130));
 sg13g2_buf_8 fanout4131 (.A(net4134),
    .X(net4131));
 sg13g2_buf_8 fanout4132 (.A(net4133),
    .X(net4132));
 sg13g2_buf_8 fanout4133 (.A(net4134),
    .X(net4133));
 sg13g2_buf_8 fanout4134 (.A(net4189),
    .X(net4134));
 sg13g2_buf_8 fanout4135 (.A(net4139),
    .X(net4135));
 sg13g2_buf_1 fanout4136 (.A(net4139),
    .X(net4136));
 sg13g2_buf_8 fanout4137 (.A(net4138),
    .X(net4137));
 sg13g2_buf_8 fanout4138 (.A(net4139),
    .X(net4138));
 sg13g2_buf_8 fanout4139 (.A(net4189),
    .X(net4139));
 sg13g2_buf_8 fanout4140 (.A(net4151),
    .X(net4140));
 sg13g2_buf_1 fanout4141 (.A(net4151),
    .X(net4141));
 sg13g2_buf_8 fanout4142 (.A(net4144),
    .X(net4142));
 sg13g2_buf_8 fanout4143 (.A(net4144),
    .X(net4143));
 sg13g2_buf_8 fanout4144 (.A(net4151),
    .X(net4144));
 sg13g2_buf_8 fanout4145 (.A(net4151),
    .X(net4145));
 sg13g2_buf_2 fanout4146 (.A(net4151),
    .X(net4146));
 sg13g2_buf_8 fanout4147 (.A(net4148),
    .X(net4147));
 sg13g2_buf_8 fanout4148 (.A(net4150),
    .X(net4148));
 sg13g2_buf_8 fanout4149 (.A(net4150),
    .X(net4149));
 sg13g2_buf_8 fanout4150 (.A(net4151),
    .X(net4150));
 sg13g2_buf_8 fanout4151 (.A(net4189),
    .X(net4151));
 sg13g2_buf_8 fanout4152 (.A(net4156),
    .X(net4152));
 sg13g2_buf_8 fanout4153 (.A(net4156),
    .X(net4153));
 sg13g2_buf_8 fanout4154 (.A(net4156),
    .X(net4154));
 sg13g2_buf_1 fanout4155 (.A(net4156),
    .X(net4155));
 sg13g2_buf_8 fanout4156 (.A(net4188),
    .X(net4156));
 sg13g2_buf_8 fanout4157 (.A(net4158),
    .X(net4157));
 sg13g2_buf_8 fanout4158 (.A(net4163),
    .X(net4158));
 sg13g2_buf_8 fanout4159 (.A(net4163),
    .X(net4159));
 sg13g2_buf_1 fanout4160 (.A(net4163),
    .X(net4160));
 sg13g2_buf_8 fanout4161 (.A(net4162),
    .X(net4161));
 sg13g2_buf_8 fanout4162 (.A(net4163),
    .X(net4162));
 sg13g2_buf_8 fanout4163 (.A(net4188),
    .X(net4163));
 sg13g2_buf_8 fanout4164 (.A(net4169),
    .X(net4164));
 sg13g2_buf_8 fanout4165 (.A(net4168),
    .X(net4165));
 sg13g2_buf_8 fanout4166 (.A(net4167),
    .X(net4166));
 sg13g2_buf_8 fanout4167 (.A(net4168),
    .X(net4167));
 sg13g2_buf_8 fanout4168 (.A(net4169),
    .X(net4168));
 sg13g2_buf_8 fanout4169 (.A(net4188),
    .X(net4169));
 sg13g2_buf_8 fanout4170 (.A(net4171),
    .X(net4170));
 sg13g2_buf_8 fanout4171 (.A(net4187),
    .X(net4171));
 sg13g2_buf_8 fanout4172 (.A(net4187),
    .X(net4172));
 sg13g2_buf_8 fanout4173 (.A(net4187),
    .X(net4173));
 sg13g2_buf_8 fanout4174 (.A(net4179),
    .X(net4174));
 sg13g2_buf_8 fanout4175 (.A(net4176),
    .X(net4175));
 sg13g2_buf_2 fanout4176 (.A(net4179),
    .X(net4176));
 sg13g2_buf_8 fanout4177 (.A(net4178),
    .X(net4177));
 sg13g2_buf_8 fanout4178 (.A(net4179),
    .X(net4178));
 sg13g2_buf_8 fanout4179 (.A(net4187),
    .X(net4179));
 sg13g2_buf_8 fanout4180 (.A(net4181),
    .X(net4180));
 sg13g2_buf_8 fanout4181 (.A(net4186),
    .X(net4181));
 sg13g2_buf_8 fanout4182 (.A(net4186),
    .X(net4182));
 sg13g2_buf_1 fanout4183 (.A(net4186),
    .X(net4183));
 sg13g2_buf_8 fanout4184 (.A(net4185),
    .X(net4184));
 sg13g2_buf_8 fanout4185 (.A(net4186),
    .X(net4185));
 sg13g2_buf_8 fanout4186 (.A(net4187),
    .X(net4186));
 sg13g2_buf_8 fanout4187 (.A(net4188),
    .X(net4187));
 sg13g2_buf_8 fanout4188 (.A(net4189),
    .X(net4188));
 sg13g2_buf_8 fanout4189 (.A(net4259),
    .X(net4189));
 sg13g2_buf_8 fanout4190 (.A(net4191),
    .X(net4190));
 sg13g2_buf_8 fanout4191 (.A(net4194),
    .X(net4191));
 sg13g2_buf_8 fanout4192 (.A(net4193),
    .X(net4192));
 sg13g2_buf_8 fanout4193 (.A(net4194),
    .X(net4193));
 sg13g2_buf_8 fanout4194 (.A(net4224),
    .X(net4194));
 sg13g2_buf_8 fanout4195 (.A(net4196),
    .X(net4195));
 sg13g2_buf_8 fanout4196 (.A(net4207),
    .X(net4196));
 sg13g2_buf_8 fanout4197 (.A(net4201),
    .X(net4197));
 sg13g2_buf_1 fanout4198 (.A(net4201),
    .X(net4198));
 sg13g2_buf_8 fanout4199 (.A(net4201),
    .X(net4199));
 sg13g2_buf_2 fanout4200 (.A(net4201),
    .X(net4200));
 sg13g2_buf_8 fanout4201 (.A(net4207),
    .X(net4201));
 sg13g2_buf_8 fanout4202 (.A(net4203),
    .X(net4202));
 sg13g2_buf_1 fanout4203 (.A(net4207),
    .X(net4203));
 sg13g2_buf_8 fanout4204 (.A(net4205),
    .X(net4204));
 sg13g2_buf_2 fanout4205 (.A(net4206),
    .X(net4205));
 sg13g2_buf_8 fanout4206 (.A(net4207),
    .X(net4206));
 sg13g2_buf_8 fanout4207 (.A(net4224),
    .X(net4207));
 sg13g2_buf_8 fanout4208 (.A(net4213),
    .X(net4208));
 sg13g2_buf_1 fanout4209 (.A(net4210),
    .X(net4209));
 sg13g2_buf_8 fanout4210 (.A(net4213),
    .X(net4210));
 sg13g2_buf_8 fanout4211 (.A(net4213),
    .X(net4211));
 sg13g2_buf_2 fanout4212 (.A(net4213),
    .X(net4212));
 sg13g2_buf_8 fanout4213 (.A(net4224),
    .X(net4213));
 sg13g2_buf_8 fanout4214 (.A(net4218),
    .X(net4214));
 sg13g2_buf_2 fanout4215 (.A(net4218),
    .X(net4215));
 sg13g2_buf_8 fanout4216 (.A(net4217),
    .X(net4216));
 sg13g2_buf_8 fanout4217 (.A(net4218),
    .X(net4217));
 sg13g2_buf_8 fanout4218 (.A(net4224),
    .X(net4218));
 sg13g2_buf_8 fanout4219 (.A(net4223),
    .X(net4219));
 sg13g2_buf_8 fanout4220 (.A(net4222),
    .X(net4220));
 sg13g2_buf_8 fanout4221 (.A(net4222),
    .X(net4221));
 sg13g2_buf_8 fanout4222 (.A(net4223),
    .X(net4222));
 sg13g2_buf_8 fanout4223 (.A(net4224),
    .X(net4223));
 sg13g2_buf_8 fanout4224 (.A(net4259),
    .X(net4224));
 sg13g2_buf_8 fanout4225 (.A(net4227),
    .X(net4225));
 sg13g2_buf_8 fanout4226 (.A(net4227),
    .X(net4226));
 sg13g2_buf_8 fanout4227 (.A(net4241),
    .X(net4227));
 sg13g2_buf_8 fanout4228 (.A(net4241),
    .X(net4228));
 sg13g2_buf_8 fanout4229 (.A(net4241),
    .X(net4229));
 sg13g2_buf_8 fanout4230 (.A(net4232),
    .X(net4230));
 sg13g2_buf_8 fanout4231 (.A(net4232),
    .X(net4231));
 sg13g2_buf_8 fanout4232 (.A(net4240),
    .X(net4232));
 sg13g2_buf_8 fanout4233 (.A(net4240),
    .X(net4233));
 sg13g2_buf_8 fanout4234 (.A(net4240),
    .X(net4234));
 sg13g2_buf_1 fanout4235 (.A(net4240),
    .X(net4235));
 sg13g2_buf_8 fanout4236 (.A(net4239),
    .X(net4236));
 sg13g2_buf_1 fanout4237 (.A(net4239),
    .X(net4237));
 sg13g2_buf_8 fanout4238 (.A(net4239),
    .X(net4238));
 sg13g2_buf_8 fanout4239 (.A(net4240),
    .X(net4239));
 sg13g2_buf_8 fanout4240 (.A(net4241),
    .X(net4240));
 sg13g2_buf_8 fanout4241 (.A(net4259),
    .X(net4241));
 sg13g2_buf_8 fanout4242 (.A(net4243),
    .X(net4242));
 sg13g2_buf_8 fanout4243 (.A(net4247),
    .X(net4243));
 sg13g2_buf_8 fanout4244 (.A(net4245),
    .X(net4244));
 sg13g2_buf_8 fanout4245 (.A(net4246),
    .X(net4245));
 sg13g2_buf_8 fanout4246 (.A(net4247),
    .X(net4246));
 sg13g2_buf_8 fanout4247 (.A(net4258),
    .X(net4247));
 sg13g2_buf_8 fanout4248 (.A(net4251),
    .X(net4248));
 sg13g2_buf_1 fanout4249 (.A(net4251),
    .X(net4249));
 sg13g2_buf_8 fanout4250 (.A(net4251),
    .X(net4250));
 sg13g2_buf_8 fanout4251 (.A(net4258),
    .X(net4251));
 sg13g2_buf_8 fanout4252 (.A(net4253),
    .X(net4252));
 sg13g2_buf_8 fanout4253 (.A(net4257),
    .X(net4253));
 sg13g2_buf_8 fanout4254 (.A(net4255),
    .X(net4254));
 sg13g2_buf_8 fanout4255 (.A(net4257),
    .X(net4255));
 sg13g2_buf_1 fanout4256 (.A(net4257),
    .X(net4256));
 sg13g2_buf_2 fanout4257 (.A(net4258),
    .X(net4257));
 sg13g2_buf_8 fanout4258 (.A(net4259),
    .X(net4258));
 sg13g2_buf_8 fanout4259 (.A(_19029_),
    .X(net4259));
 sg13g2_buf_8 fanout4260 (.A(_19032_),
    .X(net4260));
 sg13g2_buf_8 fanout4261 (.A(net4270),
    .X(net4261));
 sg13g2_buf_1 fanout4262 (.A(net4270),
    .X(net4262));
 sg13g2_buf_8 fanout4263 (.A(net4270),
    .X(net4263));
 sg13g2_buf_8 fanout4264 (.A(net4265),
    .X(net4264));
 sg13g2_buf_8 fanout4265 (.A(net4269),
    .X(net4265));
 sg13g2_buf_8 fanout4266 (.A(net4268),
    .X(net4266));
 sg13g2_buf_1 fanout4267 (.A(net4268),
    .X(net4267));
 sg13g2_buf_8 fanout4268 (.A(net4269),
    .X(net4268));
 sg13g2_buf_8 fanout4269 (.A(net4270),
    .X(net4269));
 sg13g2_buf_8 fanout4270 (.A(net4303),
    .X(net4270));
 sg13g2_buf_8 fanout4271 (.A(net4282),
    .X(net4271));
 sg13g2_buf_1 fanout4272 (.A(net4273),
    .X(net4272));
 sg13g2_buf_8 fanout4273 (.A(net4282),
    .X(net4273));
 sg13g2_buf_8 fanout4274 (.A(net4276),
    .X(net4274));
 sg13g2_buf_1 fanout4275 (.A(net4276),
    .X(net4275));
 sg13g2_buf_8 fanout4276 (.A(net4282),
    .X(net4276));
 sg13g2_buf_8 fanout4277 (.A(net4278),
    .X(net4277));
 sg13g2_buf_8 fanout4278 (.A(net4281),
    .X(net4278));
 sg13g2_buf_8 fanout4279 (.A(net4280),
    .X(net4279));
 sg13g2_buf_8 fanout4280 (.A(net4281),
    .X(net4280));
 sg13g2_buf_8 fanout4281 (.A(net4282),
    .X(net4281));
 sg13g2_buf_8 fanout4282 (.A(net4303),
    .X(net4282));
 sg13g2_buf_8 fanout4283 (.A(net4284),
    .X(net4283));
 sg13g2_buf_8 fanout4284 (.A(net4285),
    .X(net4284));
 sg13g2_buf_8 fanout4285 (.A(net4292),
    .X(net4285));
 sg13g2_buf_8 fanout4286 (.A(net4292),
    .X(net4286));
 sg13g2_buf_8 fanout4287 (.A(net4292),
    .X(net4287));
 sg13g2_buf_8 fanout4288 (.A(net4289),
    .X(net4288));
 sg13g2_buf_8 fanout4289 (.A(net4292),
    .X(net4289));
 sg13g2_buf_8 fanout4290 (.A(net4291),
    .X(net4290));
 sg13g2_buf_8 fanout4291 (.A(net4292),
    .X(net4291));
 sg13g2_buf_8 fanout4292 (.A(net4303),
    .X(net4292));
 sg13g2_buf_8 fanout4293 (.A(net4302),
    .X(net4293));
 sg13g2_buf_1 fanout4294 (.A(net4302),
    .X(net4294));
 sg13g2_buf_8 fanout4295 (.A(net4296),
    .X(net4295));
 sg13g2_buf_8 fanout4296 (.A(net4302),
    .X(net4296));
 sg13g2_buf_8 fanout4297 (.A(net4298),
    .X(net4297));
 sg13g2_buf_1 fanout4298 (.A(net4302),
    .X(net4298));
 sg13g2_buf_8 fanout4299 (.A(net4302),
    .X(net4299));
 sg13g2_buf_1 fanout4300 (.A(net4301),
    .X(net4300));
 sg13g2_buf_8 fanout4301 (.A(net4302),
    .X(net4301));
 sg13g2_buf_8 fanout4302 (.A(net4303),
    .X(net4302));
 sg13g2_buf_8 fanout4303 (.A(_19011_),
    .X(net4303));
 sg13g2_buf_8 fanout4304 (.A(net4305),
    .X(net4304));
 sg13g2_buf_8 fanout4305 (.A(net4313),
    .X(net4305));
 sg13g2_buf_8 fanout4306 (.A(net4313),
    .X(net4306));
 sg13g2_buf_1 fanout4307 (.A(net4313),
    .X(net4307));
 sg13g2_buf_8 fanout4308 (.A(net4309),
    .X(net4308));
 sg13g2_buf_8 fanout4309 (.A(net4313),
    .X(net4309));
 sg13g2_buf_8 fanout4310 (.A(net4312),
    .X(net4310));
 sg13g2_buf_1 fanout4311 (.A(net4312),
    .X(net4311));
 sg13g2_buf_8 fanout4312 (.A(net4313),
    .X(net4312));
 sg13g2_buf_8 fanout4313 (.A(net4347),
    .X(net4313));
 sg13g2_buf_8 fanout4314 (.A(net4320),
    .X(net4314));
 sg13g2_buf_1 fanout4315 (.A(net4320),
    .X(net4315));
 sg13g2_buf_8 fanout4316 (.A(net4320),
    .X(net4316));
 sg13g2_buf_8 fanout4317 (.A(net4319),
    .X(net4317));
 sg13g2_buf_1 fanout4318 (.A(net4319),
    .X(net4318));
 sg13g2_buf_8 fanout4319 (.A(net4320),
    .X(net4319));
 sg13g2_buf_8 fanout4320 (.A(net4347),
    .X(net4320));
 sg13g2_buf_8 fanout4321 (.A(net4323),
    .X(net4321));
 sg13g2_buf_1 fanout4322 (.A(net4323),
    .X(net4322));
 sg13g2_buf_8 fanout4323 (.A(net4326),
    .X(net4323));
 sg13g2_buf_8 fanout4324 (.A(net4325),
    .X(net4324));
 sg13g2_buf_8 fanout4325 (.A(net4326),
    .X(net4325));
 sg13g2_buf_8 fanout4326 (.A(net4347),
    .X(net4326));
 sg13g2_buf_8 fanout4327 (.A(net4329),
    .X(net4327));
 sg13g2_buf_1 fanout4328 (.A(net4329),
    .X(net4328));
 sg13g2_buf_8 fanout4329 (.A(net4336),
    .X(net4329));
 sg13g2_buf_8 fanout4330 (.A(net4331),
    .X(net4330));
 sg13g2_buf_8 fanout4331 (.A(net4336),
    .X(net4331));
 sg13g2_buf_8 fanout4332 (.A(net4333),
    .X(net4332));
 sg13g2_buf_8 fanout4333 (.A(net4336),
    .X(net4333));
 sg13g2_buf_8 fanout4334 (.A(net4335),
    .X(net4334));
 sg13g2_buf_8 fanout4335 (.A(net4336),
    .X(net4335));
 sg13g2_buf_8 fanout4336 (.A(net4347),
    .X(net4336));
 sg13g2_buf_8 fanout4337 (.A(net4346),
    .X(net4337));
 sg13g2_buf_1 fanout4338 (.A(net4346),
    .X(net4338));
 sg13g2_buf_8 fanout4339 (.A(net4340),
    .X(net4339));
 sg13g2_buf_8 fanout4340 (.A(net4346),
    .X(net4340));
 sg13g2_buf_8 fanout4341 (.A(net4342),
    .X(net4341));
 sg13g2_buf_1 fanout4342 (.A(net4346),
    .X(net4342));
 sg13g2_buf_8 fanout4343 (.A(net4346),
    .X(net4343));
 sg13g2_buf_1 fanout4344 (.A(net4345),
    .X(net4344));
 sg13g2_buf_8 fanout4345 (.A(net4346),
    .X(net4345));
 sg13g2_buf_8 fanout4346 (.A(net4347),
    .X(net4346));
 sg13g2_buf_8 fanout4347 (.A(_19031_),
    .X(net4347));
 sg13g2_buf_8 fanout4348 (.A(_19012_),
    .X(net4348));
 sg13g2_buf_8 fanout4349 (.A(_19012_),
    .X(net4349));
 sg13g2_buf_8 fanout4350 (.A(net4351),
    .X(net4350));
 sg13g2_buf_8 fanout4351 (.A(net4352),
    .X(net4351));
 sg13g2_buf_8 fanout4352 (.A(net4353),
    .X(net4352));
 sg13g2_buf_8 fanout4353 (.A(net4362),
    .X(net4353));
 sg13g2_buf_8 fanout4354 (.A(net4362),
    .X(net4354));
 sg13g2_buf_8 fanout4355 (.A(net4362),
    .X(net4355));
 sg13g2_buf_8 fanout4356 (.A(net4357),
    .X(net4356));
 sg13g2_buf_8 fanout4357 (.A(net4362),
    .X(net4357));
 sg13g2_buf_8 fanout4358 (.A(net4361),
    .X(net4358));
 sg13g2_buf_1 fanout4359 (.A(net4361),
    .X(net4359));
 sg13g2_buf_8 fanout4360 (.A(net4361),
    .X(net4360));
 sg13g2_buf_8 fanout4361 (.A(net4362),
    .X(net4361));
 sg13g2_buf_8 fanout4362 (.A(_19010_),
    .X(net4362));
 sg13g2_buf_8 fanout4363 (.A(net4367),
    .X(net4363));
 sg13g2_buf_8 fanout4364 (.A(net4367),
    .X(net4364));
 sg13g2_buf_8 fanout4365 (.A(net4367),
    .X(net4365));
 sg13g2_buf_8 fanout4366 (.A(net4367),
    .X(net4366));
 sg13g2_buf_8 fanout4367 (.A(net4373),
    .X(net4367));
 sg13g2_buf_8 fanout4368 (.A(net4369),
    .X(net4368));
 sg13g2_buf_8 fanout4369 (.A(net4373),
    .X(net4369));
 sg13g2_buf_8 fanout4370 (.A(net4371),
    .X(net4370));
 sg13g2_buf_8 fanout4371 (.A(net4372),
    .X(net4371));
 sg13g2_buf_8 fanout4372 (.A(net4373),
    .X(net4372));
 sg13g2_buf_8 fanout4373 (.A(_19010_),
    .X(net4373));
 sg13g2_buf_8 fanout4374 (.A(net4375),
    .X(net4374));
 sg13g2_buf_8 fanout4375 (.A(net4377),
    .X(net4375));
 sg13g2_buf_8 fanout4376 (.A(net4377),
    .X(net4376));
 sg13g2_buf_8 fanout4377 (.A(_03302_),
    .X(net4377));
 sg13g2_buf_8 fanout4378 (.A(net4379),
    .X(net4378));
 sg13g2_buf_8 fanout4379 (.A(_03302_),
    .X(net4379));
 sg13g2_buf_8 fanout4380 (.A(net4388),
    .X(net4380));
 sg13g2_buf_1 fanout4381 (.A(net4388),
    .X(net4381));
 sg13g2_buf_8 fanout4382 (.A(net4383),
    .X(net4382));
 sg13g2_buf_8 fanout4383 (.A(net4388),
    .X(net4383));
 sg13g2_buf_8 fanout4384 (.A(net4387),
    .X(net4384));
 sg13g2_buf_1 fanout4385 (.A(net4387),
    .X(net4385));
 sg13g2_buf_8 fanout4386 (.A(net4387),
    .X(net4386));
 sg13g2_buf_8 fanout4387 (.A(net4388),
    .X(net4387));
 sg13g2_buf_8 fanout4388 (.A(net4389),
    .X(net4388));
 sg13g2_buf_8 fanout4389 (.A(net4409),
    .X(net4389));
 sg13g2_buf_8 fanout4390 (.A(net4391),
    .X(net4390));
 sg13g2_buf_8 fanout4391 (.A(net4409),
    .X(net4391));
 sg13g2_buf_8 fanout4392 (.A(net4396),
    .X(net4392));
 sg13g2_buf_1 fanout4393 (.A(net4396),
    .X(net4393));
 sg13g2_buf_8 fanout4394 (.A(net4396),
    .X(net4394));
 sg13g2_buf_1 fanout4395 (.A(net4396),
    .X(net4395));
 sg13g2_buf_8 fanout4396 (.A(net4409),
    .X(net4396));
 sg13g2_buf_8 fanout4397 (.A(net4399),
    .X(net4397));
 sg13g2_buf_8 fanout4398 (.A(net4399),
    .X(net4398));
 sg13g2_buf_8 fanout4399 (.A(net4408),
    .X(net4399));
 sg13g2_buf_8 fanout4400 (.A(net4402),
    .X(net4400));
 sg13g2_buf_8 fanout4401 (.A(net4408),
    .X(net4401));
 sg13g2_buf_1 fanout4402 (.A(net4408),
    .X(net4402));
 sg13g2_buf_8 fanout4403 (.A(net4404),
    .X(net4403));
 sg13g2_buf_8 fanout4404 (.A(net4408),
    .X(net4404));
 sg13g2_buf_8 fanout4405 (.A(net4407),
    .X(net4405));
 sg13g2_buf_8 fanout4406 (.A(net4407),
    .X(net4406));
 sg13g2_buf_8 fanout4407 (.A(net4408),
    .X(net4407));
 sg13g2_buf_8 fanout4408 (.A(net4409),
    .X(net4408));
 sg13g2_buf_8 fanout4409 (.A(_19009_),
    .X(net4409));
 sg13g2_buf_8 fanout4410 (.A(net4414),
    .X(net4410));
 sg13g2_buf_1 fanout4411 (.A(net4414),
    .X(net4411));
 sg13g2_buf_8 fanout4412 (.A(net4414),
    .X(net4412));
 sg13g2_buf_1 fanout4413 (.A(net4414),
    .X(net4413));
 sg13g2_buf_8 fanout4414 (.A(net4417),
    .X(net4414));
 sg13g2_buf_8 fanout4415 (.A(net4416),
    .X(net4415));
 sg13g2_buf_8 fanout4416 (.A(net4417),
    .X(net4416));
 sg13g2_buf_2 fanout4417 (.A(net4449),
    .X(net4417));
 sg13g2_buf_8 fanout4418 (.A(net4427),
    .X(net4418));
 sg13g2_buf_1 fanout4419 (.A(net4427),
    .X(net4419));
 sg13g2_buf_8 fanout4420 (.A(net4423),
    .X(net4420));
 sg13g2_buf_8 fanout4421 (.A(net4423),
    .X(net4421));
 sg13g2_buf_1 fanout4422 (.A(net4423),
    .X(net4422));
 sg13g2_buf_8 fanout4423 (.A(net4427),
    .X(net4423));
 sg13g2_buf_8 fanout4424 (.A(net4427),
    .X(net4424));
 sg13g2_buf_1 fanout4425 (.A(net4427),
    .X(net4425));
 sg13g2_buf_8 fanout4426 (.A(net4427),
    .X(net4426));
 sg13g2_buf_8 fanout4427 (.A(net4449),
    .X(net4427));
 sg13g2_buf_8 fanout4428 (.A(net4429),
    .X(net4428));
 sg13g2_buf_8 fanout4429 (.A(net4431),
    .X(net4429));
 sg13g2_buf_8 fanout4430 (.A(net4431),
    .X(net4430));
 sg13g2_buf_8 fanout4431 (.A(net4438),
    .X(net4431));
 sg13g2_buf_8 fanout4432 (.A(net4438),
    .X(net4432));
 sg13g2_buf_1 fanout4433 (.A(net4438),
    .X(net4433));
 sg13g2_buf_8 fanout4434 (.A(net4437),
    .X(net4434));
 sg13g2_buf_8 fanout4435 (.A(net4436),
    .X(net4435));
 sg13g2_buf_2 fanout4436 (.A(net4437),
    .X(net4436));
 sg13g2_buf_2 fanout4437 (.A(net4438),
    .X(net4437));
 sg13g2_buf_8 fanout4438 (.A(net4449),
    .X(net4438));
 sg13g2_buf_8 fanout4439 (.A(net4440),
    .X(net4439));
 sg13g2_buf_8 fanout4440 (.A(net4447),
    .X(net4440));
 sg13g2_buf_8 fanout4441 (.A(net4442),
    .X(net4441));
 sg13g2_buf_2 fanout4442 (.A(net4443),
    .X(net4442));
 sg13g2_buf_8 fanout4443 (.A(net4447),
    .X(net4443));
 sg13g2_buf_8 fanout4444 (.A(net4446),
    .X(net4444));
 sg13g2_buf_1 fanout4445 (.A(net4446),
    .X(net4445));
 sg13g2_buf_8 fanout4446 (.A(net4447),
    .X(net4446));
 sg13g2_buf_8 fanout4447 (.A(net4448),
    .X(net4447));
 sg13g2_buf_8 fanout4448 (.A(net4449),
    .X(net4448));
 sg13g2_buf_8 fanout4449 (.A(_19009_),
    .X(net4449));
 sg13g2_buf_8 fanout4450 (.A(_19004_),
    .X(net4450));
 sg13g2_buf_1 fanout4451 (.A(_19004_),
    .X(net4451));
 sg13g2_buf_8 fanout4452 (.A(_03380_),
    .X(net4452));
 sg13g2_buf_1 fanout4453 (.A(_03380_),
    .X(net4453));
 sg13g2_buf_8 fanout4454 (.A(net4455),
    .X(net4454));
 sg13g2_buf_8 fanout4455 (.A(net4459),
    .X(net4455));
 sg13g2_buf_8 fanout4456 (.A(net4459),
    .X(net4456));
 sg13g2_buf_8 fanout4457 (.A(net4458),
    .X(net4457));
 sg13g2_buf_8 fanout4458 (.A(net4459),
    .X(net4458));
 sg13g2_buf_8 fanout4459 (.A(_03301_),
    .X(net4459));
 sg13g2_buf_8 fanout4460 (.A(net4461),
    .X(net4460));
 sg13g2_buf_8 fanout4461 (.A(net4462),
    .X(net4461));
 sg13g2_buf_8 fanout4462 (.A(net4469),
    .X(net4462));
 sg13g2_buf_8 fanout4463 (.A(net4465),
    .X(net4463));
 sg13g2_buf_8 fanout4464 (.A(net4465),
    .X(net4464));
 sg13g2_buf_8 fanout4465 (.A(net4469),
    .X(net4465));
 sg13g2_buf_8 fanout4466 (.A(net4467),
    .X(net4466));
 sg13g2_buf_8 fanout4467 (.A(net4468),
    .X(net4467));
 sg13g2_buf_8 fanout4468 (.A(net4469),
    .X(net4468));
 sg13g2_buf_8 fanout4469 (.A(_03301_),
    .X(net4469));
 sg13g2_buf_8 fanout4470 (.A(_03297_),
    .X(net4470));
 sg13g2_buf_8 fanout4471 (.A(_03297_),
    .X(net4471));
 sg13g2_buf_8 fanout4472 (.A(net4473),
    .X(net4472));
 sg13g2_buf_8 fanout4473 (.A(net1065),
    .X(net4473));
 sg13g2_buf_8 fanout4474 (.A(net4475),
    .X(net4474));
 sg13g2_buf_8 fanout4475 (.A(net4476),
    .X(net4475));
 sg13g2_buf_8 fanout4476 (.A(net1066),
    .X(net4476));
 sg13g2_buf_8 fanout4477 (.A(net4479),
    .X(net4477));
 sg13g2_buf_8 fanout4478 (.A(net4479),
    .X(net4478));
 sg13g2_buf_8 fanout4479 (.A(net4482),
    .X(net4479));
 sg13g2_buf_8 fanout4480 (.A(net4481),
    .X(net4480));
 sg13g2_buf_8 fanout4481 (.A(net4482),
    .X(net4481));
 sg13g2_buf_8 fanout4482 (.A(net1066),
    .X(net4482));
 sg13g2_buf_8 fanout4483 (.A(net4484),
    .X(net4483));
 sg13g2_buf_2 fanout4484 (.A(net4485),
    .X(net4484));
 sg13g2_buf_8 fanout4485 (.A(net4486),
    .X(net4485));
 sg13g2_buf_8 fanout4486 (.A(net4492),
    .X(net4486));
 sg13g2_buf_8 fanout4487 (.A(net4492),
    .X(net4487));
 sg13g2_buf_2 fanout4488 (.A(net4492),
    .X(net4488));
 sg13g2_buf_8 fanout4489 (.A(net4491),
    .X(net4489));
 sg13g2_buf_8 fanout4490 (.A(net4491),
    .X(net4490));
 sg13g2_buf_8 fanout4491 (.A(net4492),
    .X(net4491));
 sg13g2_buf_8 fanout4492 (.A(net1068),
    .X(net4492));
 sg13g2_buf_8 fanout4493 (.A(net4497),
    .X(net4493));
 sg13g2_buf_8 fanout4494 (.A(net4497),
    .X(net4494));
 sg13g2_buf_8 fanout4495 (.A(net4497),
    .X(net4495));
 sg13g2_buf_8 fanout4496 (.A(net4497),
    .X(net4496));
 sg13g2_buf_8 fanout4497 (.A(net1069),
    .X(net4497));
 sg13g2_buf_8 fanout4498 (.A(net4499),
    .X(net4498));
 sg13g2_buf_2 fanout4499 (.A(net4500),
    .X(net4499));
 sg13g2_buf_1 fanout4500 (.A(net4501),
    .X(net4500));
 sg13g2_buf_8 fanout4501 (.A(net4505),
    .X(net4501));
 sg13g2_buf_8 fanout4502 (.A(net4503),
    .X(net4502));
 sg13g2_buf_8 fanout4503 (.A(net4505),
    .X(net4503));
 sg13g2_buf_8 fanout4504 (.A(net4505),
    .X(net4504));
 sg13g2_buf_8 fanout4505 (.A(net4529),
    .X(net4505));
 sg13g2_buf_8 fanout4506 (.A(net4507),
    .X(net4506));
 sg13g2_buf_8 fanout4507 (.A(net4529),
    .X(net4507));
 sg13g2_buf_8 fanout4508 (.A(net4512),
    .X(net4508));
 sg13g2_buf_8 fanout4509 (.A(net4511),
    .X(net4509));
 sg13g2_buf_1 fanout4510 (.A(net4511),
    .X(net4510));
 sg13g2_buf_1 fanout4511 (.A(net4512),
    .X(net4511));
 sg13g2_buf_8 fanout4512 (.A(net4529),
    .X(net4512));
 sg13g2_buf_8 fanout4513 (.A(net4514),
    .X(net4513));
 sg13g2_buf_1 fanout4514 (.A(net4518),
    .X(net4514));
 sg13g2_buf_8 fanout4515 (.A(net4518),
    .X(net4515));
 sg13g2_buf_8 fanout4516 (.A(net4518),
    .X(net4516));
 sg13g2_buf_8 fanout4517 (.A(net4518),
    .X(net4517));
 sg13g2_buf_8 fanout4518 (.A(net4529),
    .X(net4518));
 sg13g2_buf_8 fanout4519 (.A(net4520),
    .X(net4519));
 sg13g2_buf_8 fanout4520 (.A(net4528),
    .X(net4520));
 sg13g2_buf_8 fanout4521 (.A(net4528),
    .X(net4521));
 sg13g2_buf_8 fanout4522 (.A(net4528),
    .X(net4522));
 sg13g2_buf_1 fanout4523 (.A(net4528),
    .X(net4523));
 sg13g2_buf_8 fanout4524 (.A(net4527),
    .X(net4524));
 sg13g2_buf_8 fanout4525 (.A(net4526),
    .X(net4525));
 sg13g2_buf_8 fanout4526 (.A(net4527),
    .X(net4526));
 sg13g2_buf_2 fanout4527 (.A(net4528),
    .X(net4527));
 sg13g2_buf_8 fanout4528 (.A(net4529),
    .X(net4528));
 sg13g2_buf_8 fanout4529 (.A(_02559_),
    .X(net4529));
 sg13g2_buf_8 fanout4530 (.A(net4534),
    .X(net4530));
 sg13g2_buf_8 fanout4531 (.A(net4533),
    .X(net4531));
 sg13g2_buf_1 fanout4532 (.A(net4533),
    .X(net4532));
 sg13g2_buf_8 fanout4533 (.A(net4534),
    .X(net4533));
 sg13g2_buf_8 fanout4534 (.A(net4540),
    .X(net4534));
 sg13g2_buf_8 fanout4535 (.A(net4536),
    .X(net4535));
 sg13g2_buf_8 fanout4536 (.A(net4540),
    .X(net4536));
 sg13g2_buf_8 fanout4537 (.A(net4538),
    .X(net4537));
 sg13g2_buf_8 fanout4538 (.A(net4539),
    .X(net4538));
 sg13g2_buf_8 fanout4539 (.A(net4540),
    .X(net4539));
 sg13g2_buf_8 fanout4540 (.A(net4574),
    .X(net4540));
 sg13g2_buf_8 fanout4541 (.A(net4544),
    .X(net4541));
 sg13g2_buf_2 fanout4542 (.A(net4544),
    .X(net4542));
 sg13g2_buf_8 fanout4543 (.A(net4544),
    .X(net4543));
 sg13g2_buf_8 fanout4544 (.A(net4574),
    .X(net4544));
 sg13g2_buf_8 fanout4545 (.A(net4549),
    .X(net4545));
 sg13g2_buf_8 fanout4546 (.A(net4549),
    .X(net4546));
 sg13g2_buf_8 fanout4547 (.A(net4549),
    .X(net4547));
 sg13g2_buf_1 fanout4548 (.A(net4549),
    .X(net4548));
 sg13g2_buf_8 fanout4549 (.A(net4574),
    .X(net4549));
 sg13g2_buf_8 fanout4550 (.A(net4552),
    .X(net4550));
 sg13g2_buf_8 fanout4551 (.A(net4552),
    .X(net4551));
 sg13g2_buf_8 fanout4552 (.A(net4555),
    .X(net4552));
 sg13g2_buf_8 fanout4553 (.A(net4554),
    .X(net4553));
 sg13g2_buf_8 fanout4554 (.A(net4555),
    .X(net4554));
 sg13g2_buf_8 fanout4555 (.A(net4573),
    .X(net4555));
 sg13g2_buf_8 fanout4556 (.A(net4558),
    .X(net4556));
 sg13g2_buf_8 fanout4557 (.A(net4558),
    .X(net4557));
 sg13g2_buf_8 fanout4558 (.A(net4573),
    .X(net4558));
 sg13g2_buf_8 fanout4559 (.A(net4560),
    .X(net4559));
 sg13g2_buf_8 fanout4560 (.A(net4573),
    .X(net4560));
 sg13g2_buf_8 fanout4561 (.A(net4563),
    .X(net4561));
 sg13g2_buf_8 fanout4562 (.A(net4572),
    .X(net4562));
 sg13g2_buf_1 fanout4563 (.A(net4572),
    .X(net4563));
 sg13g2_buf_8 fanout4564 (.A(net4566),
    .X(net4564));
 sg13g2_buf_2 fanout4565 (.A(net4566),
    .X(net4565));
 sg13g2_buf_8 fanout4566 (.A(net4572),
    .X(net4566));
 sg13g2_buf_8 fanout4567 (.A(net4568),
    .X(net4567));
 sg13g2_buf_8 fanout4568 (.A(net4571),
    .X(net4568));
 sg13g2_buf_8 fanout4569 (.A(net4570),
    .X(net4569));
 sg13g2_buf_8 fanout4570 (.A(net4571),
    .X(net4570));
 sg13g2_buf_8 fanout4571 (.A(net4572),
    .X(net4571));
 sg13g2_buf_8 fanout4572 (.A(net4573),
    .X(net4572));
 sg13g2_buf_8 fanout4573 (.A(net4574),
    .X(net4573));
 sg13g2_buf_8 fanout4574 (.A(_09674_),
    .X(net4574));
 sg13g2_buf_8 fanout4575 (.A(net4576),
    .X(net4575));
 sg13g2_buf_8 fanout4576 (.A(net4581),
    .X(net4576));
 sg13g2_buf_8 fanout4577 (.A(net4578),
    .X(net4577));
 sg13g2_buf_8 fanout4578 (.A(net4581),
    .X(net4578));
 sg13g2_buf_8 fanout4579 (.A(net4580),
    .X(net4579));
 sg13g2_buf_8 fanout4580 (.A(net4581),
    .X(net4580));
 sg13g2_buf_8 fanout4581 (.A(net4599),
    .X(net4581));
 sg13g2_buf_8 fanout4582 (.A(net4583),
    .X(net4582));
 sg13g2_buf_8 fanout4583 (.A(net4599),
    .X(net4583));
 sg13g2_buf_8 fanout4584 (.A(net4586),
    .X(net4584));
 sg13g2_buf_8 fanout4585 (.A(net4586),
    .X(net4585));
 sg13g2_buf_8 fanout4586 (.A(net4599),
    .X(net4586));
 sg13g2_buf_8 fanout4587 (.A(net4588),
    .X(net4587));
 sg13g2_buf_1 fanout4588 (.A(net4589),
    .X(net4588));
 sg13g2_buf_1 fanout4589 (.A(net4590),
    .X(net4589));
 sg13g2_buf_8 fanout4590 (.A(net4593),
    .X(net4590));
 sg13g2_buf_8 fanout4591 (.A(net4593),
    .X(net4591));
 sg13g2_buf_8 fanout4592 (.A(net4593),
    .X(net4592));
 sg13g2_buf_8 fanout4593 (.A(net4599),
    .X(net4593));
 sg13g2_buf_8 fanout4594 (.A(net4595),
    .X(net4594));
 sg13g2_buf_8 fanout4595 (.A(net4598),
    .X(net4595));
 sg13g2_buf_8 fanout4596 (.A(net4597),
    .X(net4596));
 sg13g2_buf_8 fanout4597 (.A(net4598),
    .X(net4597));
 sg13g2_buf_8 fanout4598 (.A(net4599),
    .X(net4598));
 sg13g2_buf_8 fanout4599 (.A(_09673_),
    .X(net4599));
 sg13g2_buf_8 fanout4600 (.A(net4601),
    .X(net4600));
 sg13g2_buf_8 fanout4601 (.A(net4604),
    .X(net4601));
 sg13g2_buf_8 fanout4602 (.A(net4604),
    .X(net4602));
 sg13g2_buf_8 fanout4603 (.A(net4604),
    .X(net4603));
 sg13g2_buf_8 fanout4604 (.A(net4627),
    .X(net4604));
 sg13g2_buf_8 fanout4605 (.A(net4609),
    .X(net4605));
 sg13g2_buf_2 fanout4606 (.A(net4609),
    .X(net4606));
 sg13g2_buf_8 fanout4607 (.A(net4609),
    .X(net4607));
 sg13g2_buf_2 fanout4608 (.A(net4609),
    .X(net4608));
 sg13g2_buf_8 fanout4609 (.A(net4627),
    .X(net4609));
 sg13g2_buf_8 fanout4610 (.A(net4611),
    .X(net4610));
 sg13g2_buf_8 fanout4611 (.A(net4612),
    .X(net4611));
 sg13g2_buf_8 fanout4612 (.A(net4627),
    .X(net4612));
 sg13g2_buf_8 fanout4613 (.A(net4626),
    .X(net4613));
 sg13g2_buf_8 fanout4614 (.A(net4626),
    .X(net4614));
 sg13g2_buf_8 fanout4615 (.A(net4616),
    .X(net4615));
 sg13g2_buf_8 fanout4616 (.A(net4617),
    .X(net4616));
 sg13g2_buf_8 fanout4617 (.A(net4626),
    .X(net4617));
 sg13g2_buf_8 fanout4618 (.A(net4619),
    .X(net4618));
 sg13g2_buf_8 fanout4619 (.A(net4622),
    .X(net4619));
 sg13g2_buf_8 fanout4620 (.A(net4621),
    .X(net4620));
 sg13g2_buf_2 fanout4621 (.A(net4622),
    .X(net4621));
 sg13g2_buf_8 fanout4622 (.A(net4626),
    .X(net4622));
 sg13g2_buf_8 fanout4623 (.A(net4624),
    .X(net4623));
 sg13g2_buf_8 fanout4624 (.A(net4625),
    .X(net4624));
 sg13g2_buf_8 fanout4625 (.A(net4626),
    .X(net4625));
 sg13g2_buf_8 fanout4626 (.A(net4627),
    .X(net4626));
 sg13g2_buf_8 fanout4627 (.A(_09673_),
    .X(net4627));
 sg13g2_buf_8 fanout4628 (.A(net4630),
    .X(net4628));
 sg13g2_buf_8 fanout4629 (.A(net4630),
    .X(net4629));
 sg13g2_buf_8 fanout4630 (.A(net1071),
    .X(net4630));
 sg13g2_buf_8 fanout4631 (.A(net1072),
    .X(net4631));
 sg13g2_buf_1 fanout4632 (.A(net4633),
    .X(net4632));
 sg13g2_buf_8 fanout4633 (.A(net1072),
    .X(net4633));
 sg13g2_buf_8 fanout4634 (.A(_09669_),
    .X(net4634));
 sg13g2_buf_8 fanout4635 (.A(_09672_),
    .X(net4635));
 sg13g2_buf_8 fanout4636 (.A(net4638),
    .X(net4636));
 sg13g2_buf_8 fanout4637 (.A(net4638),
    .X(net4637));
 sg13g2_buf_8 fanout4638 (.A(_09671_),
    .X(net4638));
 sg13g2_buf_8 fanout4639 (.A(_09671_),
    .X(net4639));
 sg13g2_buf_1 fanout4640 (.A(net4641),
    .X(net4640));
 sg13g2_buf_8 fanout4641 (.A(_09671_),
    .X(net4641));
 sg13g2_buf_8 fanout4642 (.A(net4645),
    .X(net4642));
 sg13g2_buf_8 fanout4643 (.A(net4644),
    .X(net4643));
 sg13g2_buf_8 fanout4644 (.A(net4645),
    .X(net4644));
 sg13g2_buf_8 fanout4645 (.A(net4651),
    .X(net4645));
 sg13g2_buf_8 fanout4646 (.A(net4651),
    .X(net4646));
 sg13g2_buf_8 fanout4647 (.A(net4650),
    .X(net4647));
 sg13g2_buf_8 fanout4648 (.A(net4649),
    .X(net4648));
 sg13g2_buf_8 fanout4649 (.A(net4650),
    .X(net4649));
 sg13g2_buf_8 fanout4650 (.A(net4651),
    .X(net4650));
 sg13g2_buf_8 fanout4651 (.A(net4664),
    .X(net4651));
 sg13g2_buf_8 fanout4652 (.A(net4653),
    .X(net4652));
 sg13g2_buf_8 fanout4653 (.A(net4664),
    .X(net4653));
 sg13g2_buf_8 fanout4654 (.A(net4656),
    .X(net4654));
 sg13g2_buf_1 fanout4655 (.A(net4656),
    .X(net4655));
 sg13g2_buf_8 fanout4656 (.A(net4664),
    .X(net4656));
 sg13g2_buf_8 fanout4657 (.A(net4660),
    .X(net4657));
 sg13g2_buf_8 fanout4658 (.A(net4660),
    .X(net4658));
 sg13g2_buf_1 fanout4659 (.A(net4660),
    .X(net4659));
 sg13g2_buf_8 fanout4660 (.A(net4663),
    .X(net4660));
 sg13g2_buf_8 fanout4661 (.A(net4662),
    .X(net4661));
 sg13g2_buf_8 fanout4662 (.A(net4663),
    .X(net4662));
 sg13g2_buf_8 fanout4663 (.A(net4664),
    .X(net4663));
 sg13g2_buf_8 fanout4664 (.A(net4685),
    .X(net4664));
 sg13g2_buf_8 fanout4665 (.A(net4666),
    .X(net4665));
 sg13g2_buf_8 fanout4666 (.A(net4669),
    .X(net4666));
 sg13g2_buf_1 fanout4667 (.A(net4669),
    .X(net4667));
 sg13g2_buf_8 fanout4668 (.A(net4669),
    .X(net4668));
 sg13g2_buf_8 fanout4669 (.A(net4685),
    .X(net4669));
 sg13g2_buf_8 fanout4670 (.A(net4671),
    .X(net4670));
 sg13g2_buf_8 fanout4671 (.A(net4674),
    .X(net4671));
 sg13g2_buf_8 fanout4672 (.A(net4673),
    .X(net4672));
 sg13g2_buf_8 fanout4673 (.A(net4674),
    .X(net4673));
 sg13g2_buf_8 fanout4674 (.A(net4685),
    .X(net4674));
 sg13g2_buf_8 fanout4675 (.A(net4684),
    .X(net4675));
 sg13g2_buf_8 fanout4676 (.A(net4684),
    .X(net4676));
 sg13g2_buf_8 fanout4677 (.A(net4678),
    .X(net4677));
 sg13g2_buf_8 fanout4678 (.A(net4684),
    .X(net4678));
 sg13g2_buf_8 fanout4679 (.A(net4681),
    .X(net4679));
 sg13g2_buf_1 fanout4680 (.A(net4681),
    .X(net4680));
 sg13g2_buf_8 fanout4681 (.A(net4684),
    .X(net4681));
 sg13g2_buf_8 fanout4682 (.A(net4683),
    .X(net4682));
 sg13g2_buf_8 fanout4683 (.A(net4684),
    .X(net4683));
 sg13g2_buf_8 fanout4684 (.A(net4685),
    .X(net4684));
 sg13g2_buf_8 fanout4685 (.A(_06456_),
    .X(net4685));
 sg13g2_buf_8 fanout4686 (.A(net4690),
    .X(net4686));
 sg13g2_buf_8 fanout4687 (.A(net4690),
    .X(net4687));
 sg13g2_buf_8 fanout4688 (.A(net4690),
    .X(net4688));
 sg13g2_buf_8 fanout4689 (.A(net4690),
    .X(net4689));
 sg13g2_buf_8 fanout4690 (.A(net4691),
    .X(net4690));
 sg13g2_buf_8 fanout4691 (.A(net4695),
    .X(net4691));
 sg13g2_buf_8 fanout4692 (.A(net4695),
    .X(net4692));
 sg13g2_buf_1 fanout4693 (.A(net4695),
    .X(net4693));
 sg13g2_buf_8 fanout4694 (.A(net4695),
    .X(net4694));
 sg13g2_buf_8 fanout4695 (.A(_06455_),
    .X(net4695));
 sg13g2_buf_8 fanout4696 (.A(net4697),
    .X(net4696));
 sg13g2_buf_8 fanout4697 (.A(net4703),
    .X(net4697));
 sg13g2_buf_8 fanout4698 (.A(net4703),
    .X(net4698));
 sg13g2_buf_1 fanout4699 (.A(net4703),
    .X(net4699));
 sg13g2_buf_8 fanout4700 (.A(net4702),
    .X(net4700));
 sg13g2_buf_8 fanout4701 (.A(net4702),
    .X(net4701));
 sg13g2_buf_8 fanout4702 (.A(net4703),
    .X(net4702));
 sg13g2_buf_8 fanout4703 (.A(_06455_),
    .X(net4703));
 sg13g2_buf_8 fanout4704 (.A(net4705),
    .X(net4704));
 sg13g2_buf_8 fanout4705 (.A(net4707),
    .X(net4705));
 sg13g2_buf_8 fanout4706 (.A(net4707),
    .X(net4706));
 sg13g2_buf_8 fanout4707 (.A(net4729),
    .X(net4707));
 sg13g2_buf_8 fanout4708 (.A(net4712),
    .X(net4708));
 sg13g2_buf_1 fanout4709 (.A(net4712),
    .X(net4709));
 sg13g2_buf_8 fanout4710 (.A(net4712),
    .X(net4710));
 sg13g2_buf_1 fanout4711 (.A(net4712),
    .X(net4711));
 sg13g2_buf_8 fanout4712 (.A(net4729),
    .X(net4712));
 sg13g2_buf_8 fanout4713 (.A(net4714),
    .X(net4713));
 sg13g2_buf_8 fanout4714 (.A(net4729),
    .X(net4714));
 sg13g2_buf_8 fanout4715 (.A(net4721),
    .X(net4715));
 sg13g2_buf_2 fanout4716 (.A(net4721),
    .X(net4716));
 sg13g2_buf_8 fanout4717 (.A(net4721),
    .X(net4717));
 sg13g2_buf_1 fanout4718 (.A(net4721),
    .X(net4718));
 sg13g2_buf_8 fanout4719 (.A(net4720),
    .X(net4719));
 sg13g2_buf_8 fanout4720 (.A(net4721),
    .X(net4720));
 sg13g2_buf_8 fanout4721 (.A(net4728),
    .X(net4721));
 sg13g2_buf_8 fanout4722 (.A(net4725),
    .X(net4722));
 sg13g2_buf_8 fanout4723 (.A(net4725),
    .X(net4723));
 sg13g2_buf_8 fanout4724 (.A(net4725),
    .X(net4724));
 sg13g2_buf_8 fanout4725 (.A(net4728),
    .X(net4725));
 sg13g2_buf_8 fanout4726 (.A(net4727),
    .X(net4726));
 sg13g2_buf_8 fanout4727 (.A(net4728),
    .X(net4727));
 sg13g2_buf_8 fanout4728 (.A(net4729),
    .X(net4728));
 sg13g2_buf_8 fanout4729 (.A(_06455_),
    .X(net4729));
 sg13g2_buf_8 fanout4730 (.A(net4731),
    .X(net4730));
 sg13g2_buf_8 fanout4731 (.A(net4734),
    .X(net4731));
 sg13g2_buf_8 fanout4732 (.A(net4733),
    .X(net4732));
 sg13g2_buf_8 fanout4733 (.A(net4734),
    .X(net4733));
 sg13g2_buf_8 fanout4734 (.A(net4754),
    .X(net4734));
 sg13g2_buf_8 fanout4735 (.A(net4737),
    .X(net4735));
 sg13g2_buf_1 fanout4736 (.A(net4737),
    .X(net4736));
 sg13g2_buf_8 fanout4737 (.A(net4754),
    .X(net4737));
 sg13g2_buf_8 fanout4738 (.A(net4739),
    .X(net4738));
 sg13g2_buf_8 fanout4739 (.A(net4740),
    .X(net4739));
 sg13g2_buf_8 fanout4740 (.A(net4741),
    .X(net4740));
 sg13g2_buf_8 fanout4741 (.A(net4754),
    .X(net4741));
 sg13g2_buf_8 fanout4742 (.A(net4743),
    .X(net4742));
 sg13g2_buf_8 fanout4743 (.A(net4753),
    .X(net4743));
 sg13g2_buf_8 fanout4744 (.A(net4746),
    .X(net4744));
 sg13g2_buf_8 fanout4745 (.A(net4746),
    .X(net4745));
 sg13g2_buf_8 fanout4746 (.A(net4753),
    .X(net4746));
 sg13g2_buf_8 fanout4747 (.A(net4753),
    .X(net4747));
 sg13g2_buf_8 fanout4748 (.A(net4753),
    .X(net4748));
 sg13g2_buf_8 fanout4749 (.A(net4752),
    .X(net4749));
 sg13g2_buf_8 fanout4750 (.A(net4751),
    .X(net4750));
 sg13g2_buf_1 fanout4751 (.A(net4752),
    .X(net4751));
 sg13g2_buf_8 fanout4752 (.A(net4753),
    .X(net4752));
 sg13g2_buf_8 fanout4753 (.A(net4754),
    .X(net4753));
 sg13g2_buf_8 fanout4754 (.A(_06443_),
    .X(net4754));
 sg13g2_buf_8 fanout4755 (.A(net4768),
    .X(net4755));
 sg13g2_buf_1 fanout4756 (.A(net4757),
    .X(net4756));
 sg13g2_buf_8 fanout4757 (.A(net4768),
    .X(net4757));
 sg13g2_buf_8 fanout4758 (.A(net4759),
    .X(net4758));
 sg13g2_buf_8 fanout4759 (.A(net4768),
    .X(net4759));
 sg13g2_buf_8 fanout4760 (.A(net4762),
    .X(net4760));
 sg13g2_buf_8 fanout4761 (.A(net4762),
    .X(net4761));
 sg13g2_buf_8 fanout4762 (.A(net4763),
    .X(net4762));
 sg13g2_buf_8 fanout4763 (.A(net4768),
    .X(net4763));
 sg13g2_buf_8 fanout4764 (.A(net4767),
    .X(net4764));
 sg13g2_buf_1 fanout4765 (.A(net4767),
    .X(net4765));
 sg13g2_buf_8 fanout4766 (.A(net4767),
    .X(net4766));
 sg13g2_buf_8 fanout4767 (.A(net4768),
    .X(net4767));
 sg13g2_buf_8 fanout4768 (.A(net4786),
    .X(net4768));
 sg13g2_buf_8 fanout4769 (.A(net4772),
    .X(net4769));
 sg13g2_buf_8 fanout4770 (.A(net4771),
    .X(net4770));
 sg13g2_buf_8 fanout4771 (.A(net4772),
    .X(net4771));
 sg13g2_buf_8 fanout4772 (.A(net4786),
    .X(net4772));
 sg13g2_buf_8 fanout4773 (.A(net4775),
    .X(net4773));
 sg13g2_buf_1 fanout4774 (.A(net4775),
    .X(net4774));
 sg13g2_buf_8 fanout4775 (.A(net4776),
    .X(net4775));
 sg13g2_buf_8 fanout4776 (.A(net4786),
    .X(net4776));
 sg13g2_buf_8 fanout4777 (.A(net4778),
    .X(net4777));
 sg13g2_buf_8 fanout4778 (.A(net4785),
    .X(net4778));
 sg13g2_buf_8 fanout4779 (.A(net4780),
    .X(net4779));
 sg13g2_buf_8 fanout4780 (.A(net4781),
    .X(net4780));
 sg13g2_buf_8 fanout4781 (.A(net4785),
    .X(net4781));
 sg13g2_buf_8 fanout4782 (.A(net4784),
    .X(net4782));
 sg13g2_buf_1 fanout4783 (.A(net4784),
    .X(net4783));
 sg13g2_buf_8 fanout4784 (.A(net4785),
    .X(net4784));
 sg13g2_buf_8 fanout4785 (.A(net4786),
    .X(net4785));
 sg13g2_buf_8 fanout4786 (.A(_06443_),
    .X(net4786));
 sg13g2_buf_8 fanout4787 (.A(net4790),
    .X(net4787));
 sg13g2_buf_8 fanout4788 (.A(net4790),
    .X(net4788));
 sg13g2_buf_8 fanout4789 (.A(net4790),
    .X(net4789));
 sg13g2_buf_8 fanout4790 (.A(net4798),
    .X(net4790));
 sg13g2_buf_8 fanout4791 (.A(net4798),
    .X(net4791));
 sg13g2_buf_2 fanout4792 (.A(net4798),
    .X(net4792));
 sg13g2_buf_8 fanout4793 (.A(net4794),
    .X(net4793));
 sg13g2_buf_1 fanout4794 (.A(net4797),
    .X(net4794));
 sg13g2_buf_8 fanout4795 (.A(net4796),
    .X(net4795));
 sg13g2_buf_8 fanout4796 (.A(net4797),
    .X(net4796));
 sg13g2_buf_8 fanout4797 (.A(net4798),
    .X(net4797));
 sg13g2_buf_8 fanout4798 (.A(net4830),
    .X(net4798));
 sg13g2_buf_8 fanout4799 (.A(net4802),
    .X(net4799));
 sg13g2_buf_8 fanout4800 (.A(net4801),
    .X(net4800));
 sg13g2_buf_8 fanout4801 (.A(net4802),
    .X(net4801));
 sg13g2_buf_8 fanout4802 (.A(net4807),
    .X(net4802));
 sg13g2_buf_8 fanout4803 (.A(net4804),
    .X(net4803));
 sg13g2_buf_8 fanout4804 (.A(net4807),
    .X(net4804));
 sg13g2_buf_8 fanout4805 (.A(net4807),
    .X(net4805));
 sg13g2_buf_8 fanout4806 (.A(net4807),
    .X(net4806));
 sg13g2_buf_8 fanout4807 (.A(net4830),
    .X(net4807));
 sg13g2_buf_8 fanout4808 (.A(net4809),
    .X(net4808));
 sg13g2_buf_1 fanout4809 (.A(net4813),
    .X(net4809));
 sg13g2_buf_8 fanout4810 (.A(net4813),
    .X(net4810));
 sg13g2_buf_8 fanout4811 (.A(net4812),
    .X(net4811));
 sg13g2_buf_8 fanout4812 (.A(net4813),
    .X(net4812));
 sg13g2_buf_8 fanout4813 (.A(net4830),
    .X(net4813));
 sg13g2_buf_8 fanout4814 (.A(net4815),
    .X(net4814));
 sg13g2_buf_8 fanout4815 (.A(net4818),
    .X(net4815));
 sg13g2_buf_8 fanout4816 (.A(net4817),
    .X(net4816));
 sg13g2_buf_8 fanout4817 (.A(net4818),
    .X(net4817));
 sg13g2_buf_8 fanout4818 (.A(net4830),
    .X(net4818));
 sg13g2_buf_8 fanout4819 (.A(net4820),
    .X(net4819));
 sg13g2_buf_8 fanout4820 (.A(net4829),
    .X(net4820));
 sg13g2_buf_8 fanout4821 (.A(net4829),
    .X(net4821));
 sg13g2_buf_8 fanout4822 (.A(net4829),
    .X(net4822));
 sg13g2_buf_8 fanout4823 (.A(net4824),
    .X(net4823));
 sg13g2_buf_8 fanout4824 (.A(net4829),
    .X(net4824));
 sg13g2_buf_8 fanout4825 (.A(net4829),
    .X(net4825));
 sg13g2_buf_8 fanout4826 (.A(net4828),
    .X(net4826));
 sg13g2_buf_8 fanout4827 (.A(net4828),
    .X(net4827));
 sg13g2_buf_8 fanout4828 (.A(net4829),
    .X(net4828));
 sg13g2_buf_8 fanout4829 (.A(net4830),
    .X(net4829));
 sg13g2_buf_8 fanout4830 (.A(_06442_),
    .X(net4830));
 sg13g2_buf_8 fanout4831 (.A(net4836),
    .X(net4831));
 sg13g2_buf_8 fanout4832 (.A(net4836),
    .X(net4832));
 sg13g2_buf_8 fanout4833 (.A(net4835),
    .X(net4833));
 sg13g2_buf_8 fanout4834 (.A(net4835),
    .X(net4834));
 sg13g2_buf_8 fanout4835 (.A(net4836),
    .X(net4835));
 sg13g2_buf_8 fanout4836 (.A(net4851),
    .X(net4836));
 sg13g2_buf_8 fanout4837 (.A(net4839),
    .X(net4837));
 sg13g2_buf_8 fanout4838 (.A(net4839),
    .X(net4838));
 sg13g2_buf_8 fanout4839 (.A(net4851),
    .X(net4839));
 sg13g2_buf_8 fanout4840 (.A(net4844),
    .X(net4840));
 sg13g2_buf_8 fanout4841 (.A(net4844),
    .X(net4841));
 sg13g2_buf_8 fanout4842 (.A(net4843),
    .X(net4842));
 sg13g2_buf_8 fanout4843 (.A(net4844),
    .X(net4843));
 sg13g2_buf_8 fanout4844 (.A(net4851),
    .X(net4844));
 sg13g2_buf_8 fanout4845 (.A(net4847),
    .X(net4845));
 sg13g2_buf_8 fanout4846 (.A(net4847),
    .X(net4846));
 sg13g2_buf_8 fanout4847 (.A(net4851),
    .X(net4847));
 sg13g2_buf_8 fanout4848 (.A(net4850),
    .X(net4848));
 sg13g2_buf_2 fanout4849 (.A(net4850),
    .X(net4849));
 sg13g2_buf_8 fanout4850 (.A(net4851),
    .X(net4850));
 sg13g2_buf_8 fanout4851 (.A(net4918),
    .X(net4851));
 sg13g2_buf_8 fanout4852 (.A(net4862),
    .X(net4852));
 sg13g2_buf_8 fanout4853 (.A(net4862),
    .X(net4853));
 sg13g2_buf_8 fanout4854 (.A(net4855),
    .X(net4854));
 sg13g2_buf_8 fanout4855 (.A(net4862),
    .X(net4855));
 sg13g2_buf_8 fanout4856 (.A(net4857),
    .X(net4856));
 sg13g2_buf_8 fanout4857 (.A(net4861),
    .X(net4857));
 sg13g2_buf_8 fanout4858 (.A(net4860),
    .X(net4858));
 sg13g2_buf_1 fanout4859 (.A(net4860),
    .X(net4859));
 sg13g2_buf_8 fanout4860 (.A(net4861),
    .X(net4860));
 sg13g2_buf_8 fanout4861 (.A(net4862),
    .X(net4861));
 sg13g2_buf_8 fanout4862 (.A(net4874),
    .X(net4862));
 sg13g2_buf_8 fanout4863 (.A(net4867),
    .X(net4863));
 sg13g2_buf_1 fanout4864 (.A(net4867),
    .X(net4864));
 sg13g2_buf_8 fanout4865 (.A(net4867),
    .X(net4865));
 sg13g2_buf_2 fanout4866 (.A(net4867),
    .X(net4866));
 sg13g2_buf_2 fanout4867 (.A(net4874),
    .X(net4867));
 sg13g2_buf_8 fanout4868 (.A(net4870),
    .X(net4868));
 sg13g2_buf_1 fanout4869 (.A(net4870),
    .X(net4869));
 sg13g2_buf_8 fanout4870 (.A(net4874),
    .X(net4870));
 sg13g2_buf_8 fanout4871 (.A(net4873),
    .X(net4871));
 sg13g2_buf_8 fanout4872 (.A(net4873),
    .X(net4872));
 sg13g2_buf_8 fanout4873 (.A(net4874),
    .X(net4873));
 sg13g2_buf_8 fanout4874 (.A(net4918),
    .X(net4874));
 sg13g2_buf_8 fanout4875 (.A(net4876),
    .X(net4875));
 sg13g2_buf_8 fanout4876 (.A(net4879),
    .X(net4876));
 sg13g2_buf_8 fanout4877 (.A(net4879),
    .X(net4877));
 sg13g2_buf_8 fanout4878 (.A(net4879),
    .X(net4878));
 sg13g2_buf_8 fanout4879 (.A(net4896),
    .X(net4879));
 sg13g2_buf_8 fanout4880 (.A(net4881),
    .X(net4880));
 sg13g2_buf_8 fanout4881 (.A(net4885),
    .X(net4881));
 sg13g2_buf_8 fanout4882 (.A(net4884),
    .X(net4882));
 sg13g2_buf_8 fanout4883 (.A(net4885),
    .X(net4883));
 sg13g2_buf_2 fanout4884 (.A(net4885),
    .X(net4884));
 sg13g2_buf_8 fanout4885 (.A(net4896),
    .X(net4885));
 sg13g2_buf_8 fanout4886 (.A(net4891),
    .X(net4886));
 sg13g2_buf_1 fanout4887 (.A(net4888),
    .X(net4887));
 sg13g2_buf_8 fanout4888 (.A(net4891),
    .X(net4888));
 sg13g2_buf_8 fanout4889 (.A(net4890),
    .X(net4889));
 sg13g2_buf_8 fanout4890 (.A(net4891),
    .X(net4890));
 sg13g2_buf_8 fanout4891 (.A(net4896),
    .X(net4891));
 sg13g2_buf_8 fanout4892 (.A(net4893),
    .X(net4892));
 sg13g2_buf_8 fanout4893 (.A(net4896),
    .X(net4893));
 sg13g2_buf_8 fanout4894 (.A(net4895),
    .X(net4894));
 sg13g2_buf_8 fanout4895 (.A(net4896),
    .X(net4895));
 sg13g2_buf_8 fanout4896 (.A(net4918),
    .X(net4896));
 sg13g2_buf_8 fanout4897 (.A(net4899),
    .X(net4897));
 sg13g2_buf_1 fanout4898 (.A(net4899),
    .X(net4898));
 sg13g2_buf_8 fanout4899 (.A(net4901),
    .X(net4899));
 sg13g2_buf_8 fanout4900 (.A(net4901),
    .X(net4900));
 sg13g2_buf_8 fanout4901 (.A(net4917),
    .X(net4901));
 sg13g2_buf_8 fanout4902 (.A(net4903),
    .X(net4902));
 sg13g2_buf_8 fanout4903 (.A(net4917),
    .X(net4903));
 sg13g2_buf_8 fanout4904 (.A(net4906),
    .X(net4904));
 sg13g2_buf_8 fanout4905 (.A(net4906),
    .X(net4905));
 sg13g2_buf_8 fanout4906 (.A(net4917),
    .X(net4906));
 sg13g2_buf_8 fanout4907 (.A(net4908),
    .X(net4907));
 sg13g2_buf_8 fanout4908 (.A(net4911),
    .X(net4908));
 sg13g2_buf_8 fanout4909 (.A(net4911),
    .X(net4909));
 sg13g2_buf_2 fanout4910 (.A(net4911),
    .X(net4910));
 sg13g2_buf_8 fanout4911 (.A(net4917),
    .X(net4911));
 sg13g2_buf_8 fanout4912 (.A(net4913),
    .X(net4912));
 sg13g2_buf_8 fanout4913 (.A(net4916),
    .X(net4913));
 sg13g2_buf_8 fanout4914 (.A(net4915),
    .X(net4914));
 sg13g2_buf_8 fanout4915 (.A(net4916),
    .X(net4915));
 sg13g2_buf_8 fanout4916 (.A(net4917),
    .X(net4916));
 sg13g2_buf_8 fanout4917 (.A(net4918),
    .X(net4917));
 sg13g2_buf_8 fanout4918 (.A(_13511_),
    .X(net4918));
 sg13g2_buf_8 fanout4919 (.A(net4921),
    .X(net4919));
 sg13g2_buf_8 fanout4920 (.A(net4921),
    .X(net4920));
 sg13g2_buf_8 fanout4921 (.A(net4926),
    .X(net4921));
 sg13g2_buf_8 fanout4922 (.A(net4926),
    .X(net4922));
 sg13g2_buf_1 fanout4923 (.A(net4926),
    .X(net4923));
 sg13g2_buf_8 fanout4924 (.A(net4926),
    .X(net4924));
 sg13g2_buf_8 fanout4925 (.A(net4926),
    .X(net4925));
 sg13g2_buf_8 fanout4926 (.A(net4944),
    .X(net4926));
 sg13g2_buf_8 fanout4927 (.A(net4928),
    .X(net4927));
 sg13g2_buf_8 fanout4928 (.A(net4944),
    .X(net4928));
 sg13g2_buf_1 fanout4929 (.A(net4944),
    .X(net4929));
 sg13g2_buf_8 fanout4930 (.A(net4932),
    .X(net4930));
 sg13g2_buf_1 fanout4931 (.A(net4932),
    .X(net4931));
 sg13g2_buf_8 fanout4932 (.A(net4937),
    .X(net4932));
 sg13g2_buf_8 fanout4933 (.A(net4936),
    .X(net4933));
 sg13g2_buf_1 fanout4934 (.A(net4936),
    .X(net4934));
 sg13g2_buf_8 fanout4935 (.A(net4936),
    .X(net4935));
 sg13g2_buf_8 fanout4936 (.A(net4937),
    .X(net4936));
 sg13g2_buf_8 fanout4937 (.A(net4944),
    .X(net4937));
 sg13g2_buf_8 fanout4938 (.A(net4940),
    .X(net4938));
 sg13g2_buf_1 fanout4939 (.A(net4940),
    .X(net4939));
 sg13g2_buf_8 fanout4940 (.A(net4944),
    .X(net4940));
 sg13g2_buf_8 fanout4941 (.A(net4943),
    .X(net4941));
 sg13g2_buf_8 fanout4942 (.A(net4943),
    .X(net4942));
 sg13g2_buf_8 fanout4943 (.A(net4944),
    .X(net4943));
 sg13g2_buf_8 fanout4944 (.A(net5017),
    .X(net4944));
 sg13g2_buf_8 fanout4945 (.A(net4946),
    .X(net4945));
 sg13g2_buf_8 fanout4946 (.A(net4950),
    .X(net4946));
 sg13g2_buf_8 fanout4947 (.A(net4949),
    .X(net4947));
 sg13g2_buf_8 fanout4948 (.A(net4949),
    .X(net4948));
 sg13g2_buf_8 fanout4949 (.A(net4950),
    .X(net4949));
 sg13g2_buf_8 fanout4950 (.A(net4956),
    .X(net4950));
 sg13g2_buf_8 fanout4951 (.A(net4956),
    .X(net4951));
 sg13g2_buf_8 fanout4952 (.A(net4956),
    .X(net4952));
 sg13g2_buf_8 fanout4953 (.A(net4955),
    .X(net4953));
 sg13g2_buf_1 fanout4954 (.A(net4955),
    .X(net4954));
 sg13g2_buf_8 fanout4955 (.A(net4956),
    .X(net4955));
 sg13g2_buf_8 fanout4956 (.A(net5017),
    .X(net4956));
 sg13g2_buf_8 fanout4957 (.A(net4958),
    .X(net4957));
 sg13g2_buf_8 fanout4958 (.A(net4966),
    .X(net4958));
 sg13g2_buf_8 fanout4959 (.A(net4966),
    .X(net4959));
 sg13g2_buf_8 fanout4960 (.A(net4966),
    .X(net4960));
 sg13g2_buf_8 fanout4961 (.A(net4965),
    .X(net4961));
 sg13g2_buf_8 fanout4962 (.A(net4965),
    .X(net4962));
 sg13g2_buf_1 fanout4963 (.A(net4964),
    .X(net4963));
 sg13g2_buf_8 fanout4964 (.A(net4965),
    .X(net4964));
 sg13g2_buf_8 fanout4965 (.A(net4966),
    .X(net4965));
 sg13g2_buf_8 fanout4966 (.A(net5017),
    .X(net4966));
 sg13g2_buf_8 fanout4967 (.A(net4968),
    .X(net4967));
 sg13g2_buf_1 fanout4968 (.A(net4973),
    .X(net4968));
 sg13g2_buf_8 fanout4969 (.A(net4973),
    .X(net4969));
 sg13g2_buf_8 fanout4970 (.A(net4972),
    .X(net4970));
 sg13g2_buf_8 fanout4971 (.A(net4972),
    .X(net4971));
 sg13g2_buf_8 fanout4972 (.A(net4973),
    .X(net4972));
 sg13g2_buf_8 fanout4973 (.A(net5016),
    .X(net4973));
 sg13g2_buf_8 fanout4974 (.A(net4980),
    .X(net4974));
 sg13g2_buf_8 fanout4975 (.A(net4976),
    .X(net4975));
 sg13g2_buf_8 fanout4976 (.A(net4980),
    .X(net4976));
 sg13g2_buf_8 fanout4977 (.A(net4978),
    .X(net4977));
 sg13g2_buf_8 fanout4978 (.A(net4979),
    .X(net4978));
 sg13g2_buf_8 fanout4979 (.A(net4980),
    .X(net4979));
 sg13g2_buf_8 fanout4980 (.A(net5016),
    .X(net4980));
 sg13g2_buf_8 fanout4981 (.A(net4983),
    .X(net4981));
 sg13g2_buf_8 fanout4982 (.A(net4983),
    .X(net4982));
 sg13g2_buf_8 fanout4983 (.A(net4987),
    .X(net4983));
 sg13g2_buf_8 fanout4984 (.A(net4985),
    .X(net4984));
 sg13g2_buf_8 fanout4985 (.A(net4986),
    .X(net4985));
 sg13g2_buf_8 fanout4986 (.A(net4987),
    .X(net4986));
 sg13g2_buf_8 fanout4987 (.A(net4992),
    .X(net4987));
 sg13g2_buf_8 fanout4988 (.A(net4989),
    .X(net4988));
 sg13g2_buf_8 fanout4989 (.A(net4992),
    .X(net4989));
 sg13g2_buf_8 fanout4990 (.A(net4992),
    .X(net4990));
 sg13g2_buf_8 fanout4991 (.A(net4992),
    .X(net4991));
 sg13g2_buf_8 fanout4992 (.A(net5016),
    .X(net4992));
 sg13g2_buf_8 fanout4993 (.A(net4999),
    .X(net4993));
 sg13g2_buf_8 fanout4994 (.A(net4995),
    .X(net4994));
 sg13g2_buf_8 fanout4995 (.A(net4999),
    .X(net4995));
 sg13g2_buf_8 fanout4996 (.A(net4998),
    .X(net4996));
 sg13g2_buf_8 fanout4997 (.A(net4998),
    .X(net4997));
 sg13g2_buf_8 fanout4998 (.A(net4999),
    .X(net4998));
 sg13g2_buf_8 fanout4999 (.A(net5015),
    .X(net4999));
 sg13g2_buf_8 fanout5000 (.A(net5004),
    .X(net5000));
 sg13g2_buf_1 fanout5001 (.A(net5004),
    .X(net5001));
 sg13g2_buf_8 fanout5002 (.A(net5004),
    .X(net5002));
 sg13g2_buf_1 fanout5003 (.A(net5004),
    .X(net5003));
 sg13g2_buf_8 fanout5004 (.A(net5015),
    .X(net5004));
 sg13g2_buf_8 fanout5005 (.A(net5006),
    .X(net5005));
 sg13g2_buf_8 fanout5006 (.A(net5010),
    .X(net5006));
 sg13g2_buf_8 fanout5007 (.A(net5008),
    .X(net5007));
 sg13g2_buf_8 fanout5008 (.A(net5009),
    .X(net5008));
 sg13g2_buf_8 fanout5009 (.A(net5010),
    .X(net5009));
 sg13g2_buf_8 fanout5010 (.A(net5015),
    .X(net5010));
 sg13g2_buf_8 fanout5011 (.A(net5012),
    .X(net5011));
 sg13g2_buf_1 fanout5012 (.A(net5014),
    .X(net5012));
 sg13g2_buf_8 fanout5013 (.A(net5014),
    .X(net5013));
 sg13g2_buf_2 fanout5014 (.A(net5015),
    .X(net5014));
 sg13g2_buf_8 fanout5015 (.A(net5016),
    .X(net5015));
 sg13g2_buf_8 fanout5016 (.A(net5017),
    .X(net5016));
 sg13g2_buf_8 fanout5017 (.A(_15969_),
    .X(net5017));
 sg13g2_buf_8 fanout5018 (.A(net5022),
    .X(net5018));
 sg13g2_buf_2 fanout5019 (.A(net5022),
    .X(net5019));
 sg13g2_buf_8 fanout5020 (.A(net5022),
    .X(net5020));
 sg13g2_buf_1 fanout5021 (.A(net5022),
    .X(net5021));
 sg13g2_buf_8 fanout5022 (.A(net5027),
    .X(net5022));
 sg13g2_buf_8 fanout5023 (.A(net5024),
    .X(net5023));
 sg13g2_buf_8 fanout5024 (.A(net5027),
    .X(net5024));
 sg13g2_buf_8 fanout5025 (.A(net5026),
    .X(net5025));
 sg13g2_buf_8 fanout5026 (.A(net5027),
    .X(net5026));
 sg13g2_buf_8 fanout5027 (.A(net5059),
    .X(net5027));
 sg13g2_buf_8 fanout5028 (.A(net5029),
    .X(net5028));
 sg13g2_buf_8 fanout5029 (.A(net5030),
    .X(net5029));
 sg13g2_buf_8 fanout5030 (.A(net5059),
    .X(net5030));
 sg13g2_buf_8 fanout5031 (.A(net5032),
    .X(net5031));
 sg13g2_buf_8 fanout5032 (.A(net5037),
    .X(net5032));
 sg13g2_buf_8 fanout5033 (.A(net5037),
    .X(net5033));
 sg13g2_buf_8 fanout5034 (.A(net5035),
    .X(net5034));
 sg13g2_buf_8 fanout5035 (.A(net5036),
    .X(net5035));
 sg13g2_buf_8 fanout5036 (.A(net5037),
    .X(net5036));
 sg13g2_buf_8 fanout5037 (.A(net5059),
    .X(net5037));
 sg13g2_buf_8 fanout5038 (.A(net5040),
    .X(net5038));
 sg13g2_buf_8 fanout5039 (.A(net5040),
    .X(net5039));
 sg13g2_buf_8 fanout5040 (.A(net5058),
    .X(net5040));
 sg13g2_buf_8 fanout5041 (.A(net5047),
    .X(net5041));
 sg13g2_buf_8 fanout5042 (.A(net5047),
    .X(net5042));
 sg13g2_buf_8 fanout5043 (.A(net5047),
    .X(net5043));
 sg13g2_buf_8 fanout5044 (.A(net5046),
    .X(net5044));
 sg13g2_buf_8 fanout5045 (.A(net5046),
    .X(net5045));
 sg13g2_buf_8 fanout5046 (.A(net5047),
    .X(net5046));
 sg13g2_buf_8 fanout5047 (.A(net5058),
    .X(net5047));
 sg13g2_buf_8 fanout5048 (.A(net5051),
    .X(net5048));
 sg13g2_buf_8 fanout5049 (.A(net5050),
    .X(net5049));
 sg13g2_buf_8 fanout5050 (.A(net5051),
    .X(net5050));
 sg13g2_buf_8 fanout5051 (.A(net5058),
    .X(net5051));
 sg13g2_buf_8 fanout5052 (.A(net5053),
    .X(net5052));
 sg13g2_buf_8 fanout5053 (.A(net5054),
    .X(net5053));
 sg13g2_buf_8 fanout5054 (.A(net5058),
    .X(net5054));
 sg13g2_buf_8 fanout5055 (.A(net5057),
    .X(net5055));
 sg13g2_buf_1 fanout5056 (.A(net5057),
    .X(net5056));
 sg13g2_buf_8 fanout5057 (.A(net5058),
    .X(net5057));
 sg13g2_buf_8 fanout5058 (.A(net5059),
    .X(net5058));
 sg13g2_buf_8 fanout5059 (.A(_15968_),
    .X(net5059));
 sg13g2_buf_8 fanout5060 (.A(net5064),
    .X(net5060));
 sg13g2_buf_1 fanout5061 (.A(net5064),
    .X(net5061));
 sg13g2_buf_8 fanout5062 (.A(net5064),
    .X(net5062));
 sg13g2_buf_1 fanout5063 (.A(net5064),
    .X(net5063));
 sg13g2_buf_2 fanout5064 (.A(net5080),
    .X(net5064));
 sg13g2_buf_8 fanout5065 (.A(net5069),
    .X(net5065));
 sg13g2_buf_2 fanout5066 (.A(net5069),
    .X(net5066));
 sg13g2_buf_8 fanout5067 (.A(net5068),
    .X(net5067));
 sg13g2_buf_8 fanout5068 (.A(net5069),
    .X(net5068));
 sg13g2_buf_8 fanout5069 (.A(net5080),
    .X(net5069));
 sg13g2_buf_8 fanout5070 (.A(net5073),
    .X(net5070));
 sg13g2_buf_8 fanout5071 (.A(net5072),
    .X(net5071));
 sg13g2_buf_8 fanout5072 (.A(net5073),
    .X(net5072));
 sg13g2_buf_8 fanout5073 (.A(net5080),
    .X(net5073));
 sg13g2_buf_8 fanout5074 (.A(net5076),
    .X(net5074));
 sg13g2_buf_1 fanout5075 (.A(net5076),
    .X(net5075));
 sg13g2_buf_8 fanout5076 (.A(net5080),
    .X(net5076));
 sg13g2_buf_8 fanout5077 (.A(net5078),
    .X(net5077));
 sg13g2_buf_8 fanout5078 (.A(net5079),
    .X(net5078));
 sg13g2_buf_2 fanout5079 (.A(net5080),
    .X(net5079));
 sg13g2_buf_8 fanout5080 (.A(net5103),
    .X(net5080));
 sg13g2_buf_8 fanout5081 (.A(net5084),
    .X(net5081));
 sg13g2_buf_8 fanout5082 (.A(net5083),
    .X(net5082));
 sg13g2_buf_8 fanout5083 (.A(net5084),
    .X(net5083));
 sg13g2_buf_8 fanout5084 (.A(net5103),
    .X(net5084));
 sg13g2_buf_8 fanout5085 (.A(net5090),
    .X(net5085));
 sg13g2_buf_8 fanout5086 (.A(net5087),
    .X(net5086));
 sg13g2_buf_1 fanout5087 (.A(net5088),
    .X(net5087));
 sg13g2_buf_2 fanout5088 (.A(net5089),
    .X(net5088));
 sg13g2_buf_8 fanout5089 (.A(net5090),
    .X(net5089));
 sg13g2_buf_8 fanout5090 (.A(net5103),
    .X(net5090));
 sg13g2_buf_8 fanout5091 (.A(net5093),
    .X(net5091));
 sg13g2_buf_2 fanout5092 (.A(net5093),
    .X(net5092));
 sg13g2_buf_8 fanout5093 (.A(net5102),
    .X(net5093));
 sg13g2_buf_8 fanout5094 (.A(net5102),
    .X(net5094));
 sg13g2_buf_8 fanout5095 (.A(net5102),
    .X(net5095));
 sg13g2_buf_8 fanout5096 (.A(net5102),
    .X(net5096));
 sg13g2_buf_8 fanout5097 (.A(net5102),
    .X(net5097));
 sg13g2_buf_8 fanout5098 (.A(net5099),
    .X(net5098));
 sg13g2_buf_8 fanout5099 (.A(net5101),
    .X(net5099));
 sg13g2_buf_8 fanout5100 (.A(net5101),
    .X(net5100));
 sg13g2_buf_8 fanout5101 (.A(net5102),
    .X(net5101));
 sg13g2_buf_8 fanout5102 (.A(net5103),
    .X(net5102));
 sg13g2_buf_8 fanout5103 (.A(_15968_),
    .X(net5103));
 sg13g2_buf_8 fanout5104 (.A(net5106),
    .X(net5104));
 sg13g2_buf_1 fanout5105 (.A(net5106),
    .X(net5105));
 sg13g2_buf_8 fanout5106 (.A(net5107),
    .X(net5106));
 sg13g2_buf_8 fanout5107 (.A(net5108),
    .X(net5107));
 sg13g2_buf_8 fanout5108 (.A(net5117),
    .X(net5108));
 sg13g2_buf_8 fanout5109 (.A(net5112),
    .X(net5109));
 sg13g2_buf_1 fanout5110 (.A(net5112),
    .X(net5110));
 sg13g2_buf_8 fanout5111 (.A(net5112),
    .X(net5111));
 sg13g2_buf_8 fanout5112 (.A(net5117),
    .X(net5112));
 sg13g2_buf_8 fanout5113 (.A(net5115),
    .X(net5113));
 sg13g2_buf_8 fanout5114 (.A(net5115),
    .X(net5114));
 sg13g2_buf_8 fanout5115 (.A(net5117),
    .X(net5115));
 sg13g2_buf_8 fanout5116 (.A(net5117),
    .X(net5116));
 sg13g2_buf_8 fanout5117 (.A(_02383_),
    .X(net5117));
 sg13g2_buf_8 fanout5118 (.A(net5119),
    .X(net5118));
 sg13g2_buf_8 fanout5119 (.A(net5123),
    .X(net5119));
 sg13g2_buf_8 fanout5120 (.A(net5123),
    .X(net5120));
 sg13g2_buf_8 fanout5121 (.A(net5122),
    .X(net5121));
 sg13g2_buf_8 fanout5122 (.A(net5123),
    .X(net5122));
 sg13g2_buf_8 fanout5123 (.A(_02383_),
    .X(net5123));
 sg13g2_buf_8 fanout5124 (.A(net5125),
    .X(net5124));
 sg13g2_buf_8 fanout5125 (.A(net5126),
    .X(net5125));
 sg13g2_buf_8 fanout5126 (.A(net5133),
    .X(net5126));
 sg13g2_buf_8 fanout5127 (.A(net5133),
    .X(net5127));
 sg13g2_buf_8 fanout5128 (.A(net5131),
    .X(net5128));
 sg13g2_buf_2 fanout5129 (.A(net5131),
    .X(net5129));
 sg13g2_buf_8 fanout5130 (.A(net5131),
    .X(net5130));
 sg13g2_buf_8 fanout5131 (.A(net5132),
    .X(net5131));
 sg13g2_buf_8 fanout5132 (.A(net5133),
    .X(net5132));
 sg13g2_buf_8 fanout5133 (.A(_02383_),
    .X(net5133));
 sg13g2_buf_8 fanout5134 (.A(net5135),
    .X(net5134));
 sg13g2_buf_1 fanout5135 (.A(net5137),
    .X(net5135));
 sg13g2_buf_8 fanout5136 (.A(net5137),
    .X(net5136));
 sg13g2_buf_1 fanout5137 (.A(net5146),
    .X(net5137));
 sg13g2_buf_8 fanout5138 (.A(net5139),
    .X(net5138));
 sg13g2_buf_8 fanout5139 (.A(net5146),
    .X(net5139));
 sg13g2_buf_8 fanout5140 (.A(net5141),
    .X(net5140));
 sg13g2_buf_1 fanout5141 (.A(net5142),
    .X(net5141));
 sg13g2_buf_8 fanout5142 (.A(net5146),
    .X(net5142));
 sg13g2_buf_8 fanout5143 (.A(net5144),
    .X(net5143));
 sg13g2_buf_2 fanout5144 (.A(net5145),
    .X(net5144));
 sg13g2_buf_1 fanout5145 (.A(net5146),
    .X(net5145));
 sg13g2_buf_2 fanout5146 (.A(net5163),
    .X(net5146));
 sg13g2_buf_8 fanout5147 (.A(net5149),
    .X(net5147));
 sg13g2_buf_1 fanout5148 (.A(net5149),
    .X(net5148));
 sg13g2_buf_8 fanout5149 (.A(net5150),
    .X(net5149));
 sg13g2_buf_2 fanout5150 (.A(net5163),
    .X(net5150));
 sg13g2_buf_8 fanout5151 (.A(net5152),
    .X(net5151));
 sg13g2_buf_8 fanout5152 (.A(net5158),
    .X(net5152));
 sg13g2_buf_8 fanout5153 (.A(net5154),
    .X(net5153));
 sg13g2_buf_2 fanout5154 (.A(net5155),
    .X(net5154));
 sg13g2_buf_1 fanout5155 (.A(net5158),
    .X(net5155));
 sg13g2_buf_8 fanout5156 (.A(net5157),
    .X(net5156));
 sg13g2_buf_8 fanout5157 (.A(net5158),
    .X(net5157));
 sg13g2_buf_2 fanout5158 (.A(net5163),
    .X(net5158));
 sg13g2_buf_8 fanout5159 (.A(net5162),
    .X(net5159));
 sg13g2_buf_8 fanout5160 (.A(net5161),
    .X(net5160));
 sg13g2_buf_8 fanout5161 (.A(net5162),
    .X(net5161));
 sg13g2_buf_8 fanout5162 (.A(net5163),
    .X(net5162));
 sg13g2_buf_8 fanout5163 (.A(net11),
    .X(net5163));
 sg13g2_buf_8 fanout5164 (.A(net5165),
    .X(net5164));
 sg13g2_buf_8 fanout5165 (.A(net5169),
    .X(net5165));
 sg13g2_buf_1 fanout5166 (.A(net5169),
    .X(net5166));
 sg13g2_buf_8 fanout5167 (.A(net5169),
    .X(net5167));
 sg13g2_buf_2 fanout5168 (.A(net5169),
    .X(net5168));
 sg13g2_buf_8 fanout5169 (.A(net5186),
    .X(net5169));
 sg13g2_buf_8 fanout5170 (.A(net5173),
    .X(net5170));
 sg13g2_buf_1 fanout5171 (.A(net5173),
    .X(net5171));
 sg13g2_buf_8 fanout5172 (.A(net5173),
    .X(net5172));
 sg13g2_buf_8 fanout5173 (.A(net5186),
    .X(net5173));
 sg13g2_buf_8 fanout5174 (.A(net5179),
    .X(net5174));
 sg13g2_buf_8 fanout5175 (.A(net5176),
    .X(net5175));
 sg13g2_buf_8 fanout5176 (.A(net5179),
    .X(net5176));
 sg13g2_buf_8 fanout5177 (.A(net5178),
    .X(net5177));
 sg13g2_buf_8 fanout5178 (.A(net5179),
    .X(net5178));
 sg13g2_buf_8 fanout5179 (.A(net5185),
    .X(net5179));
 sg13g2_buf_8 fanout5180 (.A(net5182),
    .X(net5180));
 sg13g2_buf_8 fanout5181 (.A(net5182),
    .X(net5181));
 sg13g2_buf_8 fanout5182 (.A(net5185),
    .X(net5182));
 sg13g2_buf_8 fanout5183 (.A(net5185),
    .X(net5183));
 sg13g2_buf_1 fanout5184 (.A(net5185),
    .X(net5184));
 sg13g2_buf_8 fanout5185 (.A(net5186),
    .X(net5185));
 sg13g2_buf_8 fanout5186 (.A(net11),
    .X(net5186));
 sg13g2_buf_8 fanout5187 (.A(net5190),
    .X(net5187));
 sg13g2_buf_8 fanout5188 (.A(net5189),
    .X(net5188));
 sg13g2_buf_1 fanout5189 (.A(net5190),
    .X(net5189));
 sg13g2_buf_1 fanout5190 (.A(net5191),
    .X(net5190));
 sg13g2_buf_8 fanout5191 (.A(net5196),
    .X(net5191));
 sg13g2_buf_8 fanout5192 (.A(net5196),
    .X(net5192));
 sg13g2_buf_8 fanout5193 (.A(net5195),
    .X(net5193));
 sg13g2_buf_1 fanout5194 (.A(net5195),
    .X(net5194));
 sg13g2_buf_8 fanout5195 (.A(net5196),
    .X(net5195));
 sg13g2_buf_8 fanout5196 (.A(net5229),
    .X(net5196));
 sg13g2_buf_8 fanout5197 (.A(net5201),
    .X(net5197));
 sg13g2_buf_8 fanout5198 (.A(net5201),
    .X(net5198));
 sg13g2_buf_2 fanout5199 (.A(net5200),
    .X(net5199));
 sg13g2_buf_2 fanout5200 (.A(net5201),
    .X(net5200));
 sg13g2_buf_8 fanout5201 (.A(net5229),
    .X(net5201));
 sg13g2_buf_2 fanout5202 (.A(net5204),
    .X(net5202));
 sg13g2_buf_8 fanout5203 (.A(net5204),
    .X(net5203));
 sg13g2_buf_2 fanout5204 (.A(net5205),
    .X(net5204));
 sg13g2_buf_8 fanout5205 (.A(net5229),
    .X(net5205));
 sg13g2_buf_8 fanout5206 (.A(net5210),
    .X(net5206));
 sg13g2_buf_8 fanout5207 (.A(net5209),
    .X(net5207));
 sg13g2_buf_1 fanout5208 (.A(net5209),
    .X(net5208));
 sg13g2_buf_8 fanout5209 (.A(net5210),
    .X(net5209));
 sg13g2_buf_8 fanout5210 (.A(net5229),
    .X(net5210));
 sg13g2_buf_8 fanout5211 (.A(net5213),
    .X(net5211));
 sg13g2_buf_1 fanout5212 (.A(net5213),
    .X(net5212));
 sg13g2_buf_8 fanout5213 (.A(net5214),
    .X(net5213));
 sg13g2_buf_8 fanout5214 (.A(net5229),
    .X(net5214));
 sg13g2_buf_8 fanout5215 (.A(net5218),
    .X(net5215));
 sg13g2_buf_2 fanout5216 (.A(net5218),
    .X(net5216));
 sg13g2_buf_8 fanout5217 (.A(net5218),
    .X(net5217));
 sg13g2_buf_8 fanout5218 (.A(net5228),
    .X(net5218));
 sg13g2_buf_8 fanout5219 (.A(net5223),
    .X(net5219));
 sg13g2_buf_1 fanout5220 (.A(net5223),
    .X(net5220));
 sg13g2_buf_8 fanout5221 (.A(net5222),
    .X(net5221));
 sg13g2_buf_8 fanout5222 (.A(net5223),
    .X(net5222));
 sg13g2_buf_8 fanout5223 (.A(net5228),
    .X(net5223));
 sg13g2_buf_8 fanout5224 (.A(net5226),
    .X(net5224));
 sg13g2_buf_1 fanout5225 (.A(net5226),
    .X(net5225));
 sg13g2_buf_2 fanout5226 (.A(net5228),
    .X(net5226));
 sg13g2_buf_2 fanout5227 (.A(net5228),
    .X(net5227));
 sg13g2_buf_8 fanout5228 (.A(net5229),
    .X(net5228));
 sg13g2_buf_8 fanout5229 (.A(net11),
    .X(net5229));
 sg13g2_buf_8 fanout5230 (.A(_19507_),
    .X(net5230));
 sg13g2_buf_8 fanout5231 (.A(net5232),
    .X(net5231));
 sg13g2_buf_8 fanout5232 (.A(net5239),
    .X(net5232));
 sg13g2_buf_8 fanout5233 (.A(net5238),
    .X(net5233));
 sg13g2_buf_8 fanout5234 (.A(net5238),
    .X(net5234));
 sg13g2_buf_8 fanout5235 (.A(net5237),
    .X(net5235));
 sg13g2_buf_1 fanout5236 (.A(net5237),
    .X(net5236));
 sg13g2_buf_8 fanout5237 (.A(net5238),
    .X(net5237));
 sg13g2_buf_8 fanout5238 (.A(net5239),
    .X(net5238));
 sg13g2_buf_8 fanout5239 (.A(net5266),
    .X(net5239));
 sg13g2_buf_8 fanout5240 (.A(net5241),
    .X(net5240));
 sg13g2_buf_8 fanout5241 (.A(net5242),
    .X(net5241));
 sg13g2_buf_8 fanout5242 (.A(net5249),
    .X(net5242));
 sg13g2_buf_8 fanout5243 (.A(net5249),
    .X(net5243));
 sg13g2_buf_1 fanout5244 (.A(net5249),
    .X(net5244));
 sg13g2_buf_8 fanout5245 (.A(net5248),
    .X(net5245));
 sg13g2_buf_1 fanout5246 (.A(net5248),
    .X(net5246));
 sg13g2_buf_8 fanout5247 (.A(net5248),
    .X(net5247));
 sg13g2_buf_8 fanout5248 (.A(net5249),
    .X(net5248));
 sg13g2_buf_8 fanout5249 (.A(net5266),
    .X(net5249));
 sg13g2_buf_8 fanout5250 (.A(net5252),
    .X(net5250));
 sg13g2_buf_8 fanout5251 (.A(net5252),
    .X(net5251));
 sg13g2_buf_8 fanout5252 (.A(net5253),
    .X(net5252));
 sg13g2_buf_8 fanout5253 (.A(net5266),
    .X(net5253));
 sg13g2_buf_8 fanout5254 (.A(net5256),
    .X(net5254));
 sg13g2_buf_1 fanout5255 (.A(net5256),
    .X(net5255));
 sg13g2_buf_8 fanout5256 (.A(net5266),
    .X(net5256));
 sg13g2_buf_8 fanout5257 (.A(net5259),
    .X(net5257));
 sg13g2_buf_8 fanout5258 (.A(net5259),
    .X(net5258));
 sg13g2_buf_8 fanout5259 (.A(net5265),
    .X(net5259));
 sg13g2_buf_8 fanout5260 (.A(net5261),
    .X(net5260));
 sg13g2_buf_8 fanout5261 (.A(net5264),
    .X(net5261));
 sg13g2_buf_8 fanout5262 (.A(net5264),
    .X(net5262));
 sg13g2_buf_1 fanout5263 (.A(net5264),
    .X(net5263));
 sg13g2_buf_8 fanout5264 (.A(net5265),
    .X(net5264));
 sg13g2_buf_8 fanout5265 (.A(net5266),
    .X(net5265));
 sg13g2_buf_8 fanout5266 (.A(_02382_),
    .X(net5266));
 sg13g2_buf_8 fanout5267 (.A(net5273),
    .X(net5267));
 sg13g2_buf_8 fanout5268 (.A(net5273),
    .X(net5268));
 sg13g2_buf_1 fanout5269 (.A(net5273),
    .X(net5269));
 sg13g2_buf_8 fanout5270 (.A(net5272),
    .X(net5270));
 sg13g2_buf_8 fanout5271 (.A(net5272),
    .X(net5271));
 sg13g2_buf_8 fanout5272 (.A(net5273),
    .X(net5272));
 sg13g2_buf_8 fanout5273 (.A(net5280),
    .X(net5273));
 sg13g2_buf_8 fanout5274 (.A(net5280),
    .X(net5274));
 sg13g2_buf_1 fanout5275 (.A(net5280),
    .X(net5275));
 sg13g2_buf_8 fanout5276 (.A(net5277),
    .X(net5276));
 sg13g2_buf_1 fanout5277 (.A(net5278),
    .X(net5277));
 sg13g2_buf_2 fanout5278 (.A(net5279),
    .X(net5278));
 sg13g2_buf_8 fanout5279 (.A(net5280),
    .X(net5279));
 sg13g2_buf_8 fanout5280 (.A(net5295),
    .X(net5280));
 sg13g2_buf_8 fanout5281 (.A(net5286),
    .X(net5281));
 sg13g2_buf_8 fanout5282 (.A(net5283),
    .X(net5282));
 sg13g2_buf_1 fanout5283 (.A(net5286),
    .X(net5283));
 sg13g2_buf_8 fanout5284 (.A(net5285),
    .X(net5284));
 sg13g2_buf_2 fanout5285 (.A(net5286),
    .X(net5285));
 sg13g2_buf_1 fanout5286 (.A(net5295),
    .X(net5286));
 sg13g2_buf_8 fanout5287 (.A(net5288),
    .X(net5287));
 sg13g2_buf_8 fanout5288 (.A(net5295),
    .X(net5288));
 sg13g2_buf_8 fanout5289 (.A(net5294),
    .X(net5289));
 sg13g2_buf_1 fanout5290 (.A(net5291),
    .X(net5290));
 sg13g2_buf_8 fanout5291 (.A(net5294),
    .X(net5291));
 sg13g2_buf_8 fanout5292 (.A(net5294),
    .X(net5292));
 sg13g2_buf_1 fanout5293 (.A(net5294),
    .X(net5293));
 sg13g2_buf_8 fanout5294 (.A(net5295),
    .X(net5294));
 sg13g2_buf_8 fanout5295 (.A(_02382_),
    .X(net5295));
 sg13g2_buf_8 fanout5296 (.A(_19504_),
    .X(net5296));
 sg13g2_buf_8 fanout5297 (.A(net5299),
    .X(net5297));
 sg13g2_buf_1 fanout5298 (.A(net5299),
    .X(net5298));
 sg13g2_buf_2 fanout5299 (.A(net5308),
    .X(net5299));
 sg13g2_buf_8 fanout5300 (.A(net5301),
    .X(net5300));
 sg13g2_buf_8 fanout5301 (.A(net5302),
    .X(net5301));
 sg13g2_buf_8 fanout5302 (.A(net5308),
    .X(net5302));
 sg13g2_buf_8 fanout5303 (.A(net5305),
    .X(net5303));
 sg13g2_buf_8 fanout5304 (.A(net5305),
    .X(net5304));
 sg13g2_buf_8 fanout5305 (.A(net5308),
    .X(net5305));
 sg13g2_buf_8 fanout5306 (.A(net5307),
    .X(net5306));
 sg13g2_buf_8 fanout5307 (.A(net5308),
    .X(net5307));
 sg13g2_buf_8 fanout5308 (.A(_13845_),
    .X(net5308));
 sg13g2_buf_8 fanout5309 (.A(net5311),
    .X(net5309));
 sg13g2_buf_8 fanout5310 (.A(net5320),
    .X(net5310));
 sg13g2_buf_8 fanout5311 (.A(net5320),
    .X(net5311));
 sg13g2_buf_8 fanout5312 (.A(net5314),
    .X(net5312));
 sg13g2_buf_8 fanout5313 (.A(net5314),
    .X(net5313));
 sg13g2_buf_8 fanout5314 (.A(net5320),
    .X(net5314));
 sg13g2_buf_8 fanout5315 (.A(net5317),
    .X(net5315));
 sg13g2_buf_2 fanout5316 (.A(net5317),
    .X(net5316));
 sg13g2_buf_8 fanout5317 (.A(net5320),
    .X(net5317));
 sg13g2_buf_8 fanout5318 (.A(net5319),
    .X(net5318));
 sg13g2_buf_8 fanout5319 (.A(net5320),
    .X(net5319));
 sg13g2_buf_8 fanout5320 (.A(_13845_),
    .X(net5320));
 sg13g2_buf_8 fanout5321 (.A(net5323),
    .X(net5321));
 sg13g2_buf_8 fanout5322 (.A(net5323),
    .X(net5322));
 sg13g2_buf_8 fanout5323 (.A(net5325),
    .X(net5323));
 sg13g2_buf_8 fanout5324 (.A(net5325),
    .X(net5324));
 sg13g2_buf_8 fanout5325 (.A(net5331),
    .X(net5325));
 sg13g2_buf_8 fanout5326 (.A(net5331),
    .X(net5326));
 sg13g2_buf_8 fanout5327 (.A(net5331),
    .X(net5327));
 sg13g2_buf_8 fanout5328 (.A(net5330),
    .X(net5328));
 sg13g2_buf_1 fanout5329 (.A(net5330),
    .X(net5329));
 sg13g2_buf_8 fanout5330 (.A(net5331),
    .X(net5330));
 sg13g2_buf_8 fanout5331 (.A(net5342),
    .X(net5331));
 sg13g2_buf_8 fanout5332 (.A(net5333),
    .X(net5332));
 sg13g2_buf_8 fanout5333 (.A(net5342),
    .X(net5333));
 sg13g2_buf_8 fanout5334 (.A(net5335),
    .X(net5334));
 sg13g2_buf_8 fanout5335 (.A(net5342),
    .X(net5335));
 sg13g2_buf_8 fanout5336 (.A(net5337),
    .X(net5336));
 sg13g2_buf_8 fanout5337 (.A(net5341),
    .X(net5337));
 sg13g2_buf_8 fanout5338 (.A(net5341),
    .X(net5338));
 sg13g2_buf_8 fanout5339 (.A(net5341),
    .X(net5339));
 sg13g2_buf_8 fanout5340 (.A(net5341),
    .X(net5340));
 sg13g2_buf_8 fanout5341 (.A(net5342),
    .X(net5341));
 sg13g2_buf_8 fanout5342 (.A(_13845_),
    .X(net5342));
 sg13g2_buf_8 fanout5343 (.A(net5344),
    .X(net5343));
 sg13g2_buf_1 fanout5344 (.A(net5347),
    .X(net5344));
 sg13g2_buf_8 fanout5345 (.A(net5347),
    .X(net5345));
 sg13g2_buf_1 fanout5346 (.A(net5347),
    .X(net5346));
 sg13g2_buf_8 fanout5347 (.A(net5353),
    .X(net5347));
 sg13g2_buf_8 fanout5348 (.A(net5349),
    .X(net5348));
 sg13g2_buf_8 fanout5349 (.A(net5353),
    .X(net5349));
 sg13g2_buf_8 fanout5350 (.A(net5353),
    .X(net5350));
 sg13g2_buf_8 fanout5351 (.A(net5352),
    .X(net5351));
 sg13g2_buf_8 fanout5352 (.A(net5353),
    .X(net5352));
 sg13g2_buf_8 fanout5353 (.A(_06451_),
    .X(net5353));
 sg13g2_buf_8 fanout5354 (.A(net5358),
    .X(net5354));
 sg13g2_buf_2 fanout5355 (.A(net5358),
    .X(net5355));
 sg13g2_buf_8 fanout5356 (.A(net5357),
    .X(net5356));
 sg13g2_buf_8 fanout5357 (.A(net5358),
    .X(net5357));
 sg13g2_buf_8 fanout5358 (.A(net5364),
    .X(net5358));
 sg13g2_buf_8 fanout5359 (.A(net5364),
    .X(net5359));
 sg13g2_buf_1 fanout5360 (.A(net5364),
    .X(net5360));
 sg13g2_buf_8 fanout5361 (.A(net5363),
    .X(net5361));
 sg13g2_buf_1 fanout5362 (.A(net5363),
    .X(net5362));
 sg13g2_buf_8 fanout5363 (.A(net5364),
    .X(net5363));
 sg13g2_buf_8 fanout5364 (.A(_06451_),
    .X(net5364));
 sg13g2_buf_8 fanout5365 (.A(net5366),
    .X(net5365));
 sg13g2_buf_8 fanout5366 (.A(net5368),
    .X(net5366));
 sg13g2_buf_8 fanout5367 (.A(net5368),
    .X(net5367));
 sg13g2_buf_8 fanout5368 (.A(net5386),
    .X(net5368));
 sg13g2_buf_8 fanout5369 (.A(net5372),
    .X(net5369));
 sg13g2_buf_8 fanout5370 (.A(net5372),
    .X(net5370));
 sg13g2_buf_1 fanout5371 (.A(net5372),
    .X(net5371));
 sg13g2_buf_8 fanout5372 (.A(net5386),
    .X(net5372));
 sg13g2_buf_8 fanout5373 (.A(net5375),
    .X(net5373));
 sg13g2_buf_8 fanout5374 (.A(net5375),
    .X(net5374));
 sg13g2_buf_8 fanout5375 (.A(net5386),
    .X(net5375));
 sg13g2_buf_8 fanout5376 (.A(net5379),
    .X(net5376));
 sg13g2_buf_8 fanout5377 (.A(net5379),
    .X(net5377));
 sg13g2_buf_8 fanout5378 (.A(net5379),
    .X(net5378));
 sg13g2_buf_8 fanout5379 (.A(net5385),
    .X(net5379));
 sg13g2_buf_8 fanout5380 (.A(net5381),
    .X(net5380));
 sg13g2_buf_2 fanout5381 (.A(net5382),
    .X(net5381));
 sg13g2_buf_1 fanout5382 (.A(net5385),
    .X(net5382));
 sg13g2_buf_8 fanout5383 (.A(net5385),
    .X(net5383));
 sg13g2_buf_1 fanout5384 (.A(net5385),
    .X(net5384));
 sg13g2_buf_8 fanout5385 (.A(net5386),
    .X(net5385));
 sg13g2_buf_8 fanout5386 (.A(_06451_),
    .X(net5386));
 sg13g2_buf_8 fanout5387 (.A(net5389),
    .X(net5387));
 sg13g2_buf_8 fanout5388 (.A(net5389),
    .X(net5388));
 sg13g2_buf_8 fanout5389 (.A(net5407),
    .X(net5389));
 sg13g2_buf_8 fanout5390 (.A(net5391),
    .X(net5390));
 sg13g2_buf_8 fanout5391 (.A(net5392),
    .X(net5391));
 sg13g2_buf_8 fanout5392 (.A(net5407),
    .X(net5392));
 sg13g2_buf_8 fanout5393 (.A(net5396),
    .X(net5393));
 sg13g2_buf_8 fanout5394 (.A(net5395),
    .X(net5394));
 sg13g2_buf_8 fanout5395 (.A(net5396),
    .X(net5395));
 sg13g2_buf_8 fanout5396 (.A(net5407),
    .X(net5396));
 sg13g2_buf_8 fanout5397 (.A(net5400),
    .X(net5397));
 sg13g2_buf_8 fanout5398 (.A(net5400),
    .X(net5398));
 sg13g2_buf_1 fanout5399 (.A(net5400),
    .X(net5399));
 sg13g2_buf_8 fanout5400 (.A(net5407),
    .X(net5400));
 sg13g2_buf_8 fanout5401 (.A(net5402),
    .X(net5401));
 sg13g2_buf_8 fanout5402 (.A(net5406),
    .X(net5402));
 sg13g2_buf_8 fanout5403 (.A(net5404),
    .X(net5403));
 sg13g2_buf_2 fanout5404 (.A(net5405),
    .X(net5404));
 sg13g2_buf_8 fanout5405 (.A(net5406),
    .X(net5405));
 sg13g2_buf_8 fanout5406 (.A(net5407),
    .X(net5406));
 sg13g2_buf_8 fanout5407 (.A(net5431),
    .X(net5407));
 sg13g2_buf_8 fanout5408 (.A(net5409),
    .X(net5408));
 sg13g2_buf_8 fanout5409 (.A(net5416),
    .X(net5409));
 sg13g2_buf_8 fanout5410 (.A(net5416),
    .X(net5410));
 sg13g2_buf_8 fanout5411 (.A(net5413),
    .X(net5411));
 sg13g2_buf_8 fanout5412 (.A(net5413),
    .X(net5412));
 sg13g2_buf_8 fanout5413 (.A(net5415),
    .X(net5413));
 sg13g2_buf_8 fanout5414 (.A(net5415),
    .X(net5414));
 sg13g2_buf_8 fanout5415 (.A(net5416),
    .X(net5415));
 sg13g2_buf_8 fanout5416 (.A(net5431),
    .X(net5416));
 sg13g2_buf_8 fanout5417 (.A(net5423),
    .X(net5417));
 sg13g2_buf_1 fanout5418 (.A(net5423),
    .X(net5418));
 sg13g2_buf_8 fanout5419 (.A(net5423),
    .X(net5419));
 sg13g2_buf_8 fanout5420 (.A(net5421),
    .X(net5420));
 sg13g2_buf_8 fanout5421 (.A(net5422),
    .X(net5421));
 sg13g2_buf_8 fanout5422 (.A(net5423),
    .X(net5422));
 sg13g2_buf_8 fanout5423 (.A(net5431),
    .X(net5423));
 sg13g2_buf_8 fanout5424 (.A(net5430),
    .X(net5424));
 sg13g2_buf_8 fanout5425 (.A(net5426),
    .X(net5425));
 sg13g2_buf_8 fanout5426 (.A(net5430),
    .X(net5426));
 sg13g2_buf_8 fanout5427 (.A(net5428),
    .X(net5427));
 sg13g2_buf_8 fanout5428 (.A(net5429),
    .X(net5428));
 sg13g2_buf_8 fanout5429 (.A(net5430),
    .X(net5429));
 sg13g2_buf_8 fanout5430 (.A(net5431),
    .X(net5430));
 sg13g2_buf_8 fanout5431 (.A(_06450_),
    .X(net5431));
 sg13g2_buf_2 fanout5432 (.A(net5434),
    .X(net5432));
 sg13g2_buf_2 fanout5433 (.A(net5434),
    .X(net5433));
 sg13g2_buf_8 fanout5434 (.A(net5435),
    .X(net5434));
 sg13g2_buf_8 fanout5435 (.A(net5442),
    .X(net5435));
 sg13g2_buf_1 fanout5436 (.A(net5437),
    .X(net5436));
 sg13g2_buf_8 fanout5437 (.A(net5438),
    .X(net5437));
 sg13g2_buf_8 fanout5438 (.A(net5439),
    .X(net5438));
 sg13g2_buf_8 fanout5439 (.A(net5442),
    .X(net5439));
 sg13g2_buf_8 fanout5440 (.A(net5441),
    .X(net5440));
 sg13g2_buf_8 fanout5441 (.A(net5442),
    .X(net5441));
 sg13g2_buf_8 fanout5442 (.A(_19503_),
    .X(net5442));
 sg13g2_buf_8 fanout5443 (.A(net5444),
    .X(net5443));
 sg13g2_buf_8 fanout5444 (.A(net5447),
    .X(net5444));
 sg13g2_buf_8 fanout5445 (.A(net5446),
    .X(net5445));
 sg13g2_buf_8 fanout5446 (.A(net5447),
    .X(net5446));
 sg13g2_buf_8 fanout5447 (.A(net5453),
    .X(net5447));
 sg13g2_buf_2 fanout5448 (.A(net5449),
    .X(net5448));
 sg13g2_buf_1 fanout5449 (.A(net5450),
    .X(net5449));
 sg13g2_buf_2 fanout5450 (.A(net5453),
    .X(net5450));
 sg13g2_buf_8 fanout5451 (.A(net5453),
    .X(net5451));
 sg13g2_buf_1 fanout5452 (.A(net5453),
    .X(net5452));
 sg13g2_buf_8 fanout5453 (.A(_19503_),
    .X(net5453));
 sg13g2_buf_2 fanout5454 (.A(net5455),
    .X(net5454));
 sg13g2_buf_8 fanout5455 (.A(net5459),
    .X(net5455));
 sg13g2_buf_2 fanout5456 (.A(net5459),
    .X(net5456));
 sg13g2_buf_1 fanout5457 (.A(net5459),
    .X(net5457));
 sg13g2_buf_8 fanout5458 (.A(net5459),
    .X(net5458));
 sg13g2_buf_8 fanout5459 (.A(net5476),
    .X(net5459));
 sg13g2_buf_8 fanout5460 (.A(net5463),
    .X(net5460));
 sg13g2_buf_8 fanout5461 (.A(net5462),
    .X(net5461));
 sg13g2_buf_8 fanout5462 (.A(net5463),
    .X(net5462));
 sg13g2_buf_8 fanout5463 (.A(net5476),
    .X(net5463));
 sg13g2_buf_8 fanout5464 (.A(net5466),
    .X(net5464));
 sg13g2_buf_1 fanout5465 (.A(net5466),
    .X(net5465));
 sg13g2_buf_8 fanout5466 (.A(net5476),
    .X(net5466));
 sg13g2_buf_8 fanout5467 (.A(net5468),
    .X(net5467));
 sg13g2_buf_8 fanout5468 (.A(net5476),
    .X(net5468));
 sg13g2_buf_2 fanout5469 (.A(net5475),
    .X(net5469));
 sg13g2_buf_1 fanout5470 (.A(net5475),
    .X(net5470));
 sg13g2_buf_8 fanout5471 (.A(net5472),
    .X(net5471));
 sg13g2_buf_1 fanout5472 (.A(net5473),
    .X(net5472));
 sg13g2_buf_1 fanout5473 (.A(net5475),
    .X(net5473));
 sg13g2_buf_2 fanout5474 (.A(net5475),
    .X(net5474));
 sg13g2_buf_8 fanout5475 (.A(net5476),
    .X(net5475));
 sg13g2_buf_8 fanout5476 (.A(_19503_),
    .X(net5476));
 sg13g2_buf_8 fanout5477 (.A(net5478),
    .X(net5477));
 sg13g2_buf_1 fanout5478 (.A(net5480),
    .X(net5478));
 sg13g2_buf_8 fanout5479 (.A(net5480),
    .X(net5479));
 sg13g2_buf_2 fanout5480 (.A(net5492),
    .X(net5480));
 sg13g2_buf_8 fanout5481 (.A(net5482),
    .X(net5481));
 sg13g2_buf_8 fanout5482 (.A(net5492),
    .X(net5482));
 sg13g2_buf_8 fanout5483 (.A(net5484),
    .X(net5483));
 sg13g2_buf_8 fanout5484 (.A(net5492),
    .X(net5484));
 sg13g2_buf_8 fanout5485 (.A(net5487),
    .X(net5485));
 sg13g2_buf_1 fanout5486 (.A(net5487),
    .X(net5486));
 sg13g2_buf_8 fanout5487 (.A(net5488),
    .X(net5487));
 sg13g2_buf_2 fanout5488 (.A(net5491),
    .X(net5488));
 sg13g2_buf_8 fanout5489 (.A(net5490),
    .X(net5489));
 sg13g2_buf_8 fanout5490 (.A(net5491),
    .X(net5490));
 sg13g2_buf_8 fanout5491 (.A(net5492),
    .X(net5491));
 sg13g2_buf_8 fanout5492 (.A(net5526),
    .X(net5492));
 sg13g2_buf_8 fanout5493 (.A(net5494),
    .X(net5493));
 sg13g2_buf_8 fanout5494 (.A(net5502),
    .X(net5494));
 sg13g2_buf_8 fanout5495 (.A(net5496),
    .X(net5495));
 sg13g2_buf_8 fanout5496 (.A(net5502),
    .X(net5496));
 sg13g2_buf_8 fanout5497 (.A(net5498),
    .X(net5497));
 sg13g2_buf_8 fanout5498 (.A(net5499),
    .X(net5498));
 sg13g2_buf_2 fanout5499 (.A(net5502),
    .X(net5499));
 sg13g2_buf_8 fanout5500 (.A(net5501),
    .X(net5500));
 sg13g2_buf_8 fanout5501 (.A(net5502),
    .X(net5501));
 sg13g2_buf_8 fanout5502 (.A(net5526),
    .X(net5502));
 sg13g2_buf_8 fanout5503 (.A(net5512),
    .X(net5503));
 sg13g2_buf_1 fanout5504 (.A(net5512),
    .X(net5504));
 sg13g2_buf_8 fanout5505 (.A(net5507),
    .X(net5505));
 sg13g2_buf_1 fanout5506 (.A(net5507),
    .X(net5506));
 sg13g2_buf_8 fanout5507 (.A(net5512),
    .X(net5507));
 sg13g2_buf_8 fanout5508 (.A(net5509),
    .X(net5508));
 sg13g2_buf_8 fanout5509 (.A(net5512),
    .X(net5509));
 sg13g2_buf_8 fanout5510 (.A(net5512),
    .X(net5510));
 sg13g2_buf_1 fanout5511 (.A(net5512),
    .X(net5511));
 sg13g2_buf_8 fanout5512 (.A(net5526),
    .X(net5512));
 sg13g2_buf_8 fanout5513 (.A(net5515),
    .X(net5513));
 sg13g2_buf_1 fanout5514 (.A(net5515),
    .X(net5514));
 sg13g2_buf_8 fanout5515 (.A(net5525),
    .X(net5515));
 sg13g2_buf_8 fanout5516 (.A(net5525),
    .X(net5516));
 sg13g2_buf_1 fanout5517 (.A(net5525),
    .X(net5517));
 sg13g2_buf_8 fanout5518 (.A(net5525),
    .X(net5518));
 sg13g2_buf_1 fanout5519 (.A(net5525),
    .X(net5519));
 sg13g2_buf_8 fanout5520 (.A(net5521),
    .X(net5520));
 sg13g2_buf_2 fanout5521 (.A(net5522),
    .X(net5521));
 sg13g2_buf_1 fanout5522 (.A(net5524),
    .X(net5522));
 sg13g2_buf_8 fanout5523 (.A(net5524),
    .X(net5523));
 sg13g2_buf_2 fanout5524 (.A(net5525),
    .X(net5524));
 sg13g2_buf_8 fanout5525 (.A(net5526),
    .X(net5525));
 sg13g2_buf_8 fanout5526 (.A(_19502_),
    .X(net5526));
 sg13g2_buf_8 fanout5527 (.A(net5528),
    .X(net5527));
 sg13g2_buf_8 fanout5528 (.A(net5537),
    .X(net5528));
 sg13g2_buf_8 fanout5529 (.A(net5536),
    .X(net5529));
 sg13g2_buf_2 fanout5530 (.A(net5536),
    .X(net5530));
 sg13g2_buf_8 fanout5531 (.A(net5532),
    .X(net5531));
 sg13g2_buf_2 fanout5532 (.A(net5536),
    .X(net5532));
 sg13g2_buf_8 fanout5533 (.A(net5535),
    .X(net5533));
 sg13g2_buf_1 fanout5534 (.A(net5535),
    .X(net5534));
 sg13g2_buf_8 fanout5535 (.A(net5536),
    .X(net5535));
 sg13g2_buf_8 fanout5536 (.A(net5537),
    .X(net5536));
 sg13g2_buf_8 fanout5537 (.A(net5587),
    .X(net5537));
 sg13g2_buf_8 fanout5538 (.A(net5546),
    .X(net5538));
 sg13g2_buf_8 fanout5539 (.A(net5546),
    .X(net5539));
 sg13g2_buf_8 fanout5540 (.A(net5546),
    .X(net5540));
 sg13g2_buf_1 fanout5541 (.A(net5542),
    .X(net5541));
 sg13g2_buf_8 fanout5542 (.A(net5546),
    .X(net5542));
 sg13g2_buf_8 fanout5543 (.A(net5544),
    .X(net5543));
 sg13g2_buf_8 fanout5544 (.A(net5545),
    .X(net5544));
 sg13g2_buf_8 fanout5545 (.A(net5546),
    .X(net5545));
 sg13g2_buf_8 fanout5546 (.A(net5587),
    .X(net5546));
 sg13g2_buf_8 fanout5547 (.A(net5549),
    .X(net5547));
 sg13g2_buf_1 fanout5548 (.A(net5549),
    .X(net5548));
 sg13g2_buf_8 fanout5549 (.A(net5556),
    .X(net5549));
 sg13g2_buf_8 fanout5550 (.A(net5552),
    .X(net5550));
 sg13g2_buf_1 fanout5551 (.A(net5552),
    .X(net5551));
 sg13g2_buf_8 fanout5552 (.A(net5556),
    .X(net5552));
 sg13g2_buf_8 fanout5553 (.A(net5556),
    .X(net5553));
 sg13g2_buf_1 fanout5554 (.A(net5555),
    .X(net5554));
 sg13g2_buf_8 fanout5555 (.A(net5556),
    .X(net5555));
 sg13g2_buf_8 fanout5556 (.A(net5587),
    .X(net5556));
 sg13g2_buf_8 fanout5557 (.A(net5558),
    .X(net5557));
 sg13g2_buf_8 fanout5558 (.A(net5570),
    .X(net5558));
 sg13g2_buf_8 fanout5559 (.A(net5561),
    .X(net5559));
 sg13g2_buf_1 fanout5560 (.A(net5561),
    .X(net5560));
 sg13g2_buf_8 fanout5561 (.A(net5570),
    .X(net5561));
 sg13g2_buf_8 fanout5562 (.A(net5563),
    .X(net5562));
 sg13g2_buf_8 fanout5563 (.A(net5570),
    .X(net5563));
 sg13g2_buf_8 fanout5564 (.A(net5569),
    .X(net5564));
 sg13g2_buf_8 fanout5565 (.A(net5566),
    .X(net5565));
 sg13g2_buf_8 fanout5566 (.A(net5569),
    .X(net5566));
 sg13g2_buf_8 fanout5567 (.A(net5568),
    .X(net5567));
 sg13g2_buf_8 fanout5568 (.A(net5569),
    .X(net5568));
 sg13g2_buf_8 fanout5569 (.A(net5570),
    .X(net5569));
 sg13g2_buf_8 fanout5570 (.A(net5587),
    .X(net5570));
 sg13g2_buf_8 fanout5571 (.A(net5572),
    .X(net5571));
 sg13g2_buf_8 fanout5572 (.A(net5586),
    .X(net5572));
 sg13g2_buf_8 fanout5573 (.A(net5574),
    .X(net5573));
 sg13g2_buf_8 fanout5574 (.A(net5586),
    .X(net5574));
 sg13g2_buf_8 fanout5575 (.A(net5577),
    .X(net5575));
 sg13g2_buf_1 fanout5576 (.A(net5577),
    .X(net5576));
 sg13g2_buf_8 fanout5577 (.A(net5586),
    .X(net5577));
 sg13g2_buf_8 fanout5578 (.A(net5585),
    .X(net5578));
 sg13g2_buf_8 fanout5579 (.A(net5585),
    .X(net5579));
 sg13g2_buf_8 fanout5580 (.A(net5581),
    .X(net5580));
 sg13g2_buf_8 fanout5581 (.A(net5585),
    .X(net5581));
 sg13g2_buf_8 fanout5582 (.A(net5584),
    .X(net5582));
 sg13g2_buf_8 fanout5583 (.A(net5584),
    .X(net5583));
 sg13g2_buf_8 fanout5584 (.A(net5585),
    .X(net5584));
 sg13g2_buf_8 fanout5585 (.A(net5586),
    .X(net5585));
 sg13g2_buf_8 fanout5586 (.A(net5587),
    .X(net5586));
 sg13g2_buf_8 fanout5587 (.A(_19027_),
    .X(net5587));
 sg13g2_buf_8 fanout5588 (.A(net5592),
    .X(net5588));
 sg13g2_buf_8 fanout5589 (.A(net5592),
    .X(net5589));
 sg13g2_buf_8 fanout5590 (.A(net5592),
    .X(net5590));
 sg13g2_buf_1 fanout5591 (.A(net5592),
    .X(net5591));
 sg13g2_buf_8 fanout5592 (.A(net5599),
    .X(net5592));
 sg13g2_buf_8 fanout5593 (.A(net5594),
    .X(net5593));
 sg13g2_buf_8 fanout5594 (.A(net5599),
    .X(net5594));
 sg13g2_buf_8 fanout5595 (.A(net5599),
    .X(net5595));
 sg13g2_buf_8 fanout5596 (.A(net5599),
    .X(net5596));
 sg13g2_buf_8 fanout5597 (.A(net5598),
    .X(net5597));
 sg13g2_buf_8 fanout5598 (.A(net5599),
    .X(net5598));
 sg13g2_buf_8 fanout5599 (.A(net5615),
    .X(net5599));
 sg13g2_buf_8 fanout5600 (.A(net5601),
    .X(net5600));
 sg13g2_buf_8 fanout5601 (.A(net5615),
    .X(net5601));
 sg13g2_buf_8 fanout5602 (.A(net5603),
    .X(net5602));
 sg13g2_buf_8 fanout5603 (.A(net5605),
    .X(net5603));
 sg13g2_buf_8 fanout5604 (.A(net5605),
    .X(net5604));
 sg13g2_buf_8 fanout5605 (.A(net5615),
    .X(net5605));
 sg13g2_buf_8 fanout5606 (.A(net5607),
    .X(net5606));
 sg13g2_buf_8 fanout5607 (.A(net5614),
    .X(net5607));
 sg13g2_buf_8 fanout5608 (.A(net5614),
    .X(net5608));
 sg13g2_buf_1 fanout5609 (.A(net5614),
    .X(net5609));
 sg13g2_buf_8 fanout5610 (.A(net5613),
    .X(net5610));
 sg13g2_buf_1 fanout5611 (.A(net5613),
    .X(net5611));
 sg13g2_buf_8 fanout5612 (.A(net5613),
    .X(net5612));
 sg13g2_buf_8 fanout5613 (.A(net5614),
    .X(net5613));
 sg13g2_buf_8 fanout5614 (.A(net5615),
    .X(net5614));
 sg13g2_buf_8 fanout5615 (.A(_19026_),
    .X(net5615));
 sg13g2_buf_8 fanout5616 (.A(_05559_),
    .X(net5616));
 sg13g2_buf_8 fanout5617 (.A(_05266_),
    .X(net5617));
 sg13g2_buf_8 fanout5618 (.A(_05222_),
    .X(net5618));
 sg13g2_buf_2 fanout5619 (.A(_04882_),
    .X(net5619));
 sg13g2_buf_8 fanout5620 (.A(_15407_),
    .X(net5620));
 sg13g2_buf_8 fanout5621 (.A(_15325_),
    .X(net5621));
 sg13g2_buf_8 fanout5622 (.A(_14927_),
    .X(net5622));
 sg13g2_buf_2 fanout5623 (.A(_14926_),
    .X(net5623));
 sg13g2_buf_8 fanout5624 (.A(net5626),
    .X(net5624));
 sg13g2_buf_1 fanout5625 (.A(net5626),
    .X(net5625));
 sg13g2_buf_8 fanout5626 (.A(net5631),
    .X(net5626));
 sg13g2_buf_8 fanout5627 (.A(net5628),
    .X(net5627));
 sg13g2_buf_2 fanout5628 (.A(net5631),
    .X(net5628));
 sg13g2_buf_8 fanout5629 (.A(net5631),
    .X(net5629));
 sg13g2_buf_8 fanout5630 (.A(net5631),
    .X(net5630));
 sg13g2_buf_8 fanout5631 (.A(net3379),
    .X(net5631));
 sg13g2_buf_8 fanout5632 (.A(net5633),
    .X(net5632));
 sg13g2_buf_1 fanout5633 (.A(net5634),
    .X(net5633));
 sg13g2_buf_8 fanout5634 (.A(_14827_),
    .X(net5634));
 sg13g2_buf_8 fanout5635 (.A(net5637),
    .X(net5635));
 sg13g2_buf_1 fanout5636 (.A(net5637),
    .X(net5636));
 sg13g2_buf_8 fanout5637 (.A(net5639),
    .X(net5637));
 sg13g2_buf_8 fanout5638 (.A(net5639),
    .X(net5638));
 sg13g2_buf_8 fanout5639 (.A(net5648),
    .X(net5639));
 sg13g2_buf_8 fanout5640 (.A(net5642),
    .X(net5640));
 sg13g2_buf_8 fanout5641 (.A(net5642),
    .X(net5641));
 sg13g2_buf_8 fanout5642 (.A(net5648),
    .X(net5642));
 sg13g2_buf_8 fanout5643 (.A(net5644),
    .X(net5643));
 sg13g2_buf_1 fanout5644 (.A(net5645),
    .X(net5644));
 sg13g2_buf_8 fanout5645 (.A(net5646),
    .X(net5645));
 sg13g2_buf_8 fanout5646 (.A(net5648),
    .X(net5646));
 sg13g2_buf_8 fanout5647 (.A(net5648),
    .X(net5647));
 sg13g2_buf_8 fanout5648 (.A(_14510_),
    .X(net5648));
 sg13g2_buf_8 fanout5649 (.A(net5653),
    .X(net5649));
 sg13g2_buf_8 fanout5650 (.A(net5653),
    .X(net5650));
 sg13g2_buf_8 fanout5651 (.A(net5653),
    .X(net5651));
 sg13g2_buf_1 fanout5652 (.A(net5653),
    .X(net5652));
 sg13g2_buf_8 fanout5653 (.A(net5655),
    .X(net5653));
 sg13g2_buf_8 fanout5654 (.A(net5655),
    .X(net5654));
 sg13g2_buf_8 fanout5655 (.A(net5667),
    .X(net5655));
 sg13g2_buf_8 fanout5656 (.A(net5667),
    .X(net5656));
 sg13g2_buf_8 fanout5657 (.A(net5658),
    .X(net5657));
 sg13g2_buf_8 fanout5658 (.A(net5662),
    .X(net5658));
 sg13g2_buf_8 fanout5659 (.A(net5662),
    .X(net5659));
 sg13g2_buf_1 fanout5660 (.A(net5662),
    .X(net5660));
 sg13g2_buf_8 fanout5661 (.A(net5662),
    .X(net5661));
 sg13g2_buf_8 fanout5662 (.A(net5667),
    .X(net5662));
 sg13g2_buf_8 fanout5663 (.A(net5664),
    .X(net5663));
 sg13g2_buf_8 fanout5664 (.A(net5667),
    .X(net5664));
 sg13g2_buf_8 fanout5665 (.A(net5666),
    .X(net5665));
 sg13g2_buf_8 fanout5666 (.A(net5667),
    .X(net5666));
 sg13g2_buf_8 fanout5667 (.A(net5683),
    .X(net5667));
 sg13g2_buf_8 fanout5668 (.A(net5671),
    .X(net5668));
 sg13g2_buf_8 fanout5669 (.A(net5670),
    .X(net5669));
 sg13g2_buf_8 fanout5670 (.A(net5671),
    .X(net5670));
 sg13g2_buf_8 fanout5671 (.A(net5683),
    .X(net5671));
 sg13g2_buf_8 fanout5672 (.A(net5673),
    .X(net5672));
 sg13g2_buf_8 fanout5673 (.A(net5674),
    .X(net5673));
 sg13g2_buf_8 fanout5674 (.A(net5683),
    .X(net5674));
 sg13g2_buf_8 fanout5675 (.A(net5679),
    .X(net5675));
 sg13g2_buf_1 fanout5676 (.A(net5679),
    .X(net5676));
 sg13g2_buf_8 fanout5677 (.A(net5679),
    .X(net5677));
 sg13g2_buf_8 fanout5678 (.A(net5679),
    .X(net5678));
 sg13g2_buf_8 fanout5679 (.A(net5682),
    .X(net5679));
 sg13g2_buf_8 fanout5680 (.A(net5681),
    .X(net5680));
 sg13g2_buf_8 fanout5681 (.A(net5682),
    .X(net5681));
 sg13g2_buf_8 fanout5682 (.A(net5683),
    .X(net5682));
 sg13g2_buf_8 fanout5683 (.A(_14171_),
    .X(net5683));
 sg13g2_buf_8 fanout5684 (.A(net5688),
    .X(net5684));
 sg13g2_buf_2 fanout5685 (.A(net5688),
    .X(net5685));
 sg13g2_buf_8 fanout5686 (.A(net5687),
    .X(net5686));
 sg13g2_buf_8 fanout5687 (.A(net5688),
    .X(net5687));
 sg13g2_buf_8 fanout5688 (.A(net5717),
    .X(net5688));
 sg13g2_buf_8 fanout5689 (.A(net5692),
    .X(net5689));
 sg13g2_buf_8 fanout5690 (.A(net5692),
    .X(net5690));
 sg13g2_buf_1 fanout5691 (.A(net5692),
    .X(net5691));
 sg13g2_buf_8 fanout5692 (.A(net5717),
    .X(net5692));
 sg13g2_buf_8 fanout5693 (.A(net5699),
    .X(net5693));
 sg13g2_buf_1 fanout5694 (.A(net5699),
    .X(net5694));
 sg13g2_buf_8 fanout5695 (.A(net5696),
    .X(net5695));
 sg13g2_buf_8 fanout5696 (.A(net5699),
    .X(net5696));
 sg13g2_buf_8 fanout5697 (.A(net5698),
    .X(net5697));
 sg13g2_buf_8 fanout5698 (.A(net5699),
    .X(net5698));
 sg13g2_buf_8 fanout5699 (.A(net5717),
    .X(net5699));
 sg13g2_buf_8 fanout5700 (.A(net5701),
    .X(net5700));
 sg13g2_buf_8 fanout5701 (.A(net5705),
    .X(net5701));
 sg13g2_buf_8 fanout5702 (.A(net5704),
    .X(net5702));
 sg13g2_buf_8 fanout5703 (.A(net5705),
    .X(net5703));
 sg13g2_buf_1 fanout5704 (.A(net5705),
    .X(net5704));
 sg13g2_buf_8 fanout5705 (.A(net5708),
    .X(net5705));
 sg13g2_buf_8 fanout5706 (.A(net5707),
    .X(net5706));
 sg13g2_buf_8 fanout5707 (.A(net5708),
    .X(net5707));
 sg13g2_buf_8 fanout5708 (.A(net5716),
    .X(net5708));
 sg13g2_buf_8 fanout5709 (.A(net5711),
    .X(net5709));
 sg13g2_buf_1 fanout5710 (.A(net5711),
    .X(net5710));
 sg13g2_buf_8 fanout5711 (.A(net5715),
    .X(net5711));
 sg13g2_buf_8 fanout5712 (.A(net5714),
    .X(net5712));
 sg13g2_buf_1 fanout5713 (.A(net5714),
    .X(net5713));
 sg13g2_buf_8 fanout5714 (.A(net5715),
    .X(net5714));
 sg13g2_buf_8 fanout5715 (.A(net5716),
    .X(net5715));
 sg13g2_buf_8 fanout5716 (.A(net5717),
    .X(net5716));
 sg13g2_buf_8 fanout5717 (.A(_14171_),
    .X(net5717));
 sg13g2_buf_8 fanout5718 (.A(net5719),
    .X(net5718));
 sg13g2_buf_8 fanout5719 (.A(net5723),
    .X(net5719));
 sg13g2_buf_8 fanout5720 (.A(net5722),
    .X(net5720));
 sg13g2_buf_1 fanout5721 (.A(net5722),
    .X(net5721));
 sg13g2_buf_8 fanout5722 (.A(net5723),
    .X(net5722));
 sg13g2_buf_8 fanout5723 (.A(net5743),
    .X(net5723));
 sg13g2_buf_8 fanout5724 (.A(net5726),
    .X(net5724));
 sg13g2_buf_8 fanout5725 (.A(net5726),
    .X(net5725));
 sg13g2_buf_8 fanout5726 (.A(net5743),
    .X(net5726));
 sg13g2_buf_8 fanout5727 (.A(net5729),
    .X(net5727));
 sg13g2_buf_2 fanout5728 (.A(net5729),
    .X(net5728));
 sg13g2_buf_8 fanout5729 (.A(net5730),
    .X(net5729));
 sg13g2_buf_8 fanout5730 (.A(net5743),
    .X(net5730));
 sg13g2_buf_8 fanout5731 (.A(net5742),
    .X(net5731));
 sg13g2_buf_1 fanout5732 (.A(net5742),
    .X(net5732));
 sg13g2_buf_8 fanout5733 (.A(net5742),
    .X(net5733));
 sg13g2_buf_8 fanout5734 (.A(net5737),
    .X(net5734));
 sg13g2_buf_8 fanout5735 (.A(net5737),
    .X(net5735));
 sg13g2_buf_8 fanout5736 (.A(net5737),
    .X(net5736));
 sg13g2_buf_8 fanout5737 (.A(net5741),
    .X(net5737));
 sg13g2_buf_8 fanout5738 (.A(net5739),
    .X(net5738));
 sg13g2_buf_8 fanout5739 (.A(net5741),
    .X(net5739));
 sg13g2_buf_8 fanout5740 (.A(net5741),
    .X(net5740));
 sg13g2_buf_8 fanout5741 (.A(net5742),
    .X(net5741));
 sg13g2_buf_8 fanout5742 (.A(net5743),
    .X(net5742));
 sg13g2_buf_8 fanout5743 (.A(net5771),
    .X(net5743));
 sg13g2_buf_8 fanout5744 (.A(net5745),
    .X(net5744));
 sg13g2_buf_8 fanout5745 (.A(net5748),
    .X(net5745));
 sg13g2_buf_8 fanout5746 (.A(net5748),
    .X(net5746));
 sg13g2_buf_8 fanout5747 (.A(net5748),
    .X(net5747));
 sg13g2_buf_8 fanout5748 (.A(net5771),
    .X(net5748));
 sg13g2_buf_8 fanout5749 (.A(net5757),
    .X(net5749));
 sg13g2_buf_1 fanout5750 (.A(net5757),
    .X(net5750));
 sg13g2_buf_8 fanout5751 (.A(net5752),
    .X(net5751));
 sg13g2_buf_8 fanout5752 (.A(net5757),
    .X(net5752));
 sg13g2_buf_8 fanout5753 (.A(net5756),
    .X(net5753));
 sg13g2_buf_8 fanout5754 (.A(net5755),
    .X(net5754));
 sg13g2_buf_8 fanout5755 (.A(net5756),
    .X(net5755));
 sg13g2_buf_8 fanout5756 (.A(net5757),
    .X(net5756));
 sg13g2_buf_8 fanout5757 (.A(net5771),
    .X(net5757));
 sg13g2_buf_8 fanout5758 (.A(net5759),
    .X(net5758));
 sg13g2_buf_2 fanout5759 (.A(net5770),
    .X(net5759));
 sg13g2_buf_8 fanout5760 (.A(net5770),
    .X(net5760));
 sg13g2_buf_8 fanout5761 (.A(net5770),
    .X(net5761));
 sg13g2_buf_8 fanout5762 (.A(net5764),
    .X(net5762));
 sg13g2_buf_8 fanout5763 (.A(net5764),
    .X(net5763));
 sg13g2_buf_8 fanout5764 (.A(net5769),
    .X(net5764));
 sg13g2_buf_8 fanout5765 (.A(net5769),
    .X(net5765));
 sg13g2_buf_8 fanout5766 (.A(net5769),
    .X(net5766));
 sg13g2_buf_8 fanout5767 (.A(net5769),
    .X(net5767));
 sg13g2_buf_8 fanout5768 (.A(net5769),
    .X(net5768));
 sg13g2_buf_8 fanout5769 (.A(net5770),
    .X(net5769));
 sg13g2_buf_8 fanout5770 (.A(net5771),
    .X(net5770));
 sg13g2_buf_8 fanout5771 (.A(\u_inv.f_next[0] ),
    .X(net5771));
 sg13g2_buf_8 fanout5772 (.A(net5773),
    .X(net5772));
 sg13g2_buf_8 fanout5773 (.A(net5799),
    .X(net5773));
 sg13g2_buf_8 fanout5774 (.A(net5776),
    .X(net5774));
 sg13g2_buf_8 fanout5775 (.A(net5776),
    .X(net5775));
 sg13g2_buf_8 fanout5776 (.A(net5799),
    .X(net5776));
 sg13g2_buf_8 fanout5777 (.A(net5778),
    .X(net5777));
 sg13g2_buf_8 fanout5778 (.A(net5785),
    .X(net5778));
 sg13g2_buf_1 fanout5779 (.A(net5785),
    .X(net5779));
 sg13g2_buf_8 fanout5780 (.A(net5785),
    .X(net5780));
 sg13g2_buf_8 fanout5781 (.A(net5784),
    .X(net5781));
 sg13g2_buf_8 fanout5782 (.A(net5784),
    .X(net5782));
 sg13g2_buf_1 fanout5783 (.A(net5784),
    .X(net5783));
 sg13g2_buf_8 fanout5784 (.A(net5785),
    .X(net5784));
 sg13g2_buf_8 fanout5785 (.A(net5799),
    .X(net5785));
 sg13g2_buf_8 fanout5786 (.A(net5787),
    .X(net5786));
 sg13g2_buf_8 fanout5787 (.A(net5799),
    .X(net5787));
 sg13g2_buf_8 fanout5788 (.A(net5789),
    .X(net5788));
 sg13g2_buf_8 fanout5789 (.A(net5790),
    .X(net5789));
 sg13g2_buf_8 fanout5790 (.A(net5799),
    .X(net5790));
 sg13g2_buf_8 fanout5791 (.A(net5798),
    .X(net5791));
 sg13g2_buf_8 fanout5792 (.A(net5798),
    .X(net5792));
 sg13g2_buf_8 fanout5793 (.A(net5798),
    .X(net5793));
 sg13g2_buf_8 fanout5794 (.A(net5796),
    .X(net5794));
 sg13g2_buf_1 fanout5795 (.A(net5796),
    .X(net5795));
 sg13g2_buf_8 fanout5796 (.A(net5797),
    .X(net5796));
 sg13g2_buf_8 fanout5797 (.A(net5798),
    .X(net5797));
 sg13g2_buf_8 fanout5798 (.A(net5799),
    .X(net5798));
 sg13g2_buf_8 fanout5799 (.A(\u_inv.f_next[0] ),
    .X(net5799));
 sg13g2_buf_8 fanout5800 (.A(net5804),
    .X(net5800));
 sg13g2_buf_8 fanout5801 (.A(net5804),
    .X(net5801));
 sg13g2_buf_8 fanout5802 (.A(net5804),
    .X(net5802));
 sg13g2_buf_1 fanout5803 (.A(net5804),
    .X(net5803));
 sg13g2_buf_8 fanout5804 (.A(net5811),
    .X(net5804));
 sg13g2_buf_8 fanout5805 (.A(net5806),
    .X(net5805));
 sg13g2_buf_8 fanout5806 (.A(net5811),
    .X(net5806));
 sg13g2_buf_8 fanout5807 (.A(net5808),
    .X(net5807));
 sg13g2_buf_1 fanout5808 (.A(net5809),
    .X(net5808));
 sg13g2_buf_8 fanout5809 (.A(net5811),
    .X(net5809));
 sg13g2_buf_8 fanout5810 (.A(net5811),
    .X(net5810));
 sg13g2_buf_8 fanout5811 (.A(net5828),
    .X(net5811));
 sg13g2_buf_8 fanout5812 (.A(net5814),
    .X(net5812));
 sg13g2_buf_2 fanout5813 (.A(net5814),
    .X(net5813));
 sg13g2_buf_8 fanout5814 (.A(net5828),
    .X(net5814));
 sg13g2_buf_8 fanout5815 (.A(net5817),
    .X(net5815));
 sg13g2_buf_2 fanout5816 (.A(net5817),
    .X(net5816));
 sg13g2_buf_8 fanout5817 (.A(net5828),
    .X(net5817));
 sg13g2_buf_8 fanout5818 (.A(net5827),
    .X(net5818));
 sg13g2_buf_1 fanout5819 (.A(net5827),
    .X(net5819));
 sg13g2_buf_8 fanout5820 (.A(net5827),
    .X(net5820));
 sg13g2_buf_8 fanout5821 (.A(net5823),
    .X(net5821));
 sg13g2_buf_1 fanout5822 (.A(net5823),
    .X(net5822));
 sg13g2_buf_8 fanout5823 (.A(net5827),
    .X(net5823));
 sg13g2_buf_8 fanout5824 (.A(net5826),
    .X(net5824));
 sg13g2_buf_1 fanout5825 (.A(net5826),
    .X(net5825));
 sg13g2_buf_8 fanout5826 (.A(net5827),
    .X(net5826));
 sg13g2_buf_8 fanout5827 (.A(net5828),
    .X(net5827));
 sg13g2_buf_8 fanout5828 (.A(\u_inv.f_next[0] ),
    .X(net5828));
 sg13g2_buf_8 fanout5829 (.A(net3432),
    .X(net5829));
 sg13g2_buf_8 fanout5830 (.A(net5831),
    .X(net5830));
 sg13g2_buf_8 fanout5831 (.A(net5832),
    .X(net5831));
 sg13g2_buf_8 fanout5832 (.A(net5833),
    .X(net5832));
 sg13g2_buf_8 fanout5833 (.A(net5847),
    .X(net5833));
 sg13g2_buf_8 fanout5834 (.A(net5838),
    .X(net5834));
 sg13g2_buf_1 fanout5835 (.A(net5838),
    .X(net5835));
 sg13g2_buf_8 fanout5836 (.A(net5838),
    .X(net5836));
 sg13g2_buf_1 fanout5837 (.A(net5838),
    .X(net5837));
 sg13g2_buf_8 fanout5838 (.A(net5839),
    .X(net5838));
 sg13g2_buf_8 fanout5839 (.A(net5847),
    .X(net5839));
 sg13g2_buf_8 fanout5840 (.A(net5843),
    .X(net5840));
 sg13g2_buf_8 fanout5841 (.A(net5842),
    .X(net5841));
 sg13g2_buf_8 fanout5842 (.A(net5843),
    .X(net5842));
 sg13g2_buf_8 fanout5843 (.A(net5847),
    .X(net5843));
 sg13g2_buf_8 fanout5844 (.A(net5845),
    .X(net5844));
 sg13g2_buf_2 fanout5845 (.A(net5846),
    .X(net5845));
 sg13g2_buf_8 fanout5846 (.A(net5847),
    .X(net5846));
 sg13g2_buf_8 fanout5847 (.A(net5864),
    .X(net5847));
 sg13g2_buf_8 fanout5848 (.A(net5850),
    .X(net5848));
 sg13g2_buf_8 fanout5849 (.A(net5850),
    .X(net5849));
 sg13g2_buf_8 fanout5850 (.A(net5855),
    .X(net5850));
 sg13g2_buf_8 fanout5851 (.A(net5852),
    .X(net5851));
 sg13g2_buf_8 fanout5852 (.A(net5854),
    .X(net5852));
 sg13g2_buf_8 fanout5853 (.A(net5854),
    .X(net5853));
 sg13g2_buf_8 fanout5854 (.A(net5855),
    .X(net5854));
 sg13g2_buf_8 fanout5855 (.A(net5864),
    .X(net5855));
 sg13g2_buf_8 fanout5856 (.A(net5858),
    .X(net5856));
 sg13g2_buf_1 fanout5857 (.A(net5858),
    .X(net5857));
 sg13g2_buf_8 fanout5858 (.A(net5859),
    .X(net5858));
 sg13g2_buf_8 fanout5859 (.A(net5864),
    .X(net5859));
 sg13g2_buf_8 fanout5860 (.A(net5863),
    .X(net5860));
 sg13g2_buf_8 fanout5861 (.A(net5863),
    .X(net5861));
 sg13g2_buf_8 fanout5862 (.A(net5863),
    .X(net5862));
 sg13g2_buf_8 fanout5863 (.A(net5864),
    .X(net5863));
 sg13g2_buf_8 fanout5864 (.A(\u_inv.f_reg[256] ),
    .X(net5864));
 sg13g2_buf_8 fanout5865 (.A(net2898),
    .X(net5865));
 sg13g2_buf_8 fanout5866 (.A(\u_inv.d_reg[184] ),
    .X(net5866));
 sg13g2_buf_8 fanout5867 (.A(\u_inv.d_reg[164] ),
    .X(net5867));
 sg13g2_buf_8 fanout5868 (.A(net2782),
    .X(net5868));
 sg13g2_buf_8 fanout5869 (.A(\u_inv.d_reg[140] ),
    .X(net5869));
 sg13g2_buf_8 fanout5870 (.A(\u_inv.d_reg[98] ),
    .X(net5870));
 sg13g2_buf_8 fanout5871 (.A(net3153),
    .X(net5871));
 sg13g2_buf_8 fanout5872 (.A(\u_inv.d_reg[77] ),
    .X(net5872));
 sg13g2_buf_8 fanout5873 (.A(\u_inv.d_reg[16] ),
    .X(net5873));
 sg13g2_buf_8 fanout5874 (.A(\u_inv.d_reg[11] ),
    .X(net5874));
 sg13g2_buf_8 fanout5875 (.A(net1331),
    .X(net5875));
 sg13g2_buf_8 fanout5876 (.A(net1222),
    .X(net5876));
 sg13g2_buf_8 fanout5877 (.A(net1359),
    .X(net5877));
 sg13g2_buf_8 fanout5878 (.A(net3418),
    .X(net5878));
 sg13g2_buf_8 fanout5879 (.A(net1406),
    .X(net5879));
 sg13g2_buf_8 fanout5880 (.A(net1260),
    .X(net5880));
 sg13g2_buf_8 fanout5881 (.A(net3427),
    .X(net5881));
 sg13g2_buf_8 fanout5882 (.A(net3435),
    .X(net5882));
 sg13g2_buf_8 fanout5883 (.A(net5884),
    .X(net5883));
 sg13g2_buf_8 fanout5884 (.A(net5928),
    .X(net5884));
 sg13g2_buf_8 fanout5885 (.A(net5886),
    .X(net5885));
 sg13g2_buf_8 fanout5886 (.A(net5887),
    .X(net5886));
 sg13g2_buf_8 fanout5887 (.A(net5928),
    .X(net5887));
 sg13g2_buf_8 fanout5888 (.A(net5892),
    .X(net5888));
 sg13g2_buf_8 fanout5889 (.A(net5891),
    .X(net5889));
 sg13g2_buf_2 fanout5890 (.A(net5891),
    .X(net5890));
 sg13g2_buf_8 fanout5891 (.A(net5892),
    .X(net5891));
 sg13g2_buf_8 fanout5892 (.A(net5906),
    .X(net5892));
 sg13g2_buf_8 fanout5893 (.A(net5895),
    .X(net5893));
 sg13g2_buf_8 fanout5894 (.A(net5895),
    .X(net5894));
 sg13g2_buf_8 fanout5895 (.A(net5899),
    .X(net5895));
 sg13g2_buf_8 fanout5896 (.A(net5899),
    .X(net5896));
 sg13g2_buf_8 fanout5897 (.A(net5898),
    .X(net5897));
 sg13g2_buf_8 fanout5898 (.A(net5899),
    .X(net5898));
 sg13g2_buf_8 fanout5899 (.A(net5906),
    .X(net5899));
 sg13g2_buf_8 fanout5900 (.A(net5901),
    .X(net5900));
 sg13g2_buf_8 fanout5901 (.A(net5902),
    .X(net5901));
 sg13g2_buf_8 fanout5902 (.A(net5906),
    .X(net5902));
 sg13g2_buf_8 fanout5903 (.A(net5905),
    .X(net5903));
 sg13g2_buf_8 fanout5904 (.A(net5905),
    .X(net5904));
 sg13g2_buf_8 fanout5905 (.A(net5906),
    .X(net5905));
 sg13g2_buf_8 fanout5906 (.A(net5928),
    .X(net5906));
 sg13g2_buf_8 fanout5907 (.A(net5915),
    .X(net5907));
 sg13g2_buf_1 fanout5908 (.A(net5915),
    .X(net5908));
 sg13g2_buf_8 fanout5909 (.A(net5910),
    .X(net5909));
 sg13g2_buf_8 fanout5910 (.A(net5912),
    .X(net5910));
 sg13g2_buf_8 fanout5911 (.A(net5912),
    .X(net5911));
 sg13g2_buf_8 fanout5912 (.A(net5915),
    .X(net5912));
 sg13g2_buf_8 fanout5913 (.A(net5914),
    .X(net5913));
 sg13g2_buf_8 fanout5914 (.A(net5915),
    .X(net5914));
 sg13g2_buf_8 fanout5915 (.A(net5928),
    .X(net5915));
 sg13g2_buf_8 fanout5916 (.A(net5927),
    .X(net5916));
 sg13g2_buf_8 fanout5917 (.A(net5927),
    .X(net5917));
 sg13g2_buf_8 fanout5918 (.A(net5920),
    .X(net5918));
 sg13g2_buf_2 fanout5919 (.A(net5920),
    .X(net5919));
 sg13g2_buf_8 fanout5920 (.A(net5927),
    .X(net5920));
 sg13g2_buf_8 fanout5921 (.A(net5922),
    .X(net5921));
 sg13g2_buf_8 fanout5922 (.A(net5926),
    .X(net5922));
 sg13g2_buf_8 fanout5923 (.A(net5926),
    .X(net5923));
 sg13g2_buf_2 fanout5924 (.A(net5925),
    .X(net5924));
 sg13g2_buf_8 fanout5925 (.A(net5926),
    .X(net5925));
 sg13g2_buf_8 fanout5926 (.A(net5927),
    .X(net5926));
 sg13g2_buf_8 fanout5927 (.A(net5928),
    .X(net5927));
 sg13g2_buf_8 fanout5928 (.A(rst_n),
    .X(net5928));
 sg13g2_buf_8 fanout5929 (.A(net5931),
    .X(net5929));
 sg13g2_buf_8 fanout5930 (.A(net5931),
    .X(net5930));
 sg13g2_buf_8 fanout5931 (.A(net5932),
    .X(net5931));
 sg13g2_buf_8 fanout5932 (.A(net5945),
    .X(net5932));
 sg13g2_buf_8 fanout5933 (.A(net5935),
    .X(net5933));
 sg13g2_buf_8 fanout5934 (.A(net5935),
    .X(net5934));
 sg13g2_buf_8 fanout5935 (.A(net5945),
    .X(net5935));
 sg13g2_buf_8 fanout5936 (.A(net5937),
    .X(net5936));
 sg13g2_buf_8 fanout5937 (.A(net5945),
    .X(net5937));
 sg13g2_buf_8 fanout5938 (.A(net5939),
    .X(net5938));
 sg13g2_buf_8 fanout5939 (.A(net5945),
    .X(net5939));
 sg13g2_buf_8 fanout5940 (.A(net5944),
    .X(net5940));
 sg13g2_buf_8 fanout5941 (.A(net5944),
    .X(net5941));
 sg13g2_buf_8 fanout5942 (.A(net5944),
    .X(net5942));
 sg13g2_buf_8 fanout5943 (.A(net5944),
    .X(net5943));
 sg13g2_buf_8 fanout5944 (.A(net5945),
    .X(net5944));
 sg13g2_buf_8 fanout5945 (.A(net5965),
    .X(net5945));
 sg13g2_buf_8 fanout5946 (.A(net5947),
    .X(net5946));
 sg13g2_buf_8 fanout5947 (.A(net5949),
    .X(net5947));
 sg13g2_buf_8 fanout5948 (.A(net5949),
    .X(net5948));
 sg13g2_buf_8 fanout5949 (.A(net5952),
    .X(net5949));
 sg13g2_buf_8 fanout5950 (.A(net5951),
    .X(net5950));
 sg13g2_buf_2 fanout5951 (.A(net5952),
    .X(net5951));
 sg13g2_buf_2 fanout5952 (.A(net5965),
    .X(net5952));
 sg13g2_buf_8 fanout5953 (.A(net5959),
    .X(net5953));
 sg13g2_buf_8 fanout5954 (.A(net5959),
    .X(net5954));
 sg13g2_buf_8 fanout5955 (.A(net5958),
    .X(net5955));
 sg13g2_buf_8 fanout5956 (.A(net5958),
    .X(net5956));
 sg13g2_buf_2 fanout5957 (.A(net5958),
    .X(net5957));
 sg13g2_buf_8 fanout5958 (.A(net5959),
    .X(net5958));
 sg13g2_buf_8 fanout5959 (.A(net5965),
    .X(net5959));
 sg13g2_buf_8 fanout5960 (.A(net5961),
    .X(net5960));
 sg13g2_buf_8 fanout5961 (.A(net5964),
    .X(net5961));
 sg13g2_buf_8 fanout5962 (.A(net5963),
    .X(net5962));
 sg13g2_buf_8 fanout5963 (.A(net5964),
    .X(net5963));
 sg13g2_buf_8 fanout5964 (.A(net5965),
    .X(net5964));
 sg13g2_buf_8 fanout5965 (.A(rst_n),
    .X(net5965));
 sg13g2_buf_8 fanout5966 (.A(net5967),
    .X(net5966));
 sg13g2_buf_8 fanout5967 (.A(net5968),
    .X(net5967));
 sg13g2_buf_8 fanout5968 (.A(net5981),
    .X(net5968));
 sg13g2_buf_8 fanout5969 (.A(net5970),
    .X(net5969));
 sg13g2_buf_8 fanout5970 (.A(net5974),
    .X(net5970));
 sg13g2_buf_8 fanout5971 (.A(net5973),
    .X(net5971));
 sg13g2_buf_2 fanout5972 (.A(net5973),
    .X(net5972));
 sg13g2_buf_8 fanout5973 (.A(net5974),
    .X(net5973));
 sg13g2_buf_8 fanout5974 (.A(net5980),
    .X(net5974));
 sg13g2_buf_8 fanout5975 (.A(net5976),
    .X(net5975));
 sg13g2_buf_8 fanout5976 (.A(net5977),
    .X(net5976));
 sg13g2_buf_8 fanout5977 (.A(net5979),
    .X(net5977));
 sg13g2_buf_2 fanout5978 (.A(net5979),
    .X(net5978));
 sg13g2_buf_8 fanout5979 (.A(net5980),
    .X(net5979));
 sg13g2_buf_8 fanout5980 (.A(net5981),
    .X(net5980));
 sg13g2_buf_8 fanout5981 (.A(net6031),
    .X(net5981));
 sg13g2_buf_8 fanout5982 (.A(net5983),
    .X(net5982));
 sg13g2_buf_8 fanout5983 (.A(net5986),
    .X(net5983));
 sg13g2_buf_8 fanout5984 (.A(net5986),
    .X(net5984));
 sg13g2_buf_2 fanout5985 (.A(net5986),
    .X(net5985));
 sg13g2_buf_8 fanout5986 (.A(net6031),
    .X(net5986));
 sg13g2_buf_8 fanout5987 (.A(net5988),
    .X(net5987));
 sg13g2_buf_8 fanout5988 (.A(net5989),
    .X(net5988));
 sg13g2_buf_8 fanout5989 (.A(net5990),
    .X(net5989));
 sg13g2_buf_8 fanout5990 (.A(net5995),
    .X(net5990));
 sg13g2_buf_8 fanout5991 (.A(net5993),
    .X(net5991));
 sg13g2_buf_8 fanout5992 (.A(net5993),
    .X(net5992));
 sg13g2_buf_8 fanout5993 (.A(net5994),
    .X(net5993));
 sg13g2_buf_8 fanout5994 (.A(net5995),
    .X(net5994));
 sg13g2_buf_8 fanout5995 (.A(net6031),
    .X(net5995));
 sg13g2_buf_8 fanout5996 (.A(net5997),
    .X(net5996));
 sg13g2_buf_8 fanout5997 (.A(net6012),
    .X(net5997));
 sg13g2_buf_8 fanout5998 (.A(net6000),
    .X(net5998));
 sg13g2_buf_8 fanout5999 (.A(net6000),
    .X(net5999));
 sg13g2_buf_8 fanout6000 (.A(net6002),
    .X(net6000));
 sg13g2_buf_8 fanout6001 (.A(net6002),
    .X(net6001));
 sg13g2_buf_8 fanout6002 (.A(net6011),
    .X(net6002));
 sg13g2_buf_8 fanout6003 (.A(net6011),
    .X(net6003));
 sg13g2_buf_2 fanout6004 (.A(net6011),
    .X(net6004));
 sg13g2_buf_8 fanout6005 (.A(net6009),
    .X(net6005));
 sg13g2_buf_2 fanout6006 (.A(net6009),
    .X(net6006));
 sg13g2_buf_8 fanout6007 (.A(net6009),
    .X(net6007));
 sg13g2_buf_8 fanout6008 (.A(net6009),
    .X(net6008));
 sg13g2_buf_8 fanout6009 (.A(net6010),
    .X(net6009));
 sg13g2_buf_8 fanout6010 (.A(net6011),
    .X(net6010));
 sg13g2_buf_8 fanout6011 (.A(net6012),
    .X(net6011));
 sg13g2_buf_8 fanout6012 (.A(net6031),
    .X(net6012));
 sg13g2_buf_8 fanout6013 (.A(net6015),
    .X(net6013));
 sg13g2_buf_8 fanout6014 (.A(net6015),
    .X(net6014));
 sg13g2_buf_8 fanout6015 (.A(net6016),
    .X(net6015));
 sg13g2_buf_8 fanout6016 (.A(net6031),
    .X(net6016));
 sg13g2_buf_8 fanout6017 (.A(net6022),
    .X(net6017));
 sg13g2_buf_8 fanout6018 (.A(net6022),
    .X(net6018));
 sg13g2_buf_8 fanout6019 (.A(net6022),
    .X(net6019));
 sg13g2_buf_8 fanout6020 (.A(net6021),
    .X(net6020));
 sg13g2_buf_8 fanout6021 (.A(net6022),
    .X(net6021));
 sg13g2_buf_8 fanout6022 (.A(net6030),
    .X(net6022));
 sg13g2_buf_8 fanout6023 (.A(net6026),
    .X(net6023));
 sg13g2_buf_8 fanout6024 (.A(net6026),
    .X(net6024));
 sg13g2_buf_8 fanout6025 (.A(net6026),
    .X(net6025));
 sg13g2_buf_8 fanout6026 (.A(net6029),
    .X(net6026));
 sg13g2_buf_8 fanout6027 (.A(net6029),
    .X(net6027));
 sg13g2_buf_8 fanout6028 (.A(net6029),
    .X(net6028));
 sg13g2_buf_8 fanout6029 (.A(net6030),
    .X(net6029));
 sg13g2_buf_8 fanout6030 (.A(net6031),
    .X(net6030));
 sg13g2_buf_8 fanout6031 (.A(rst_n),
    .X(net6031));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_8 wire11 (.A(_19522_),
    .X(net11));
 sg13g2_tielo tt_um_corey_12 (.L_LO(net12));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sg13g2_buf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sg13g2_buf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sg13g2_buf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sg13g2_buf_8 clkbuf_5_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0_0_clk));
 sg13g2_buf_8 clkbuf_5_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1_0_clk));
 sg13g2_buf_8 clkbuf_5_2_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2_0_clk));
 sg13g2_buf_8 clkbuf_5_3_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3_0_clk));
 sg13g2_buf_8 clkbuf_5_4_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4_0_clk));
 sg13g2_buf_8 clkbuf_5_5_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5_0_clk));
 sg13g2_buf_8 clkbuf_5_6_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6_0_clk));
 sg13g2_buf_8 clkbuf_5_7_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7_0_clk));
 sg13g2_buf_8 clkbuf_5_8_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8_0_clk));
 sg13g2_buf_8 clkbuf_5_9_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9_0_clk));
 sg13g2_buf_8 clkbuf_5_10_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10_0_clk));
 sg13g2_buf_8 clkbuf_5_11_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11_0_clk));
 sg13g2_buf_8 clkbuf_5_12_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12_0_clk));
 sg13g2_buf_8 clkbuf_5_13_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13_0_clk));
 sg13g2_buf_8 clkbuf_5_14_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14_0_clk));
 sg13g2_buf_8 clkbuf_5_15_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15_0_clk));
 sg13g2_buf_8 clkbuf_5_16_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16_0_clk));
 sg13g2_buf_8 clkbuf_5_17_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17_0_clk));
 sg13g2_buf_8 clkbuf_5_18_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18_0_clk));
 sg13g2_buf_8 clkbuf_5_19_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19_0_clk));
 sg13g2_buf_8 clkbuf_5_20_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20_0_clk));
 sg13g2_buf_8 clkbuf_5_21_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21_0_clk));
 sg13g2_buf_8 clkbuf_5_22_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22_0_clk));
 sg13g2_buf_8 clkbuf_5_23_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23_0_clk));
 sg13g2_buf_8 clkbuf_5_24_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24_0_clk));
 sg13g2_buf_8 clkbuf_5_25_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25_0_clk));
 sg13g2_buf_8 clkbuf_5_26_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26_0_clk));
 sg13g2_buf_8 clkbuf_5_27_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27_0_clk));
 sg13g2_buf_8 clkbuf_5_28_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28_0_clk));
 sg13g2_buf_8 clkbuf_5_29_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29_0_clk));
 sg13g2_buf_8 clkbuf_5_30_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30_0_clk));
 sg13g2_buf_8 clkbuf_5_31_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31_0_clk));
 sg13g2_buf_8 clkbuf_6_0__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_8 clkbuf_6_1__f_clk (.A(clknet_5_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkbuf_6_2__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_8 clkbuf_6_3__f_clk (.A(clknet_5_1_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkbuf_6_4__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_8 clkbuf_6_5__f_clk (.A(clknet_5_2_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkbuf_6_6__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_8 clkbuf_6_7__f_clk (.A(clknet_5_3_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkbuf_6_8__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_8 clkbuf_6_9__f_clk (.A(clknet_5_4_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkbuf_6_10__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_8 clkbuf_6_11__f_clk (.A(clknet_5_5_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkbuf_6_12__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_8 clkbuf_6_13__f_clk (.A(clknet_5_6_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkbuf_6_14__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_8 clkbuf_6_15__f_clk (.A(clknet_5_7_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkbuf_6_16__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_8 clkbuf_6_17__f_clk (.A(clknet_5_8_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkbuf_6_18__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_8 clkbuf_6_19__f_clk (.A(clknet_5_9_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkbuf_6_20__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_8 clkbuf_6_21__f_clk (.A(clknet_5_10_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkbuf_6_22__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_8 clkbuf_6_23__f_clk (.A(clknet_5_11_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkbuf_6_24__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_8 clkbuf_6_25__f_clk (.A(clknet_5_12_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkbuf_6_26__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_8 clkbuf_6_27__f_clk (.A(clknet_5_13_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkbuf_6_28__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_8 clkbuf_6_29__f_clk (.A(clknet_5_14_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkbuf_6_30__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_8 clkbuf_6_31__f_clk (.A(clknet_5_15_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkbuf_6_32__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_8 clkbuf_6_33__f_clk (.A(clknet_5_16_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkbuf_6_34__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_8 clkbuf_6_35__f_clk (.A(clknet_5_17_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkbuf_6_36__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_8 clkbuf_6_37__f_clk (.A(clknet_5_18_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkbuf_6_38__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_8 clkbuf_6_39__f_clk (.A(clknet_5_19_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkbuf_6_40__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_8 clkbuf_6_41__f_clk (.A(clknet_5_20_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkbuf_6_42__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_8 clkbuf_6_43__f_clk (.A(clknet_5_21_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkbuf_6_44__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_8 clkbuf_6_45__f_clk (.A(clknet_5_22_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkbuf_6_46__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_8 clkbuf_6_47__f_clk (.A(clknet_5_23_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkbuf_6_48__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_8 clkbuf_6_49__f_clk (.A(clknet_5_24_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkbuf_6_50__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_8 clkbuf_6_51__f_clk (.A(clknet_5_25_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkbuf_6_52__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_8 clkbuf_6_53__f_clk (.A(clknet_5_26_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkbuf_6_54__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_8 clkbuf_6_55__f_clk (.A(clknet_5_27_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkbuf_6_56__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_8 clkbuf_6_57__f_clk (.A(clknet_5_28_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_8 clkbuf_6_58__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_8 clkbuf_6_59__f_clk (.A(clknet_5_29_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkbuf_6_60__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_8 clkbuf_6_61__f_clk (.A(clknet_5_30_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_8 clkbuf_6_62__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_8 clkbuf_6_63__f_clk (.A(clknet_5_31_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_6_61__leaf_clk));
 sg13g2_buf_8 clkload18 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_17_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_223_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_13_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_230_clk));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_79_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_236_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_232_clk));
 sg13g2_buf_8 clkload26 (.A(clknet_leaf_135_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_199_clk));
 sg13g2_buf_8 clkload28 (.A(clknet_leaf_198_clk));
 sg13g2_inv_2 clkload29 (.A(clknet_leaf_203_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_195_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_187_clk));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_212_clk));
 sg13g2_inv_1 clkload33 (.A(clknet_leaf_213_clk));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_208_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_209_clk));
 sg13g2_buf_8 clkload36 (.A(clknet_leaf_214_clk));
 sg13g2_inv_1 clkload37 (.A(clknet_leaf_129_clk));
 sg13g2_buf_8 rebuffer1 (.A(_09601_),
    .X(net1064));
 sg13g2_buf_8 rebuffer2 (.A(_03296_),
    .X(net1065));
 sg13g2_buf_1 rebuffer3 (.A(net1065),
    .X(net1066));
 sg13g2_buf_8 rebuffer4 (.A(_11595_),
    .X(net1067));
 sg13g2_buf_8 rebuffer5 (.A(_02560_),
    .X(net1068));
 sg13g2_buf_1 rebuffer6 (.A(net1068),
    .X(net1069));
 sg13g2_buf_8 rebuffer7 (.A(_06247_),
    .X(net1070));
 sg13g2_buf_8 rebuffer8 (.A(_09670_),
    .X(net1071));
 sg13g2_buf_1 rebuffer9 (.A(net1071),
    .X(net1072));
 sg13g2_buf_8 rebuffer10 (.A(_02486_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_inv.load_input ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold12 (.A(_00227_),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold13 (.A(\inv_result[18] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold14 (.A(\inv_result[34] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold15 (.A(\inv_result[30] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold16 (.A(\inv_result[32] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold17 (.A(\inv_result[12] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold18 (.A(\inv_result[67] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold19 (.A(\inv_result[246] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold20 (.A(\inv_result[65] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold21 (.A(\inv_result[58] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold22 (.A(\inv_result[10] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold23 (.A(\inv_result[60] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold24 (.A(\inv_result[16] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold25 (.A(\inv_result[160] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold26 (.A(\inv_result[250] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold27 (.A(\inv_result[56] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold28 (.A(\inv_result[57] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold29 (.A(\inv_result[70] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold30 (.A(\inv_result[61] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold31 (.A(\inv_result[193] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold32 (.A(\inv_result[91] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold33 (.A(\inv_result[59] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold34 (.A(\inv_result[80] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold35 (.A(\inv_result[238] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold36 (.A(\inv_result[229] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold37 (.A(\inv_result[224] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold38 (.A(\inv_result[165] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold39 (.A(\inv_result[153] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold40 (.A(\inv_result[211] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold41 (.A(\inv_result[213] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold42 (.A(\inv_result[66] ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold43 (.A(\inv_result[227] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold44 (.A(\inv_result[152] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold45 (.A(\inv_result[177] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold46 (.A(\inv_result[163] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold47 (.A(\inv_result[92] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold48 (.A(\inv_result[7] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold49 (.A(\inv_result[99] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold50 (.A(\shift_reg[264] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold51 (.A(_00499_),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold52 (.A(\shift_reg[270] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold53 (.A(_00505_),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold54 (.A(\shift_reg[271] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold55 (.A(_00506_),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold56 (.A(\inv_result[251] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold57 (.A(\inv_result[245] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold58 (.A(\inv_result[88] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold59 (.A(\inv_result[226] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold60 (.A(\inv_result[215] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold61 (.A(\inv_cycles[3] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold62 (.A(_01550_),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold63 (.A(\inv_result[72] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold64 (.A(\inv_result[217] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold65 (.A(\inv_result[68] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold66 (.A(\inv_result[204] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold67 (.A(\shift_reg[266] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold68 (.A(_00501_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold69 (.A(\inv_cycles[8] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold70 (.A(_01555_),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold71 (.A(\inv_result[225] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold72 (.A(\inv_result[168] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold73 (.A(\inv_result[207] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold74 (.A(\inv_result[184] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold75 (.A(\inv_result[111] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold76 (.A(\inv_result[100] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold77 (.A(_00618_),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold78 (.A(\shift_reg[256] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold79 (.A(_00491_),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold80 (.A(\inv_result[76] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold81 (.A(\inv_result[35] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_inv.d_next[205] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold83 (.A(_01236_),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold84 (.A(\inv_result[51] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold85 (.A(\u_inv.input_reg[11] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold86 (.A(_01579_),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold87 (.A(\shift_reg[263] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold88 (.A(_00498_),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold89 (.A(\inv_result[84] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold90 (.A(\byte_cnt[4] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold91 (.A(_00234_),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold92 (.A(\inv_result[21] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold93 (.A(\inv_result[162] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold94 (.A(\inv_result[181] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_inv.input_reg[12] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold96 (.A(_01580_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold97 (.A(\inv_result[98] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold98 (.A(\u_inv.input_reg[13] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold99 (.A(_01581_),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold100 (.A(\shift_reg[267] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold101 (.A(_00502_),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold102 (.A(\inv_result[147] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold103 (.A(\inv_result[49] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold104 (.A(\inv_result[54] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold105 (.A(\inv_result[71] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold106 (.A(\inv_result[113] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold107 (.A(\inv_result[252] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold108 (.A(\inv_result[36] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold109 (.A(\inv_cycles[0] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold110 (.A(_01547_),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold111 (.A(\inv_result[244] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold112 (.A(\inv_result[26] ),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold113 (.A(\inv_result[38] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold114 (.A(\inv_result[15] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold115 (.A(\inv_result[45] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold116 (.A(\inv_result[55] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold117 (.A(\inv_result[202] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold118 (.A(\byte_cnt[1] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold119 (.A(_19510_),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold120 (.A(_00231_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold121 (.A(\inv_result[94] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold122 (.A(\inv_result[89] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold123 (.A(\inv_result[46] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold124 (.A(\inv_result[120] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold125 (.A(\inv_result[39] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold126 (.A(\inv_result[140] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold127 (.A(\inv_result[144] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold128 (.A(\inv_result[112] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold129 (.A(\shift_reg[259] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold130 (.A(_00494_),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold131 (.A(\shift_reg[260] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold132 (.A(_00495_),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold133 (.A(\u_inv.f_reg[0] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold134 (.A(\inv_result[40] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold135 (.A(\inv_result[124] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold136 (.A(_00642_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold137 (.A(\inv_result[208] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold138 (.A(\inv_result[110] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold139 (.A(\inv_result[146] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold140 (.A(\inv_result[79] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold141 (.A(\shift_reg[261] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold142 (.A(_00496_),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold143 (.A(\inv_result[6] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold144 (.A(\inv_result[78] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold145 (.A(\inv_result[234] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold146 (.A(\inv_result[221] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold147 (.A(\shift_reg[268] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold148 (.A(\inv_result[249] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold149 (.A(\inv_result[248] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold150 (.A(\inv_result[103] ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold151 (.A(\u_inv.input_reg[10] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold152 (.A(_01578_),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold153 (.A(\inv_result[47] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold154 (.A(\shift_reg[269] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold155 (.A(_00504_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold156 (.A(\inv_result[62] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold157 (.A(\inv_result[150] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold158 (.A(\inv_result[154] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_inv.d_next[145] ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold160 (.A(_01176_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold161 (.A(\u_inv.delta_reg[9] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold162 (.A(_01566_),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold163 (.A(\inv_result[196] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold164 (.A(\inv_result[240] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold165 (.A(\inv_result[23] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold166 (.A(\inv_result[164] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold167 (.A(\shift_reg[258] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold168 (.A(_00493_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold169 (.A(\inv_result[161] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold170 (.A(\inv_result[167] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold171 (.A(\inv_result[206] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold172 (.A(\inv_result[197] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold173 (.A(\inv_result[145] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold174 (.A(\inv_cycles[7] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold175 (.A(_01554_),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold176 (.A(\inv_result[186] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold177 (.A(\shift_reg[265] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold178 (.A(_00500_),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold179 (.A(\shift_reg[257] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold180 (.A(_00492_),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_inv.f_next[8] ),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold182 (.A(_01296_),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold183 (.A(\inv_result[41] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold184 (.A(\u_inv.delta_reg[7] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold185 (.A(\inv_result[216] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold186 (.A(\inv_result[0] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold187 (.A(_00518_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold188 (.A(\inv_result[233] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold189 (.A(\inv_result[115] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold190 (.A(\inv_result[75] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold191 (.A(\inv_result[158] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold192 (.A(\inv_result[166] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold193 (.A(\inv_result[156] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold194 (.A(\inv_result[8] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold195 (.A(\inv_result[133] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold196 (.A(\inv_result[25] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_inv.d_next[66] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold198 (.A(_01097_),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold199 (.A(\inv_result[24] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold200 (.A(\inv_result[64] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold201 (.A(\inv_result[9] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold202 (.A(\inv_result[33] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold203 (.A(\inv_result[86] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold204 (.A(\inv_result[242] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold205 (.A(\inv_result[102] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold206 (.A(\inv_result[173] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold207 (.A(\inv_cycles[5] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold208 (.A(_01552_),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold209 (.A(\inv_result[96] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold210 (.A(\inv_cycles[1] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold211 (.A(_01548_),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold212 (.A(\inv_result[212] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold213 (.A(\inv_result[171] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold214 (.A(\inv_result[114] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold215 (.A(\inv_result[170] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold216 (.A(\inv_result[48] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold217 (.A(\inv_result[93] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold218 (.A(\inv_result[239] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold219 (.A(\inv_result[82] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold220 (.A(\inv_result[220] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold221 (.A(\inv_result[218] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold222 (.A(\inv_result[214] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold223 (.A(\inv_result[195] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold224 (.A(\shift_reg[3] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold225 (.A(_00246_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold226 (.A(\inv_result[178] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold227 (.A(\inv_result[44] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold228 (.A(\u_inv.input_reg[15] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold229 (.A(_01583_),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold230 (.A(\inv_result[228] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold231 (.A(\inv_result[105] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_inv.input_reg[14] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold233 (.A(_01582_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold234 (.A(\u_inv.f_reg[108] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold235 (.A(_01396_),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold236 (.A(\inv_result[50] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold237 (.A(\inv_result[101] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold238 (.A(_00619_),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold239 (.A(\inv_result[210] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold240 (.A(\inv_result[63] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold241 (.A(\inv_result[104] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold242 (.A(\inv_result[143] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold243 (.A(\inv_result[43] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold244 (.A(\shift_reg[163] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold245 (.A(_00398_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold246 (.A(\inv_result[69] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold247 (.A(\shift_reg[49] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold248 (.A(_00284_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold249 (.A(\shift_reg[2] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold250 (.A(_00245_),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold251 (.A(\inv_result[199] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold252 (.A(\inv_result[97] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold253 (.A(\inv_result[106] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold254 (.A(\inv_result[125] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold255 (.A(\inv_result[232] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold256 (.A(\inv_result[149] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold257 (.A(\inv_result[180] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold258 (.A(\inv_result[230] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold259 (.A(\inv_result[159] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold260 (.A(\shift_reg[262] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold261 (.A(_00497_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold262 (.A(\inv_result[5] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold263 (.A(\shift_reg[4] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold264 (.A(_00247_),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold265 (.A(\inv_result[188] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold266 (.A(\shift_reg[67] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00302_),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold268 (.A(\u_inv.d_next[225] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold269 (.A(_01256_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold270 (.A(\inv_result[118] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold271 (.A(\inv_result[231] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold272 (.A(\inv_result[151] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold273 (.A(\inv_result[169] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold274 (.A(\inv_result[190] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold275 (.A(\inv_result[142] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold276 (.A(\inv_result[29] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold277 (.A(\inv_result[176] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold278 (.A(\inv_result[247] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold279 (.A(\inv_result[172] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold280 (.A(\u_inv.d_next[191] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold281 (.A(_01222_),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold282 (.A(\shift_reg[243] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold283 (.A(_00478_),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold284 (.A(\inv_result[189] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold285 (.A(\inv_result[183] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold286 (.A(\inv_result[179] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold287 (.A(\inv_result[117] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold288 (.A(\inv_result[222] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold289 (.A(\inv_result[37] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold290 (.A(\inv_result[13] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold291 (.A(\shift_reg[38] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold292 (.A(_00273_),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold293 (.A(\inv_result[31] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold294 (.A(\inv_result[223] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold295 (.A(\inv_result[42] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold296 (.A(\u_inv.d_next[74] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold297 (.A(_01105_),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold298 (.A(\shift_reg[144] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold299 (.A(_00379_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold300 (.A(\inv_result[192] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold301 (.A(\inv_cycles[6] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold302 (.A(_01553_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold303 (.A(\inv_result[254] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold304 (.A(\inv_result[90] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold305 (.A(\u_inv.f_reg[137] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold306 (.A(_01425_),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold307 (.A(\shift_reg[178] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold308 (.A(_00413_),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold309 (.A(\inv_result[14] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold310 (.A(\inv_result[108] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold311 (.A(\shift_reg[102] ),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold312 (.A(_00337_),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold313 (.A(\shift_reg[84] ),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold314 (.A(_00319_),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold315 (.A(\shift_reg[34] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold316 (.A(_00269_),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold317 (.A(\inv_result[11] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold318 (.A(\inv_result[243] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold319 (.A(\inv_result[129] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold320 (.A(_00647_),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold321 (.A(\u_inv.d_next[0] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold322 (.A(_01031_),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold323 (.A(\inv_result[22] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold324 (.A(\inv_result[85] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold325 (.A(\inv_result[28] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold326 (.A(\shift_reg[127] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold327 (.A(_00362_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold328 (.A(\shift_reg[166] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold329 (.A(_00401_),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold330 (.A(\shift_reg[184] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold331 (.A(_00419_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold332 (.A(\shift_reg[87] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold333 (.A(_00322_),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold334 (.A(\shift_reg[0] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold335 (.A(\shift_reg[134] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold336 (.A(_00369_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold337 (.A(\shift_reg[159] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold338 (.A(_00394_),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold339 (.A(\shift_reg[254] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold340 (.A(_00489_),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold341 (.A(\shift_reg[244] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold342 (.A(_00479_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold343 (.A(\u_inv.d_next[70] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold344 (.A(_01101_),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold345 (.A(\shift_reg[162] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold346 (.A(_00397_),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold347 (.A(\inv_result[116] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold348 (.A(\inv_cycles[4] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold349 (.A(_01551_),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold350 (.A(\shift_reg[125] ),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold351 (.A(_00360_),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold352 (.A(\inv_result[87] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold353 (.A(\shift_reg[51] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold354 (.A(_00286_),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold355 (.A(\inv_result[119] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold356 (.A(\u_inv.d_next[253] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold357 (.A(_01284_),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold358 (.A(\u_inv.d_next[109] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold359 (.A(_01140_),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold360 (.A(\u_inv.d_next[175] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold361 (.A(_01206_),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold362 (.A(\shift_reg[215] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold363 (.A(_00450_),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold364 (.A(\shift_reg[239] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold365 (.A(_00474_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold366 (.A(\shift_reg[229] ),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold367 (.A(_00464_),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold368 (.A(\shift_reg[226] ),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold369 (.A(_00461_),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold370 (.A(\inv_result[95] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold371 (.A(\shift_reg[222] ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold372 (.A(_00457_),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold373 (.A(\u_inv.input_reg[60] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold374 (.A(_01628_),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold375 (.A(\u_inv.input_reg[8] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold376 (.A(_01576_),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold377 (.A(\u_inv.input_reg[174] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold378 (.A(_01742_),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold379 (.A(\inv_cycles[9] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold380 (.A(_01556_),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold381 (.A(\inv_result[174] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold382 (.A(\shift_reg[157] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold383 (.A(_00392_),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold384 (.A(\u_inv.input_reg[107] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold385 (.A(_01675_),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold386 (.A(\shift_reg[37] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold387 (.A(_00272_),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold388 (.A(\shift_reg[221] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold389 (.A(_00456_),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold390 (.A(\shift_reg[198] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold391 (.A(_00433_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold392 (.A(\u_inv.input_reg[52] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold393 (.A(_01620_),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold394 (.A(\u_inv.input_reg[63] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold395 (.A(_01631_),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold396 (.A(\u_inv.input_reg[155] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold397 (.A(_01723_),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold398 (.A(\u_inv.input_reg[79] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold399 (.A(_01647_),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold400 (.A(\shift_reg[65] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold401 (.A(_00300_),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold402 (.A(\shift_reg[23] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold403 (.A(_00258_),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold404 (.A(\u_inv.input_reg[224] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold405 (.A(_01792_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold406 (.A(\u_inv.input_reg[228] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold407 (.A(_01796_),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold408 (.A(\shift_reg[124] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold409 (.A(_00359_),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold410 (.A(\u_inv.input_reg[240] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold411 (.A(_01808_),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold412 (.A(\u_inv.input_reg[134] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold413 (.A(\inv_result[255] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold414 (.A(\shift_reg[123] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold415 (.A(_00358_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold416 (.A(\shift_reg[64] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold417 (.A(_00299_),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold418 (.A(\u_inv.input_reg[192] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold419 (.A(_01760_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold420 (.A(\u_inv.input_reg[55] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold421 (.A(_01623_),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold422 (.A(\u_inv.input_reg[103] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold423 (.A(_01671_),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold424 (.A(\shift_reg[237] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold425 (.A(\u_inv.input_reg[62] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold426 (.A(_01630_),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold427 (.A(\u_inv.input_reg[251] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold428 (.A(_01819_),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold429 (.A(\shift_reg[86] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold430 (.A(_00321_),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold431 (.A(\u_inv.input_reg[95] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold432 (.A(_01663_),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold433 (.A(\inv_result[175] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold434 (.A(\inv_result[122] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold435 (.A(\u_inv.input_reg[241] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold436 (.A(_01809_),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold437 (.A(\shift_reg[26] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold438 (.A(_00261_),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold439 (.A(\shift_reg[242] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold440 (.A(_00477_),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold441 (.A(\u_inv.f_next[220] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold442 (.A(_01508_),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold443 (.A(\u_inv.input_reg[139] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold444 (.A(_01707_),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold445 (.A(\u_inv.input_reg[54] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold446 (.A(_01622_),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold447 (.A(\shift_reg[70] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold448 (.A(_00305_),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold449 (.A(\u_inv.input_reg[99] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold450 (.A(_01667_),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold451 (.A(\u_inv.input_reg[71] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold452 (.A(_01639_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold453 (.A(\shift_reg[50] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold454 (.A(_00285_),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold455 (.A(\shift_reg[211] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold456 (.A(_00446_),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold457 (.A(\u_inv.input_reg[218] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold458 (.A(_01786_),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold459 (.A(\u_inv.input_reg[83] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold460 (.A(_01651_),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold461 (.A(\u_inv.d_next[87] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold462 (.A(_01118_),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold463 (.A(\inv_result[73] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold464 (.A(\u_inv.input_reg[115] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold465 (.A(_01683_),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold466 (.A(\u_inv.input_reg[36] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold467 (.A(_01604_),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold468 (.A(\u_inv.input_reg[114] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold469 (.A(_01682_),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold470 (.A(\shift_reg[59] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold471 (.A(\u_inv.d_next[110] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold472 (.A(_01141_),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold473 (.A(\u_inv.input_reg[181] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold474 (.A(_01749_),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold475 (.A(\u_inv.input_reg[61] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold476 (.A(_01629_),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold477 (.A(\u_inv.input_reg[219] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold478 (.A(_01787_),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold479 (.A(\u_inv.input_reg[65] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold480 (.A(\shift_reg[210] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold481 (.A(_00445_),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold482 (.A(\inv_result[209] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold483 (.A(\u_inv.input_reg[0] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold484 (.A(\u_inv.input_reg[69] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold485 (.A(_01637_),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold486 (.A(\u_inv.input_reg[111] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold487 (.A(_01679_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold488 (.A(\u_inv.input_reg[231] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold489 (.A(_01799_),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold490 (.A(\u_inv.input_reg[243] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold491 (.A(\u_inv.f_next[21] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold492 (.A(_01309_),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold493 (.A(\u_inv.input_reg[137] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold494 (.A(_01705_),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold495 (.A(\shift_reg[33] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold496 (.A(_00268_),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold497 (.A(\u_inv.input_reg[217] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold498 (.A(_01785_),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold499 (.A(\u_inv.input_reg[77] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold500 (.A(_01645_),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold501 (.A(\u_inv.input_reg[193] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold502 (.A(_01761_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold503 (.A(\shift_reg[146] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold504 (.A(_00381_),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold505 (.A(\u_inv.input_reg[242] ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold506 (.A(\u_inv.input_reg[76] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold507 (.A(_01644_),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold508 (.A(\u_inv.input_reg[177] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold509 (.A(_01745_),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold510 (.A(\u_inv.input_reg[48] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold511 (.A(_01616_),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold512 (.A(\u_inv.input_reg[87] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold513 (.A(\u_inv.input_reg[92] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold514 (.A(_01660_),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold515 (.A(\u_inv.input_reg[81] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold516 (.A(_01649_),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold517 (.A(\u_inv.input_reg[244] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold518 (.A(\u_inv.d_next[171] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold519 (.A(\u_inv.d_next[62] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold520 (.A(_01093_),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold521 (.A(\shift_reg[116] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold522 (.A(_00351_),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold523 (.A(\u_inv.input_reg[229] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold524 (.A(\u_inv.input_reg[132] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold525 (.A(_01700_),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold526 (.A(\u_inv.input_reg[80] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold527 (.A(_01648_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold528 (.A(\u_inv.input_reg[75] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold529 (.A(_01643_),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold530 (.A(\u_inv.input_reg[234] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold531 (.A(_01802_),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold532 (.A(\u_inv.input_reg[160] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold533 (.A(_01728_),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold534 (.A(\u_inv.d_next[28] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold535 (.A(_01059_),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold536 (.A(\u_inv.input_reg[91] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold537 (.A(_01659_),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold538 (.A(\shift_reg[183] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold539 (.A(_00418_),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold540 (.A(\u_inv.input_reg[208] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold541 (.A(_01776_),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold542 (.A(\u_inv.input_reg[255] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold543 (.A(_01823_),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold544 (.A(\u_inv.input_reg[164] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold545 (.A(_01732_),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold546 (.A(\inv_result[253] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold547 (.A(_00771_),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold548 (.A(\shift_reg[247] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold549 (.A(\u_inv.d_next[25] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold550 (.A(_01056_),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold551 (.A(\shift_reg[180] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold552 (.A(_00415_),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold553 (.A(\inv_result[205] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold555 (.A(\u_inv.input_reg[216] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold556 (.A(_01784_),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold557 (.A(\u_inv.input_reg[161] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold558 (.A(_01729_),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold559 (.A(\u_inv.input_reg[130] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold560 (.A(_01698_),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold561 (.A(\inv_result[123] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold562 (.A(_00641_),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold563 (.A(\u_inv.input_reg[72] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold564 (.A(_01640_),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold565 (.A(\inv_result[134] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold566 (.A(\shift_reg[5] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold567 (.A(_00248_),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold568 (.A(\inv_result[194] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold569 (.A(\u_inv.input_reg[116] ),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold570 (.A(\u_inv.input_reg[106] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold571 (.A(_01674_),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold572 (.A(\u_inv.input_reg[252] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold573 (.A(_01820_),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold574 (.A(\u_inv.input_reg[236] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold575 (.A(_01804_),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold576 (.A(\u_inv.input_reg[222] ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold577 (.A(\u_inv.d_next[103] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold578 (.A(_01134_),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold579 (.A(\u_inv.input_reg[248] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold580 (.A(_01816_),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold581 (.A(\shift_reg[7] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold582 (.A(\inv_result[135] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold583 (.A(\u_inv.input_reg[119] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold584 (.A(_01687_),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold585 (.A(\u_inv.input_reg[250] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold586 (.A(_01818_),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold587 (.A(\u_inv.input_reg[74] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold588 (.A(_01642_),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold589 (.A(\u_inv.input_reg[143] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold590 (.A(_01711_),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold591 (.A(\u_inv.input_reg[58] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold592 (.A(_01626_),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold593 (.A(\inv_cycles[2] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold594 (.A(_01549_),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold595 (.A(\shift_reg[194] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold596 (.A(_00429_),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold597 (.A(\shift_reg[58] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold598 (.A(\u_inv.d_next[179] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold599 (.A(\u_inv.input_reg[221] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold600 (.A(\u_inv.input_reg[53] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold601 (.A(_01621_),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold602 (.A(\u_inv.input_reg[135] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold603 (.A(_01703_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold604 (.A(\u_inv.input_reg[64] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold605 (.A(\shift_reg[217] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold606 (.A(_00452_),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold607 (.A(\shift_reg[145] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold608 (.A(_00380_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold609 (.A(\u_inv.input_reg[47] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold610 (.A(_01615_),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold611 (.A(\u_inv.d_next[212] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold612 (.A(\u_inv.input_reg[204] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold613 (.A(_01772_),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold614 (.A(\u_inv.input_reg[38] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold615 (.A(\u_inv.f_reg[222] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold616 (.A(_01510_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold617 (.A(\u_inv.input_reg[180] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold618 (.A(\u_inv.input_reg[121] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold619 (.A(_01689_),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold620 (.A(\u_inv.input_reg[191] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold621 (.A(_01759_),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold622 (.A(\u_inv.input_reg[226] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold623 (.A(\u_inv.input_reg[128] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold624 (.A(_01696_),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold625 (.A(\u_inv.input_reg[183] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold626 (.A(\u_inv.input_reg[159] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold627 (.A(\u_inv.input_reg[43] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold628 (.A(_01611_),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold629 (.A(\shift_reg[202] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold630 (.A(\u_inv.input_reg[133] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold631 (.A(_01701_),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold632 (.A(\u_inv.input_reg[175] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold633 (.A(_01743_),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold634 (.A(\u_inv.input_reg[6] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold635 (.A(_01574_),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold636 (.A(\u_inv.input_reg[57] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold637 (.A(_01625_),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold638 (.A(\shift_reg[135] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold639 (.A(\u_inv.input_reg[90] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold640 (.A(_01658_),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold641 (.A(\u_inv.input_reg[167] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold642 (.A(_01735_),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold643 (.A(\u_inv.input_reg[239] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold644 (.A(\u_inv.input_reg[94] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold645 (.A(_01662_),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold646 (.A(\shift_reg[99] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold647 (.A(_00334_),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold648 (.A(\u_inv.d_next[201] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold649 (.A(_01232_),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold650 (.A(\shift_reg[192] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold651 (.A(\u_inv.input_reg[184] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold652 (.A(\u_inv.input_reg[129] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold653 (.A(_01697_),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold654 (.A(\u_inv.input_reg[109] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold655 (.A(_01677_),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold656 (.A(\shift_reg[203] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold657 (.A(_00438_),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold658 (.A(\shift_reg[46] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold659 (.A(\shift_reg[42] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold660 (.A(\u_inv.input_reg[168] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold661 (.A(_01736_),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold662 (.A(\u_inv.d_next[192] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold663 (.A(\u_inv.d_next[54] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold664 (.A(_01085_),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold665 (.A(\u_inv.input_reg[97] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold666 (.A(_01665_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold667 (.A(\inv_result[136] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold668 (.A(\shift_reg[24] ),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold669 (.A(_00259_),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold670 (.A(\shift_reg[114] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold671 (.A(_00349_),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold672 (.A(\u_inv.input_reg[170] ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold673 (.A(_01738_),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold674 (.A(\shift_reg[60] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold675 (.A(_00295_),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold676 (.A(\u_inv.input_reg[44] ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold677 (.A(_01612_),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold678 (.A(\u_inv.input_reg[34] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold679 (.A(\u_inv.input_reg[42] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold680 (.A(\u_inv.f_next[32] ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold681 (.A(_01320_),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold682 (.A(\u_inv.input_reg[30] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold683 (.A(_01598_),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold684 (.A(\u_inv.input_reg[209] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold685 (.A(_01777_),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold686 (.A(\u_inv.input_reg[166] ),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold687 (.A(\u_inv.input_reg[51] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold688 (.A(\shift_reg[177] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold689 (.A(_00412_),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold690 (.A(\u_inv.input_reg[35] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold691 (.A(_01603_),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold692 (.A(\u_inv.input_reg[37] ),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold693 (.A(\u_inv.input_reg[96] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold694 (.A(_01664_),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold695 (.A(\u_inv.input_reg[194] ),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold696 (.A(\u_inv.input_reg[148] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold697 (.A(_01716_),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold698 (.A(\inv_result[148] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold699 (.A(\shift_reg[176] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold700 (.A(_00411_),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold701 (.A(\u_inv.input_reg[199] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold702 (.A(_01767_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold703 (.A(\shift_reg[155] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold704 (.A(_00390_),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold705 (.A(\inv_result[19] ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold706 (.A(\u_inv.input_reg[66] ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold707 (.A(_01634_),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold708 (.A(\u_inv.input_reg[202] ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold709 (.A(\inv_result[132] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold710 (.A(\u_inv.input_reg[25] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold711 (.A(_01593_),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold712 (.A(\shift_reg[95] ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold713 (.A(\u_inv.input_reg[147] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold714 (.A(_01715_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold715 (.A(\u_inv.input_reg[40] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold716 (.A(_01608_),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold717 (.A(\u_inv.input_reg[189] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold718 (.A(_01757_),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold719 (.A(\u_inv.input_reg[86] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold720 (.A(\u_inv.input_reg[211] ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold721 (.A(\shift_reg[118] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold722 (.A(_00353_),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold723 (.A(\shift_reg[209] ),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold724 (.A(_00444_),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold725 (.A(\shift_reg[223] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold726 (.A(\u_inv.input_reg[198] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold727 (.A(\shift_reg[130] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold728 (.A(_00365_),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold729 (.A(\u_inv.input_reg[32] ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold730 (.A(_01600_),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold731 (.A(\u_inv.input_reg[246] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold732 (.A(_01814_),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold733 (.A(\shift_reg[186] ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold734 (.A(\u_inv.input_reg[45] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold735 (.A(_01613_),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold736 (.A(\shift_reg[15] ),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold737 (.A(\shift_reg[120] ),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold738 (.A(_00355_),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold739 (.A(\u_inv.input_reg[67] ),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold740 (.A(\u_inv.input_reg[138] ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold741 (.A(_01706_),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold742 (.A(\u_inv.input_reg[108] ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold743 (.A(_01676_),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold744 (.A(\u_inv.input_reg[50] ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold745 (.A(\shift_reg[228] ),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold746 (.A(_00463_),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold747 (.A(\shift_reg[71] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold748 (.A(_00306_),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold749 (.A(\u_inv.d_reg[171] ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold750 (.A(\u_inv.input_reg[46] ),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold751 (.A(\u_inv.input_reg[233] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold752 (.A(_01801_),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold753 (.A(\u_inv.input_reg[156] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold754 (.A(_01724_),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold755 (.A(\u_inv.f_reg[166] ),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold756 (.A(_01454_),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold757 (.A(\u_inv.f_next[82] ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold758 (.A(_01370_),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold759 (.A(\u_inv.input_reg[88] ),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold760 (.A(_01656_),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold761 (.A(\u_inv.input_reg[220] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold762 (.A(_01788_),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold763 (.A(\u_inv.input_reg[185] ),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold764 (.A(_01753_),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold765 (.A(\shift_reg[240] ),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold766 (.A(_00475_),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold767 (.A(wr_prev),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold768 (.A(\inv_result[127] ),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold769 (.A(\inv_result[81] ),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold770 (.A(\u_inv.input_reg[245] ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold771 (.A(_01813_),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold772 (.A(\shift_reg[201] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold773 (.A(_00436_),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold774 (.A(\inv_result[3] ),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold775 (.A(\u_inv.input_reg[31] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold776 (.A(_01599_),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold777 (.A(\u_inv.input_reg[9] ),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold778 (.A(_01577_),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold779 (.A(\u_inv.input_reg[254] ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold780 (.A(_00225_),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold781 (.A(\u_inv.input_reg[215] ),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold782 (.A(\shift_reg[212] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold783 (.A(_00447_),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold784 (.A(\shift_reg[204] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold785 (.A(_00439_),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold786 (.A(\u_inv.f_next[148] ),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold787 (.A(_01436_),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold788 (.A(\u_inv.input_reg[150] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold789 (.A(_01718_),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold790 (.A(\shift_reg[69] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold791 (.A(_00304_),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold792 (.A(\u_inv.input_reg[120] ),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold793 (.A(\u_inv.input_reg[82] ),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold794 (.A(_01650_),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold795 (.A(\u_inv.input_reg[178] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold796 (.A(\u_inv.input_reg[153] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold797 (.A(_01721_),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold798 (.A(\u_inv.input_reg[145] ),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold799 (.A(\shift_reg[193] ),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold800 (.A(_00428_),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold801 (.A(\u_inv.delta_reg[8] ),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold802 (.A(\shift_reg[44] ),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold803 (.A(_00279_),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold804 (.A(\shift_reg[164] ),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold805 (.A(_00399_),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold806 (.A(\u_inv.f_reg[242] ),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold807 (.A(_01530_),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold808 (.A(\shift_reg[149] ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold809 (.A(_00384_),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold810 (.A(\u_inv.input_reg[206] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold811 (.A(_01774_),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold812 (.A(\u_inv.input_reg[187] ),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold813 (.A(_01755_),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold814 (.A(\u_inv.f_reg[62] ),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold815 (.A(_01350_),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold816 (.A(\u_inv.input_reg[101] ),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold817 (.A(_01669_),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold818 (.A(\shift_reg[189] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold819 (.A(_00424_),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold820 (.A(\u_inv.input_reg[144] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold821 (.A(\u_inv.input_reg[127] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold822 (.A(\u_inv.input_reg[210] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold823 (.A(\u_inv.input_reg[154] ),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold824 (.A(_01722_),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold825 (.A(\u_inv.input_reg[78] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold826 (.A(_01646_),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold827 (.A(\shift_reg[119] ),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold828 (.A(_00354_),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold829 (.A(\u_inv.input_reg[113] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold830 (.A(_01681_),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold831 (.A(\u_inv.input_reg[176] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold832 (.A(\u_inv.input_reg[182] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold833 (.A(_01750_),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold834 (.A(\u_inv.input_reg[163] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold835 (.A(\shift_reg[153] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold836 (.A(_00388_),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold837 (.A(\shift_reg[27] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold838 (.A(_00262_),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold839 (.A(\shift_reg[172] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold840 (.A(\shift_reg[80] ),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold841 (.A(_00315_),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold842 (.A(\u_inv.input_reg[227] ),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold843 (.A(_01795_),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold844 (.A(\u_inv.input_reg[85] ),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold845 (.A(_01653_),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold846 (.A(\u_inv.input_reg[223] ),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold847 (.A(\shift_reg[19] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold848 (.A(_00254_),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold849 (.A(\u_inv.input_reg[123] ),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold850 (.A(\u_inv.input_reg[112] ),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold851 (.A(_01680_),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold852 (.A(\shift_reg[61] ),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold853 (.A(_00296_),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold854 (.A(\u_inv.input_reg[110] ),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold855 (.A(_01678_),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold856 (.A(\u_inv.input_reg[232] ),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold857 (.A(_01800_),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold858 (.A(\shift_reg[205] ),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold859 (.A(_00440_),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold860 (.A(\shift_reg[77] ),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold861 (.A(\u_inv.input_reg[26] ),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold862 (.A(\u_inv.f_next[150] ),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold863 (.A(_01438_),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold864 (.A(\u_inv.input_reg[205] ),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold865 (.A(\u_inv.input_reg[39] ),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold866 (.A(_01607_),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold867 (.A(\u_inv.input_reg[104] ),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold868 (.A(_01672_),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold869 (.A(\u_inv.input_reg[151] ),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold870 (.A(_01719_),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold871 (.A(\u_inv.input_reg[24] ),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold872 (.A(\u_inv.input_reg[162] ),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold873 (.A(\shift_reg[109] ),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold874 (.A(_00344_),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold875 (.A(\shift_reg[136] ),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold876 (.A(_00371_),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold877 (.A(\u_inv.input_reg[158] ),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold878 (.A(_01726_),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold879 (.A(\shift_reg[213] ),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold880 (.A(\u_inv.input_reg[186] ),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold881 (.A(\u_inv.input_reg[190] ),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold882 (.A(_01758_),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold883 (.A(\shift_reg[147] ),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold884 (.A(_00382_),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold885 (.A(\shift_reg[233] ),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold886 (.A(_00468_),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold887 (.A(\shift_reg[104] ),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold888 (.A(_00339_),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold889 (.A(\shift_reg[63] ),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold890 (.A(_00298_),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold891 (.A(\u_inv.d_next[75] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold892 (.A(_01106_),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold893 (.A(\u_inv.d_next[244] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold894 (.A(_01275_),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold895 (.A(\u_inv.input_reg[70] ),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold896 (.A(\shift_reg[132] ),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold897 (.A(\u_inv.input_reg[196] ),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold898 (.A(_01764_),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold899 (.A(\shift_reg[20] ),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold900 (.A(_00255_),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold901 (.A(\shift_reg[126] ),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold902 (.A(pipe_pending),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold903 (.A(_01824_),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold904 (.A(\shift_reg[48] ),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold905 (.A(_00283_),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold906 (.A(\u_inv.d_next[138] ),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold907 (.A(\u_inv.input_reg[188] ),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold908 (.A(_01756_),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold909 (.A(\shift_reg[185] ),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold910 (.A(\shift_reg[225] ),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold911 (.A(\u_inv.input_reg[122] ),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold912 (.A(_01690_),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold913 (.A(\shift_reg[249] ),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold914 (.A(_00484_),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold915 (.A(\u_inv.input_reg[197] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold916 (.A(_01765_),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold917 (.A(\shift_reg[238] ),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold918 (.A(_00473_),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold919 (.A(\u_inv.d_next[177] ),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold920 (.A(_01208_),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold921 (.A(\u_inv.input_reg[102] ),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold922 (.A(\u_inv.input_reg[225] ),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold923 (.A(\u_inv.input_reg[214] ),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold924 (.A(_01782_),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold925 (.A(\shift_reg[108] ),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold926 (.A(_00343_),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold927 (.A(\u_inv.input_reg[28] ),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold928 (.A(_01596_),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold929 (.A(\u_inv.input_reg[200] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold930 (.A(_01768_),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold931 (.A(\shift_reg[98] ),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold932 (.A(_00333_),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold933 (.A(\inv_result[74] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold934 (.A(\shift_reg[218] ),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold935 (.A(\shift_reg[165] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold936 (.A(\u_inv.d_next[185] ),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold937 (.A(\shift_reg[236] ),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold938 (.A(\u_inv.input_reg[203] ),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold939 (.A(\u_inv.f_next[85] ),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold940 (.A(_01373_),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold941 (.A(\shift_reg[115] ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold942 (.A(_00350_),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold943 (.A(\u_inv.input_reg[195] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold944 (.A(_01763_),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold945 (.A(\shift_reg[179] ),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold946 (.A(_00414_),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold947 (.A(\shift_reg[113] ),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold948 (.A(_00348_),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold949 (.A(\shift_reg[171] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold950 (.A(_00406_),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold951 (.A(\u_inv.input_reg[146] ),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold952 (.A(\u_inv.input_reg[105] ),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold953 (.A(_01673_),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold954 (.A(\shift_reg[197] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold955 (.A(\u_inv.d_next[255] ),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold956 (.A(_01286_),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold957 (.A(\shift_reg[106] ),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold958 (.A(\u_inv.d_next[189] ),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold959 (.A(_01220_),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold960 (.A(\shift_reg[111] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold961 (.A(_00346_),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold962 (.A(\u_inv.input_reg[140] ),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold963 (.A(_01708_),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold964 (.A(\inv_result[27] ),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold965 (.A(\shift_reg[22] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold966 (.A(_00257_),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold967 (.A(\u_inv.f_reg[182] ),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold968 (.A(_01470_),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold969 (.A(\inv_result[128] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold970 (.A(\u_inv.f_reg[234] ),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold971 (.A(_01522_),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold972 (.A(\u_inv.input_reg[1] ),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold973 (.A(_01569_),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold974 (.A(\shift_reg[85] ),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold975 (.A(\u_inv.f_reg[122] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold976 (.A(_01410_),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold977 (.A(\inv_result[107] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold978 (.A(\shift_reg[231] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold979 (.A(\u_inv.d_reg[185] ),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold980 (.A(\inv_result[138] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold981 (.A(\shift_reg[137] ),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold982 (.A(_00372_),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold983 (.A(\u_inv.input_reg[149] ),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold984 (.A(\shift_reg[230] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold985 (.A(\u_inv.input_reg[41] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold986 (.A(_01609_),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold987 (.A(\u_inv.f_reg[118] ),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold988 (.A(_01406_),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold989 (.A(\inv_result[137] ),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold990 (.A(\shift_reg[158] ),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold991 (.A(_00393_),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold992 (.A(\u_inv.d_next[30] ),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold993 (.A(\shift_reg[224] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold994 (.A(_00459_),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold995 (.A(\shift_reg[174] ),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold996 (.A(\u_inv.input_reg[230] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold997 (.A(\u_inv.d_next[217] ),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold998 (.A(_01248_),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold999 (.A(\u_inv.d_next[155] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold1000 (.A(_01186_),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\u_inv.input_reg[125] ),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\u_inv.input_reg[201] ),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\shift_reg[1] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\u_inv.input_reg[131] ),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold1005 (.A(_01699_),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\u_inv.f_next[240] ),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold1007 (.A(_01528_),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\u_inv.input_reg[21] ),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold1009 (.A(_01589_),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\shift_reg[68] ),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold1011 (.A(_00303_),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\shift_reg[36] ),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold1013 (.A(_00271_),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\u_inv.input_reg[89] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold1015 (.A(_01657_),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\u_inv.input_reg[73] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold1017 (.A(_01641_),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\shift_reg[169] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold1019 (.A(_00404_),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\u_inv.delta_reg[1] ),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold1021 (.A(_01558_),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\u_inv.input_reg[124] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\u_inv.input_reg[173] ),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold1024 (.A(_01741_),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\u_inv.input_reg[171] ),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\u_inv.input_reg[237] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\u_inv.input_reg[141] ),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold1028 (.A(_01709_),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\u_inv.d_next[127] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold1030 (.A(_01158_),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\shift_reg[105] ),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_00340_),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\u_inv.f_next[253] ),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold1034 (.A(_01541_),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\u_inv.input_reg[179] ),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\u_inv.d_next[210] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\shift_reg[112] ),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\shift_reg[219] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold1039 (.A(_00454_),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\shift_reg[35] ),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\u_inv.d_next[45] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_01076_),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\shift_reg[227] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\shift_reg[195] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold1045 (.A(_00430_),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\u_inv.input_reg[169] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\u_inv.d_next[204] ),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_01235_),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\inv_result[198] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\shift_reg[122] ),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\u_inv.input_reg[23] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\shift_reg[89] ),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_00324_),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\u_inv.d_next[59] ),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_01090_),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\u_inv.input_reg[29] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold1057 (.A(_01597_),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\shift_reg[208] ),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold1059 (.A(_00443_),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\inv_result[130] ),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\shift_reg[196] ),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold1062 (.A(_00431_),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\shift_reg[21] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold1064 (.A(_00256_),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\shift_reg[141] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold1066 (.A(_00376_),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\u_inv.d_next[31] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold1068 (.A(_01062_),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\inv_result[157] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\u_inv.input_reg[207] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold1071 (.A(_01775_),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\u_inv.input_reg[136] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\shift_reg[78] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\u_inv.d_next[122] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\shift_reg[66] ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\u_inv.input_reg[5] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\u_inv.d_next[176] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\inv_result[126] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\shift_reg[148] ),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold1080 (.A(_00383_),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\shift_reg[43] ),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\u_inv.d_next[136] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold1083 (.A(_01167_),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\shift_reg[182] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\u_inv.d_next[202] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\shift_reg[246] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\u_inv.d_next[245] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold1088 (.A(_01276_),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\u_inv.input_reg[213] ),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\u_inv.d_reg[212] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\u_inv.input_reg[22] ),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\shift_reg[133] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\u_inv.input_reg[165] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\u_inv.input_reg[117] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold1095 (.A(_01685_),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\u_inv.f_next[65] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold1097 (.A(_01353_),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\shift_reg[25] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold1099 (.A(_00260_),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\u_inv.f_reg[6] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold1101 (.A(_01294_),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\shift_reg[121] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\u_inv.input_reg[157] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\shift_reg[167] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\shift_reg[75] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\shift_reg[28] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\shift_reg[214] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold1108 (.A(_00449_),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\inv_result[200] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\u_inv.d_reg[179] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\shift_reg[250] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\inv_result[17] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold1113 (.A(_00535_),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\u_inv.d_next[56] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold1115 (.A(_01087_),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\u_inv.input_reg[235] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold1117 (.A(_01803_),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\inv_result[20] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\u_inv.input_reg[84] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\u_inv.input_reg[212] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\shift_reg[140] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\u_inv.d_reg[98] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold1123 (.A(_01129_),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\u_inv.input_reg[49] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\shift_reg[161] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\u_inv.d_next[226] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\shift_reg[187] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\u_inv.input_reg[126] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\u_inv.input_reg[238] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\shift_reg[241] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\shift_reg[160] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold1132 (.A(_00395_),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\u_inv.f_reg[254] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_01542_),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\u_inv.delta_reg[3] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold1136 (.A(_01560_),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\shift_reg[129] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\u_inv.f_reg[248] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold1139 (.A(_01536_),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\shift_reg[220] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\u_inv.input_reg[3] ),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\u_inv.d_next[186] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold1143 (.A(_01217_),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\shift_reg[76] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\u_inv.input_reg[172] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\u_inv.input_reg[17] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold1147 (.A(_01585_),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\shift_reg[18] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold1149 (.A(_00253_),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\u_inv.d_next[43] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold1151 (.A(_01074_),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\u_inv.input_reg[247] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\u_inv.d_next[206] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold1154 (.A(_01237_),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\shift_reg[53] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold1156 (.A(_00288_),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\u_inv.f_reg[68] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold1158 (.A(_01356_),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\shift_reg[131] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\shift_reg[103] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\shift_reg[101] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold1162 (.A(_00336_),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\shift_reg[156] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\u_inv.d_reg[226] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\shift_reg[17] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold1166 (.A(_00252_),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\shift_reg[96] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold1168 (.A(_00331_),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\shift_reg[150] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold1170 (.A(_00385_),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\u_inv.f_reg[123] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold1172 (.A(_01411_),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\u_inv.d_next[241] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold1174 (.A(_01272_),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\u_inv.d_next[196] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold1176 (.A(_01227_),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\u_inv.input_reg[59] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\shift_reg[232] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\u_inv.f_reg[46] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold1180 (.A(_01334_),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\shift_reg[188] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\shift_reg[54] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\u_inv.d_next[172] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold1184 (.A(_01203_),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\u_inv.d_reg[210] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\u_inv.d_next[143] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_01174_),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\u_inv.f_next[255] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold1189 (.A(_01543_),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\u_inv.f_reg[2] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold1191 (.A(_01290_),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\u_inv.f_reg[203] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold1193 (.A(_01491_),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\u_inv.d_next[197] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_01228_),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\shift_reg[100] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold1197 (.A(_00335_),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\u_inv.d_next[39] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_01070_),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\u_inv.input_reg[142] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold1201 (.A(_01710_),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\u_inv.d_next[249] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold1203 (.A(_01280_),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\shift_reg[117] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\u_inv.d_next[38] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_01069_),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\u_inv.f_reg[188] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold1208 (.A(_01476_),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\shift_reg[168] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\u_inv.d_next[29] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold1211 (.A(_01060_),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\shift_reg[110] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\u_inv.d_next[86] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold1214 (.A(_01117_),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\u_inv.d_next[198] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\u_inv.d_next[194] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold1217 (.A(_01225_),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\u_inv.f_next[204] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_01492_),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\u_inv.input_reg[118] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\u_inv.d_next[170] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\u_inv.input_reg[2] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\u_inv.input_reg[33] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\inv_result[53] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\u_inv.input_reg[253] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold1226 (.A(_01821_),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\u_inv.d_reg[198] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\shift_reg[142] ),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\u_inv.d_next[190] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold1230 (.A(_01221_),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\u_inv.d_next[238] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\u_inv.f_next[89] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold1233 (.A(_01377_),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\u_inv.f_reg[212] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold1235 (.A(_01500_),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\u_inv.d_next[21] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold1237 (.A(_01052_),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\u_inv.f_reg[52] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold1239 (.A(_01340_),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\shift_reg[253] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold1241 (.A(_00488_),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\u_inv.d_next[195] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\u_inv.d_next[78] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold1244 (.A(_01109_),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\u_inv.d_next[22] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\shift_reg[190] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\shift_reg[82] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold1248 (.A(_00317_),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\shift_reg[47] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold1250 (.A(_00282_),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\u_inv.input_reg[93] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold1252 (.A(_01661_),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\u_inv.f_next[256] ),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\u_inv.d_next[130] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_01161_),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\shift_reg[6] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold1257 (.A(_00249_),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\u_inv.d_next[104] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_01135_),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\shift_reg[181] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold1261 (.A(_00416_),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\u_inv.d_next[46] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold1263 (.A(_01077_),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\u_inv.d_next[102] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold1265 (.A(_01133_),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\inv_result[83] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\u_inv.d_reg[192] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\u_inv.input_reg[56] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold1269 (.A(_01624_),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\shift_reg[107] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\u_inv.d_next[65] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold1272 (.A(_01096_),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\shift_reg[216] ),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\u_inv.d_next[100] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold1275 (.A(_01131_),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\shift_reg[170] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\shift_reg[173] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\u_inv.d_next[188] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold1279 (.A(_01219_),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\u_inv.d_next[42] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold1281 (.A(_01073_),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\u_inv.input_reg[19] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\u_inv.d_reg[176] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\u_inv.d_next[60] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold1285 (.A(_01091_),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\u_inv.d_next[256] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\shift_reg[31] ),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\u_inv.f_next[205] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold1289 (.A(_01493_),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\u_inv.f_reg[186] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold1291 (.A(_01474_),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\u_inv.f_next[4] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold1293 (.A(_01292_),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\shift_reg[175] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\shift_reg[199] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold1296 (.A(_00434_),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\u_inv.f_reg[1] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold1298 (.A(_01289_),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\shift_reg[128] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\u_inv.d_reg[122] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\u_inv.f_next[23] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\u_inv.f_reg[236] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold1303 (.A(_01524_),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\shift_reg[139] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\u_inv.f_next[252] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_01540_),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\u_inv.d_next[115] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold1308 (.A(_01146_),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\u_inv.d_next[114] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold1310 (.A(_01145_),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\shift_reg[91] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold1312 (.A(_00326_),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\u_inv.input_reg[152] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold1314 (.A(_01720_),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\u_inv.d_next[234] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold1316 (.A(_01265_),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\shift_reg[152] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\u_inv.d_next[152] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold1319 (.A(_01183_),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\u_inv.d_next[156] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\u_inv.input_reg[27] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\u_inv.d_next[182] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\shift_reg[143] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\u_inv.input_reg[100] ),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\u_inv.d_next[92] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold1326 (.A(_01123_),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\u_inv.d_reg[195] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\u_inv.f_next[94] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_01382_),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold1330 (.A(next_loaded),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold1331 (.A(_02336_),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\shift_reg[191] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\u_inv.d_next[200] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\inv_result[109] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\u_inv.d_next[1] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold1336 (.A(_01032_),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\shift_reg[93] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold1338 (.A(_00328_),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\u_inv.d_reg[202] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\shift_reg[234] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\shift_reg[40] ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold1342 (.A(_00275_),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\u_inv.d_next[154] ),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\u_inv.d_next[44] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold1345 (.A(_01075_),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\u_inv.f_reg[42] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold1347 (.A(_01330_),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\shift_reg[207] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold1349 (.A(_00442_),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\u_inv.f_next[208] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold1351 (.A(_01496_),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\u_inv.d_next[41] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_01072_),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\u_inv.d_reg[22] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\u_inv.d_next[178] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold1356 (.A(_01209_),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\u_inv.d_next[99] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold1358 (.A(_01130_),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\inv_result[182] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold1360 (.A(_00700_),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\u_inv.f_reg[145] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold1362 (.A(_01433_),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\u_inv.d_next[7] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold1364 (.A(_01038_),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\u_inv.d_reg[138] ),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\u_inv.d_reg[154] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\u_inv.d_next[2] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold1368 (.A(_01033_),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\shift_reg[138] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\u_inv.d_next[153] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\shift_reg[39] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\u_inv.input_reg[68] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\u_inv.input_reg[98] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\u_inv.d_next[112] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\u_inv.d_next[53] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold1376 (.A(_01084_),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\shift_reg[45] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\u_inv.d_next[14] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold1379 (.A(_01045_),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\u_inv.d_next[126] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold1381 (.A(_01157_),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\shift_reg[32] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\u_inv.d_next[250] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\u_inv.input_reg[20] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\u_inv.d_next[82] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold1386 (.A(_01113_),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\u_inv.f_next[241] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold1388 (.A(_01529_),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\shift_reg[206] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\shift_reg[9] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\shift_reg[90] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\u_inv.f_reg[133] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold1393 (.A(_01421_),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\u_inv.d_next[203] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold1395 (.A(_01234_),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\shift_reg[200] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\shift_reg[16] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold1398 (.A(_00251_),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\u_inv.d_next[193] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold1400 (.A(_01224_),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\u_inv.f_reg[26] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold1402 (.A(_01314_),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\u_inv.f_reg[70] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold1404 (.A(_01358_),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\u_inv.d_next[85] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold1406 (.A(_01116_),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\u_inv.d_next[132] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\u_inv.f_reg[130] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold1409 (.A(_01418_),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\u_inv.d_next[24] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold1411 (.A(_01055_),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\shift_reg[88] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\u_inv.d_next[242] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold1414 (.A(_01273_),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\u_inv.d_next[246] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\u_inv.d_next[47] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold1417 (.A(_01078_),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\u_inv.f_next[210] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold1419 (.A(_01498_),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\u_inv.f_reg[226] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold1421 (.A(_01514_),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\u_inv.d_next[235] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\u_inv.d_reg[182] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\inv_result[131] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\u_inv.input_reg[18] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\u_inv.f_reg[110] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold1427 (.A(_01398_),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\u_inv.f_next[100] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold1429 (.A(_01388_),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\u_inv.f_next[199] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold1431 (.A(_01487_),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\u_inv.d_reg[200] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\u_inv.d_next[211] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold1434 (.A(_01242_),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\u_inv.d_reg[170] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\u_inv.f_reg[131] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold1437 (.A(_01419_),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\u_inv.f_reg[15] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold1439 (.A(_01303_),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\u_inv.d_next[9] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold1441 (.A(_01040_),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\inv_result[4] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\u_inv.d_next[252] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold1444 (.A(_01283_),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\u_inv.d_next[13] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold1446 (.A(_01044_),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\u_inv.input_reg[4] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\u_inv.d_reg[250] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\u_inv.f_next[50] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold1450 (.A(_01338_),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\u_inv.d_next[105] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold1452 (.A(_01136_),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\u_inv.d_next[108] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold1454 (.A(_01139_),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\shift_reg[154] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\u_inv.d_next[141] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold1457 (.A(_01172_),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\inv_result[235] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\u_inv.input_reg[7] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\u_inv.d_next[12] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold1461 (.A(_01043_),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\u_inv.d_reg[30] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\u_inv.f_next[9] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold1464 (.A(_01297_),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\u_inv.d_next[222] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold1466 (.A(_01253_),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\u_inv.d_next[218] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold1468 (.A(_01249_),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\u_inv.f_next[211] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold1470 (.A(_01499_),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\shift_reg[30] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\u_inv.d_reg[153] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\u_inv.d_next[71] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold1474 (.A(_01102_),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\u_inv.d_next[173] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\shift_reg[97] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\u_inv.f_next[213] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold1478 (.A(_01501_),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\shift_reg[248] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\u_inv.d_next[6] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold1481 (.A(_01037_),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\shift_reg[8] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\u_inv.f_next[56] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_01344_),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\byte_cnt[0] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold1486 (.A(_00230_),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\inv_result[52] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\shift_reg[79] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\u_inv.d_next[142] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold1490 (.A(_01173_),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\u_inv.f_next[117] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold1492 (.A(_01405_),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\shift_reg[62] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\u_inv.d_reg[140] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold1495 (.A(_01171_),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\u_inv.f_next[51] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold1497 (.A(_01339_),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\u_inv.d_next[168] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold1499 (.A(_01199_),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\u_inv.d_next[3] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold1501 (.A(_01034_),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\u_inv.f_next[136] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold1503 (.A(_01424_),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\shift_reg[245] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\shift_reg[151] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\u_inv.d_next[113] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold1507 (.A(_01144_),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\u_inv.d_next[233] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold1509 (.A(_01264_),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\u_inv.d_next[231] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold1511 (.A(_01262_),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\u_inv.d_next[216] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold1513 (.A(_01247_),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\u_inv.f_next[223] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold1515 (.A(_01511_),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\u_inv.f_next[197] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold1517 (.A(_01485_),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\u_inv.d_next[35] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold1519 (.A(_01066_),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\u_inv.f_next[190] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold1521 (.A(_01478_),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\u_inv.f_reg[95] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold1523 (.A(_01383_),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\u_inv.d_next[169] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\u_inv.d_next[34] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold1526 (.A(_01065_),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\u_inv.d_next[55] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold1528 (.A(_01086_),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\inv_result[236] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\u_inv.f_reg[20] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold1531 (.A(_01308_),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\u_inv.d_reg[256] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\u_inv.d_next[20] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_01051_),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\u_inv.f_reg[156] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold1536 (.A(_01444_),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\u_inv.d_next[61] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold1538 (.A(_01092_),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\inv_result[2] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\u_inv.d_next[237] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\u_inv.d_next[8] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold1542 (.A(_01039_),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\u_inv.d_next[58] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_01089_),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\u_inv.f_next[7] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold1546 (.A(_01295_),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\u_inv.d_next[129] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold1548 (.A(_01160_),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\u_inv.d_next[101] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold1550 (.A(_01132_),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\u_inv.f_next[97] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_01385_),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\u_inv.d_reg[169] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\u_inv.f_next[229] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold1555 (.A(_01517_),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\u_inv.d_next[15] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold1557 (.A(_01046_),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\u_inv.d_next[123] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold1559 (.A(_01154_),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\shift_reg[83] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\u_inv.d_next[57] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold1562 (.A(_01088_),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\u_inv.d_next[94] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold1564 (.A(_01125_),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\u_inv.d_next[229] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold1566 (.A(_01260_),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\u_inv.f_next[221] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\shift_reg[29] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\u_inv.d_next[134] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\u_inv.counter[9] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold1571 (.A(_02379_),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold1572 (.A(_00517_),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\u_inv.d_next[83] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold1574 (.A(_01114_),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\u_inv.d_next[118] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_01149_),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\inv_result[187] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\u_inv.d_next[64] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold1579 (.A(_01095_),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\shift_reg[235] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_00470_),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\u_inv.d_next[51] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold1583 (.A(_01082_),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\u_inv.f_reg[91] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold1585 (.A(_01379_),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\u_inv.d_next[228] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold1587 (.A(_01259_),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\shift_reg[74] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\u_inv.f_reg[198] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold1590 (.A(_01486_),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\u_inv.f_next[161] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold1592 (.A(_01449_),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\u_inv.f_reg[238] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold1594 (.A(_01526_),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\u_inv.d_next[251] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold1596 (.A(_01282_),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\shift_reg[255] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\u_inv.f_reg[132] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_01420_),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\u_inv.d_next[181] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold1601 (.A(_01212_),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\u_inv.f_next[129] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold1603 (.A(_01417_),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\u_inv.d_next[91] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold1605 (.A(_01122_),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\u_inv.d_next[240] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\u_inv.f_reg[22] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold1608 (.A(_01310_),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\inv_result[185] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\u_inv.f_next[84] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_01372_),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\shift_reg[92] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\u_inv.f_next[187] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold1614 (.A(_01475_),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\u_inv.d_next[63] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold1616 (.A(_01094_),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\u_inv.d_reg[235] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\u_inv.f_next[152] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\u_inv.d_next[144] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold1620 (.A(_01175_),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\u_inv.f_reg[45] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold1622 (.A(_01333_),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\shift_reg[94] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\u_inv.f_reg[101] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold1625 (.A(_01389_),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\u_inv.d_next[32] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold1627 (.A(_01063_),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\u_inv.d_next[207] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold1629 (.A(_01238_),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\u_inv.d_next[131] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold1631 (.A(_01162_),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\u_inv.f_reg[78] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold1633 (.A(_01366_),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\u_inv.d_next[124] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\u_inv.f_next[43] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold1636 (.A(_01331_),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\u_inv.f_reg[143] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold1638 (.A(_01431_),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\u_inv.f_next[149] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\u_inv.d_reg[132] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\u_inv.d_next[18] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold1642 (.A(_01049_),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\u_inv.d_reg[112] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\u_inv.d_next[174] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold1645 (.A(_01205_),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\u_inv.f_next[63] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold1647 (.A(_01351_),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\u_inv.f_next[249] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold1649 (.A(_01537_),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\u_inv.f_next[212] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\u_inv.f_reg[179] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold1652 (.A(_01467_),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\inv_result[139] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\u_inv.f_reg[244] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold1655 (.A(_01532_),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\u_inv.f_reg[162] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold1657 (.A(_01450_),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\shift_reg[41] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\u_inv.d_next[161] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold1660 (.A(_01192_),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\u_inv.d_reg[238] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\u_inv.d_reg[164] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold1663 (.A(_01195_),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\u_inv.input_reg[16] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\inv_result[155] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\u_inv.f_next[225] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold1667 (.A(_01513_),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\shift_reg[55] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\u_inv.d_next[160] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\u_inv.f_reg[231] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold1671 (.A(_01519_),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\u_inv.f_next[183] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold1673 (.A(_01471_),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\u_inv.d_next[209] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold1675 (.A(_01240_),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\u_inv.d_next[140] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\u_inv.d_next[52] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold1678 (.A(_01083_),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\shift_reg[81] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold1680 (.A(_00316_),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\u_inv.f_next[163] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold1682 (.A(_01451_),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\u_inv.f_reg[126] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold1684 (.A(_01414_),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\u_inv.f_reg[170] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold1686 (.A(_01458_),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\inv_result[1] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\u_inv.d_reg[237] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\u_inv.f_reg[66] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold1690 (.A(_01354_),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\u_inv.f_next[251] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold1692 (.A(_01539_),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\u_inv.d_next[146] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold1694 (.A(_01177_),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\u_inv.f_next[69] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold1696 (.A(_01357_),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\u_inv.f_reg[27] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold1698 (.A(_01315_),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\inv_result[141] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\u_inv.f_reg[221] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\u_inv.f_reg[206] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold1702 (.A(_01494_),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\u_inv.f_reg[38] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold1704 (.A(_01326_),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\u_inv.f_reg[250] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold1706 (.A(_01538_),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\inv_result[77] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\u_inv.f_reg[80] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold1709 (.A(_01368_),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\u_inv.f_next[181] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold1711 (.A(_01469_),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\inv_result[219] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\u_inv.f_reg[230] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_01518_),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\u_inv.f_next[47] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold1716 (.A(_01335_),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\u_inv.input_reg[249] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\u_inv.d_next[4] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\u_inv.d_reg[160] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\u_inv.f_next[128] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold1721 (.A(_01416_),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\u_inv.f_reg[224] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold1723 (.A(_01512_),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\u_inv.d_next[17] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold1725 (.A(_01048_),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\u_inv.f_reg[104] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold1727 (.A(_01392_),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\u_inv.d_next[232] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold1729 (.A(_01263_),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\u_inv.f_reg[194] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold1731 (.A(_01482_),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\shift_reg[251] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\u_inv.f_next[185] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold1734 (.A(_01473_),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\u_inv.f_reg[147] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold1736 (.A(_01435_),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\u_inv.f_next[245] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold1738 (.A(_01533_),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\u_inv.d_next[183] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\u_inv.f_reg[202] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold1741 (.A(_01490_),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\u_inv.f_reg[144] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold1743 (.A(_01432_),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\u_inv.f_reg[174] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold1745 (.A(_01462_),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\u_inv.d_reg[183] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\u_inv.d_next[84] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold1748 (.A(_01115_),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\u_inv.f_reg[86] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold1750 (.A(_01374_),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\u_inv.d_next[139] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold1752 (.A(_01170_),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\inv_result[237] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\u_inv.f_reg[14] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold1755 (.A(_01302_),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\shift_reg[56] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\u_inv.f_reg[140] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold1758 (.A(_01428_),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\u_inv.d_reg[124] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\u_inv.f_next[66] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\u_inv.d_reg[246] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\u_inv.f_next[81] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold1763 (.A(_01369_),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\u_inv.f_reg[196] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold1765 (.A(_01484_),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\u_inv.f_reg[114] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold1767 (.A(_01402_),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\byte_cnt[3] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold1769 (.A(_19517_),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\u_inv.f_reg[3] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold1771 (.A(_01291_),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\u_inv.d_reg[156] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\u_inv.d_next[180] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold1774 (.A(_01211_),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\u_inv.f_reg[83] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold1776 (.A(_01371_),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\u_inv.d_next[26] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold1778 (.A(_01057_),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\u_inv.delta_reg[2] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold1780 (.A(_01559_),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\u_inv.counter[4] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold1782 (.A(_02351_),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\u_inv.f_next[125] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold1784 (.A(_01413_),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\u_inv.f_next[57] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\u_inv.d_next[80] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold1787 (.A(_01111_),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\u_inv.f_next[24] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold1789 (.A(_01312_),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\u_inv.d_next[90] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\u_inv.f_reg[165] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold1792 (.A(_01453_),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\u_inv.f_reg[5] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold1794 (.A(_01293_),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\u_inv.f_next[90] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\shift_reg[72] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\u_inv.f_reg[11] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold1798 (.A(_01299_),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\u_inv.d_next[5] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold1800 (.A(_01036_),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\u_inv.d_next[37] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold1802 (.A(_01068_),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\u_inv.delta_reg[4] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\u_inv.f_reg[23] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\shift_reg[252] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\u_inv.f_reg[164] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold1807 (.A(_01452_),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\u_inv.d_next[68] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold1809 (.A(_01099_),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\u_inv.f_next[246] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold1811 (.A(_01534_),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\u_inv.d_next[166] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold1813 (.A(_01197_),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\u_inv.f_reg[58] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold1815 (.A(_01346_),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\u_inv.d_next[67] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold1817 (.A(_01098_),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\u_inv.d_next[48] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold1819 (.A(_01079_),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\u_inv.d_next[119] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold1821 (.A(_01150_),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\u_inv.d_next[40] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold1823 (.A(_01071_),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\u_inv.d_next[223] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\u_inv.delta_reg[5] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold1826 (.A(_13816_),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\u_inv.f_reg[40] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold1828 (.A(_01328_),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\u_inv.f_reg[34] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold1830 (.A(_01322_),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\u_inv.f_reg[76] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold1832 (.A(_01364_),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\shift_reg[52] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\shift_reg[73] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\u_inv.d_reg[240] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\u_inv.f_reg[44] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold1837 (.A(_01332_),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\u_inv.d_next[230] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\u_inv.d_next[248] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold1840 (.A(_01279_),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\u_inv.d_next[19] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold1842 (.A(_01050_),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\u_inv.d_next[116] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold1844 (.A(_01147_),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\u_inv.d_next[163] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\u_inv.d_next[184] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold1847 (.A(_01215_),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\u_inv.f_next[88] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold1849 (.A(_01376_),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\u_inv.f_reg[61] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold1851 (.A(_01349_),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\u_inv.f_reg[106] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold1853 (.A(_01394_),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\u_inv.d_next[243] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold1855 (.A(_01274_),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\u_inv.d_next[111] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold1857 (.A(_01142_),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\u_inv.d_next[208] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold1859 (.A(_01239_),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\u_inv.d_reg[230] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\u_inv.f_reg[10] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold1862 (.A(_01298_),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\u_inv.d_next[49] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold1864 (.A(_01080_),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\u_inv.d_next[81] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold1866 (.A(_01112_),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\u_inv.f_reg[120] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold1868 (.A(_01408_),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\u_inv.d_next[149] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold1870 (.A(_01180_),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\u_inv.d_next[16] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold1872 (.A(_01047_),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\u_inv.d_next[167] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold1874 (.A(_01198_),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\u_inv.d_next[199] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\u_inv.f_reg[36] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold1877 (.A(_01324_),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\shift_reg[57] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\u_inv.d_next[148] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold1880 (.A(_01179_),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\u_inv.d_next[95] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold1882 (.A(_01126_),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\u_inv.f_next[146] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold1884 (.A(_01434_),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\inv_result[203] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\u_inv.d_next[224] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold1887 (.A(_01255_),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\u_inv.f_next[86] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\u_inv.d_next[69] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold1890 (.A(_01100_),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\u_inv.f_next[201] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\u_inv.d_reg[4] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\u_inv.f_reg[215] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold1894 (.A(_01503_),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\u_inv.f_reg[134] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold1896 (.A(_01422_),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\u_inv.f_next[44] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\u_inv.f_next[214] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\u_inv.d_next[254] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\u_inv.d_next[73] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold1901 (.A(_01104_),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\u_inv.d_reg[134] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\u_inv.d_reg[254] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\u_inv.f_reg[64] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold1905 (.A(_01352_),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\u_inv.d_reg[199] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\u_inv.d_next[27] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold1908 (.A(_01058_),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\u_inv.f_next[52] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\u_inv.d_next[147] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\u_inv.d_next[76] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold1912 (.A(_01107_),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\u_inv.d_next[128] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold1914 (.A(_01159_),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\u_inv.f_next[96] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\inv_result[201] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\u_inv.f_next[19] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold1918 (.A(_01307_),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\u_inv.f_reg[158] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold1920 (.A(_01446_),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\u_inv.d_next[33] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold1922 (.A(_01064_),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\u_inv.f_next[115] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold1924 (.A(_01403_),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\u_inv.d_next[220] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold1926 (.A(_01251_),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\u_inv.delta_reg[6] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\u_inv.f_next[224] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\u_inv.f_next[235] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold1930 (.A(_01523_),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\u_inv.f_reg[243] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold1932 (.A(_01531_),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\u_inv.d_next[135] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold1934 (.A(_01166_),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\u_inv.f_next[25] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold1936 (.A(_01313_),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\u_inv.f_next[182] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\u_inv.f_next[73] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold1939 (.A(_01361_),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\u_inv.d_next[150] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold1941 (.A(_01181_),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\u_inv.f_next[45] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\u_inv.f_next[200] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold1944 (.A(_01488_),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\u_inv.f_next[15] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\u_inv.d_reg[147] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\u_inv.f_reg[178] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold1948 (.A(_01466_),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\u_inv.d_next[247] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold1950 (.A(_01278_),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\u_inv.f_reg[154] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold1952 (.A(_01442_),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\u_inv.f_reg[184] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold1954 (.A(_01472_),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\u_inv.f_reg[180] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold1956 (.A(_01468_),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\u_inv.f_next[68] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\u_inv.d_reg[223] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\u_inv.d_next[239] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold1960 (.A(_01270_),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\u_inv.f_next[132] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\u_inv.f_next[177] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold1963 (.A(_01465_),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\u_inv.d_next[79] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold1965 (.A(_01110_),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\u_inv.d_next[157] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\u_inv.f_reg[116] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold1968 (.A(_01404_),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\u_inv.f_reg[218] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold1970 (.A(_01506_),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\u_inv.f_reg[18] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold1972 (.A(_01306_),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\u_inv.f_next[243] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\u_inv.f_next[75] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold1975 (.A(_01363_),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\u_inv.f_reg[30] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold1977 (.A(_01318_),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\u_inv.f_next[48] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold1979 (.A(_01336_),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\u_inv.f_next[70] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\u_inv.d_next[96] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold1982 (.A(_01127_),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\u_inv.f_reg[90] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\u_inv.d_next[89] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold1985 (.A(_01120_),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\u_inv.f_reg[228] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold1987 (.A(_01516_),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\u_inv.f_reg[149] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\u_inv.f_next[113] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\u_inv.f_next[33] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold1991 (.A(_01321_),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\u_inv.d_next[23] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold1993 (.A(_01054_),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\u_inv.f_reg[74] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold1995 (.A(_01362_),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\u_inv.f_next[191] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\u_inv.f_next[143] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\u_inv.f_next[137] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\u_inv.f_reg[172] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold2000 (.A(_01460_),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\u_inv.f_next[64] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\u_inv.f_next[49] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\u_inv.d_next[117] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold2004 (.A(_01148_),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\u_inv.d_next[120] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold2006 (.A(_01151_),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\u_inv.f_next[41] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold2008 (.A(_01329_),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\u_inv.counter[5] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold2010 (.A(_00513_),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\u_inv.d_next[133] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold2012 (.A(_01164_),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\u_inv.d_next[187] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold2014 (.A(_01218_),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\u_inv.f_next[184] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\u_inv.f_next[164] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\u_inv.f_next[67] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold2018 (.A(_01355_),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\u_inv.d_next[162] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold2020 (.A(_01193_),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\inv_result[191] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\u_inv.f_next[193] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold2023 (.A(_01481_),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\u_inv.d_next[77] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold2025 (.A(_01108_),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\u_inv.f_reg[16] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold2027 (.A(_01304_),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\u_inv.d_next[219] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold2029 (.A(_01250_),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\u_inv.d_next[10] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold2031 (.A(_01041_),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\u_inv.d_next[215] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold2033 (.A(_01246_),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\u_inv.d_next[106] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold2035 (.A(_01137_),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\u_inv.f_next[186] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\u_inv.f_next[159] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold2038 (.A(_01447_),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\u_inv.f_next[79] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold2040 (.A(_01367_),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\u_inv.d_next[97] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold2042 (.A(_01128_),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold2043 (.A(\u_inv.d_next[214] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\u_inv.f_reg[112] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold2045 (.A(_01400_),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\u_inv.f_next[59] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold2047 (.A(_01347_),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\u_inv.f_next[111] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold2049 (.A(_01399_),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\u_inv.f_reg[124] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold2051 (.A(_01412_),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\u_inv.f_reg[237] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold2053 (.A(_01525_),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\u_inv.f_next[17] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold2055 (.A(_01305_),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\u_inv.f_reg[227] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold2057 (.A(_01515_),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\u_inv.f_reg[217] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold2059 (.A(_01505_),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\u_inv.f_reg[54] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold2061 (.A(_01342_),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\u_inv.d_reg[173] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\u_inv.d_reg[157] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\u_inv.f_reg[219] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold2065 (.A(_01507_),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\u_inv.f_next[99] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\u_inv.d_next[165] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold2068 (.A(_01196_),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\u_inv.f_reg[55] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold2070 (.A(_01343_),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\u_inv.f_reg[102] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold2072 (.A(_01390_),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\u_inv.f_next[42] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\u_inv.f_next[131] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\u_inv.f_next[133] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\u_inv.f_next[206] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\u_inv.f_next[61] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\u_inv.f_next[155] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold2079 (.A(_01443_),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\u_inv.f_next[160] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold2081 (.A(_01448_),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\u_inv.f_next[77] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold2083 (.A(_01365_),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\u_inv.f_next[29] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold2085 (.A(_01317_),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\u_inv.d_reg[163] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\u_inv.f_reg[109] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold2088 (.A(_01397_),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\u_inv.f_next[238] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\u_inv.d_reg[90] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\u_inv.f_next[167] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold2092 (.A(_01455_),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\u_inv.f_next[123] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\u_inv.f_next[233] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold2095 (.A(_01521_),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\u_inv.f_reg[232] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold2097 (.A(_01520_),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\u_inv.f_reg[28] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold2099 (.A(_01316_),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\u_inv.f_reg[135] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold2101 (.A(_01423_),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\inv_result[121] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold2103 (.A(\u_inv.f_reg[72] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold2104 (.A(_01360_),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\u_inv.f_next[156] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\u_inv.f_next[12] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold2107 (.A(_01300_),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\u_inv.f_next[138] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\u_inv.f_reg[216] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold2110 (.A(_01504_),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\u_inv.f_reg[96] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\u_inv.f_next[127] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold2113 (.A(_01415_),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\u_inv.d_next[213] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold2115 (.A(_01244_),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\u_inv.f_reg[53] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold2117 (.A(_01341_),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\u_inv.f_next[151] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold2119 (.A(_01439_),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\u_inv.f_reg[192] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold2121 (.A(_01480_),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\u_inv.f_next[130] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\u_inv.f_next[87] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\u_inv.d_next[221] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold2125 (.A(_01252_),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\u_inv.f_next[46] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\u_inv.f_reg[176] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold2128 (.A(_01464_),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\u_inv.f_next[31] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold2130 (.A(_01319_),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold2131 (.A(\u_inv.f_reg[169] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold2132 (.A(_01457_),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\u_inv.f_next[95] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold2134 (.A(\u_inv.f_reg[195] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold2135 (.A(_01483_),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\u_inv.f_next[78] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\u_inv.f_next[11] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\u_inv.f_next[126] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\u_inv.f_reg[121] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold2140 (.A(_01409_),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\u_inv.f_reg[105] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold2142 (.A(_01393_),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\u_inv.f_next[139] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\u_inv.f_next[10] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\u_inv.f_reg[98] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold2146 (.A(_01386_),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\u_inv.d_next[236] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold2148 (.A(\u_inv.f_next[116] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\u_inv.f_reg[141] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold2150 (.A(_01429_),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\u_inv.f_reg[49] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold2152 (.A(\u_inv.d_next[11] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold2153 (.A(_01042_),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\u_inv.d_next[36] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold2155 (.A(_01067_),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold2156 (.A(\u_inv.f_next[122] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\u_inv.d_next[151] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold2158 (.A(_01182_),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\u_inv.d_next[125] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold2160 (.A(_01156_),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\u_inv.f_next[40] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\u_inv.f_next[227] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\u_inv.d_next[227] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold2164 (.A(_01258_),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\u_inv.f_reg[207] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold2166 (.A(_01495_),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\u_inv.d_reg[214] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\u_inv.d_next[107] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold2169 (.A(_01138_),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\u_inv.f_next[60] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\u_inv.f_next[27] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold2172 (.A(\u_inv.d_next[137] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold2173 (.A(_01168_),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\u_inv.f_reg[71] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold2175 (.A(_01359_),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\u_inv.f_reg[209] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold2177 (.A(_01497_),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\u_inv.counter[6] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\u_inv.f_next[103] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold2180 (.A(_01391_),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\u_inv.f_reg[175] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold2182 (.A(_01463_),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\u_inv.f_next[58] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\u_inv.f_next[76] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\u_inv.f_reg[152] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\u_inv.f_next[112] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\u_inv.f_next[178] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\u_inv.f_next[35] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\u_inv.f_next[108] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\u_inv.f_next[83] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\u_inv.d_next[158] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold2192 (.A(_01189_),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\u_inv.f_next[162] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold2194 (.A(\u_inv.f_reg[60] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold2195 (.A(\u_inv.f_next[231] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\u_inv.f_next[34] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\u_inv.f_reg[93] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold2198 (.A(_01381_),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\u_inv.f_next[104] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold2200 (.A(\u_inv.f_next[38] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\u_inv.f_reg[247] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold2202 (.A(_01535_),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\u_inv.f_next[192] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\u_inv.f_next[195] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\u_inv.f_reg[142] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold2206 (.A(_01430_),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\u_inv.d_next[88] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold2208 (.A(_01119_),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\u_inv.f_next[6] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\u_inv.f_next[13] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\u_inv.f_reg[201] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold2212 (.A(\u_inv.f_next[158] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold2213 (.A(\u_inv.f_next[118] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\u_inv.f_reg[153] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold2215 (.A(_01441_),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold2216 (.A(\u_inv.f_reg[138] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\u_inv.f_reg[157] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold2218 (.A(_01445_),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\u_inv.f_next[170] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\u_inv.f_next[222] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\u_inv.f_reg[37] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold2222 (.A(_01325_),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold2223 (.A(\u_inv.f_next[74] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\u_inv.d_next[121] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold2225 (.A(_01152_),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\u_inv.d_reg[236] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold2227 (.A(\u_inv.f_reg[214] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\u_inv.f_next[26] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\u_inv.f_next[250] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\u_inv.f_next[179] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold2231 (.A(\u_inv.f_reg[57] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\u_inv.f_next[37] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\u_inv.f_next[145] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\u_inv.f_reg[139] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\u_inv.f_next[247] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\u_inv.f_reg[35] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\u_inv.f_next[202] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold2238 (.A(_00173_),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\u_inv.f_reg[39] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold2240 (.A(_01327_),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\u_inv.d_next[50] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold2242 (.A(_01081_),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\u_inv.f_next[30] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\u_inv.f_next[72] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\u_inv.f_next[92] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold2246 (.A(_01380_),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\u_inv.f_next[230] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\u_inv.f_next[55] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\u_inv.f_next[237] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\byte_cnt[2] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\u_inv.f_next[198] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\u_inv.d_next[93] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold2253 (.A(_01124_),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\u_inv.f_next[105] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\u_inv.f_next[180] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\u_inv.f_reg[113] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\u_inv.f_next[32] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\u_inv.f_reg[189] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold2259 (.A(_01477_),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold2260 (.A(\u_inv.f_next[166] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold2261 (.A(\u_inv.f_reg[173] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold2262 (.A(_01461_),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\u_inv.f_next[110] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold2264 (.A(\u_inv.f_next[154] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\u_inv.f_next[226] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\u_inv.f_next[28] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\u_inv.f_next[174] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold2268 (.A(\u_inv.state[1] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold2269 (.A(_19016_),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold2270 (.A(_00000_),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\u_inv.f_next[188] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold2272 (.A(\u_inv.f_next[54] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold2273 (.A(\u_inv.f_next[236] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\u_inv.f_next[242] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\u_inv.f_next[175] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\u_inv.f_next[165] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\u_inv.f_next[18] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold2278 (.A(\u_inv.f_next[157] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\u_inv.f_next[101] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold2280 (.A(\u_inv.counter[8] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\u_inv.f_reg[107] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold2282 (.A(_01395_),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold2283 (.A(\u_inv.f_next[22] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\u_inv.f_reg[239] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold2285 (.A(_01527_),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\u_inv.f_reg[13] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold2287 (.A(\u_inv.f_next[91] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\u_inv.f_next[71] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold2289 (.A(\u_inv.f_next[5] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\u_inv.f_reg[119] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold2291 (.A(_01407_),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\u_inv.f_reg[168] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold2293 (.A(_01456_),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold2294 (.A(\u_inv.f_next[203] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold2295 (.A(\u_inv.f_next[39] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold2296 (.A(\u_inv.f_next[228] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\u_inv.f_next[1] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\u_inv.f_next[140] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\u_inv.f_next[80] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\u_inv.f_next[239] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold2301 (.A(\u_inv.f_next[248] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\u_inv.f_next[234] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\u_inv.f_next[189] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold2304 (.A(\u_inv.f_next[196] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold2305 (.A(\u_inv.delta_double[0] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\u_inv.f_next[53] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold2307 (.A(\u_inv.f_reg[99] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold2308 (.A(\u_inv.counter[3] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\u_inv.f_reg[191] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold2310 (.A(\u_inv.f_next[215] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\u_inv.f_next[98] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\u_inv.f_next[244] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\u_inv.f_reg[171] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold2314 (.A(_01459_),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold2315 (.A(\u_inv.state[0] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold2316 (.A(_14828_),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\u_inv.f_next[169] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold2318 (.A(\u_inv.d_next[98] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\u_inv.f_next[93] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold2320 (.A(\u_inv.f_next[141] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold2321 (.A(\u_inv.d_next[164] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\u_inv.f_next[62] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\u_inv.f_next[119] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\u_inv.f_next[121] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\u_inv.f_next[217] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\u_inv.counter[1] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold2327 (.A(_00509_),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold2328 (.A(\u_inv.f_next[219] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold2329 (.A(\u_inv.f_next[20] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold2330 (.A(\u_inv.f_next[3] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\u_inv.f_next[194] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\u_inv.f_next[16] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold2333 (.A(\u_inv.f_next[218] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold2334 (.A(\u_inv.f_next[171] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\u_inv.f_next[173] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold2336 (.A(\u_inv.f_reg[87] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold2337 (.A(\u_inv.d_next[159] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold2338 (.A(\u_inv.f_next[153] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold2339 (.A(\u_inv.f_next[36] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold2340 (.A(\u_inv.f_next[144] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\u_inv.f_next[114] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\u_inv.f_next[135] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\u_inv.f_next[207] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold2344 (.A(\u_inv.f_next[106] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\u_inv.f_next[209] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold2346 (.A(\u_inv.f_next[134] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold2347 (.A(\u_inv.f_next[2] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\inv_result[241] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\u_inv.d_reg[159] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\u_inv.f_next[232] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold2351 (.A(\u_inv.f_next[172] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\u_inv.f_next[142] ),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\u_inv.f_next[102] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold2354 (.A(inv_done),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\u_inv.d_next[72] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold2356 (.A(_01103_),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\u_inv.f_next[109] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\u_inv.f_next[168] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold2359 (.A(\u_inv.f_next[107] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\u_inv.f_next[176] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\u_inv.f_next[216] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold2362 (.A(\u_inv.f_next[14] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold2363 (.A(\u_inv.f_next[120] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold2364 (.A(\u_inv.counter[2] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold2365 (.A(_00510_),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\u_inv.f_next[124] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold2367 (.A(\u_inv.f_next[147] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold2368 (.A(\u_inv.counter[7] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold2369 (.A(\u_inv.counter[0] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold2370 (.A(\state[1] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold2371 (.A(_14821_),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\state[0] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold2373 (.A(\u_inv.input_valid ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\state[1] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold2375 (.A(\u_inv.d_reg[205] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold2376 (.A(\u_inv.counter[1] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\u_inv.counter[3] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\u_inv.delta_reg[6] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold2379 (.A(\u_inv.d_reg[240] ),
    .X(net3442));
 sg13g2_antennanp ANTENNA_1 (.A(_03302_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(_17242_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_fill_2 FILLER_0_679 ();
 sg13g2_fill_1 FILLER_0_681 ();
 sg13g2_fill_2 FILLER_0_694 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_730 ();
 sg13g2_fill_1 FILLER_0_737 ();
 sg13g2_fill_1 FILLER_0_746 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_4 FILLER_0_759 ();
 sg13g2_fill_2 FILLER_0_763 ();
 sg13g2_decap_4 FILLER_0_773 ();
 sg13g2_fill_2 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_4 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_fill_1 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_4 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_988 ();
 sg13g2_decap_8 FILLER_0_995 ();
 sg13g2_decap_8 FILLER_0_1002 ();
 sg13g2_decap_8 FILLER_0_1009 ();
 sg13g2_decap_8 FILLER_0_1016 ();
 sg13g2_decap_8 FILLER_0_1023 ();
 sg13g2_decap_8 FILLER_0_1030 ();
 sg13g2_decap_8 FILLER_0_1037 ();
 sg13g2_decap_8 FILLER_0_1044 ();
 sg13g2_decap_8 FILLER_0_1051 ();
 sg13g2_decap_8 FILLER_0_1058 ();
 sg13g2_decap_8 FILLER_0_1065 ();
 sg13g2_decap_8 FILLER_0_1072 ();
 sg13g2_decap_8 FILLER_0_1079 ();
 sg13g2_decap_8 FILLER_0_1086 ();
 sg13g2_decap_4 FILLER_0_1093 ();
 sg13g2_decap_8 FILLER_0_1102 ();
 sg13g2_decap_8 FILLER_0_1109 ();
 sg13g2_decap_8 FILLER_0_1126 ();
 sg13g2_decap_4 FILLER_0_1133 ();
 sg13g2_fill_1 FILLER_0_1137 ();
 sg13g2_decap_8 FILLER_0_1159 ();
 sg13g2_decap_8 FILLER_0_1166 ();
 sg13g2_decap_8 FILLER_0_1173 ();
 sg13g2_decap_8 FILLER_0_1180 ();
 sg13g2_fill_2 FILLER_0_1187 ();
 sg13g2_fill_1 FILLER_0_1189 ();
 sg13g2_fill_1 FILLER_0_1195 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_decap_8 FILLER_0_1211 ();
 sg13g2_decap_8 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1225 ();
 sg13g2_decap_8 FILLER_0_1232 ();
 sg13g2_decap_8 FILLER_0_1239 ();
 sg13g2_decap_8 FILLER_0_1246 ();
 sg13g2_decap_8 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1260 ();
 sg13g2_decap_8 FILLER_0_1267 ();
 sg13g2_decap_8 FILLER_0_1274 ();
 sg13g2_decap_8 FILLER_0_1281 ();
 sg13g2_decap_8 FILLER_0_1288 ();
 sg13g2_decap_8 FILLER_0_1295 ();
 sg13g2_decap_8 FILLER_0_1302 ();
 sg13g2_decap_8 FILLER_0_1309 ();
 sg13g2_decap_8 FILLER_0_1316 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1337 ();
 sg13g2_decap_8 FILLER_0_1344 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_8 FILLER_0_1365 ();
 sg13g2_decap_8 FILLER_0_1372 ();
 sg13g2_decap_8 FILLER_0_1379 ();
 sg13g2_decap_8 FILLER_0_1386 ();
 sg13g2_decap_8 FILLER_0_1393 ();
 sg13g2_decap_8 FILLER_0_1400 ();
 sg13g2_decap_8 FILLER_0_1407 ();
 sg13g2_decap_8 FILLER_0_1414 ();
 sg13g2_decap_8 FILLER_0_1421 ();
 sg13g2_decap_8 FILLER_0_1428 ();
 sg13g2_decap_8 FILLER_0_1435 ();
 sg13g2_decap_8 FILLER_0_1442 ();
 sg13g2_decap_8 FILLER_0_1449 ();
 sg13g2_decap_8 FILLER_0_1456 ();
 sg13g2_decap_8 FILLER_0_1463 ();
 sg13g2_decap_8 FILLER_0_1470 ();
 sg13g2_decap_8 FILLER_0_1477 ();
 sg13g2_decap_8 FILLER_0_1484 ();
 sg13g2_decap_8 FILLER_0_1491 ();
 sg13g2_decap_8 FILLER_0_1498 ();
 sg13g2_decap_8 FILLER_0_1505 ();
 sg13g2_decap_8 FILLER_0_1512 ();
 sg13g2_decap_8 FILLER_0_1519 ();
 sg13g2_decap_8 FILLER_0_1526 ();
 sg13g2_decap_8 FILLER_0_1533 ();
 sg13g2_decap_8 FILLER_0_1540 ();
 sg13g2_fill_1 FILLER_0_1547 ();
 sg13g2_decap_8 FILLER_0_1564 ();
 sg13g2_decap_8 FILLER_0_1571 ();
 sg13g2_fill_2 FILLER_0_1578 ();
 sg13g2_fill_2 FILLER_0_1585 ();
 sg13g2_fill_1 FILLER_0_1587 ();
 sg13g2_decap_8 FILLER_0_1601 ();
 sg13g2_decap_8 FILLER_0_1608 ();
 sg13g2_decap_4 FILLER_0_1615 ();
 sg13g2_fill_1 FILLER_0_1623 ();
 sg13g2_decap_8 FILLER_0_1629 ();
 sg13g2_decap_8 FILLER_0_1636 ();
 sg13g2_decap_8 FILLER_0_1643 ();
 sg13g2_decap_8 FILLER_0_1650 ();
 sg13g2_decap_8 FILLER_0_1657 ();
 sg13g2_decap_8 FILLER_0_1664 ();
 sg13g2_decap_8 FILLER_0_1671 ();
 sg13g2_decap_8 FILLER_0_1678 ();
 sg13g2_decap_8 FILLER_0_1685 ();
 sg13g2_decap_8 FILLER_0_1692 ();
 sg13g2_decap_8 FILLER_0_1699 ();
 sg13g2_decap_8 FILLER_0_1706 ();
 sg13g2_decap_8 FILLER_0_1713 ();
 sg13g2_decap_8 FILLER_0_1720 ();
 sg13g2_decap_8 FILLER_0_1727 ();
 sg13g2_decap_8 FILLER_0_1734 ();
 sg13g2_decap_8 FILLER_0_1741 ();
 sg13g2_decap_8 FILLER_0_1748 ();
 sg13g2_fill_2 FILLER_0_1755 ();
 sg13g2_fill_2 FILLER_0_1770 ();
 sg13g2_fill_1 FILLER_0_1772 ();
 sg13g2_fill_1 FILLER_0_1780 ();
 sg13g2_decap_8 FILLER_0_1794 ();
 sg13g2_decap_8 FILLER_0_1801 ();
 sg13g2_decap_8 FILLER_0_1821 ();
 sg13g2_decap_8 FILLER_0_1828 ();
 sg13g2_decap_8 FILLER_0_1835 ();
 sg13g2_decap_8 FILLER_0_1846 ();
 sg13g2_decap_8 FILLER_0_1853 ();
 sg13g2_decap_8 FILLER_0_1860 ();
 sg13g2_decap_8 FILLER_0_1867 ();
 sg13g2_decap_8 FILLER_0_1874 ();
 sg13g2_decap_8 FILLER_0_1881 ();
 sg13g2_decap_8 FILLER_0_1888 ();
 sg13g2_decap_8 FILLER_0_1895 ();
 sg13g2_decap_8 FILLER_0_1902 ();
 sg13g2_decap_8 FILLER_0_1909 ();
 sg13g2_decap_8 FILLER_0_1916 ();
 sg13g2_decap_4 FILLER_0_1923 ();
 sg13g2_fill_2 FILLER_0_1927 ();
 sg13g2_decap_8 FILLER_0_1957 ();
 sg13g2_decap_8 FILLER_0_1964 ();
 sg13g2_decap_8 FILLER_0_1971 ();
 sg13g2_decap_8 FILLER_0_1978 ();
 sg13g2_fill_1 FILLER_0_1985 ();
 sg13g2_fill_2 FILLER_0_1999 ();
 sg13g2_decap_8 FILLER_0_2014 ();
 sg13g2_decap_8 FILLER_0_2021 ();
 sg13g2_decap_8 FILLER_0_2028 ();
 sg13g2_decap_8 FILLER_0_2035 ();
 sg13g2_decap_8 FILLER_0_2042 ();
 sg13g2_decap_8 FILLER_0_2049 ();
 sg13g2_decap_8 FILLER_0_2056 ();
 sg13g2_decap_8 FILLER_0_2063 ();
 sg13g2_decap_8 FILLER_0_2070 ();
 sg13g2_decap_8 FILLER_0_2077 ();
 sg13g2_decap_8 FILLER_0_2084 ();
 sg13g2_decap_8 FILLER_0_2091 ();
 sg13g2_decap_8 FILLER_0_2098 ();
 sg13g2_decap_8 FILLER_0_2105 ();
 sg13g2_decap_8 FILLER_0_2112 ();
 sg13g2_decap_8 FILLER_0_2119 ();
 sg13g2_decap_8 FILLER_0_2126 ();
 sg13g2_decap_8 FILLER_0_2133 ();
 sg13g2_decap_8 FILLER_0_2140 ();
 sg13g2_decap_8 FILLER_0_2147 ();
 sg13g2_decap_4 FILLER_0_2154 ();
 sg13g2_fill_1 FILLER_0_2158 ();
 sg13g2_decap_8 FILLER_0_2185 ();
 sg13g2_decap_8 FILLER_0_2192 ();
 sg13g2_decap_8 FILLER_0_2199 ();
 sg13g2_fill_1 FILLER_0_2206 ();
 sg13g2_decap_8 FILLER_0_2212 ();
 sg13g2_decap_8 FILLER_0_2219 ();
 sg13g2_fill_2 FILLER_0_2226 ();
 sg13g2_fill_1 FILLER_0_2240 ();
 sg13g2_fill_2 FILLER_0_2246 ();
 sg13g2_decap_4 FILLER_0_2253 ();
 sg13g2_fill_2 FILLER_0_2257 ();
 sg13g2_decap_4 FILLER_0_2264 ();
 sg13g2_decap_8 FILLER_0_2276 ();
 sg13g2_decap_4 FILLER_0_2283 ();
 sg13g2_fill_1 FILLER_0_2287 ();
 sg13g2_decap_8 FILLER_0_2309 ();
 sg13g2_decap_8 FILLER_0_2316 ();
 sg13g2_decap_8 FILLER_0_2323 ();
 sg13g2_decap_8 FILLER_0_2330 ();
 sg13g2_decap_8 FILLER_0_2337 ();
 sg13g2_decap_8 FILLER_0_2344 ();
 sg13g2_decap_8 FILLER_0_2351 ();
 sg13g2_decap_8 FILLER_0_2358 ();
 sg13g2_decap_8 FILLER_0_2365 ();
 sg13g2_fill_1 FILLER_0_2372 ();
 sg13g2_decap_8 FILLER_0_2381 ();
 sg13g2_decap_8 FILLER_0_2388 ();
 sg13g2_decap_8 FILLER_0_2395 ();
 sg13g2_decap_8 FILLER_0_2402 ();
 sg13g2_decap_8 FILLER_0_2409 ();
 sg13g2_decap_8 FILLER_0_2416 ();
 sg13g2_decap_8 FILLER_0_2423 ();
 sg13g2_decap_4 FILLER_0_2447 ();
 sg13g2_fill_2 FILLER_0_2463 ();
 sg13g2_fill_1 FILLER_0_2465 ();
 sg13g2_decap_8 FILLER_0_2472 ();
 sg13g2_decap_8 FILLER_0_2479 ();
 sg13g2_fill_2 FILLER_0_2486 ();
 sg13g2_decap_8 FILLER_0_2493 ();
 sg13g2_decap_8 FILLER_0_2500 ();
 sg13g2_decap_8 FILLER_0_2507 ();
 sg13g2_decap_8 FILLER_0_2514 ();
 sg13g2_decap_8 FILLER_0_2521 ();
 sg13g2_decap_8 FILLER_0_2528 ();
 sg13g2_decap_8 FILLER_0_2535 ();
 sg13g2_decap_8 FILLER_0_2542 ();
 sg13g2_decap_8 FILLER_0_2549 ();
 sg13g2_decap_8 FILLER_0_2556 ();
 sg13g2_decap_8 FILLER_0_2563 ();
 sg13g2_decap_4 FILLER_0_2570 ();
 sg13g2_fill_1 FILLER_0_2574 ();
 sg13g2_fill_2 FILLER_0_2583 ();
 sg13g2_decap_8 FILLER_0_2590 ();
 sg13g2_fill_2 FILLER_0_2597 ();
 sg13g2_fill_1 FILLER_0_2599 ();
 sg13g2_fill_1 FILLER_0_2608 ();
 sg13g2_decap_8 FILLER_0_2614 ();
 sg13g2_fill_2 FILLER_0_2621 ();
 sg13g2_fill_2 FILLER_0_2632 ();
 sg13g2_fill_1 FILLER_0_2639 ();
 sg13g2_decap_8 FILLER_0_2644 ();
 sg13g2_decap_8 FILLER_0_2651 ();
 sg13g2_decap_8 FILLER_0_2671 ();
 sg13g2_decap_8 FILLER_0_2678 ();
 sg13g2_decap_8 FILLER_0_2685 ();
 sg13g2_decap_8 FILLER_0_2692 ();
 sg13g2_decap_8 FILLER_0_2699 ();
 sg13g2_decap_8 FILLER_0_2706 ();
 sg13g2_decap_8 FILLER_0_2713 ();
 sg13g2_decap_8 FILLER_0_2720 ();
 sg13g2_decap_8 FILLER_0_2727 ();
 sg13g2_decap_8 FILLER_0_2734 ();
 sg13g2_fill_1 FILLER_0_2749 ();
 sg13g2_decap_8 FILLER_0_2755 ();
 sg13g2_fill_2 FILLER_0_2762 ();
 sg13g2_decap_8 FILLER_0_2775 ();
 sg13g2_decap_8 FILLER_0_2782 ();
 sg13g2_decap_8 FILLER_0_2789 ();
 sg13g2_decap_8 FILLER_0_2796 ();
 sg13g2_decap_8 FILLER_0_2803 ();
 sg13g2_decap_8 FILLER_0_2810 ();
 sg13g2_decap_8 FILLER_0_2817 ();
 sg13g2_decap_8 FILLER_0_2824 ();
 sg13g2_decap_8 FILLER_0_2831 ();
 sg13g2_decap_8 FILLER_0_2838 ();
 sg13g2_decap_8 FILLER_0_2845 ();
 sg13g2_decap_8 FILLER_0_2852 ();
 sg13g2_decap_8 FILLER_0_2859 ();
 sg13g2_decap_4 FILLER_0_2866 ();
 sg13g2_fill_1 FILLER_0_2879 ();
 sg13g2_decap_8 FILLER_0_2885 ();
 sg13g2_decap_4 FILLER_0_2892 ();
 sg13g2_fill_1 FILLER_0_2896 ();
 sg13g2_decap_8 FILLER_0_2915 ();
 sg13g2_decap_8 FILLER_0_2922 ();
 sg13g2_decap_8 FILLER_0_2929 ();
 sg13g2_decap_8 FILLER_0_2936 ();
 sg13g2_decap_8 FILLER_0_2943 ();
 sg13g2_decap_8 FILLER_0_2950 ();
 sg13g2_decap_8 FILLER_0_2957 ();
 sg13g2_decap_8 FILLER_0_2964 ();
 sg13g2_decap_4 FILLER_0_2971 ();
 sg13g2_fill_2 FILLER_0_2975 ();
 sg13g2_decap_8 FILLER_0_2985 ();
 sg13g2_decap_8 FILLER_0_2992 ();
 sg13g2_decap_8 FILLER_0_2999 ();
 sg13g2_decap_8 FILLER_0_3006 ();
 sg13g2_decap_8 FILLER_0_3013 ();
 sg13g2_decap_8 FILLER_0_3020 ();
 sg13g2_fill_2 FILLER_0_3027 ();
 sg13g2_decap_4 FILLER_0_3033 ();
 sg13g2_decap_8 FILLER_0_3042 ();
 sg13g2_decap_4 FILLER_0_3049 ();
 sg13g2_decap_8 FILLER_0_3069 ();
 sg13g2_decap_8 FILLER_0_3076 ();
 sg13g2_decap_8 FILLER_0_3083 ();
 sg13g2_decap_8 FILLER_0_3090 ();
 sg13g2_decap_8 FILLER_0_3097 ();
 sg13g2_decap_8 FILLER_0_3104 ();
 sg13g2_decap_8 FILLER_0_3111 ();
 sg13g2_decap_8 FILLER_0_3118 ();
 sg13g2_decap_8 FILLER_0_3125 ();
 sg13g2_decap_8 FILLER_0_3132 ();
 sg13g2_decap_8 FILLER_0_3139 ();
 sg13g2_decap_8 FILLER_0_3146 ();
 sg13g2_decap_8 FILLER_0_3153 ();
 sg13g2_decap_8 FILLER_0_3160 ();
 sg13g2_decap_8 FILLER_0_3167 ();
 sg13g2_decap_8 FILLER_0_3174 ();
 sg13g2_decap_8 FILLER_0_3181 ();
 sg13g2_decap_8 FILLER_0_3188 ();
 sg13g2_decap_8 FILLER_0_3195 ();
 sg13g2_decap_8 FILLER_0_3202 ();
 sg13g2_decap_8 FILLER_0_3209 ();
 sg13g2_decap_8 FILLER_0_3216 ();
 sg13g2_decap_8 FILLER_0_3223 ();
 sg13g2_decap_8 FILLER_0_3230 ();
 sg13g2_decap_8 FILLER_0_3237 ();
 sg13g2_decap_8 FILLER_0_3244 ();
 sg13g2_decap_8 FILLER_0_3251 ();
 sg13g2_decap_8 FILLER_0_3258 ();
 sg13g2_decap_8 FILLER_0_3265 ();
 sg13g2_decap_8 FILLER_0_3272 ();
 sg13g2_decap_8 FILLER_0_3279 ();
 sg13g2_decap_8 FILLER_0_3286 ();
 sg13g2_decap_8 FILLER_0_3293 ();
 sg13g2_decap_8 FILLER_0_3300 ();
 sg13g2_decap_8 FILLER_0_3307 ();
 sg13g2_decap_8 FILLER_0_3314 ();
 sg13g2_decap_8 FILLER_0_3321 ();
 sg13g2_decap_8 FILLER_0_3328 ();
 sg13g2_decap_8 FILLER_0_3335 ();
 sg13g2_decap_8 FILLER_0_3342 ();
 sg13g2_decap_8 FILLER_0_3349 ();
 sg13g2_decap_8 FILLER_0_3356 ();
 sg13g2_decap_8 FILLER_0_3363 ();
 sg13g2_decap_8 FILLER_0_3370 ();
 sg13g2_decap_8 FILLER_0_3377 ();
 sg13g2_decap_8 FILLER_0_3384 ();
 sg13g2_decap_8 FILLER_0_3391 ();
 sg13g2_decap_8 FILLER_0_3398 ();
 sg13g2_decap_8 FILLER_0_3405 ();
 sg13g2_decap_8 FILLER_0_3412 ();
 sg13g2_decap_8 FILLER_0_3419 ();
 sg13g2_decap_8 FILLER_0_3426 ();
 sg13g2_decap_8 FILLER_0_3433 ();
 sg13g2_decap_8 FILLER_0_3440 ();
 sg13g2_decap_8 FILLER_0_3447 ();
 sg13g2_decap_8 FILLER_0_3454 ();
 sg13g2_decap_8 FILLER_0_3461 ();
 sg13g2_decap_8 FILLER_0_3468 ();
 sg13g2_decap_8 FILLER_0_3475 ();
 sg13g2_decap_8 FILLER_0_3482 ();
 sg13g2_decap_8 FILLER_0_3489 ();
 sg13g2_decap_8 FILLER_0_3496 ();
 sg13g2_decap_8 FILLER_0_3503 ();
 sg13g2_decap_8 FILLER_0_3510 ();
 sg13g2_decap_8 FILLER_0_3517 ();
 sg13g2_decap_8 FILLER_0_3524 ();
 sg13g2_decap_8 FILLER_0_3531 ();
 sg13g2_decap_8 FILLER_0_3538 ();
 sg13g2_decap_8 FILLER_0_3545 ();
 sg13g2_decap_8 FILLER_0_3552 ();
 sg13g2_decap_8 FILLER_0_3559 ();
 sg13g2_decap_8 FILLER_0_3566 ();
 sg13g2_decap_8 FILLER_0_3573 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_4 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_225 ();
 sg13g2_decap_4 FILLER_1_241 ();
 sg13g2_fill_1 FILLER_1_245 ();
 sg13g2_fill_2 FILLER_1_251 ();
 sg13g2_fill_1 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_decap_4 FILLER_1_289 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_8 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_1_412 ();
 sg13g2_decap_8 FILLER_1_419 ();
 sg13g2_decap_8 FILLER_1_426 ();
 sg13g2_decap_8 FILLER_1_433 ();
 sg13g2_decap_8 FILLER_1_440 ();
 sg13g2_decap_8 FILLER_1_447 ();
 sg13g2_decap_8 FILLER_1_454 ();
 sg13g2_decap_8 FILLER_1_461 ();
 sg13g2_decap_8 FILLER_1_468 ();
 sg13g2_decap_8 FILLER_1_475 ();
 sg13g2_decap_8 FILLER_1_482 ();
 sg13g2_decap_8 FILLER_1_489 ();
 sg13g2_decap_8 FILLER_1_496 ();
 sg13g2_decap_8 FILLER_1_503 ();
 sg13g2_decap_8 FILLER_1_510 ();
 sg13g2_decap_8 FILLER_1_517 ();
 sg13g2_decap_8 FILLER_1_524 ();
 sg13g2_decap_8 FILLER_1_531 ();
 sg13g2_decap_8 FILLER_1_538 ();
 sg13g2_decap_8 FILLER_1_545 ();
 sg13g2_decap_8 FILLER_1_552 ();
 sg13g2_decap_8 FILLER_1_559 ();
 sg13g2_decap_8 FILLER_1_566 ();
 sg13g2_decap_8 FILLER_1_573 ();
 sg13g2_decap_8 FILLER_1_580 ();
 sg13g2_decap_8 FILLER_1_587 ();
 sg13g2_decap_8 FILLER_1_594 ();
 sg13g2_decap_8 FILLER_1_601 ();
 sg13g2_decap_8 FILLER_1_612 ();
 sg13g2_decap_8 FILLER_1_619 ();
 sg13g2_decap_8 FILLER_1_626 ();
 sg13g2_fill_2 FILLER_1_633 ();
 sg13g2_decap_4 FILLER_1_663 ();
 sg13g2_fill_1 FILLER_1_667 ();
 sg13g2_fill_1 FILLER_1_676 ();
 sg13g2_fill_1 FILLER_1_706 ();
 sg13g2_decap_8 FILLER_1_727 ();
 sg13g2_decap_4 FILLER_1_734 ();
 sg13g2_decap_4 FILLER_1_750 ();
 sg13g2_fill_2 FILLER_1_759 ();
 sg13g2_fill_2 FILLER_1_783 ();
 sg13g2_fill_1 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_816 ();
 sg13g2_decap_4 FILLER_1_823 ();
 sg13g2_fill_1 FILLER_1_827 ();
 sg13g2_decap_4 FILLER_1_841 ();
 sg13g2_fill_2 FILLER_1_857 ();
 sg13g2_fill_2 FILLER_1_864 ();
 sg13g2_fill_1 FILLER_1_866 ();
 sg13g2_decap_8 FILLER_1_871 ();
 sg13g2_fill_1 FILLER_1_878 ();
 sg13g2_fill_2 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_891 ();
 sg13g2_decap_8 FILLER_1_898 ();
 sg13g2_fill_1 FILLER_1_905 ();
 sg13g2_decap_8 FILLER_1_916 ();
 sg13g2_fill_1 FILLER_1_928 ();
 sg13g2_decap_8 FILLER_1_934 ();
 sg13g2_decap_8 FILLER_1_954 ();
 sg13g2_decap_8 FILLER_1_961 ();
 sg13g2_decap_8 FILLER_1_968 ();
 sg13g2_fill_1 FILLER_1_975 ();
 sg13g2_decap_8 FILLER_1_1007 ();
 sg13g2_fill_2 FILLER_1_1014 ();
 sg13g2_fill_1 FILLER_1_1016 ();
 sg13g2_decap_8 FILLER_1_1030 ();
 sg13g2_decap_8 FILLER_1_1037 ();
 sg13g2_decap_8 FILLER_1_1044 ();
 sg13g2_decap_8 FILLER_1_1051 ();
 sg13g2_decap_8 FILLER_1_1058 ();
 sg13g2_decap_4 FILLER_1_1065 ();
 sg13g2_fill_1 FILLER_1_1069 ();
 sg13g2_decap_4 FILLER_1_1083 ();
 sg13g2_decap_8 FILLER_1_1103 ();
 sg13g2_fill_1 FILLER_1_1123 ();
 sg13g2_fill_1 FILLER_1_1155 ();
 sg13g2_fill_2 FILLER_1_1179 ();
 sg13g2_fill_1 FILLER_1_1181 ();
 sg13g2_decap_8 FILLER_1_1210 ();
 sg13g2_decap_8 FILLER_1_1225 ();
 sg13g2_decap_8 FILLER_1_1232 ();
 sg13g2_decap_8 FILLER_1_1239 ();
 sg13g2_fill_1 FILLER_1_1246 ();
 sg13g2_decap_8 FILLER_1_1260 ();
 sg13g2_decap_8 FILLER_1_1267 ();
 sg13g2_decap_8 FILLER_1_1274 ();
 sg13g2_decap_8 FILLER_1_1281 ();
 sg13g2_decap_8 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1302 ();
 sg13g2_decap_4 FILLER_1_1309 ();
 sg13g2_fill_1 FILLER_1_1313 ();
 sg13g2_decap_8 FILLER_1_1319 ();
 sg13g2_decap_8 FILLER_1_1326 ();
 sg13g2_fill_2 FILLER_1_1333 ();
 sg13g2_fill_1 FILLER_1_1335 ();
 sg13g2_decap_8 FILLER_1_1341 ();
 sg13g2_decap_8 FILLER_1_1348 ();
 sg13g2_decap_8 FILLER_1_1355 ();
 sg13g2_fill_1 FILLER_1_1362 ();
 sg13g2_decap_8 FILLER_1_1368 ();
 sg13g2_decap_8 FILLER_1_1375 ();
 sg13g2_decap_4 FILLER_1_1382 ();
 sg13g2_fill_1 FILLER_1_1386 ();
 sg13g2_decap_8 FILLER_1_1404 ();
 sg13g2_fill_2 FILLER_1_1411 ();
 sg13g2_decap_8 FILLER_1_1417 ();
 sg13g2_decap_8 FILLER_1_1424 ();
 sg13g2_decap_8 FILLER_1_1444 ();
 sg13g2_decap_4 FILLER_1_1457 ();
 sg13g2_decap_8 FILLER_1_1474 ();
 sg13g2_decap_8 FILLER_1_1481 ();
 sg13g2_decap_8 FILLER_1_1488 ();
 sg13g2_decap_8 FILLER_1_1495 ();
 sg13g2_decap_4 FILLER_1_1502 ();
 sg13g2_decap_8 FILLER_1_1511 ();
 sg13g2_decap_4 FILLER_1_1518 ();
 sg13g2_decap_4 FILLER_1_1534 ();
 sg13g2_fill_1 FILLER_1_1538 ();
 sg13g2_decap_4 FILLER_1_1608 ();
 sg13g2_fill_2 FILLER_1_1612 ();
 sg13g2_decap_8 FILLER_1_1642 ();
 sg13g2_decap_8 FILLER_1_1649 ();
 sg13g2_decap_8 FILLER_1_1656 ();
 sg13g2_decap_8 FILLER_1_1663 ();
 sg13g2_fill_2 FILLER_1_1670 ();
 sg13g2_decap_8 FILLER_1_1682 ();
 sg13g2_decap_8 FILLER_1_1689 ();
 sg13g2_fill_1 FILLER_1_1696 ();
 sg13g2_decap_8 FILLER_1_1710 ();
 sg13g2_decap_8 FILLER_1_1717 ();
 sg13g2_decap_8 FILLER_1_1724 ();
 sg13g2_decap_8 FILLER_1_1731 ();
 sg13g2_decap_8 FILLER_1_1738 ();
 sg13g2_decap_8 FILLER_1_1745 ();
 sg13g2_decap_8 FILLER_1_1752 ();
 sg13g2_fill_2 FILLER_1_1759 ();
 sg13g2_decap_4 FILLER_1_1831 ();
 sg13g2_fill_2 FILLER_1_1835 ();
 sg13g2_decap_8 FILLER_1_1865 ();
 sg13g2_decap_8 FILLER_1_1885 ();
 sg13g2_decap_8 FILLER_1_1892 ();
 sg13g2_decap_8 FILLER_1_1899 ();
 sg13g2_fill_2 FILLER_1_1932 ();
 sg13g2_fill_2 FILLER_1_1938 ();
 sg13g2_decap_8 FILLER_1_1944 ();
 sg13g2_decap_8 FILLER_1_1951 ();
 sg13g2_decap_8 FILLER_1_1958 ();
 sg13g2_decap_8 FILLER_1_1965 ();
 sg13g2_fill_2 FILLER_1_1972 ();
 sg13g2_decap_8 FILLER_1_2019 ();
 sg13g2_decap_8 FILLER_1_2026 ();
 sg13g2_decap_8 FILLER_1_2033 ();
 sg13g2_decap_8 FILLER_1_2040 ();
 sg13g2_decap_4 FILLER_1_2047 ();
 sg13g2_fill_2 FILLER_1_2051 ();
 sg13g2_decap_8 FILLER_1_2057 ();
 sg13g2_decap_8 FILLER_1_2064 ();
 sg13g2_decap_8 FILLER_1_2071 ();
 sg13g2_decap_8 FILLER_1_2078 ();
 sg13g2_decap_8 FILLER_1_2085 ();
 sg13g2_decap_8 FILLER_1_2092 ();
 sg13g2_decap_8 FILLER_1_2099 ();
 sg13g2_decap_8 FILLER_1_2106 ();
 sg13g2_fill_1 FILLER_1_2113 ();
 sg13g2_decap_8 FILLER_1_2123 ();
 sg13g2_decap_4 FILLER_1_2130 ();
 sg13g2_decap_8 FILLER_1_2139 ();
 sg13g2_decap_8 FILLER_1_2146 ();
 sg13g2_decap_8 FILLER_1_2153 ();
 sg13g2_decap_4 FILLER_1_2160 ();
 sg13g2_fill_1 FILLER_1_2164 ();
 sg13g2_decap_8 FILLER_1_2170 ();
 sg13g2_decap_8 FILLER_1_2177 ();
 sg13g2_decap_8 FILLER_1_2184 ();
 sg13g2_decap_8 FILLER_1_2191 ();
 sg13g2_fill_2 FILLER_1_2198 ();
 sg13g2_fill_1 FILLER_1_2200 ();
 sg13g2_decap_8 FILLER_1_2210 ();
 sg13g2_decap_4 FILLER_1_2217 ();
 sg13g2_fill_1 FILLER_1_2221 ();
 sg13g2_fill_1 FILLER_1_2235 ();
 sg13g2_fill_2 FILLER_1_2261 ();
 sg13g2_fill_1 FILLER_1_2284 ();
 sg13g2_decap_8 FILLER_1_2312 ();
 sg13g2_decap_8 FILLER_1_2319 ();
 sg13g2_fill_2 FILLER_1_2326 ();
 sg13g2_decap_8 FILLER_1_2337 ();
 sg13g2_decap_4 FILLER_1_2344 ();
 sg13g2_decap_8 FILLER_1_2358 ();
 sg13g2_fill_1 FILLER_1_2365 ();
 sg13g2_decap_8 FILLER_1_2386 ();
 sg13g2_decap_8 FILLER_1_2393 ();
 sg13g2_decap_8 FILLER_1_2400 ();
 sg13g2_decap_8 FILLER_1_2407 ();
 sg13g2_fill_2 FILLER_1_2414 ();
 sg13g2_fill_1 FILLER_1_2421 ();
 sg13g2_fill_1 FILLER_1_2445 ();
 sg13g2_fill_2 FILLER_1_2470 ();
 sg13g2_fill_2 FILLER_1_2481 ();
 sg13g2_decap_8 FILLER_1_2504 ();
 sg13g2_fill_1 FILLER_1_2511 ();
 sg13g2_decap_4 FILLER_1_2525 ();
 sg13g2_decap_8 FILLER_1_2542 ();
 sg13g2_fill_2 FILLER_1_2549 ();
 sg13g2_decap_8 FILLER_1_2555 ();
 sg13g2_decap_4 FILLER_1_2562 ();
 sg13g2_fill_2 FILLER_1_2566 ();
 sg13g2_fill_2 FILLER_1_2576 ();
 sg13g2_fill_1 FILLER_1_2616 ();
 sg13g2_fill_1 FILLER_1_2632 ();
 sg13g2_decap_8 FILLER_1_2654 ();
 sg13g2_fill_2 FILLER_1_2661 ();
 sg13g2_decap_4 FILLER_1_2676 ();
 sg13g2_fill_1 FILLER_1_2680 ();
 sg13g2_decap_8 FILLER_1_2689 ();
 sg13g2_fill_1 FILLER_1_2696 ();
 sg13g2_decap_8 FILLER_1_2712 ();
 sg13g2_decap_4 FILLER_1_2719 ();
 sg13g2_fill_2 FILLER_1_2723 ();
 sg13g2_fill_1 FILLER_1_2746 ();
 sg13g2_decap_8 FILLER_1_2779 ();
 sg13g2_decap_8 FILLER_1_2786 ();
 sg13g2_decap_8 FILLER_1_2793 ();
 sg13g2_decap_8 FILLER_1_2800 ();
 sg13g2_decap_8 FILLER_1_2807 ();
 sg13g2_decap_8 FILLER_1_2814 ();
 sg13g2_decap_8 FILLER_1_2821 ();
 sg13g2_decap_8 FILLER_1_2828 ();
 sg13g2_decap_8 FILLER_1_2835 ();
 sg13g2_decap_8 FILLER_1_2842 ();
 sg13g2_decap_8 FILLER_1_2849 ();
 sg13g2_decap_8 FILLER_1_2856 ();
 sg13g2_decap_4 FILLER_1_2863 ();
 sg13g2_fill_2 FILLER_1_2895 ();
 sg13g2_decap_4 FILLER_1_2910 ();
 sg13g2_fill_1 FILLER_1_2932 ();
 sg13g2_decap_8 FILLER_1_2945 ();
 sg13g2_fill_2 FILLER_1_2952 ();
 sg13g2_fill_2 FILLER_1_2967 ();
 sg13g2_decap_8 FILLER_1_2994 ();
 sg13g2_fill_1 FILLER_1_3001 ();
 sg13g2_fill_2 FILLER_1_3022 ();
 sg13g2_fill_2 FILLER_1_3041 ();
 sg13g2_fill_1 FILLER_1_3043 ();
 sg13g2_fill_1 FILLER_1_3052 ();
 sg13g2_decap_4 FILLER_1_3085 ();
 sg13g2_fill_1 FILLER_1_3089 ();
 sg13g2_decap_8 FILLER_1_3095 ();
 sg13g2_decap_8 FILLER_1_3102 ();
 sg13g2_decap_8 FILLER_1_3109 ();
 sg13g2_decap_8 FILLER_1_3116 ();
 sg13g2_fill_2 FILLER_1_3123 ();
 sg13g2_decap_8 FILLER_1_3130 ();
 sg13g2_decap_8 FILLER_1_3137 ();
 sg13g2_decap_8 FILLER_1_3144 ();
 sg13g2_decap_8 FILLER_1_3151 ();
 sg13g2_decap_4 FILLER_1_3158 ();
 sg13g2_decap_8 FILLER_1_3170 ();
 sg13g2_decap_8 FILLER_1_3177 ();
 sg13g2_decap_8 FILLER_1_3184 ();
 sg13g2_decap_8 FILLER_1_3191 ();
 sg13g2_decap_8 FILLER_1_3198 ();
 sg13g2_decap_8 FILLER_1_3205 ();
 sg13g2_fill_1 FILLER_1_3212 ();
 sg13g2_decap_8 FILLER_1_3226 ();
 sg13g2_decap_8 FILLER_1_3233 ();
 sg13g2_decap_8 FILLER_1_3240 ();
 sg13g2_decap_8 FILLER_1_3247 ();
 sg13g2_decap_8 FILLER_1_3254 ();
 sg13g2_decap_8 FILLER_1_3261 ();
 sg13g2_decap_8 FILLER_1_3268 ();
 sg13g2_decap_8 FILLER_1_3275 ();
 sg13g2_decap_8 FILLER_1_3282 ();
 sg13g2_decap_8 FILLER_1_3289 ();
 sg13g2_decap_8 FILLER_1_3296 ();
 sg13g2_decap_8 FILLER_1_3303 ();
 sg13g2_decap_8 FILLER_1_3310 ();
 sg13g2_decap_8 FILLER_1_3317 ();
 sg13g2_decap_8 FILLER_1_3324 ();
 sg13g2_decap_8 FILLER_1_3331 ();
 sg13g2_decap_8 FILLER_1_3338 ();
 sg13g2_decap_8 FILLER_1_3345 ();
 sg13g2_decap_8 FILLER_1_3352 ();
 sg13g2_decap_8 FILLER_1_3359 ();
 sg13g2_decap_8 FILLER_1_3366 ();
 sg13g2_decap_8 FILLER_1_3373 ();
 sg13g2_decap_8 FILLER_1_3380 ();
 sg13g2_decap_8 FILLER_1_3387 ();
 sg13g2_decap_8 FILLER_1_3394 ();
 sg13g2_decap_8 FILLER_1_3401 ();
 sg13g2_decap_8 FILLER_1_3408 ();
 sg13g2_decap_8 FILLER_1_3415 ();
 sg13g2_decap_8 FILLER_1_3422 ();
 sg13g2_decap_8 FILLER_1_3429 ();
 sg13g2_decap_8 FILLER_1_3436 ();
 sg13g2_decap_8 FILLER_1_3443 ();
 sg13g2_decap_8 FILLER_1_3450 ();
 sg13g2_decap_8 FILLER_1_3457 ();
 sg13g2_decap_8 FILLER_1_3464 ();
 sg13g2_decap_8 FILLER_1_3471 ();
 sg13g2_decap_8 FILLER_1_3478 ();
 sg13g2_decap_8 FILLER_1_3485 ();
 sg13g2_decap_8 FILLER_1_3492 ();
 sg13g2_decap_8 FILLER_1_3499 ();
 sg13g2_decap_8 FILLER_1_3506 ();
 sg13g2_decap_8 FILLER_1_3513 ();
 sg13g2_decap_8 FILLER_1_3520 ();
 sg13g2_decap_8 FILLER_1_3527 ();
 sg13g2_decap_8 FILLER_1_3534 ();
 sg13g2_decap_8 FILLER_1_3541 ();
 sg13g2_decap_8 FILLER_1_3548 ();
 sg13g2_decap_8 FILLER_1_3555 ();
 sg13g2_decap_8 FILLER_1_3562 ();
 sg13g2_decap_8 FILLER_1_3569 ();
 sg13g2_decap_4 FILLER_1_3576 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_fill_2 FILLER_2_175 ();
 sg13g2_fill_1 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_192 ();
 sg13g2_decap_4 FILLER_2_199 ();
 sg13g2_fill_2 FILLER_2_207 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_fill_1 FILLER_2_243 ();
 sg13g2_fill_2 FILLER_2_254 ();
 sg13g2_fill_1 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_fill_2 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_4 FILLER_2_292 ();
 sg13g2_fill_2 FILLER_2_296 ();
 sg13g2_decap_8 FILLER_2_302 ();
 sg13g2_decap_4 FILLER_2_309 ();
 sg13g2_fill_2 FILLER_2_313 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_fill_2 FILLER_2_326 ();
 sg13g2_fill_1 FILLER_2_328 ();
 sg13g2_fill_1 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_4 FILLER_2_532 ();
 sg13g2_fill_2 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_547 ();
 sg13g2_decap_8 FILLER_2_554 ();
 sg13g2_decap_8 FILLER_2_561 ();
 sg13g2_decap_8 FILLER_2_568 ();
 sg13g2_decap_8 FILLER_2_575 ();
 sg13g2_fill_1 FILLER_2_582 ();
 sg13g2_decap_4 FILLER_2_631 ();
 sg13g2_fill_2 FILLER_2_635 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_fill_2 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_675 ();
 sg13g2_decap_4 FILLER_2_682 ();
 sg13g2_fill_2 FILLER_2_686 ();
 sg13g2_fill_2 FILLER_2_698 ();
 sg13g2_fill_1 FILLER_2_705 ();
 sg13g2_fill_1 FILLER_2_718 ();
 sg13g2_decap_4 FILLER_2_731 ();
 sg13g2_fill_1 FILLER_2_735 ();
 sg13g2_fill_1 FILLER_2_751 ();
 sg13g2_fill_2 FILLER_2_769 ();
 sg13g2_fill_1 FILLER_2_784 ();
 sg13g2_decap_4 FILLER_2_796 ();
 sg13g2_fill_2 FILLER_2_800 ();
 sg13g2_fill_1 FILLER_2_806 ();
 sg13g2_decap_8 FILLER_2_814 ();
 sg13g2_decap_8 FILLER_2_821 ();
 sg13g2_fill_2 FILLER_2_828 ();
 sg13g2_fill_2 FILLER_2_843 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_fill_2 FILLER_2_926 ();
 sg13g2_decap_4 FILLER_2_936 ();
 sg13g2_fill_2 FILLER_2_947 ();
 sg13g2_fill_1 FILLER_2_949 ();
 sg13g2_fill_2 FILLER_2_969 ();
 sg13g2_fill_1 FILLER_2_971 ();
 sg13g2_decap_8 FILLER_2_982 ();
 sg13g2_fill_2 FILLER_2_989 ();
 sg13g2_fill_2 FILLER_2_999 ();
 sg13g2_fill_1 FILLER_2_1001 ();
 sg13g2_fill_2 FILLER_2_1015 ();
 sg13g2_fill_1 FILLER_2_1017 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_2_1042 ();
 sg13g2_decap_8 FILLER_2_1049 ();
 sg13g2_fill_2 FILLER_2_1056 ();
 sg13g2_decap_8 FILLER_2_1065 ();
 sg13g2_decap_8 FILLER_2_1072 ();
 sg13g2_decap_4 FILLER_2_1079 ();
 sg13g2_decap_4 FILLER_2_1096 ();
 sg13g2_fill_2 FILLER_2_1112 ();
 sg13g2_fill_1 FILLER_2_1114 ();
 sg13g2_decap_8 FILLER_2_1127 ();
 sg13g2_decap_4 FILLER_2_1134 ();
 sg13g2_decap_8 FILLER_2_1161 ();
 sg13g2_decap_4 FILLER_2_1168 ();
 sg13g2_fill_2 FILLER_2_1172 ();
 sg13g2_fill_2 FILLER_2_1204 ();
 sg13g2_fill_1 FILLER_2_1206 ();
 sg13g2_decap_8 FILLER_2_1235 ();
 sg13g2_decap_8 FILLER_2_1242 ();
 sg13g2_decap_8 FILLER_2_1249 ();
 sg13g2_decap_8 FILLER_2_1256 ();
 sg13g2_decap_8 FILLER_2_1263 ();
 sg13g2_decap_8 FILLER_2_1288 ();
 sg13g2_decap_8 FILLER_2_1295 ();
 sg13g2_decap_4 FILLER_2_1327 ();
 sg13g2_fill_2 FILLER_2_1344 ();
 sg13g2_decap_8 FILLER_2_1375 ();
 sg13g2_decap_8 FILLER_2_1382 ();
 sg13g2_fill_1 FILLER_2_1389 ();
 sg13g2_decap_8 FILLER_2_1421 ();
 sg13g2_fill_2 FILLER_2_1432 ();
 sg13g2_fill_1 FILLER_2_1434 ();
 sg13g2_fill_2 FILLER_2_1440 ();
 sg13g2_fill_2 FILLER_2_1446 ();
 sg13g2_fill_1 FILLER_2_1448 ();
 sg13g2_decap_8 FILLER_2_1466 ();
 sg13g2_decap_8 FILLER_2_1473 ();
 sg13g2_decap_4 FILLER_2_1480 ();
 sg13g2_decap_8 FILLER_2_1497 ();
 sg13g2_decap_4 FILLER_2_1511 ();
 sg13g2_fill_1 FILLER_2_1515 ();
 sg13g2_decap_8 FILLER_2_1523 ();
 sg13g2_fill_2 FILLER_2_1530 ();
 sg13g2_fill_2 FILLER_2_1545 ();
 sg13g2_fill_2 FILLER_2_1552 ();
 sg13g2_decap_8 FILLER_2_1567 ();
 sg13g2_decap_4 FILLER_2_1574 ();
 sg13g2_fill_1 FILLER_2_1578 ();
 sg13g2_decap_8 FILLER_2_1597 ();
 sg13g2_decap_8 FILLER_2_1604 ();
 sg13g2_fill_1 FILLER_2_1611 ();
 sg13g2_decap_4 FILLER_2_1621 ();
 sg13g2_fill_1 FILLER_2_1637 ();
 sg13g2_decap_8 FILLER_2_1643 ();
 sg13g2_fill_2 FILLER_2_1654 ();
 sg13g2_fill_2 FILLER_2_1664 ();
 sg13g2_fill_1 FILLER_2_1666 ();
 sg13g2_decap_8 FILLER_2_1688 ();
 sg13g2_decap_4 FILLER_2_1695 ();
 sg13g2_decap_4 FILLER_2_1709 ();
 sg13g2_fill_2 FILLER_2_1713 ();
 sg13g2_fill_2 FILLER_2_1743 ();
 sg13g2_decap_8 FILLER_2_1758 ();
 sg13g2_decap_4 FILLER_2_1765 ();
 sg13g2_fill_2 FILLER_2_1787 ();
 sg13g2_fill_1 FILLER_2_1789 ();
 sg13g2_decap_8 FILLER_2_1794 ();
 sg13g2_decap_8 FILLER_2_1801 ();
 sg13g2_decap_4 FILLER_2_1830 ();
 sg13g2_fill_1 FILLER_2_1834 ();
 sg13g2_decap_4 FILLER_2_1839 ();
 sg13g2_decap_4 FILLER_2_1847 ();
 sg13g2_fill_2 FILLER_2_1879 ();
 sg13g2_decap_8 FILLER_2_1909 ();
 sg13g2_fill_1 FILLER_2_1916 ();
 sg13g2_fill_2 FILLER_2_1930 ();
 sg13g2_fill_1 FILLER_2_1943 ();
 sg13g2_decap_8 FILLER_2_1952 ();
 sg13g2_fill_1 FILLER_2_1967 ();
 sg13g2_decap_8 FILLER_2_1980 ();
 sg13g2_fill_2 FILLER_2_1987 ();
 sg13g2_fill_2 FILLER_2_1992 ();
 sg13g2_decap_8 FILLER_2_1999 ();
 sg13g2_decap_4 FILLER_2_2006 ();
 sg13g2_fill_2 FILLER_2_2010 ();
 sg13g2_decap_8 FILLER_2_2033 ();
 sg13g2_decap_4 FILLER_2_2040 ();
 sg13g2_fill_1 FILLER_2_2044 ();
 sg13g2_fill_1 FILLER_2_2055 ();
 sg13g2_decap_8 FILLER_2_2061 ();
 sg13g2_decap_8 FILLER_2_2068 ();
 sg13g2_decap_8 FILLER_2_2075 ();
 sg13g2_decap_8 FILLER_2_2082 ();
 sg13g2_decap_8 FILLER_2_2089 ();
 sg13g2_decap_8 FILLER_2_2096 ();
 sg13g2_decap_8 FILLER_2_2103 ();
 sg13g2_decap_4 FILLER_2_2110 ();
 sg13g2_decap_8 FILLER_2_2142 ();
 sg13g2_fill_2 FILLER_2_2149 ();
 sg13g2_fill_1 FILLER_2_2151 ();
 sg13g2_fill_2 FILLER_2_2160 ();
 sg13g2_fill_2 FILLER_2_2177 ();
 sg13g2_fill_1 FILLER_2_2179 ();
 sg13g2_fill_2 FILLER_2_2188 ();
 sg13g2_decap_8 FILLER_2_2215 ();
 sg13g2_decap_4 FILLER_2_2222 ();
 sg13g2_fill_1 FILLER_2_2226 ();
 sg13g2_fill_2 FILLER_2_2230 ();
 sg13g2_fill_2 FILLER_2_2237 ();
 sg13g2_decap_8 FILLER_2_2244 ();
 sg13g2_decap_4 FILLER_2_2251 ();
 sg13g2_decap_4 FILLER_2_2259 ();
 sg13g2_fill_1 FILLER_2_2263 ();
 sg13g2_decap_8 FILLER_2_2274 ();
 sg13g2_decap_4 FILLER_2_2281 ();
 sg13g2_fill_2 FILLER_2_2285 ();
 sg13g2_decap_4 FILLER_2_2312 ();
 sg13g2_fill_1 FILLER_2_2316 ();
 sg13g2_decap_8 FILLER_2_2341 ();
 sg13g2_fill_2 FILLER_2_2348 ();
 sg13g2_decap_8 FILLER_2_2362 ();
 sg13g2_fill_1 FILLER_2_2369 ();
 sg13g2_decap_8 FILLER_2_2392 ();
 sg13g2_decap_8 FILLER_2_2399 ();
 sg13g2_decap_4 FILLER_2_2406 ();
 sg13g2_fill_1 FILLER_2_2410 ();
 sg13g2_decap_8 FILLER_2_2424 ();
 sg13g2_fill_2 FILLER_2_2431 ();
 sg13g2_fill_1 FILLER_2_2433 ();
 sg13g2_fill_1 FILLER_2_2444 ();
 sg13g2_decap_8 FILLER_2_2450 ();
 sg13g2_decap_8 FILLER_2_2457 ();
 sg13g2_fill_2 FILLER_2_2464 ();
 sg13g2_fill_1 FILLER_2_2466 ();
 sg13g2_decap_8 FILLER_2_2510 ();
 sg13g2_fill_1 FILLER_2_2517 ();
 sg13g2_decap_8 FILLER_2_2525 ();
 sg13g2_decap_8 FILLER_2_2532 ();
 sg13g2_decap_4 FILLER_2_2539 ();
 sg13g2_fill_2 FILLER_2_2543 ();
 sg13g2_fill_2 FILLER_2_2551 ();
 sg13g2_fill_1 FILLER_2_2553 ();
 sg13g2_decap_8 FILLER_2_2559 ();
 sg13g2_fill_2 FILLER_2_2566 ();
 sg13g2_decap_8 FILLER_2_2589 ();
 sg13g2_decap_4 FILLER_2_2596 ();
 sg13g2_decap_8 FILLER_2_2608 ();
 sg13g2_decap_8 FILLER_2_2615 ();
 sg13g2_fill_2 FILLER_2_2622 ();
 sg13g2_fill_1 FILLER_2_2624 ();
 sg13g2_decap_4 FILLER_2_2630 ();
 sg13g2_fill_2 FILLER_2_2634 ();
 sg13g2_decap_4 FILLER_2_2641 ();
 sg13g2_fill_2 FILLER_2_2645 ();
 sg13g2_decap_4 FILLER_2_2651 ();
 sg13g2_fill_1 FILLER_2_2655 ();
 sg13g2_fill_2 FILLER_2_2659 ();
 sg13g2_fill_1 FILLER_2_2661 ();
 sg13g2_decap_4 FILLER_2_2675 ();
 sg13g2_fill_2 FILLER_2_2679 ();
 sg13g2_fill_1 FILLER_2_2720 ();
 sg13g2_fill_2 FILLER_2_2739 ();
 sg13g2_decap_8 FILLER_2_2759 ();
 sg13g2_decap_8 FILLER_2_2776 ();
 sg13g2_decap_8 FILLER_2_2783 ();
 sg13g2_decap_8 FILLER_2_2790 ();
 sg13g2_decap_8 FILLER_2_2797 ();
 sg13g2_fill_2 FILLER_2_2804 ();
 sg13g2_fill_1 FILLER_2_2806 ();
 sg13g2_decap_8 FILLER_2_2820 ();
 sg13g2_decap_4 FILLER_2_2855 ();
 sg13g2_fill_1 FILLER_2_2859 ();
 sg13g2_decap_8 FILLER_2_2869 ();
 sg13g2_fill_2 FILLER_2_2876 ();
 sg13g2_fill_2 FILLER_2_2883 ();
 sg13g2_fill_2 FILLER_2_2895 ();
 sg13g2_fill_1 FILLER_2_2897 ();
 sg13g2_decap_8 FILLER_2_2906 ();
 sg13g2_decap_4 FILLER_2_2913 ();
 sg13g2_fill_2 FILLER_2_2917 ();
 sg13g2_decap_4 FILLER_2_2933 ();
 sg13g2_decap_8 FILLER_2_2949 ();
 sg13g2_decap_8 FILLER_2_2956 ();
 sg13g2_decap_4 FILLER_2_2963 ();
 sg13g2_fill_1 FILLER_2_2967 ();
 sg13g2_decap_8 FILLER_2_2987 ();
 sg13g2_decap_8 FILLER_2_2994 ();
 sg13g2_decap_4 FILLER_2_3001 ();
 sg13g2_fill_2 FILLER_2_3005 ();
 sg13g2_decap_8 FILLER_2_3014 ();
 sg13g2_decap_8 FILLER_2_3026 ();
 sg13g2_decap_4 FILLER_2_3033 ();
 sg13g2_fill_2 FILLER_2_3037 ();
 sg13g2_decap_4 FILLER_2_3044 ();
 sg13g2_decap_8 FILLER_2_3069 ();
 sg13g2_decap_8 FILLER_2_3076 ();
 sg13g2_fill_2 FILLER_2_3083 ();
 sg13g2_fill_2 FILLER_2_3090 ();
 sg13g2_fill_1 FILLER_2_3092 ();
 sg13g2_decap_8 FILLER_2_3103 ();
 sg13g2_decap_8 FILLER_2_3110 ();
 sg13g2_fill_2 FILLER_2_3117 ();
 sg13g2_decap_8 FILLER_2_3135 ();
 sg13g2_decap_8 FILLER_2_3142 ();
 sg13g2_decap_8 FILLER_2_3149 ();
 sg13g2_decap_4 FILLER_2_3156 ();
 sg13g2_fill_2 FILLER_2_3160 ();
 sg13g2_fill_2 FILLER_2_3178 ();
 sg13g2_fill_1 FILLER_2_3180 ();
 sg13g2_decap_8 FILLER_2_3190 ();
 sg13g2_fill_2 FILLER_2_3197 ();
 sg13g2_fill_1 FILLER_2_3199 ();
 sg13g2_decap_4 FILLER_2_3207 ();
 sg13g2_decap_8 FILLER_2_3220 ();
 sg13g2_decap_8 FILLER_2_3227 ();
 sg13g2_decap_8 FILLER_2_3234 ();
 sg13g2_decap_8 FILLER_2_3241 ();
 sg13g2_decap_8 FILLER_2_3248 ();
 sg13g2_decap_8 FILLER_2_3255 ();
 sg13g2_decap_8 FILLER_2_3262 ();
 sg13g2_decap_8 FILLER_2_3269 ();
 sg13g2_decap_8 FILLER_2_3276 ();
 sg13g2_decap_8 FILLER_2_3283 ();
 sg13g2_decap_8 FILLER_2_3290 ();
 sg13g2_decap_8 FILLER_2_3297 ();
 sg13g2_decap_8 FILLER_2_3304 ();
 sg13g2_decap_8 FILLER_2_3311 ();
 sg13g2_decap_8 FILLER_2_3318 ();
 sg13g2_decap_8 FILLER_2_3325 ();
 sg13g2_decap_8 FILLER_2_3332 ();
 sg13g2_fill_2 FILLER_2_3339 ();
 sg13g2_decap_8 FILLER_2_3351 ();
 sg13g2_decap_8 FILLER_2_3358 ();
 sg13g2_decap_8 FILLER_2_3365 ();
 sg13g2_decap_8 FILLER_2_3372 ();
 sg13g2_decap_8 FILLER_2_3379 ();
 sg13g2_decap_8 FILLER_2_3386 ();
 sg13g2_decap_8 FILLER_2_3393 ();
 sg13g2_decap_8 FILLER_2_3400 ();
 sg13g2_decap_8 FILLER_2_3407 ();
 sg13g2_decap_8 FILLER_2_3414 ();
 sg13g2_decap_8 FILLER_2_3421 ();
 sg13g2_decap_8 FILLER_2_3428 ();
 sg13g2_decap_8 FILLER_2_3435 ();
 sg13g2_decap_8 FILLER_2_3442 ();
 sg13g2_decap_8 FILLER_2_3449 ();
 sg13g2_decap_8 FILLER_2_3456 ();
 sg13g2_decap_8 FILLER_2_3463 ();
 sg13g2_decap_8 FILLER_2_3470 ();
 sg13g2_decap_8 FILLER_2_3477 ();
 sg13g2_decap_8 FILLER_2_3484 ();
 sg13g2_decap_8 FILLER_2_3491 ();
 sg13g2_decap_8 FILLER_2_3498 ();
 sg13g2_decap_8 FILLER_2_3505 ();
 sg13g2_decap_8 FILLER_2_3512 ();
 sg13g2_decap_8 FILLER_2_3519 ();
 sg13g2_decap_8 FILLER_2_3526 ();
 sg13g2_decap_8 FILLER_2_3533 ();
 sg13g2_decap_8 FILLER_2_3540 ();
 sg13g2_decap_8 FILLER_2_3547 ();
 sg13g2_decap_8 FILLER_2_3554 ();
 sg13g2_decap_8 FILLER_2_3561 ();
 sg13g2_decap_8 FILLER_2_3568 ();
 sg13g2_decap_4 FILLER_2_3575 ();
 sg13g2_fill_1 FILLER_2_3579 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_140 ();
 sg13g2_fill_2 FILLER_3_144 ();
 sg13g2_decap_4 FILLER_3_158 ();
 sg13g2_fill_2 FILLER_3_194 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_fill_2 FILLER_3_224 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_fill_2 FILLER_3_240 ();
 sg13g2_fill_1 FILLER_3_250 ();
 sg13g2_decap_4 FILLER_3_263 ();
 sg13g2_fill_2 FILLER_3_267 ();
 sg13g2_fill_1 FILLER_3_289 ();
 sg13g2_fill_2 FILLER_3_295 ();
 sg13g2_fill_1 FILLER_3_297 ();
 sg13g2_fill_2 FILLER_3_314 ();
 sg13g2_fill_2 FILLER_3_321 ();
 sg13g2_fill_1 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_fill_2 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_decap_8 FILLER_3_430 ();
 sg13g2_decap_8 FILLER_3_437 ();
 sg13g2_decap_8 FILLER_3_444 ();
 sg13g2_decap_8 FILLER_3_451 ();
 sg13g2_decap_8 FILLER_3_458 ();
 sg13g2_decap_8 FILLER_3_465 ();
 sg13g2_fill_1 FILLER_3_472 ();
 sg13g2_decap_8 FILLER_3_486 ();
 sg13g2_decap_8 FILLER_3_493 ();
 sg13g2_decap_8 FILLER_3_500 ();
 sg13g2_decap_8 FILLER_3_507 ();
 sg13g2_decap_8 FILLER_3_514 ();
 sg13g2_decap_8 FILLER_3_554 ();
 sg13g2_decap_8 FILLER_3_561 ();
 sg13g2_decap_4 FILLER_3_568 ();
 sg13g2_fill_1 FILLER_3_576 ();
 sg13g2_decap_8 FILLER_3_598 ();
 sg13g2_fill_2 FILLER_3_605 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_8 FILLER_3_620 ();
 sg13g2_fill_1 FILLER_3_627 ();
 sg13g2_fill_1 FILLER_3_641 ();
 sg13g2_decap_8 FILLER_3_646 ();
 sg13g2_fill_2 FILLER_3_659 ();
 sg13g2_fill_2 FILLER_3_676 ();
 sg13g2_fill_1 FILLER_3_678 ();
 sg13g2_fill_2 FILLER_3_688 ();
 sg13g2_fill_1 FILLER_3_708 ();
 sg13g2_decap_8 FILLER_3_723 ();
 sg13g2_decap_4 FILLER_3_730 ();
 sg13g2_decap_8 FILLER_3_739 ();
 sg13g2_decap_4 FILLER_3_746 ();
 sg13g2_fill_2 FILLER_3_750 ();
 sg13g2_fill_1 FILLER_3_780 ();
 sg13g2_fill_1 FILLER_3_785 ();
 sg13g2_fill_1 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_799 ();
 sg13g2_decap_8 FILLER_3_806 ();
 sg13g2_fill_2 FILLER_3_813 ();
 sg13g2_fill_1 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_821 ();
 sg13g2_fill_2 FILLER_3_828 ();
 sg13g2_fill_1 FILLER_3_830 ();
 sg13g2_decap_4 FILLER_3_844 ();
 sg13g2_fill_2 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_856 ();
 sg13g2_decap_8 FILLER_3_866 ();
 sg13g2_decap_8 FILLER_3_873 ();
 sg13g2_decap_8 FILLER_3_880 ();
 sg13g2_decap_8 FILLER_3_887 ();
 sg13g2_decap_4 FILLER_3_894 ();
 sg13g2_fill_1 FILLER_3_898 ();
 sg13g2_fill_1 FILLER_3_904 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_decap_4 FILLER_3_921 ();
 sg13g2_fill_2 FILLER_3_925 ();
 sg13g2_fill_1 FILLER_3_932 ();
 sg13g2_decap_8 FILLER_3_937 ();
 sg13g2_decap_8 FILLER_3_944 ();
 sg13g2_decap_8 FILLER_3_951 ();
 sg13g2_decap_8 FILLER_3_958 ();
 sg13g2_decap_4 FILLER_3_965 ();
 sg13g2_fill_2 FILLER_3_969 ();
 sg13g2_fill_1 FILLER_3_986 ();
 sg13g2_fill_2 FILLER_3_1028 ();
 sg13g2_fill_1 FILLER_3_1030 ();
 sg13g2_decap_4 FILLER_3_1047 ();
 sg13g2_fill_2 FILLER_3_1051 ();
 sg13g2_fill_2 FILLER_3_1081 ();
 sg13g2_fill_1 FILLER_3_1083 ();
 sg13g2_fill_2 FILLER_3_1149 ();
 sg13g2_fill_1 FILLER_3_1151 ();
 sg13g2_fill_1 FILLER_3_1157 ();
 sg13g2_fill_1 FILLER_3_1168 ();
 sg13g2_decap_4 FILLER_3_1186 ();
 sg13g2_decap_4 FILLER_3_1204 ();
 sg13g2_fill_1 FILLER_3_1208 ();
 sg13g2_fill_1 FILLER_3_1213 ();
 sg13g2_decap_4 FILLER_3_1224 ();
 sg13g2_decap_4 FILLER_3_1237 ();
 sg13g2_fill_1 FILLER_3_1241 ();
 sg13g2_decap_4 FILLER_3_1270 ();
 sg13g2_decap_8 FILLER_3_1287 ();
 sg13g2_decap_8 FILLER_3_1294 ();
 sg13g2_fill_2 FILLER_3_1301 ();
 sg13g2_decap_8 FILLER_3_1324 ();
 sg13g2_decap_4 FILLER_3_1331 ();
 sg13g2_fill_1 FILLER_3_1335 ();
 sg13g2_decap_8 FILLER_3_1351 ();
 sg13g2_decap_4 FILLER_3_1358 ();
 sg13g2_decap_4 FILLER_3_1370 ();
 sg13g2_fill_2 FILLER_3_1374 ();
 sg13g2_decap_8 FILLER_3_1380 ();
 sg13g2_decap_4 FILLER_3_1387 ();
 sg13g2_fill_2 FILLER_3_1391 ();
 sg13g2_fill_2 FILLER_3_1406 ();
 sg13g2_fill_1 FILLER_3_1408 ();
 sg13g2_fill_2 FILLER_3_1417 ();
 sg13g2_fill_1 FILLER_3_1419 ();
 sg13g2_fill_1 FILLER_3_1455 ();
 sg13g2_decap_8 FILLER_3_1473 ();
 sg13g2_decap_4 FILLER_3_1480 ();
 sg13g2_fill_2 FILLER_3_1512 ();
 sg13g2_fill_1 FILLER_3_1542 ();
 sg13g2_fill_2 FILLER_3_1561 ();
 sg13g2_fill_1 FILLER_3_1563 ();
 sg13g2_decap_4 FILLER_3_1575 ();
 sg13g2_fill_2 FILLER_3_1579 ();
 sg13g2_fill_2 FILLER_3_1600 ();
 sg13g2_fill_1 FILLER_3_1602 ();
 sg13g2_fill_1 FILLER_3_1606 ();
 sg13g2_fill_2 FILLER_3_1627 ();
 sg13g2_decap_8 FILLER_3_1637 ();
 sg13g2_fill_1 FILLER_3_1644 ();
 sg13g2_decap_8 FILLER_3_1662 ();
 sg13g2_decap_8 FILLER_3_1669 ();
 sg13g2_fill_1 FILLER_3_1676 ();
 sg13g2_fill_2 FILLER_3_1714 ();
 sg13g2_fill_1 FILLER_3_1716 ();
 sg13g2_fill_2 FILLER_3_1724 ();
 sg13g2_decap_8 FILLER_3_1730 ();
 sg13g2_decap_8 FILLER_3_1737 ();
 sg13g2_fill_2 FILLER_3_1769 ();
 sg13g2_fill_2 FILLER_3_1788 ();
 sg13g2_decap_8 FILLER_3_1805 ();
 sg13g2_fill_1 FILLER_3_1812 ();
 sg13g2_fill_1 FILLER_3_1833 ();
 sg13g2_decap_4 FILLER_3_1839 ();
 sg13g2_fill_1 FILLER_3_1843 ();
 sg13g2_decap_8 FILLER_3_1878 ();
 sg13g2_fill_2 FILLER_3_1885 ();
 sg13g2_decap_8 FILLER_3_1891 ();
 sg13g2_decap_4 FILLER_3_1926 ();
 sg13g2_fill_2 FILLER_3_1930 ();
 sg13g2_fill_1 FILLER_3_1969 ();
 sg13g2_fill_1 FILLER_3_2018 ();
 sg13g2_fill_1 FILLER_3_2038 ();
 sg13g2_fill_2 FILLER_3_2052 ();
 sg13g2_decap_8 FILLER_3_2070 ();
 sg13g2_decap_8 FILLER_3_2077 ();
 sg13g2_decap_8 FILLER_3_2112 ();
 sg13g2_decap_8 FILLER_3_2119 ();
 sg13g2_decap_4 FILLER_3_2126 ();
 sg13g2_fill_2 FILLER_3_2140 ();
 sg13g2_fill_1 FILLER_3_2142 ();
 sg13g2_decap_8 FILLER_3_2155 ();
 sg13g2_decap_8 FILLER_3_2162 ();
 sg13g2_decap_4 FILLER_3_2169 ();
 sg13g2_fill_2 FILLER_3_2182 ();
 sg13g2_fill_1 FILLER_3_2184 ();
 sg13g2_fill_1 FILLER_3_2190 ();
 sg13g2_fill_2 FILLER_3_2201 ();
 sg13g2_decap_8 FILLER_3_2222 ();
 sg13g2_fill_1 FILLER_3_2229 ();
 sg13g2_decap_8 FILLER_3_2276 ();
 sg13g2_decap_4 FILLER_3_2283 ();
 sg13g2_fill_2 FILLER_3_2292 ();
 sg13g2_fill_1 FILLER_3_2299 ();
 sg13g2_decap_4 FILLER_3_2308 ();
 sg13g2_fill_1 FILLER_3_2312 ();
 sg13g2_fill_1 FILLER_3_2326 ();
 sg13g2_decap_4 FILLER_3_2344 ();
 sg13g2_decap_8 FILLER_3_2360 ();
 sg13g2_decap_4 FILLER_3_2367 ();
 sg13g2_fill_1 FILLER_3_2384 ();
 sg13g2_decap_4 FILLER_3_2397 ();
 sg13g2_fill_1 FILLER_3_2412 ();
 sg13g2_decap_4 FILLER_3_2429 ();
 sg13g2_fill_2 FILLER_3_2433 ();
 sg13g2_fill_1 FILLER_3_2456 ();
 sg13g2_fill_2 FILLER_3_2465 ();
 sg13g2_decap_8 FILLER_3_2471 ();
 sg13g2_fill_2 FILLER_3_2478 ();
 sg13g2_fill_2 FILLER_3_2494 ();
 sg13g2_fill_1 FILLER_3_2496 ();
 sg13g2_decap_8 FILLER_3_2502 ();
 sg13g2_fill_2 FILLER_3_2509 ();
 sg13g2_fill_1 FILLER_3_2511 ();
 sg13g2_decap_8 FILLER_3_2529 ();
 sg13g2_fill_2 FILLER_3_2567 ();
 sg13g2_fill_1 FILLER_3_2595 ();
 sg13g2_decap_4 FILLER_3_2618 ();
 sg13g2_fill_1 FILLER_3_2622 ();
 sg13g2_decap_4 FILLER_3_2632 ();
 sg13g2_fill_1 FILLER_3_2641 ();
 sg13g2_fill_1 FILLER_3_2652 ();
 sg13g2_decap_8 FILLER_3_2686 ();
 sg13g2_fill_2 FILLER_3_2707 ();
 sg13g2_fill_1 FILLER_3_2709 ();
 sg13g2_decap_8 FILLER_3_2715 ();
 sg13g2_decap_8 FILLER_3_2722 ();
 sg13g2_fill_2 FILLER_3_2729 ();
 sg13g2_decap_8 FILLER_3_2751 ();
 sg13g2_decap_8 FILLER_3_2758 ();
 sg13g2_fill_1 FILLER_3_2765 ();
 sg13g2_decap_8 FILLER_3_2771 ();
 sg13g2_decap_4 FILLER_3_2778 ();
 sg13g2_fill_2 FILLER_3_2782 ();
 sg13g2_fill_2 FILLER_3_2804 ();
 sg13g2_decap_8 FILLER_3_2837 ();
 sg13g2_decap_4 FILLER_3_2844 ();
 sg13g2_fill_2 FILLER_3_2848 ();
 sg13g2_fill_1 FILLER_3_2858 ();
 sg13g2_fill_1 FILLER_3_2868 ();
 sg13g2_decap_8 FILLER_3_2894 ();
 sg13g2_fill_1 FILLER_3_2901 ();
 sg13g2_decap_8 FILLER_3_2923 ();
 sg13g2_fill_2 FILLER_3_2930 ();
 sg13g2_fill_1 FILLER_3_2932 ();
 sg13g2_fill_2 FILLER_3_2946 ();
 sg13g2_decap_4 FILLER_3_2965 ();
 sg13g2_fill_2 FILLER_3_2969 ();
 sg13g2_fill_2 FILLER_3_2986 ();
 sg13g2_fill_1 FILLER_3_2988 ();
 sg13g2_decap_8 FILLER_3_3037 ();
 sg13g2_decap_4 FILLER_3_3044 ();
 sg13g2_fill_1 FILLER_3_3053 ();
 sg13g2_decap_4 FILLER_3_3063 ();
 sg13g2_fill_2 FILLER_3_3067 ();
 sg13g2_fill_2 FILLER_3_3089 ();
 sg13g2_decap_8 FILLER_3_3108 ();
 sg13g2_decap_8 FILLER_3_3115 ();
 sg13g2_fill_2 FILLER_3_3122 ();
 sg13g2_decap_4 FILLER_3_3190 ();
 sg13g2_fill_1 FILLER_3_3194 ();
 sg13g2_fill_2 FILLER_3_3207 ();
 sg13g2_fill_1 FILLER_3_3225 ();
 sg13g2_decap_8 FILLER_3_3230 ();
 sg13g2_decap_8 FILLER_3_3237 ();
 sg13g2_decap_8 FILLER_3_3244 ();
 sg13g2_decap_8 FILLER_3_3251 ();
 sg13g2_decap_8 FILLER_3_3258 ();
 sg13g2_decap_8 FILLER_3_3265 ();
 sg13g2_decap_8 FILLER_3_3272 ();
 sg13g2_decap_8 FILLER_3_3279 ();
 sg13g2_decap_8 FILLER_3_3286 ();
 sg13g2_decap_8 FILLER_3_3293 ();
 sg13g2_decap_4 FILLER_3_3300 ();
 sg13g2_fill_1 FILLER_3_3304 ();
 sg13g2_decap_4 FILLER_3_3309 ();
 sg13g2_fill_1 FILLER_3_3313 ();
 sg13g2_decap_8 FILLER_3_3318 ();
 sg13g2_fill_2 FILLER_3_3325 ();
 sg13g2_fill_1 FILLER_3_3327 ();
 sg13g2_decap_8 FILLER_3_3363 ();
 sg13g2_fill_2 FILLER_3_3370 ();
 sg13g2_fill_1 FILLER_3_3372 ();
 sg13g2_decap_8 FILLER_3_3429 ();
 sg13g2_decap_8 FILLER_3_3436 ();
 sg13g2_decap_8 FILLER_3_3443 ();
 sg13g2_decap_8 FILLER_3_3450 ();
 sg13g2_decap_8 FILLER_3_3457 ();
 sg13g2_decap_8 FILLER_3_3464 ();
 sg13g2_decap_8 FILLER_3_3471 ();
 sg13g2_decap_8 FILLER_3_3478 ();
 sg13g2_decap_8 FILLER_3_3485 ();
 sg13g2_decap_8 FILLER_3_3492 ();
 sg13g2_decap_8 FILLER_3_3499 ();
 sg13g2_decap_8 FILLER_3_3506 ();
 sg13g2_decap_8 FILLER_3_3513 ();
 sg13g2_decap_8 FILLER_3_3520 ();
 sg13g2_decap_8 FILLER_3_3527 ();
 sg13g2_decap_8 FILLER_3_3534 ();
 sg13g2_decap_8 FILLER_3_3541 ();
 sg13g2_decap_8 FILLER_3_3548 ();
 sg13g2_decap_8 FILLER_3_3555 ();
 sg13g2_decap_8 FILLER_3_3562 ();
 sg13g2_decap_8 FILLER_3_3569 ();
 sg13g2_decap_4 FILLER_3_3576 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_fill_2 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_163 ();
 sg13g2_fill_2 FILLER_4_174 ();
 sg13g2_decap_8 FILLER_4_190 ();
 sg13g2_fill_2 FILLER_4_197 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_218 ();
 sg13g2_fill_2 FILLER_4_225 ();
 sg13g2_fill_1 FILLER_4_227 ();
 sg13g2_fill_2 FILLER_4_241 ();
 sg13g2_fill_1 FILLER_4_243 ();
 sg13g2_fill_2 FILLER_4_265 ();
 sg13g2_fill_1 FILLER_4_267 ();
 sg13g2_fill_2 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_4 FILLER_4_333 ();
 sg13g2_fill_2 FILLER_4_337 ();
 sg13g2_decap_4 FILLER_4_344 ();
 sg13g2_fill_2 FILLER_4_348 ();
 sg13g2_fill_2 FILLER_4_368 ();
 sg13g2_fill_1 FILLER_4_370 ();
 sg13g2_decap_4 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_decap_8 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_4_415 ();
 sg13g2_decap_4 FILLER_4_422 ();
 sg13g2_fill_1 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_4_440 ();
 sg13g2_decap_8 FILLER_4_447 ();
 sg13g2_decap_8 FILLER_4_454 ();
 sg13g2_decap_8 FILLER_4_461 ();
 sg13g2_decap_8 FILLER_4_468 ();
 sg13g2_decap_8 FILLER_4_475 ();
 sg13g2_decap_8 FILLER_4_482 ();
 sg13g2_decap_8 FILLER_4_489 ();
 sg13g2_fill_2 FILLER_4_496 ();
 sg13g2_fill_2 FILLER_4_511 ();
 sg13g2_fill_1 FILLER_4_513 ();
 sg13g2_decap_8 FILLER_4_536 ();
 sg13g2_decap_8 FILLER_4_548 ();
 sg13g2_fill_1 FILLER_4_555 ();
 sg13g2_fill_2 FILLER_4_574 ();
 sg13g2_fill_1 FILLER_4_576 ();
 sg13g2_decap_8 FILLER_4_594 ();
 sg13g2_fill_2 FILLER_4_618 ();
 sg13g2_fill_1 FILLER_4_633 ();
 sg13g2_decap_8 FILLER_4_678 ();
 sg13g2_decap_8 FILLER_4_685 ();
 sg13g2_fill_2 FILLER_4_692 ();
 sg13g2_decap_8 FILLER_4_704 ();
 sg13g2_fill_1 FILLER_4_711 ();
 sg13g2_decap_4 FILLER_4_722 ();
 sg13g2_fill_2 FILLER_4_726 ();
 sg13g2_decap_4 FILLER_4_756 ();
 sg13g2_fill_1 FILLER_4_773 ();
 sg13g2_fill_1 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_829 ();
 sg13g2_fill_2 FILLER_4_836 ();
 sg13g2_fill_2 FILLER_4_866 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_fill_2 FILLER_4_882 ();
 sg13g2_fill_1 FILLER_4_884 ();
 sg13g2_decap_8 FILLER_4_900 ();
 sg13g2_fill_1 FILLER_4_907 ();
 sg13g2_decap_4 FILLER_4_918 ();
 sg13g2_decap_8 FILLER_4_927 ();
 sg13g2_decap_8 FILLER_4_934 ();
 sg13g2_fill_1 FILLER_4_941 ();
 sg13g2_fill_2 FILLER_4_987 ();
 sg13g2_decap_4 FILLER_4_1002 ();
 sg13g2_fill_1 FILLER_4_1006 ();
 sg13g2_decap_4 FILLER_4_1013 ();
 sg13g2_fill_1 FILLER_4_1017 ();
 sg13g2_decap_4 FILLER_4_1029 ();
 sg13g2_fill_2 FILLER_4_1033 ();
 sg13g2_fill_2 FILLER_4_1050 ();
 sg13g2_fill_1 FILLER_4_1052 ();
 sg13g2_decap_8 FILLER_4_1057 ();
 sg13g2_decap_8 FILLER_4_1064 ();
 sg13g2_fill_2 FILLER_4_1071 ();
 sg13g2_fill_1 FILLER_4_1073 ();
 sg13g2_fill_2 FILLER_4_1090 ();
 sg13g2_decap_4 FILLER_4_1106 ();
 sg13g2_fill_2 FILLER_4_1110 ();
 sg13g2_decap_8 FILLER_4_1126 ();
 sg13g2_decap_8 FILLER_4_1133 ();
 sg13g2_decap_8 FILLER_4_1140 ();
 sg13g2_fill_1 FILLER_4_1163 ();
 sg13g2_fill_2 FILLER_4_1192 ();
 sg13g2_fill_1 FILLER_4_1194 ();
 sg13g2_decap_4 FILLER_4_1200 ();
 sg13g2_fill_2 FILLER_4_1213 ();
 sg13g2_fill_1 FILLER_4_1215 ();
 sg13g2_fill_1 FILLER_4_1235 ();
 sg13g2_fill_2 FILLER_4_1245 ();
 sg13g2_decap_8 FILLER_4_1251 ();
 sg13g2_fill_2 FILLER_4_1266 ();
 sg13g2_fill_1 FILLER_4_1268 ();
 sg13g2_decap_8 FILLER_4_1297 ();
 sg13g2_decap_4 FILLER_4_1304 ();
 sg13g2_fill_2 FILLER_4_1321 ();
 sg13g2_fill_1 FILLER_4_1323 ();
 sg13g2_decap_8 FILLER_4_1342 ();
 sg13g2_fill_2 FILLER_4_1349 ();
 sg13g2_fill_2 FILLER_4_1369 ();
 sg13g2_decap_4 FILLER_4_1403 ();
 sg13g2_fill_1 FILLER_4_1407 ();
 sg13g2_decap_8 FILLER_4_1420 ();
 sg13g2_decap_4 FILLER_4_1427 ();
 sg13g2_decap_8 FILLER_4_1440 ();
 sg13g2_fill_1 FILLER_4_1447 ();
 sg13g2_fill_2 FILLER_4_1460 ();
 sg13g2_decap_8 FILLER_4_1474 ();
 sg13g2_decap_4 FILLER_4_1481 ();
 sg13g2_decap_8 FILLER_4_1493 ();
 sg13g2_decap_8 FILLER_4_1500 ();
 sg13g2_decap_8 FILLER_4_1507 ();
 sg13g2_fill_1 FILLER_4_1514 ();
 sg13g2_decap_8 FILLER_4_1519 ();
 sg13g2_decap_8 FILLER_4_1526 ();
 sg13g2_fill_1 FILLER_4_1570 ();
 sg13g2_decap_8 FILLER_4_1594 ();
 sg13g2_decap_4 FILLER_4_1601 ();
 sg13g2_fill_1 FILLER_4_1605 ();
 sg13g2_fill_2 FILLER_4_1619 ();
 sg13g2_fill_1 FILLER_4_1621 ();
 sg13g2_decap_4 FILLER_4_1666 ();
 sg13g2_fill_2 FILLER_4_1670 ();
 sg13g2_decap_8 FILLER_4_1689 ();
 sg13g2_decap_4 FILLER_4_1713 ();
 sg13g2_fill_2 FILLER_4_1728 ();
 sg13g2_fill_1 FILLER_4_1730 ();
 sg13g2_decap_8 FILLER_4_1739 ();
 sg13g2_fill_1 FILLER_4_1746 ();
 sg13g2_decap_8 FILLER_4_1770 ();
 sg13g2_decap_8 FILLER_4_1796 ();
 sg13g2_decap_8 FILLER_4_1803 ();
 sg13g2_fill_1 FILLER_4_1829 ();
 sg13g2_fill_2 FILLER_4_1855 ();
 sg13g2_fill_1 FILLER_4_1857 ();
 sg13g2_decap_4 FILLER_4_1893 ();
 sg13g2_fill_2 FILLER_4_1897 ();
 sg13g2_decap_8 FILLER_4_1912 ();
 sg13g2_decap_4 FILLER_4_1919 ();
 sg13g2_decap_4 FILLER_4_1930 ();
 sg13g2_fill_1 FILLER_4_1934 ();
 sg13g2_fill_2 FILLER_4_1951 ();
 sg13g2_fill_1 FILLER_4_1953 ();
 sg13g2_fill_2 FILLER_4_1969 ();
 sg13g2_decap_4 FILLER_4_1986 ();
 sg13g2_fill_2 FILLER_4_1995 ();
 sg13g2_decap_4 FILLER_4_2005 ();
 sg13g2_fill_1 FILLER_4_2009 ();
 sg13g2_fill_1 FILLER_4_2019 ();
 sg13g2_decap_8 FILLER_4_2036 ();
 sg13g2_fill_2 FILLER_4_2051 ();
 sg13g2_fill_1 FILLER_4_2053 ();
 sg13g2_fill_1 FILLER_4_2064 ();
 sg13g2_fill_2 FILLER_4_2071 ();
 sg13g2_fill_1 FILLER_4_2073 ();
 sg13g2_decap_8 FILLER_4_2095 ();
 sg13g2_decap_4 FILLER_4_2102 ();
 sg13g2_fill_1 FILLER_4_2106 ();
 sg13g2_decap_8 FILLER_4_2111 ();
 sg13g2_decap_8 FILLER_4_2118 ();
 sg13g2_fill_2 FILLER_4_2125 ();
 sg13g2_fill_1 FILLER_4_2127 ();
 sg13g2_fill_1 FILLER_4_2133 ();
 sg13g2_decap_8 FILLER_4_2154 ();
 sg13g2_decap_4 FILLER_4_2176 ();
 sg13g2_fill_2 FILLER_4_2180 ();
 sg13g2_decap_8 FILLER_4_2196 ();
 sg13g2_decap_8 FILLER_4_2203 ();
 sg13g2_fill_1 FILLER_4_2210 ();
 sg13g2_fill_1 FILLER_4_2216 ();
 sg13g2_decap_8 FILLER_4_2234 ();
 sg13g2_fill_2 FILLER_4_2241 ();
 sg13g2_decap_4 FILLER_4_2261 ();
 sg13g2_fill_2 FILLER_4_2265 ();
 sg13g2_fill_2 FILLER_4_2289 ();
 sg13g2_decap_8 FILLER_4_2304 ();
 sg13g2_decap_8 FILLER_4_2311 ();
 sg13g2_decap_4 FILLER_4_2322 ();
 sg13g2_decap_8 FILLER_4_2340 ();
 sg13g2_decap_8 FILLER_4_2347 ();
 sg13g2_fill_2 FILLER_4_2354 ();
 sg13g2_fill_1 FILLER_4_2356 ();
 sg13g2_decap_8 FILLER_4_2362 ();
 sg13g2_decap_8 FILLER_4_2369 ();
 sg13g2_decap_4 FILLER_4_2376 ();
 sg13g2_fill_1 FILLER_4_2384 ();
 sg13g2_decap_4 FILLER_4_2389 ();
 sg13g2_fill_1 FILLER_4_2393 ();
 sg13g2_decap_8 FILLER_4_2399 ();
 sg13g2_fill_2 FILLER_4_2406 ();
 sg13g2_fill_1 FILLER_4_2408 ();
 sg13g2_decap_8 FILLER_4_2423 ();
 sg13g2_decap_4 FILLER_4_2430 ();
 sg13g2_fill_1 FILLER_4_2434 ();
 sg13g2_fill_2 FILLER_4_2458 ();
 sg13g2_fill_1 FILLER_4_2460 ();
 sg13g2_decap_8 FILLER_4_2509 ();
 sg13g2_decap_4 FILLER_4_2516 ();
 sg13g2_fill_1 FILLER_4_2520 ();
 sg13g2_decap_8 FILLER_4_2538 ();
 sg13g2_fill_2 FILLER_4_2550 ();
 sg13g2_decap_4 FILLER_4_2556 ();
 sg13g2_fill_1 FILLER_4_2560 ();
 sg13g2_decap_8 FILLER_4_2587 ();
 sg13g2_decap_8 FILLER_4_2594 ();
 sg13g2_fill_2 FILLER_4_2606 ();
 sg13g2_decap_8 FILLER_4_2613 ();
 sg13g2_fill_2 FILLER_4_2620 ();
 sg13g2_fill_1 FILLER_4_2622 ();
 sg13g2_fill_1 FILLER_4_2633 ();
 sg13g2_decap_8 FILLER_4_2639 ();
 sg13g2_decap_8 FILLER_4_2646 ();
 sg13g2_fill_1 FILLER_4_2653 ();
 sg13g2_fill_2 FILLER_4_2664 ();
 sg13g2_fill_1 FILLER_4_2666 ();
 sg13g2_decap_8 FILLER_4_2672 ();
 sg13g2_decap_8 FILLER_4_2679 ();
 sg13g2_fill_2 FILLER_4_2686 ();
 sg13g2_decap_8 FILLER_4_2693 ();
 sg13g2_fill_1 FILLER_4_2700 ();
 sg13g2_decap_4 FILLER_4_2721 ();
 sg13g2_fill_1 FILLER_4_2725 ();
 sg13g2_decap_4 FILLER_4_2757 ();
 sg13g2_decap_8 FILLER_4_2806 ();
 sg13g2_decap_8 FILLER_4_2813 ();
 sg13g2_fill_1 FILLER_4_2820 ();
 sg13g2_decap_8 FILLER_4_2839 ();
 sg13g2_fill_1 FILLER_4_2846 ();
 sg13g2_decap_4 FILLER_4_2867 ();
 sg13g2_fill_2 FILLER_4_2886 ();
 sg13g2_decap_8 FILLER_4_2896 ();
 sg13g2_fill_1 FILLER_4_2903 ();
 sg13g2_decap_4 FILLER_4_2917 ();
 sg13g2_fill_1 FILLER_4_2921 ();
 sg13g2_decap_8 FILLER_4_2927 ();
 sg13g2_decap_8 FILLER_4_2934 ();
 sg13g2_fill_2 FILLER_4_2941 ();
 sg13g2_fill_1 FILLER_4_2943 ();
 sg13g2_fill_2 FILLER_4_2972 ();
 sg13g2_fill_1 FILLER_4_2974 ();
 sg13g2_decap_4 FILLER_4_2979 ();
 sg13g2_fill_2 FILLER_4_2992 ();
 sg13g2_fill_1 FILLER_4_2994 ();
 sg13g2_fill_2 FILLER_4_2999 ();
 sg13g2_decap_8 FILLER_4_3006 ();
 sg13g2_decap_8 FILLER_4_3013 ();
 sg13g2_decap_4 FILLER_4_3020 ();
 sg13g2_fill_2 FILLER_4_3024 ();
 sg13g2_fill_2 FILLER_4_3049 ();
 sg13g2_fill_2 FILLER_4_3064 ();
 sg13g2_fill_1 FILLER_4_3066 ();
 sg13g2_fill_1 FILLER_4_3072 ();
 sg13g2_decap_8 FILLER_4_3085 ();
 sg13g2_decap_8 FILLER_4_3092 ();
 sg13g2_decap_8 FILLER_4_3099 ();
 sg13g2_fill_2 FILLER_4_3106 ();
 sg13g2_fill_1 FILLER_4_3108 ();
 sg13g2_decap_4 FILLER_4_3129 ();
 sg13g2_fill_2 FILLER_4_3133 ();
 sg13g2_decap_8 FILLER_4_3150 ();
 sg13g2_decap_4 FILLER_4_3157 ();
 sg13g2_fill_1 FILLER_4_3161 ();
 sg13g2_decap_8 FILLER_4_3172 ();
 sg13g2_decap_8 FILLER_4_3179 ();
 sg13g2_fill_1 FILLER_4_3186 ();
 sg13g2_decap_8 FILLER_4_3191 ();
 sg13g2_decap_4 FILLER_4_3198 ();
 sg13g2_fill_1 FILLER_4_3212 ();
 sg13g2_decap_4 FILLER_4_3217 ();
 sg13g2_decap_8 FILLER_4_3247 ();
 sg13g2_decap_8 FILLER_4_3254 ();
 sg13g2_decap_8 FILLER_4_3261 ();
 sg13g2_decap_8 FILLER_4_3268 ();
 sg13g2_decap_8 FILLER_4_3275 ();
 sg13g2_decap_8 FILLER_4_3282 ();
 sg13g2_decap_8 FILLER_4_3289 ();
 sg13g2_decap_8 FILLER_4_3296 ();
 sg13g2_decap_8 FILLER_4_3303 ();
 sg13g2_decap_8 FILLER_4_3310 ();
 sg13g2_decap_8 FILLER_4_3317 ();
 sg13g2_fill_1 FILLER_4_3324 ();
 sg13g2_fill_2 FILLER_4_3342 ();
 sg13g2_decap_8 FILLER_4_3349 ();
 sg13g2_decap_4 FILLER_4_3361 ();
 sg13g2_fill_2 FILLER_4_3365 ();
 sg13g2_decap_8 FILLER_4_3388 ();
 sg13g2_fill_2 FILLER_4_3395 ();
 sg13g2_decap_8 FILLER_4_3408 ();
 sg13g2_decap_8 FILLER_4_3415 ();
 sg13g2_decap_8 FILLER_4_3422 ();
 sg13g2_decap_8 FILLER_4_3429 ();
 sg13g2_decap_8 FILLER_4_3436 ();
 sg13g2_decap_8 FILLER_4_3443 ();
 sg13g2_decap_8 FILLER_4_3450 ();
 sg13g2_fill_2 FILLER_4_3457 ();
 sg13g2_fill_1 FILLER_4_3459 ();
 sg13g2_decap_8 FILLER_4_3464 ();
 sg13g2_decap_8 FILLER_4_3471 ();
 sg13g2_decap_8 FILLER_4_3478 ();
 sg13g2_decap_8 FILLER_4_3485 ();
 sg13g2_decap_8 FILLER_4_3492 ();
 sg13g2_decap_8 FILLER_4_3499 ();
 sg13g2_decap_8 FILLER_4_3506 ();
 sg13g2_decap_8 FILLER_4_3513 ();
 sg13g2_decap_8 FILLER_4_3520 ();
 sg13g2_decap_8 FILLER_4_3527 ();
 sg13g2_decap_8 FILLER_4_3534 ();
 sg13g2_decap_8 FILLER_4_3541 ();
 sg13g2_decap_8 FILLER_4_3548 ();
 sg13g2_decap_8 FILLER_4_3555 ();
 sg13g2_decap_8 FILLER_4_3562 ();
 sg13g2_decap_8 FILLER_4_3569 ();
 sg13g2_decap_4 FILLER_4_3576 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_2 FILLER_5_130 ();
 sg13g2_decap_4 FILLER_5_135 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_fill_2 FILLER_5_156 ();
 sg13g2_fill_1 FILLER_5_158 ();
 sg13g2_fill_2 FILLER_5_164 ();
 sg13g2_fill_1 FILLER_5_166 ();
 sg13g2_decap_8 FILLER_5_192 ();
 sg13g2_decap_8 FILLER_5_199 ();
 sg13g2_fill_1 FILLER_5_206 ();
 sg13g2_decap_4 FILLER_5_220 ();
 sg13g2_fill_1 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_decap_4 FILLER_5_268 ();
 sg13g2_fill_1 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_289 ();
 sg13g2_decap_4 FILLER_5_296 ();
 sg13g2_fill_2 FILLER_5_300 ();
 sg13g2_fill_1 FILLER_5_306 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_4 FILLER_5_326 ();
 sg13g2_fill_2 FILLER_5_330 ();
 sg13g2_fill_2 FILLER_5_339 ();
 sg13g2_fill_1 FILLER_5_341 ();
 sg13g2_fill_2 FILLER_5_347 ();
 sg13g2_fill_1 FILLER_5_349 ();
 sg13g2_fill_2 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_decap_4 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_440 ();
 sg13g2_decap_8 FILLER_5_460 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_508 ();
 sg13g2_decap_4 FILLER_5_515 ();
 sg13g2_fill_2 FILLER_5_519 ();
 sg13g2_fill_1 FILLER_5_528 ();
 sg13g2_decap_4 FILLER_5_542 ();
 sg13g2_fill_1 FILLER_5_562 ();
 sg13g2_decap_8 FILLER_5_572 ();
 sg13g2_fill_2 FILLER_5_579 ();
 sg13g2_fill_1 FILLER_5_581 ();
 sg13g2_decap_4 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_617 ();
 sg13g2_fill_2 FILLER_5_637 ();
 sg13g2_fill_1 FILLER_5_639 ();
 sg13g2_fill_1 FILLER_5_653 ();
 sg13g2_decap_8 FILLER_5_659 ();
 sg13g2_decap_8 FILLER_5_666 ();
 sg13g2_decap_4 FILLER_5_673 ();
 sg13g2_decap_8 FILLER_5_694 ();
 sg13g2_decap_4 FILLER_5_701 ();
 sg13g2_fill_2 FILLER_5_719 ();
 sg13g2_fill_2 FILLER_5_738 ();
 sg13g2_fill_1 FILLER_5_740 ();
 sg13g2_decap_8 FILLER_5_745 ();
 sg13g2_decap_8 FILLER_5_752 ();
 sg13g2_decap_4 FILLER_5_782 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_fill_1 FILLER_5_809 ();
 sg13g2_decap_4 FILLER_5_867 ();
 sg13g2_fill_2 FILLER_5_871 ();
 sg13g2_decap_4 FILLER_5_905 ();
 sg13g2_fill_2 FILLER_5_944 ();
 sg13g2_fill_1 FILLER_5_946 ();
 sg13g2_decap_8 FILLER_5_951 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_decap_4 FILLER_5_965 ();
 sg13g2_fill_2 FILLER_5_969 ();
 sg13g2_decap_4 FILLER_5_976 ();
 sg13g2_fill_2 FILLER_5_980 ();
 sg13g2_fill_2 FILLER_5_1004 ();
 sg13g2_fill_1 FILLER_5_1006 ();
 sg13g2_fill_2 FILLER_5_1011 ();
 sg13g2_fill_1 FILLER_5_1013 ();
 sg13g2_fill_2 FILLER_5_1019 ();
 sg13g2_decap_8 FILLER_5_1025 ();
 sg13g2_decap_4 FILLER_5_1032 ();
 sg13g2_fill_1 FILLER_5_1036 ();
 sg13g2_fill_2 FILLER_5_1046 ();
 sg13g2_decap_4 FILLER_5_1076 ();
 sg13g2_decap_8 FILLER_5_1109 ();
 sg13g2_fill_1 FILLER_5_1116 ();
 sg13g2_decap_8 FILLER_5_1127 ();
 sg13g2_decap_8 FILLER_5_1146 ();
 sg13g2_fill_1 FILLER_5_1153 ();
 sg13g2_decap_4 FILLER_5_1164 ();
 sg13g2_fill_1 FILLER_5_1168 ();
 sg13g2_decap_8 FILLER_5_1173 ();
 sg13g2_decap_4 FILLER_5_1180 ();
 sg13g2_fill_1 FILLER_5_1184 ();
 sg13g2_fill_2 FILLER_5_1203 ();
 sg13g2_decap_8 FILLER_5_1215 ();
 sg13g2_fill_2 FILLER_5_1222 ();
 sg13g2_fill_1 FILLER_5_1224 ();
 sg13g2_decap_8 FILLER_5_1230 ();
 sg13g2_fill_1 FILLER_5_1237 ();
 sg13g2_decap_8 FILLER_5_1242 ();
 sg13g2_fill_2 FILLER_5_1249 ();
 sg13g2_fill_1 FILLER_5_1251 ();
 sg13g2_decap_8 FILLER_5_1269 ();
 sg13g2_decap_4 FILLER_5_1276 ();
 sg13g2_fill_1 FILLER_5_1280 ();
 sg13g2_fill_1 FILLER_5_1312 ();
 sg13g2_fill_2 FILLER_5_1319 ();
 sg13g2_fill_1 FILLER_5_1326 ();
 sg13g2_fill_2 FILLER_5_1331 ();
 sg13g2_fill_2 FILLER_5_1337 ();
 sg13g2_fill_2 FILLER_5_1376 ();
 sg13g2_fill_2 FILLER_5_1394 ();
 sg13g2_fill_1 FILLER_5_1396 ();
 sg13g2_fill_1 FILLER_5_1410 ();
 sg13g2_decap_4 FILLER_5_1442 ();
 sg13g2_fill_2 FILLER_5_1460 ();
 sg13g2_fill_2 FILLER_5_1508 ();
 sg13g2_fill_2 FILLER_5_1545 ();
 sg13g2_decap_4 FILLER_5_1552 ();
 sg13g2_fill_1 FILLER_5_1556 ();
 sg13g2_fill_1 FILLER_5_1565 ();
 sg13g2_fill_2 FILLER_5_1577 ();
 sg13g2_fill_1 FILLER_5_1579 ();
 sg13g2_fill_1 FILLER_5_1588 ();
 sg13g2_decap_8 FILLER_5_1593 ();
 sg13g2_decap_8 FILLER_5_1600 ();
 sg13g2_decap_8 FILLER_5_1607 ();
 sg13g2_decap_4 FILLER_5_1614 ();
 sg13g2_fill_2 FILLER_5_1618 ();
 sg13g2_decap_8 FILLER_5_1623 ();
 sg13g2_decap_8 FILLER_5_1634 ();
 sg13g2_decap_8 FILLER_5_1641 ();
 sg13g2_decap_4 FILLER_5_1659 ();
 sg13g2_fill_1 FILLER_5_1663 ();
 sg13g2_decap_4 FILLER_5_1669 ();
 sg13g2_fill_2 FILLER_5_1673 ();
 sg13g2_decap_8 FILLER_5_1690 ();
 sg13g2_decap_8 FILLER_5_1697 ();
 sg13g2_decap_8 FILLER_5_1704 ();
 sg13g2_decap_8 FILLER_5_1711 ();
 sg13g2_decap_4 FILLER_5_1718 ();
 sg13g2_fill_1 FILLER_5_1722 ();
 sg13g2_decap_4 FILLER_5_1741 ();
 sg13g2_fill_1 FILLER_5_1745 ();
 sg13g2_fill_2 FILLER_5_1760 ();
 sg13g2_decap_8 FILLER_5_1773 ();
 sg13g2_decap_8 FILLER_5_1780 ();
 sg13g2_decap_8 FILLER_5_1800 ();
 sg13g2_decap_4 FILLER_5_1830 ();
 sg13g2_fill_2 FILLER_5_1879 ();
 sg13g2_fill_2 FILLER_5_1929 ();
 sg13g2_fill_1 FILLER_5_1931 ();
 sg13g2_fill_1 FILLER_5_1942 ();
 sg13g2_fill_1 FILLER_5_1959 ();
 sg13g2_fill_2 FILLER_5_1966 ();
 sg13g2_fill_1 FILLER_5_1973 ();
 sg13g2_decap_8 FILLER_5_1979 ();
 sg13g2_decap_4 FILLER_5_1986 ();
 sg13g2_fill_1 FILLER_5_1990 ();
 sg13g2_fill_2 FILLER_5_1996 ();
 sg13g2_decap_4 FILLER_5_2008 ();
 sg13g2_decap_8 FILLER_5_2041 ();
 sg13g2_fill_2 FILLER_5_2048 ();
 sg13g2_fill_1 FILLER_5_2050 ();
 sg13g2_decap_4 FILLER_5_2089 ();
 sg13g2_fill_1 FILLER_5_2093 ();
 sg13g2_decap_4 FILLER_5_2097 ();
 sg13g2_fill_1 FILLER_5_2101 ();
 sg13g2_decap_8 FILLER_5_2130 ();
 sg13g2_decap_8 FILLER_5_2137 ();
 sg13g2_fill_2 FILLER_5_2144 ();
 sg13g2_fill_2 FILLER_5_2159 ();
 sg13g2_fill_1 FILLER_5_2161 ();
 sg13g2_decap_4 FILLER_5_2175 ();
 sg13g2_decap_4 FILLER_5_2204 ();
 sg13g2_fill_2 FILLER_5_2208 ();
 sg13g2_decap_4 FILLER_5_2237 ();
 sg13g2_fill_2 FILLER_5_2241 ();
 sg13g2_decap_8 FILLER_5_2283 ();
 sg13g2_decap_8 FILLER_5_2297 ();
 sg13g2_fill_2 FILLER_5_2304 ();
 sg13g2_decap_4 FILLER_5_2341 ();
 sg13g2_fill_2 FILLER_5_2345 ();
 sg13g2_decap_8 FILLER_5_2384 ();
 sg13g2_decap_4 FILLER_5_2391 ();
 sg13g2_fill_1 FILLER_5_2395 ();
 sg13g2_fill_2 FILLER_5_2400 ();
 sg13g2_fill_2 FILLER_5_2451 ();
 sg13g2_fill_1 FILLER_5_2466 ();
 sg13g2_fill_1 FILLER_5_2471 ();
 sg13g2_decap_8 FILLER_5_2476 ();
 sg13g2_decap_8 FILLER_5_2483 ();
 sg13g2_decap_8 FILLER_5_2506 ();
 sg13g2_fill_2 FILLER_5_2513 ();
 sg13g2_fill_1 FILLER_5_2515 ();
 sg13g2_decap_4 FILLER_5_2539 ();
 sg13g2_fill_2 FILLER_5_2543 ();
 sg13g2_fill_1 FILLER_5_2580 ();
 sg13g2_decap_8 FILLER_5_2589 ();
 sg13g2_fill_2 FILLER_5_2596 ();
 sg13g2_decap_8 FILLER_5_2605 ();
 sg13g2_fill_2 FILLER_5_2612 ();
 sg13g2_fill_1 FILLER_5_2614 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_4 FILLER_5_2653 ();
 sg13g2_fill_1 FILLER_5_2657 ();
 sg13g2_decap_8 FILLER_5_2662 ();
 sg13g2_decap_8 FILLER_5_2669 ();
 sg13g2_decap_8 FILLER_5_2676 ();
 sg13g2_fill_1 FILLER_5_2683 ();
 sg13g2_decap_4 FILLER_5_2702 ();
 sg13g2_fill_2 FILLER_5_2706 ();
 sg13g2_decap_8 FILLER_5_2725 ();
 sg13g2_fill_2 FILLER_5_2732 ();
 sg13g2_fill_1 FILLER_5_2738 ();
 sg13g2_fill_1 FILLER_5_2744 ();
 sg13g2_decap_8 FILLER_5_2751 ();
 sg13g2_fill_1 FILLER_5_2758 ();
 sg13g2_fill_2 FILLER_5_2764 ();
 sg13g2_fill_1 FILLER_5_2766 ();
 sg13g2_fill_2 FILLER_5_2780 ();
 sg13g2_fill_1 FILLER_5_2782 ();
 sg13g2_decap_4 FILLER_5_2792 ();
 sg13g2_fill_1 FILLER_5_2796 ();
 sg13g2_decap_4 FILLER_5_2808 ();
 sg13g2_fill_1 FILLER_5_2812 ();
 sg13g2_fill_2 FILLER_5_2826 ();
 sg13g2_fill_1 FILLER_5_2828 ();
 sg13g2_fill_2 FILLER_5_2847 ();
 sg13g2_fill_2 FILLER_5_2870 ();
 sg13g2_fill_1 FILLER_5_2882 ();
 sg13g2_decap_4 FILLER_5_2944 ();
 sg13g2_fill_1 FILLER_5_2948 ();
 sg13g2_decap_8 FILLER_5_2953 ();
 sg13g2_decap_8 FILLER_5_2960 ();
 sg13g2_decap_8 FILLER_5_2978 ();
 sg13g2_fill_1 FILLER_5_2985 ();
 sg13g2_decap_8 FILLER_5_3012 ();
 sg13g2_fill_2 FILLER_5_3055 ();
 sg13g2_fill_1 FILLER_5_3057 ();
 sg13g2_decap_8 FILLER_5_3081 ();
 sg13g2_fill_1 FILLER_5_3088 ();
 sg13g2_fill_1 FILLER_5_3097 ();
 sg13g2_decap_8 FILLER_5_3124 ();
 sg13g2_fill_1 FILLER_5_3131 ();
 sg13g2_decap_4 FILLER_5_3152 ();
 sg13g2_fill_1 FILLER_5_3156 ();
 sg13g2_decap_8 FILLER_5_3162 ();
 sg13g2_fill_2 FILLER_5_3169 ();
 sg13g2_fill_1 FILLER_5_3200 ();
 sg13g2_fill_1 FILLER_5_3262 ();
 sg13g2_decap_4 FILLER_5_3276 ();
 sg13g2_fill_2 FILLER_5_3298 ();
 sg13g2_decap_8 FILLER_5_3308 ();
 sg13g2_fill_2 FILLER_5_3315 ();
 sg13g2_fill_1 FILLER_5_3330 ();
 sg13g2_fill_1 FILLER_5_3336 ();
 sg13g2_fill_1 FILLER_5_3351 ();
 sg13g2_decap_8 FILLER_5_3359 ();
 sg13g2_decap_4 FILLER_5_3366 ();
 sg13g2_fill_2 FILLER_5_3370 ();
 sg13g2_decap_8 FILLER_5_3377 ();
 sg13g2_decap_8 FILLER_5_3384 ();
 sg13g2_fill_2 FILLER_5_3391 ();
 sg13g2_decap_8 FILLER_5_3415 ();
 sg13g2_fill_2 FILLER_5_3422 ();
 sg13g2_fill_1 FILLER_5_3424 ();
 sg13g2_decap_8 FILLER_5_3443 ();
 sg13g2_decap_4 FILLER_5_3450 ();
 sg13g2_fill_2 FILLER_5_3462 ();
 sg13g2_decap_8 FILLER_5_3472 ();
 sg13g2_decap_8 FILLER_5_3479 ();
 sg13g2_decap_8 FILLER_5_3486 ();
 sg13g2_decap_8 FILLER_5_3493 ();
 sg13g2_decap_8 FILLER_5_3500 ();
 sg13g2_decap_8 FILLER_5_3507 ();
 sg13g2_decap_8 FILLER_5_3514 ();
 sg13g2_decap_8 FILLER_5_3521 ();
 sg13g2_decap_8 FILLER_5_3528 ();
 sg13g2_decap_8 FILLER_5_3535 ();
 sg13g2_decap_8 FILLER_5_3542 ();
 sg13g2_decap_8 FILLER_5_3549 ();
 sg13g2_decap_8 FILLER_5_3556 ();
 sg13g2_decap_8 FILLER_5_3563 ();
 sg13g2_decap_8 FILLER_5_3570 ();
 sg13g2_fill_2 FILLER_5_3577 ();
 sg13g2_fill_1 FILLER_5_3579 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_126 ();
 sg13g2_decap_4 FILLER_6_156 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_fill_1 FILLER_6_172 ();
 sg13g2_fill_2 FILLER_6_181 ();
 sg13g2_fill_1 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_190 ();
 sg13g2_decap_4 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_226 ();
 sg13g2_decap_8 FILLER_6_244 ();
 sg13g2_decap_8 FILLER_6_251 ();
 sg13g2_fill_2 FILLER_6_275 ();
 sg13g2_fill_1 FILLER_6_277 ();
 sg13g2_decap_4 FILLER_6_290 ();
 sg13g2_fill_2 FILLER_6_323 ();
 sg13g2_fill_1 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_fill_1 FILLER_6_372 ();
 sg13g2_decap_4 FILLER_6_378 ();
 sg13g2_fill_2 FILLER_6_382 ();
 sg13g2_fill_1 FILLER_6_396 ();
 sg13g2_fill_1 FILLER_6_401 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_1 FILLER_6_427 ();
 sg13g2_fill_2 FILLER_6_443 ();
 sg13g2_decap_8 FILLER_6_463 ();
 sg13g2_fill_1 FILLER_6_526 ();
 sg13g2_fill_2 FILLER_6_535 ();
 sg13g2_fill_2 FILLER_6_548 ();
 sg13g2_decap_8 FILLER_6_570 ();
 sg13g2_fill_1 FILLER_6_577 ();
 sg13g2_decap_8 FILLER_6_582 ();
 sg13g2_decap_8 FILLER_6_589 ();
 sg13g2_fill_2 FILLER_6_607 ();
 sg13g2_decap_4 FILLER_6_622 ();
 sg13g2_fill_2 FILLER_6_626 ();
 sg13g2_decap_4 FILLER_6_645 ();
 sg13g2_fill_1 FILLER_6_649 ();
 sg13g2_fill_1 FILLER_6_665 ();
 sg13g2_fill_2 FILLER_6_682 ();
 sg13g2_fill_1 FILLER_6_684 ();
 sg13g2_decap_4 FILLER_6_693 ();
 sg13g2_fill_2 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_724 ();
 sg13g2_decap_4 FILLER_6_731 ();
 sg13g2_fill_1 FILLER_6_735 ();
 sg13g2_fill_2 FILLER_6_749 ();
 sg13g2_fill_2 FILLER_6_775 ();
 sg13g2_decap_4 FILLER_6_782 ();
 sg13g2_fill_2 FILLER_6_786 ();
 sg13g2_decap_4 FILLER_6_802 ();
 sg13g2_fill_1 FILLER_6_806 ();
 sg13g2_fill_2 FILLER_6_812 ();
 sg13g2_fill_2 FILLER_6_819 ();
 sg13g2_fill_1 FILLER_6_821 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_fill_1 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_849 ();
 sg13g2_decap_4 FILLER_6_856 ();
 sg13g2_fill_1 FILLER_6_860 ();
 sg13g2_decap_8 FILLER_6_873 ();
 sg13g2_decap_8 FILLER_6_880 ();
 sg13g2_decap_4 FILLER_6_887 ();
 sg13g2_fill_2 FILLER_6_903 ();
 sg13g2_fill_1 FILLER_6_905 ();
 sg13g2_fill_2 FILLER_6_931 ();
 sg13g2_fill_1 FILLER_6_933 ();
 sg13g2_decap_4 FILLER_6_946 ();
 sg13g2_fill_1 FILLER_6_950 ();
 sg13g2_fill_1 FILLER_6_959 ();
 sg13g2_decap_4 FILLER_6_981 ();
 sg13g2_fill_2 FILLER_6_1013 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_fill_2 FILLER_6_1038 ();
 sg13g2_fill_1 FILLER_6_1040 ();
 sg13g2_fill_2 FILLER_6_1070 ();
 sg13g2_decap_8 FILLER_6_1089 ();
 sg13g2_decap_4 FILLER_6_1124 ();
 sg13g2_fill_2 FILLER_6_1128 ();
 sg13g2_decap_4 FILLER_6_1155 ();
 sg13g2_fill_1 FILLER_6_1159 ();
 sg13g2_decap_8 FILLER_6_1178 ();
 sg13g2_fill_2 FILLER_6_1185 ();
 sg13g2_fill_1 FILLER_6_1187 ();
 sg13g2_fill_1 FILLER_6_1193 ();
 sg13g2_decap_8 FILLER_6_1203 ();
 sg13g2_decap_4 FILLER_6_1222 ();
 sg13g2_fill_2 FILLER_6_1226 ();
 sg13g2_fill_2 FILLER_6_1243 ();
 sg13g2_fill_1 FILLER_6_1245 ();
 sg13g2_fill_2 FILLER_6_1259 ();
 sg13g2_decap_4 FILLER_6_1279 ();
 sg13g2_fill_2 FILLER_6_1283 ();
 sg13g2_decap_8 FILLER_6_1294 ();
 sg13g2_decap_4 FILLER_6_1301 ();
 sg13g2_decap_8 FILLER_6_1328 ();
 sg13g2_fill_2 FILLER_6_1335 ();
 sg13g2_fill_1 FILLER_6_1337 ();
 sg13g2_decap_8 FILLER_6_1353 ();
 sg13g2_decap_8 FILLER_6_1360 ();
 sg13g2_fill_2 FILLER_6_1367 ();
 sg13g2_fill_2 FILLER_6_1382 ();
 sg13g2_fill_1 FILLER_6_1384 ();
 sg13g2_decap_4 FILLER_6_1406 ();
 sg13g2_decap_8 FILLER_6_1415 ();
 sg13g2_fill_2 FILLER_6_1422 ();
 sg13g2_fill_1 FILLER_6_1424 ();
 sg13g2_fill_1 FILLER_6_1430 ();
 sg13g2_fill_2 FILLER_6_1436 ();
 sg13g2_fill_1 FILLER_6_1438 ();
 sg13g2_fill_1 FILLER_6_1456 ();
 sg13g2_decap_8 FILLER_6_1462 ();
 sg13g2_fill_1 FILLER_6_1469 ();
 sg13g2_fill_2 FILLER_6_1487 ();
 sg13g2_fill_1 FILLER_6_1489 ();
 sg13g2_decap_8 FILLER_6_1493 ();
 sg13g2_decap_4 FILLER_6_1500 ();
 sg13g2_decap_8 FILLER_6_1508 ();
 sg13g2_decap_8 FILLER_6_1515 ();
 sg13g2_decap_8 FILLER_6_1522 ();
 sg13g2_decap_8 FILLER_6_1529 ();
 sg13g2_fill_2 FILLER_6_1536 ();
 sg13g2_fill_2 FILLER_6_1558 ();
 sg13g2_fill_2 FILLER_6_1587 ();
 sg13g2_fill_2 FILLER_6_1597 ();
 sg13g2_fill_1 FILLER_6_1599 ();
 sg13g2_fill_2 FILLER_6_1610 ();
 sg13g2_fill_1 FILLER_6_1627 ();
 sg13g2_decap_8 FILLER_6_1636 ();
 sg13g2_fill_1 FILLER_6_1643 ();
 sg13g2_fill_1 FILLER_6_1667 ();
 sg13g2_decap_4 FILLER_6_1678 ();
 sg13g2_fill_2 FILLER_6_1682 ();
 sg13g2_fill_1 FILLER_6_1687 ();
 sg13g2_decap_8 FILLER_6_1716 ();
 sg13g2_decap_8 FILLER_6_1723 ();
 sg13g2_fill_2 FILLER_6_1735 ();
 sg13g2_decap_8 FILLER_6_1764 ();
 sg13g2_fill_1 FILLER_6_1780 ();
 sg13g2_decap_4 FILLER_6_1788 ();
 sg13g2_decap_8 FILLER_6_1805 ();
 sg13g2_decap_8 FILLER_6_1812 ();
 sg13g2_decap_4 FILLER_6_1819 ();
 sg13g2_fill_1 FILLER_6_1823 ();
 sg13g2_decap_8 FILLER_6_1829 ();
 sg13g2_fill_2 FILLER_6_1836 ();
 sg13g2_fill_1 FILLER_6_1838 ();
 sg13g2_decap_8 FILLER_6_1843 ();
 sg13g2_fill_2 FILLER_6_1850 ();
 sg13g2_fill_1 FILLER_6_1861 ();
 sg13g2_fill_2 FILLER_6_1871 ();
 sg13g2_decap_8 FILLER_6_1909 ();
 sg13g2_decap_4 FILLER_6_1916 ();
 sg13g2_fill_1 FILLER_6_1920 ();
 sg13g2_decap_8 FILLER_6_1962 ();
 sg13g2_decap_4 FILLER_6_1969 ();
 sg13g2_fill_1 FILLER_6_1973 ();
 sg13g2_decap_4 FILLER_6_1984 ();
 sg13g2_fill_1 FILLER_6_1988 ();
 sg13g2_decap_8 FILLER_6_1994 ();
 sg13g2_fill_1 FILLER_6_2001 ();
 sg13g2_decap_4 FILLER_6_2006 ();
 sg13g2_fill_1 FILLER_6_2010 ();
 sg13g2_fill_2 FILLER_6_2028 ();
 sg13g2_decap_8 FILLER_6_2038 ();
 sg13g2_fill_2 FILLER_6_2060 ();
 sg13g2_fill_1 FILLER_6_2062 ();
 sg13g2_decap_4 FILLER_6_2076 ();
 sg13g2_fill_2 FILLER_6_2084 ();
 sg13g2_fill_1 FILLER_6_2086 ();
 sg13g2_fill_2 FILLER_6_2096 ();
 sg13g2_fill_1 FILLER_6_2101 ();
 sg13g2_fill_2 FILLER_6_2130 ();
 sg13g2_decap_8 FILLER_6_2136 ();
 sg13g2_fill_1 FILLER_6_2143 ();
 sg13g2_decap_4 FILLER_6_2151 ();
 sg13g2_decap_4 FILLER_6_2180 ();
 sg13g2_decap_8 FILLER_6_2205 ();
 sg13g2_decap_8 FILLER_6_2212 ();
 sg13g2_decap_8 FILLER_6_2232 ();
 sg13g2_decap_4 FILLER_6_2239 ();
 sg13g2_fill_2 FILLER_6_2243 ();
 sg13g2_decap_4 FILLER_6_2249 ();
 sg13g2_decap_8 FILLER_6_2267 ();
 sg13g2_decap_8 FILLER_6_2274 ();
 sg13g2_fill_2 FILLER_6_2281 ();
 sg13g2_fill_1 FILLER_6_2283 ();
 sg13g2_fill_2 FILLER_6_2312 ();
 sg13g2_fill_1 FILLER_6_2314 ();
 sg13g2_decap_8 FILLER_6_2324 ();
 sg13g2_decap_4 FILLER_6_2331 ();
 sg13g2_fill_1 FILLER_6_2335 ();
 sg13g2_fill_1 FILLER_6_2341 ();
 sg13g2_decap_4 FILLER_6_2356 ();
 sg13g2_fill_1 FILLER_6_2360 ();
 sg13g2_fill_2 FILLER_6_2365 ();
 sg13g2_fill_1 FILLER_6_2367 ();
 sg13g2_decap_4 FILLER_6_2386 ();
 sg13g2_fill_1 FILLER_6_2390 ();
 sg13g2_fill_2 FILLER_6_2460 ();
 sg13g2_fill_1 FILLER_6_2462 ();
 sg13g2_fill_1 FILLER_6_2471 ();
 sg13g2_fill_2 FILLER_6_2496 ();
 sg13g2_fill_1 FILLER_6_2498 ();
 sg13g2_decap_8 FILLER_6_2503 ();
 sg13g2_decap_8 FILLER_6_2510 ();
 sg13g2_decap_8 FILLER_6_2517 ();
 sg13g2_fill_1 FILLER_6_2524 ();
 sg13g2_decap_8 FILLER_6_2536 ();
 sg13g2_decap_8 FILLER_6_2543 ();
 sg13g2_decap_8 FILLER_6_2554 ();
 sg13g2_decap_4 FILLER_6_2561 ();
 sg13g2_fill_2 FILLER_6_2572 ();
 sg13g2_fill_1 FILLER_6_2579 ();
 sg13g2_decap_8 FILLER_6_2585 ();
 sg13g2_decap_4 FILLER_6_2592 ();
 sg13g2_fill_1 FILLER_6_2624 ();
 sg13g2_decap_4 FILLER_6_2638 ();
 sg13g2_fill_1 FILLER_6_2642 ();
 sg13g2_decap_8 FILLER_6_2697 ();
 sg13g2_fill_2 FILLER_6_2704 ();
 sg13g2_fill_1 FILLER_6_2706 ();
 sg13g2_fill_2 FILLER_6_2733 ();
 sg13g2_fill_1 FILLER_6_2735 ();
 sg13g2_fill_2 FILLER_6_2783 ();
 sg13g2_fill_1 FILLER_6_2785 ();
 sg13g2_fill_1 FILLER_6_2793 ();
 sg13g2_decap_4 FILLER_6_2822 ();
 sg13g2_decap_4 FILLER_6_2844 ();
 sg13g2_fill_2 FILLER_6_2857 ();
 sg13g2_decap_8 FILLER_6_2864 ();
 sg13g2_fill_2 FILLER_6_2871 ();
 sg13g2_decap_8 FILLER_6_2890 ();
 sg13g2_decap_8 FILLER_6_2897 ();
 sg13g2_fill_2 FILLER_6_2904 ();
 sg13g2_decap_4 FILLER_6_2910 ();
 sg13g2_fill_1 FILLER_6_2914 ();
 sg13g2_decap_8 FILLER_6_2919 ();
 sg13g2_decap_8 FILLER_6_2926 ();
 sg13g2_fill_1 FILLER_6_2933 ();
 sg13g2_fill_2 FILLER_6_2964 ();
 sg13g2_fill_1 FILLER_6_2966 ();
 sg13g2_fill_1 FILLER_6_3022 ();
 sg13g2_fill_2 FILLER_6_3034 ();
 sg13g2_fill_1 FILLER_6_3036 ();
 sg13g2_fill_1 FILLER_6_3042 ();
 sg13g2_decap_8 FILLER_6_3060 ();
 sg13g2_decap_8 FILLER_6_3067 ();
 sg13g2_decap_8 FILLER_6_3074 ();
 sg13g2_fill_2 FILLER_6_3098 ();
 sg13g2_fill_1 FILLER_6_3106 ();
 sg13g2_decap_8 FILLER_6_3118 ();
 sg13g2_fill_2 FILLER_6_3125 ();
 sg13g2_fill_2 FILLER_6_3158 ();
 sg13g2_fill_1 FILLER_6_3160 ();
 sg13g2_decap_4 FILLER_6_3166 ();
 sg13g2_fill_2 FILLER_6_3188 ();
 sg13g2_fill_1 FILLER_6_3190 ();
 sg13g2_fill_2 FILLER_6_3195 ();
 sg13g2_decap_8 FILLER_6_3213 ();
 sg13g2_fill_1 FILLER_6_3220 ();
 sg13g2_fill_1 FILLER_6_3230 ();
 sg13g2_decap_4 FILLER_6_3235 ();
 sg13g2_decap_8 FILLER_6_3243 ();
 sg13g2_decap_8 FILLER_6_3250 ();
 sg13g2_decap_4 FILLER_6_3257 ();
 sg13g2_fill_2 FILLER_6_3261 ();
 sg13g2_decap_4 FILLER_6_3273 ();
 sg13g2_fill_1 FILLER_6_3277 ();
 sg13g2_fill_2 FILLER_6_3293 ();
 sg13g2_decap_4 FILLER_6_3312 ();
 sg13g2_fill_2 FILLER_6_3316 ();
 sg13g2_decap_8 FILLER_6_3334 ();
 sg13g2_fill_2 FILLER_6_3341 ();
 sg13g2_fill_2 FILLER_6_3365 ();
 sg13g2_decap_8 FILLER_6_3390 ();
 sg13g2_fill_2 FILLER_6_3397 ();
 sg13g2_fill_2 FILLER_6_3420 ();
 sg13g2_decap_4 FILLER_6_3442 ();
 sg13g2_fill_2 FILLER_6_3471 ();
 sg13g2_fill_1 FILLER_6_3473 ();
 sg13g2_fill_1 FILLER_6_3483 ();
 sg13g2_decap_8 FILLER_6_3494 ();
 sg13g2_decap_8 FILLER_6_3529 ();
 sg13g2_decap_8 FILLER_6_3536 ();
 sg13g2_decap_8 FILLER_6_3543 ();
 sg13g2_decap_8 FILLER_6_3550 ();
 sg13g2_decap_8 FILLER_6_3557 ();
 sg13g2_decap_8 FILLER_6_3564 ();
 sg13g2_decap_8 FILLER_6_3571 ();
 sg13g2_fill_2 FILLER_6_3578 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_124 ();
 sg13g2_fill_2 FILLER_7_131 ();
 sg13g2_decap_8 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_151 ();
 sg13g2_fill_2 FILLER_7_158 ();
 sg13g2_fill_2 FILLER_7_175 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_fill_2 FILLER_7_194 ();
 sg13g2_fill_1 FILLER_7_196 ();
 sg13g2_fill_1 FILLER_7_207 ();
 sg13g2_decap_4 FILLER_7_212 ();
 sg13g2_fill_2 FILLER_7_216 ();
 sg13g2_fill_2 FILLER_7_226 ();
 sg13g2_fill_1 FILLER_7_228 ();
 sg13g2_fill_2 FILLER_7_279 ();
 sg13g2_fill_1 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_292 ();
 sg13g2_fill_2 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_fill_2 FILLER_7_333 ();
 sg13g2_fill_2 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_fill_1 FILLER_7_357 ();
 sg13g2_fill_2 FILLER_7_361 ();
 sg13g2_fill_1 FILLER_7_363 ();
 sg13g2_decap_4 FILLER_7_384 ();
 sg13g2_fill_1 FILLER_7_388 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_7_437 ();
 sg13g2_fill_1 FILLER_7_444 ();
 sg13g2_fill_1 FILLER_7_461 ();
 sg13g2_fill_1 FILLER_7_480 ();
 sg13g2_decap_4 FILLER_7_494 ();
 sg13g2_fill_1 FILLER_7_509 ();
 sg13g2_decap_4 FILLER_7_520 ();
 sg13g2_fill_2 FILLER_7_529 ();
 sg13g2_fill_1 FILLER_7_531 ();
 sg13g2_decap_8 FILLER_7_537 ();
 sg13g2_decap_4 FILLER_7_544 ();
 sg13g2_fill_1 FILLER_7_548 ();
 sg13g2_decap_8 FILLER_7_561 ();
 sg13g2_fill_1 FILLER_7_572 ();
 sg13g2_fill_1 FILLER_7_624 ();
 sg13g2_fill_2 FILLER_7_646 ();
 sg13g2_fill_1 FILLER_7_648 ();
 sg13g2_decap_4 FILLER_7_670 ();
 sg13g2_fill_2 FILLER_7_674 ();
 sg13g2_decap_4 FILLER_7_701 ();
 sg13g2_fill_1 FILLER_7_705 ();
 sg13g2_decap_8 FILLER_7_719 ();
 sg13g2_fill_2 FILLER_7_726 ();
 sg13g2_fill_1 FILLER_7_728 ();
 sg13g2_fill_1 FILLER_7_751 ();
 sg13g2_fill_1 FILLER_7_772 ();
 sg13g2_fill_1 FILLER_7_783 ();
 sg13g2_fill_1 FILLER_7_803 ();
 sg13g2_fill_1 FILLER_7_816 ();
 sg13g2_decap_8 FILLER_7_822 ();
 sg13g2_fill_2 FILLER_7_842 ();
 sg13g2_fill_1 FILLER_7_856 ();
 sg13g2_fill_1 FILLER_7_882 ();
 sg13g2_fill_1 FILLER_7_888 ();
 sg13g2_fill_2 FILLER_7_897 ();
 sg13g2_fill_1 FILLER_7_913 ();
 sg13g2_decap_4 FILLER_7_927 ();
 sg13g2_fill_1 FILLER_7_931 ();
 sg13g2_fill_2 FILLER_7_937 ();
 sg13g2_fill_1 FILLER_7_939 ();
 sg13g2_fill_2 FILLER_7_945 ();
 sg13g2_fill_1 FILLER_7_947 ();
 sg13g2_fill_1 FILLER_7_953 ();
 sg13g2_fill_1 FILLER_7_959 ();
 sg13g2_fill_2 FILLER_7_968 ();
 sg13g2_fill_1 FILLER_7_970 ();
 sg13g2_decap_8 FILLER_7_979 ();
 sg13g2_decap_4 FILLER_7_986 ();
 sg13g2_decap_8 FILLER_7_994 ();
 sg13g2_decap_8 FILLER_7_1001 ();
 sg13g2_decap_8 FILLER_7_1008 ();
 sg13g2_fill_2 FILLER_7_1015 ();
 sg13g2_fill_1 FILLER_7_1017 ();
 sg13g2_fill_1 FILLER_7_1027 ();
 sg13g2_fill_2 FILLER_7_1059 ();
 sg13g2_fill_2 FILLER_7_1078 ();
 sg13g2_decap_4 FILLER_7_1094 ();
 sg13g2_fill_2 FILLER_7_1098 ();
 sg13g2_decap_8 FILLER_7_1120 ();
 sg13g2_decap_4 FILLER_7_1127 ();
 sg13g2_fill_2 FILLER_7_1138 ();
 sg13g2_decap_8 FILLER_7_1145 ();
 sg13g2_fill_1 FILLER_7_1152 ();
 sg13g2_fill_2 FILLER_7_1176 ();
 sg13g2_fill_2 FILLER_7_1206 ();
 sg13g2_fill_1 FILLER_7_1208 ();
 sg13g2_decap_8 FILLER_7_1244 ();
 sg13g2_fill_2 FILLER_7_1251 ();
 sg13g2_decap_4 FILLER_7_1282 ();
 sg13g2_fill_2 FILLER_7_1286 ();
 sg13g2_decap_8 FILLER_7_1293 ();
 sg13g2_decap_4 FILLER_7_1300 ();
 sg13g2_fill_1 FILLER_7_1329 ();
 sg13g2_decap_4 FILLER_7_1338 ();
 sg13g2_fill_2 FILLER_7_1342 ();
 sg13g2_decap_8 FILLER_7_1359 ();
 sg13g2_decap_8 FILLER_7_1366 ();
 sg13g2_decap_4 FILLER_7_1382 ();
 sg13g2_decap_4 FILLER_7_1399 ();
 sg13g2_fill_2 FILLER_7_1403 ();
 sg13g2_decap_8 FILLER_7_1421 ();
 sg13g2_fill_2 FILLER_7_1428 ();
 sg13g2_fill_2 FILLER_7_1440 ();
 sg13g2_fill_1 FILLER_7_1442 ();
 sg13g2_decap_8 FILLER_7_1453 ();
 sg13g2_fill_2 FILLER_7_1460 ();
 sg13g2_fill_1 FILLER_7_1462 ();
 sg13g2_decap_8 FILLER_7_1527 ();
 sg13g2_decap_4 FILLER_7_1534 ();
 sg13g2_fill_2 FILLER_7_1538 ();
 sg13g2_decap_8 FILLER_7_1551 ();
 sg13g2_fill_1 FILLER_7_1571 ();
 sg13g2_decap_8 FILLER_7_1590 ();
 sg13g2_decap_4 FILLER_7_1597 ();
 sg13g2_fill_1 FILLER_7_1647 ();
 sg13g2_fill_2 FILLER_7_1672 ();
 sg13g2_decap_8 FILLER_7_1682 ();
 sg13g2_decap_4 FILLER_7_1689 ();
 sg13g2_decap_8 FILLER_7_1697 ();
 sg13g2_decap_4 FILLER_7_1704 ();
 sg13g2_fill_2 FILLER_7_1708 ();
 sg13g2_fill_2 FILLER_7_1756 ();
 sg13g2_decap_8 FILLER_7_1770 ();
 sg13g2_decap_8 FILLER_7_1777 ();
 sg13g2_fill_2 FILLER_7_1789 ();
 sg13g2_fill_1 FILLER_7_1791 ();
 sg13g2_fill_2 FILLER_7_1811 ();
 sg13g2_fill_1 FILLER_7_1833 ();
 sg13g2_fill_2 FILLER_7_1842 ();
 sg13g2_fill_1 FILLER_7_1844 ();
 sg13g2_fill_1 FILLER_7_1895 ();
 sg13g2_fill_1 FILLER_7_1908 ();
 sg13g2_decap_4 FILLER_7_1922 ();
 sg13g2_decap_8 FILLER_7_1930 ();
 sg13g2_decap_8 FILLER_7_1937 ();
 sg13g2_decap_4 FILLER_7_1944 ();
 sg13g2_fill_1 FILLER_7_1948 ();
 sg13g2_fill_2 FILLER_7_1977 ();
 sg13g2_fill_2 FILLER_7_1999 ();
 sg13g2_fill_1 FILLER_7_2001 ();
 sg13g2_decap_4 FILLER_7_2012 ();
 sg13g2_fill_1 FILLER_7_2037 ();
 sg13g2_decap_4 FILLER_7_2054 ();
 sg13g2_decap_4 FILLER_7_2071 ();
 sg13g2_fill_1 FILLER_7_2103 ();
 sg13g2_decap_8 FILLER_7_2117 ();
 sg13g2_fill_2 FILLER_7_2124 ();
 sg13g2_fill_1 FILLER_7_2126 ();
 sg13g2_decap_8 FILLER_7_2155 ();
 sg13g2_fill_2 FILLER_7_2162 ();
 sg13g2_decap_8 FILLER_7_2169 ();
 sg13g2_fill_2 FILLER_7_2176 ();
 sg13g2_fill_1 FILLER_7_2178 ();
 sg13g2_decap_4 FILLER_7_2186 ();
 sg13g2_fill_2 FILLER_7_2190 ();
 sg13g2_decap_8 FILLER_7_2201 ();
 sg13g2_decap_8 FILLER_7_2208 ();
 sg13g2_decap_4 FILLER_7_2215 ();
 sg13g2_fill_2 FILLER_7_2219 ();
 sg13g2_decap_8 FILLER_7_2235 ();
 sg13g2_fill_1 FILLER_7_2242 ();
 sg13g2_fill_2 FILLER_7_2264 ();
 sg13g2_fill_1 FILLER_7_2266 ();
 sg13g2_decap_8 FILLER_7_2277 ();
 sg13g2_decap_4 FILLER_7_2284 ();
 sg13g2_fill_1 FILLER_7_2288 ();
 sg13g2_decap_8 FILLER_7_2298 ();
 sg13g2_decap_4 FILLER_7_2305 ();
 sg13g2_fill_2 FILLER_7_2309 ();
 sg13g2_decap_8 FILLER_7_2361 ();
 sg13g2_decap_4 FILLER_7_2368 ();
 sg13g2_fill_1 FILLER_7_2372 ();
 sg13g2_decap_8 FILLER_7_2386 ();
 sg13g2_decap_8 FILLER_7_2393 ();
 sg13g2_decap_8 FILLER_7_2400 ();
 sg13g2_fill_1 FILLER_7_2407 ();
 sg13g2_decap_8 FILLER_7_2413 ();
 sg13g2_decap_8 FILLER_7_2420 ();
 sg13g2_fill_2 FILLER_7_2427 ();
 sg13g2_fill_1 FILLER_7_2429 ();
 sg13g2_fill_1 FILLER_7_2437 ();
 sg13g2_fill_2 FILLER_7_2476 ();
 sg13g2_fill_1 FILLER_7_2478 ();
 sg13g2_fill_2 FILLER_7_2484 ();
 sg13g2_fill_1 FILLER_7_2486 ();
 sg13g2_decap_4 FILLER_7_2522 ();
 sg13g2_decap_8 FILLER_7_2554 ();
 sg13g2_decap_8 FILLER_7_2561 ();
 sg13g2_decap_8 FILLER_7_2568 ();
 sg13g2_decap_4 FILLER_7_2575 ();
 sg13g2_fill_1 FILLER_7_2579 ();
 sg13g2_decap_8 FILLER_7_2593 ();
 sg13g2_fill_1 FILLER_7_2600 ();
 sg13g2_fill_2 FILLER_7_2610 ();
 sg13g2_decap_4 FILLER_7_2621 ();
 sg13g2_fill_1 FILLER_7_2625 ();
 sg13g2_fill_2 FILLER_7_2631 ();
 sg13g2_fill_1 FILLER_7_2633 ();
 sg13g2_fill_2 FILLER_7_2639 ();
 sg13g2_decap_8 FILLER_7_2652 ();
 sg13g2_decap_4 FILLER_7_2659 ();
 sg13g2_fill_1 FILLER_7_2663 ();
 sg13g2_fill_2 FILLER_7_2668 ();
 sg13g2_decap_4 FILLER_7_2675 ();
 sg13g2_fill_2 FILLER_7_2715 ();
 sg13g2_decap_8 FILLER_7_2726 ();
 sg13g2_fill_2 FILLER_7_2733 ();
 sg13g2_fill_1 FILLER_7_2735 ();
 sg13g2_decap_4 FILLER_7_2744 ();
 sg13g2_decap_8 FILLER_7_2752 ();
 sg13g2_decap_8 FILLER_7_2759 ();
 sg13g2_fill_2 FILLER_7_2766 ();
 sg13g2_decap_8 FILLER_7_2786 ();
 sg13g2_fill_2 FILLER_7_2793 ();
 sg13g2_fill_2 FILLER_7_2804 ();
 sg13g2_fill_1 FILLER_7_2806 ();
 sg13g2_decap_8 FILLER_7_2811 ();
 sg13g2_decap_4 FILLER_7_2818 ();
 sg13g2_fill_2 FILLER_7_2822 ();
 sg13g2_fill_2 FILLER_7_2855 ();
 sg13g2_fill_2 FILLER_7_2866 ();
 sg13g2_fill_1 FILLER_7_2868 ();
 sg13g2_fill_1 FILLER_7_2874 ();
 sg13g2_decap_8 FILLER_7_2885 ();
 sg13g2_decap_4 FILLER_7_2892 ();
 sg13g2_fill_2 FILLER_7_2896 ();
 sg13g2_decap_8 FILLER_7_2913 ();
 sg13g2_decap_4 FILLER_7_2920 ();
 sg13g2_fill_2 FILLER_7_2924 ();
 sg13g2_decap_4 FILLER_7_2950 ();
 sg13g2_decap_4 FILLER_7_2988 ();
 sg13g2_fill_1 FILLER_7_2992 ();
 sg13g2_decap_4 FILLER_7_2998 ();
 sg13g2_decap_4 FILLER_7_3012 ();
 sg13g2_fill_2 FILLER_7_3021 ();
 sg13g2_fill_1 FILLER_7_3023 ();
 sg13g2_decap_8 FILLER_7_3051 ();
 sg13g2_decap_8 FILLER_7_3063 ();
 sg13g2_decap_8 FILLER_7_3105 ();
 sg13g2_fill_2 FILLER_7_3112 ();
 sg13g2_decap_4 FILLER_7_3127 ();
 sg13g2_decap_8 FILLER_7_3139 ();
 sg13g2_fill_2 FILLER_7_3146 ();
 sg13g2_decap_4 FILLER_7_3153 ();
 sg13g2_fill_1 FILLER_7_3157 ();
 sg13g2_decap_8 FILLER_7_3163 ();
 sg13g2_decap_8 FILLER_7_3170 ();
 sg13g2_fill_2 FILLER_7_3181 ();
 sg13g2_decap_8 FILLER_7_3200 ();
 sg13g2_decap_8 FILLER_7_3207 ();
 sg13g2_decap_4 FILLER_7_3214 ();
 sg13g2_fill_1 FILLER_7_3218 ();
 sg13g2_decap_8 FILLER_7_3254 ();
 sg13g2_fill_1 FILLER_7_3261 ();
 sg13g2_fill_2 FILLER_7_3273 ();
 sg13g2_decap_8 FILLER_7_3278 ();
 sg13g2_fill_2 FILLER_7_3285 ();
 sg13g2_fill_1 FILLER_7_3287 ();
 sg13g2_decap_8 FILLER_7_3304 ();
 sg13g2_decap_8 FILLER_7_3311 ();
 sg13g2_fill_2 FILLER_7_3326 ();
 sg13g2_decap_8 FILLER_7_3336 ();
 sg13g2_decap_8 FILLER_7_3343 ();
 sg13g2_decap_4 FILLER_7_3366 ();
 sg13g2_decap_4 FILLER_7_3390 ();
 sg13g2_fill_1 FILLER_7_3399 ();
 sg13g2_fill_1 FILLER_7_3418 ();
 sg13g2_fill_1 FILLER_7_3428 ();
 sg13g2_decap_8 FILLER_7_3446 ();
 sg13g2_fill_2 FILLER_7_3462 ();
 sg13g2_fill_1 FILLER_7_3464 ();
 sg13g2_fill_2 FILLER_7_3473 ();
 sg13g2_fill_1 FILLER_7_3475 ();
 sg13g2_decap_4 FILLER_7_3491 ();
 sg13g2_fill_1 FILLER_7_3502 ();
 sg13g2_decap_8 FILLER_7_3511 ();
 sg13g2_decap_8 FILLER_7_3518 ();
 sg13g2_decap_8 FILLER_7_3525 ();
 sg13g2_decap_8 FILLER_7_3532 ();
 sg13g2_decap_8 FILLER_7_3539 ();
 sg13g2_decap_8 FILLER_7_3546 ();
 sg13g2_decap_8 FILLER_7_3553 ();
 sg13g2_decap_8 FILLER_7_3560 ();
 sg13g2_decap_8 FILLER_7_3567 ();
 sg13g2_decap_4 FILLER_7_3574 ();
 sg13g2_fill_2 FILLER_7_3578 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_4 FILLER_8_105 ();
 sg13g2_fill_2 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_174 ();
 sg13g2_fill_1 FILLER_8_176 ();
 sg13g2_fill_1 FILLER_8_211 ();
 sg13g2_fill_2 FILLER_8_230 ();
 sg13g2_fill_1 FILLER_8_232 ();
 sg13g2_fill_2 FILLER_8_241 ();
 sg13g2_fill_1 FILLER_8_243 ();
 sg13g2_decap_8 FILLER_8_248 ();
 sg13g2_decap_4 FILLER_8_255 ();
 sg13g2_fill_2 FILLER_8_275 ();
 sg13g2_fill_2 FILLER_8_293 ();
 sg13g2_fill_2 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_330 ();
 sg13g2_fill_1 FILLER_8_332 ();
 sg13g2_fill_2 FILLER_8_352 ();
 sg13g2_fill_1 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_fill_1 FILLER_8_391 ();
 sg13g2_fill_1 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_409 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_4 FILLER_8_423 ();
 sg13g2_fill_1 FILLER_8_440 ();
 sg13g2_fill_1 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_468 ();
 sg13g2_decap_4 FILLER_8_475 ();
 sg13g2_decap_8 FILLER_8_496 ();
 sg13g2_fill_1 FILLER_8_503 ();
 sg13g2_decap_4 FILLER_8_511 ();
 sg13g2_fill_1 FILLER_8_530 ();
 sg13g2_decap_8 FILLER_8_536 ();
 sg13g2_fill_2 FILLER_8_566 ();
 sg13g2_fill_1 FILLER_8_568 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_fill_2 FILLER_8_595 ();
 sg13g2_fill_1 FILLER_8_597 ();
 sg13g2_fill_2 FILLER_8_617 ();
 sg13g2_fill_1 FILLER_8_625 ();
 sg13g2_decap_8 FILLER_8_643 ();
 sg13g2_fill_2 FILLER_8_650 ();
 sg13g2_decap_8 FILLER_8_671 ();
 sg13g2_fill_1 FILLER_8_678 ();
 sg13g2_fill_2 FILLER_8_696 ();
 sg13g2_fill_1 FILLER_8_698 ();
 sg13g2_decap_8 FILLER_8_719 ();
 sg13g2_decap_8 FILLER_8_726 ();
 sg13g2_decap_4 FILLER_8_733 ();
 sg13g2_fill_2 FILLER_8_737 ();
 sg13g2_fill_1 FILLER_8_760 ();
 sg13g2_decap_4 FILLER_8_774 ();
 sg13g2_decap_8 FILLER_8_786 ();
 sg13g2_fill_2 FILLER_8_793 ();
 sg13g2_decap_4 FILLER_8_800 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_fill_1 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_849 ();
 sg13g2_decap_8 FILLER_8_856 ();
 sg13g2_fill_2 FILLER_8_863 ();
 sg13g2_fill_2 FILLER_8_873 ();
 sg13g2_fill_1 FILLER_8_875 ();
 sg13g2_fill_2 FILLER_8_881 ();
 sg13g2_fill_1 FILLER_8_887 ();
 sg13g2_fill_1 FILLER_8_897 ();
 sg13g2_fill_2 FILLER_8_902 ();
 sg13g2_fill_1 FILLER_8_904 ();
 sg13g2_fill_2 FILLER_8_913 ();
 sg13g2_fill_2 FILLER_8_920 ();
 sg13g2_fill_2 FILLER_8_926 ();
 sg13g2_decap_4 FILLER_8_933 ();
 sg13g2_fill_1 FILLER_8_937 ();
 sg13g2_decap_4 FILLER_8_943 ();
 sg13g2_fill_1 FILLER_8_947 ();
 sg13g2_decap_8 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_987 ();
 sg13g2_fill_1 FILLER_8_994 ();
 sg13g2_decap_8 FILLER_8_1020 ();
 sg13g2_decap_4 FILLER_8_1027 ();
 sg13g2_fill_1 FILLER_8_1031 ();
 sg13g2_decap_8 FILLER_8_1036 ();
 sg13g2_fill_2 FILLER_8_1043 ();
 sg13g2_fill_1 FILLER_8_1045 ();
 sg13g2_decap_8 FILLER_8_1058 ();
 sg13g2_decap_4 FILLER_8_1065 ();
 sg13g2_fill_2 FILLER_8_1069 ();
 sg13g2_decap_4 FILLER_8_1099 ();
 sg13g2_fill_1 FILLER_8_1107 ();
 sg13g2_fill_1 FILLER_8_1116 ();
 sg13g2_decap_8 FILLER_8_1149 ();
 sg13g2_fill_2 FILLER_8_1156 ();
 sg13g2_fill_2 FILLER_8_1170 ();
 sg13g2_fill_1 FILLER_8_1172 ();
 sg13g2_decap_4 FILLER_8_1178 ();
 sg13g2_fill_1 FILLER_8_1182 ();
 sg13g2_decap_4 FILLER_8_1190 ();
 sg13g2_fill_2 FILLER_8_1194 ();
 sg13g2_decap_8 FILLER_8_1200 ();
 sg13g2_decap_8 FILLER_8_1207 ();
 sg13g2_fill_1 FILLER_8_1214 ();
 sg13g2_decap_8 FILLER_8_1219 ();
 sg13g2_fill_1 FILLER_8_1226 ();
 sg13g2_decap_8 FILLER_8_1239 ();
 sg13g2_decap_8 FILLER_8_1246 ();
 sg13g2_decap_8 FILLER_8_1253 ();
 sg13g2_decap_4 FILLER_8_1260 ();
 sg13g2_fill_1 FILLER_8_1264 ();
 sg13g2_fill_1 FILLER_8_1275 ();
 sg13g2_fill_2 FILLER_8_1289 ();
 sg13g2_decap_8 FILLER_8_1300 ();
 sg13g2_fill_1 FILLER_8_1307 ();
 sg13g2_decap_4 FILLER_8_1334 ();
 sg13g2_fill_2 FILLER_8_1338 ();
 sg13g2_fill_2 FILLER_8_1362 ();
 sg13g2_decap_4 FILLER_8_1391 ();
 sg13g2_fill_2 FILLER_8_1395 ();
 sg13g2_fill_1 FILLER_8_1413 ();
 sg13g2_fill_2 FILLER_8_1419 ();
 sg13g2_fill_1 FILLER_8_1421 ();
 sg13g2_decap_8 FILLER_8_1455 ();
 sg13g2_decap_4 FILLER_8_1467 ();
 sg13g2_decap_8 FILLER_8_1484 ();
 sg13g2_decap_4 FILLER_8_1491 ();
 sg13g2_fill_2 FILLER_8_1495 ();
 sg13g2_fill_2 FILLER_8_1501 ();
 sg13g2_decap_8 FILLER_8_1512 ();
 sg13g2_fill_2 FILLER_8_1519 ();
 sg13g2_fill_1 FILLER_8_1521 ();
 sg13g2_fill_2 FILLER_8_1563 ();
 sg13g2_fill_1 FILLER_8_1565 ();
 sg13g2_fill_2 FILLER_8_1574 ();
 sg13g2_decap_8 FILLER_8_1600 ();
 sg13g2_fill_1 FILLER_8_1607 ();
 sg13g2_fill_1 FILLER_8_1611 ();
 sg13g2_decap_4 FILLER_8_1620 ();
 sg13g2_fill_2 FILLER_8_1629 ();
 sg13g2_fill_1 FILLER_8_1631 ();
 sg13g2_decap_8 FILLER_8_1650 ();
 sg13g2_fill_2 FILLER_8_1665 ();
 sg13g2_fill_1 FILLER_8_1667 ();
 sg13g2_decap_4 FILLER_8_1677 ();
 sg13g2_fill_2 FILLER_8_1681 ();
 sg13g2_fill_1 FILLER_8_1688 ();
 sg13g2_fill_2 FILLER_8_1694 ();
 sg13g2_decap_4 FILLER_8_1710 ();
 sg13g2_fill_1 FILLER_8_1714 ();
 sg13g2_decap_8 FILLER_8_1719 ();
 sg13g2_decap_4 FILLER_8_1733 ();
 sg13g2_fill_2 FILLER_8_1737 ();
 sg13g2_decap_4 FILLER_8_1749 ();
 sg13g2_fill_1 FILLER_8_1753 ();
 sg13g2_fill_2 FILLER_8_1775 ();
 sg13g2_fill_1 FILLER_8_1777 ();
 sg13g2_fill_2 FILLER_8_1782 ();
 sg13g2_fill_1 FILLER_8_1784 ();
 sg13g2_fill_2 FILLER_8_1801 ();
 sg13g2_fill_1 FILLER_8_1817 ();
 sg13g2_decap_8 FILLER_8_1843 ();
 sg13g2_fill_2 FILLER_8_1850 ();
 sg13g2_decap_4 FILLER_8_1861 ();
 sg13g2_fill_2 FILLER_8_1872 ();
 sg13g2_fill_1 FILLER_8_1874 ();
 sg13g2_fill_2 FILLER_8_1884 ();
 sg13g2_fill_1 FILLER_8_1886 ();
 sg13g2_fill_1 FILLER_8_1895 ();
 sg13g2_decap_8 FILLER_8_1937 ();
 sg13g2_decap_4 FILLER_8_1944 ();
 sg13g2_fill_1 FILLER_8_1948 ();
 sg13g2_decap_8 FILLER_8_1969 ();
 sg13g2_fill_2 FILLER_8_1976 ();
 sg13g2_fill_2 FILLER_8_1989 ();
 sg13g2_fill_1 FILLER_8_1991 ();
 sg13g2_decap_4 FILLER_8_2017 ();
 sg13g2_fill_2 FILLER_8_2029 ();
 sg13g2_decap_4 FILLER_8_2075 ();
 sg13g2_fill_2 FILLER_8_2079 ();
 sg13g2_decap_8 FILLER_8_2086 ();
 sg13g2_decap_4 FILLER_8_2093 ();
 sg13g2_fill_2 FILLER_8_2097 ();
 sg13g2_decap_4 FILLER_8_2127 ();
 sg13g2_decap_8 FILLER_8_2139 ();
 sg13g2_decap_8 FILLER_8_2146 ();
 sg13g2_fill_1 FILLER_8_2153 ();
 sg13g2_decap_8 FILLER_8_2186 ();
 sg13g2_fill_2 FILLER_8_2193 ();
 sg13g2_fill_2 FILLER_8_2210 ();
 sg13g2_fill_1 FILLER_8_2212 ();
 sg13g2_fill_2 FILLER_8_2238 ();
 sg13g2_fill_1 FILLER_8_2240 ();
 sg13g2_decap_4 FILLER_8_2258 ();
 sg13g2_fill_2 FILLER_8_2280 ();
 sg13g2_fill_2 FILLER_8_2286 ();
 sg13g2_fill_1 FILLER_8_2288 ();
 sg13g2_fill_2 FILLER_8_2302 ();
 sg13g2_fill_1 FILLER_8_2304 ();
 sg13g2_fill_2 FILLER_8_2335 ();
 sg13g2_fill_1 FILLER_8_2337 ();
 sg13g2_fill_2 FILLER_8_2341 ();
 sg13g2_fill_1 FILLER_8_2343 ();
 sg13g2_decap_4 FILLER_8_2357 ();
 sg13g2_fill_1 FILLER_8_2361 ();
 sg13g2_fill_2 FILLER_8_2378 ();
 sg13g2_fill_1 FILLER_8_2380 ();
 sg13g2_fill_1 FILLER_8_2397 ();
 sg13g2_fill_2 FILLER_8_2454 ();
 sg13g2_fill_1 FILLER_8_2456 ();
 sg13g2_decap_8 FILLER_8_2497 ();
 sg13g2_decap_4 FILLER_8_2504 ();
 sg13g2_fill_1 FILLER_8_2508 ();
 sg13g2_decap_8 FILLER_8_2520 ();
 sg13g2_decap_4 FILLER_8_2527 ();
 sg13g2_decap_8 FILLER_8_2535 ();
 sg13g2_fill_2 FILLER_8_2542 ();
 sg13g2_fill_1 FILLER_8_2544 ();
 sg13g2_decap_4 FILLER_8_2565 ();
 sg13g2_fill_2 FILLER_8_2569 ();
 sg13g2_fill_1 FILLER_8_2583 ();
 sg13g2_fill_1 FILLER_8_2595 ();
 sg13g2_fill_1 FILLER_8_2614 ();
 sg13g2_fill_1 FILLER_8_2624 ();
 sg13g2_decap_8 FILLER_8_2644 ();
 sg13g2_fill_2 FILLER_8_2651 ();
 sg13g2_decap_4 FILLER_8_2688 ();
 sg13g2_decap_8 FILLER_8_2696 ();
 sg13g2_decap_4 FILLER_8_2703 ();
 sg13g2_fill_2 FILLER_8_2727 ();
 sg13g2_fill_1 FILLER_8_2729 ();
 sg13g2_decap_8 FILLER_8_2754 ();
 sg13g2_fill_2 FILLER_8_2761 ();
 sg13g2_fill_1 FILLER_8_2763 ();
 sg13g2_fill_2 FILLER_8_2790 ();
 sg13g2_fill_1 FILLER_8_2792 ();
 sg13g2_fill_1 FILLER_8_2800 ();
 sg13g2_fill_2 FILLER_8_2821 ();
 sg13g2_fill_1 FILLER_8_2823 ();
 sg13g2_decap_8 FILLER_8_2828 ();
 sg13g2_fill_2 FILLER_8_2835 ();
 sg13g2_fill_1 FILLER_8_2837 ();
 sg13g2_fill_1 FILLER_8_2862 ();
 sg13g2_decap_8 FILLER_8_2881 ();
 sg13g2_fill_2 FILLER_8_2888 ();
 sg13g2_fill_1 FILLER_8_2890 ();
 sg13g2_fill_1 FILLER_8_2919 ();
 sg13g2_fill_1 FILLER_8_2930 ();
 sg13g2_fill_2 FILLER_8_2947 ();
 sg13g2_fill_2 FILLER_8_2975 ();
 sg13g2_fill_1 FILLER_8_2990 ();
 sg13g2_fill_1 FILLER_8_3001 ();
 sg13g2_decap_4 FILLER_8_3024 ();
 sg13g2_fill_1 FILLER_8_3028 ();
 sg13g2_decap_4 FILLER_8_3033 ();
 sg13g2_decap_4 FILLER_8_3041 ();
 sg13g2_fill_1 FILLER_8_3060 ();
 sg13g2_decap_4 FILLER_8_3071 ();
 sg13g2_fill_1 FILLER_8_3075 ();
 sg13g2_decap_8 FILLER_8_3091 ();
 sg13g2_decap_8 FILLER_8_3098 ();
 sg13g2_fill_2 FILLER_8_3105 ();
 sg13g2_fill_1 FILLER_8_3107 ();
 sg13g2_fill_2 FILLER_8_3121 ();
 sg13g2_fill_1 FILLER_8_3123 ();
 sg13g2_fill_1 FILLER_8_3144 ();
 sg13g2_decap_4 FILLER_8_3179 ();
 sg13g2_fill_1 FILLER_8_3183 ();
 sg13g2_decap_8 FILLER_8_3229 ();
 sg13g2_fill_2 FILLER_8_3253 ();
 sg13g2_fill_1 FILLER_8_3255 ();
 sg13g2_decap_8 FILLER_8_3263 ();
 sg13g2_decap_4 FILLER_8_3298 ();
 sg13g2_fill_1 FILLER_8_3312 ();
 sg13g2_fill_2 FILLER_8_3326 ();
 sg13g2_decap_4 FILLER_8_3340 ();
 sg13g2_fill_2 FILLER_8_3360 ();
 sg13g2_fill_1 FILLER_8_3362 ();
 sg13g2_fill_1 FILLER_8_3376 ();
 sg13g2_decap_8 FILLER_8_3446 ();
 sg13g2_fill_2 FILLER_8_3453 ();
 sg13g2_decap_8 FILLER_8_3475 ();
 sg13g2_fill_2 FILLER_8_3482 ();
 sg13g2_fill_1 FILLER_8_3484 ();
 sg13g2_decap_4 FILLER_8_3489 ();
 sg13g2_fill_1 FILLER_8_3493 ();
 sg13g2_fill_1 FILLER_8_3501 ();
 sg13g2_decap_8 FILLER_8_3530 ();
 sg13g2_decap_8 FILLER_8_3537 ();
 sg13g2_decap_8 FILLER_8_3544 ();
 sg13g2_decap_8 FILLER_8_3551 ();
 sg13g2_decap_8 FILLER_8_3558 ();
 sg13g2_decap_8 FILLER_8_3565 ();
 sg13g2_decap_8 FILLER_8_3572 ();
 sg13g2_fill_1 FILLER_8_3579 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_89 ();
 sg13g2_fill_1 FILLER_9_96 ();
 sg13g2_fill_2 FILLER_9_102 ();
 sg13g2_fill_1 FILLER_9_104 ();
 sg13g2_decap_8 FILLER_9_110 ();
 sg13g2_decap_4 FILLER_9_117 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_148 ();
 sg13g2_decap_8 FILLER_9_155 ();
 sg13g2_fill_1 FILLER_9_162 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_fill_2 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_decap_4 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_211 ();
 sg13g2_decap_4 FILLER_9_258 ();
 sg13g2_fill_1 FILLER_9_262 ();
 sg13g2_decap_4 FILLER_9_276 ();
 sg13g2_fill_1 FILLER_9_280 ();
 sg13g2_decap_4 FILLER_9_285 ();
 sg13g2_fill_2 FILLER_9_289 ();
 sg13g2_decap_4 FILLER_9_295 ();
 sg13g2_fill_2 FILLER_9_299 ();
 sg13g2_fill_2 FILLER_9_322 ();
 sg13g2_fill_1 FILLER_9_324 ();
 sg13g2_fill_1 FILLER_9_352 ();
 sg13g2_fill_1 FILLER_9_386 ();
 sg13g2_fill_1 FILLER_9_415 ();
 sg13g2_fill_1 FILLER_9_446 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_4 FILLER_9_469 ();
 sg13g2_fill_2 FILLER_9_514 ();
 sg13g2_decap_8 FILLER_9_529 ();
 sg13g2_decap_8 FILLER_9_536 ();
 sg13g2_fill_1 FILLER_9_543 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_4 FILLER_9_567 ();
 sg13g2_fill_1 FILLER_9_571 ();
 sg13g2_decap_4 FILLER_9_588 ();
 sg13g2_fill_2 FILLER_9_592 ();
 sg13g2_fill_2 FILLER_9_599 ();
 sg13g2_fill_1 FILLER_9_618 ();
 sg13g2_fill_2 FILLER_9_637 ();
 sg13g2_fill_1 FILLER_9_639 ();
 sg13g2_fill_2 FILLER_9_681 ();
 sg13g2_decap_8 FILLER_9_696 ();
 sg13g2_decap_4 FILLER_9_703 ();
 sg13g2_fill_1 FILLER_9_707 ();
 sg13g2_fill_2 FILLER_9_712 ();
 sg13g2_decap_4 FILLER_9_749 ();
 sg13g2_fill_2 FILLER_9_753 ();
 sg13g2_decap_8 FILLER_9_790 ();
 sg13g2_fill_2 FILLER_9_797 ();
 sg13g2_decap_4 FILLER_9_821 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_fill_1 FILLER_9_862 ();
 sg13g2_fill_1 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_895 ();
 sg13g2_fill_1 FILLER_9_902 ();
 sg13g2_decap_8 FILLER_9_908 ();
 sg13g2_fill_2 FILLER_9_915 ();
 sg13g2_fill_2 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_947 ();
 sg13g2_decap_4 FILLER_9_954 ();
 sg13g2_decap_8 FILLER_9_967 ();
 sg13g2_fill_2 FILLER_9_974 ();
 sg13g2_fill_2 FILLER_9_993 ();
 sg13g2_fill_2 FILLER_9_1023 ();
 sg13g2_decap_4 FILLER_9_1056 ();
 sg13g2_fill_1 FILLER_9_1073 ();
 sg13g2_fill_2 FILLER_9_1088 ();
 sg13g2_fill_1 FILLER_9_1090 ();
 sg13g2_decap_8 FILLER_9_1102 ();
 sg13g2_decap_4 FILLER_9_1109 ();
 sg13g2_fill_1 FILLER_9_1113 ();
 sg13g2_fill_2 FILLER_9_1133 ();
 sg13g2_fill_1 FILLER_9_1135 ();
 sg13g2_decap_8 FILLER_9_1145 ();
 sg13g2_fill_2 FILLER_9_1152 ();
 sg13g2_fill_1 FILLER_9_1154 ();
 sg13g2_decap_8 FILLER_9_1160 ();
 sg13g2_fill_2 FILLER_9_1173 ();
 sg13g2_fill_1 FILLER_9_1175 ();
 sg13g2_decap_8 FILLER_9_1218 ();
 sg13g2_decap_8 FILLER_9_1225 ();
 sg13g2_fill_2 FILLER_9_1249 ();
 sg13g2_fill_2 FILLER_9_1281 ();
 sg13g2_decap_8 FILLER_9_1301 ();
 sg13g2_decap_4 FILLER_9_1308 ();
 sg13g2_fill_2 FILLER_9_1312 ();
 sg13g2_decap_4 FILLER_9_1330 ();
 sg13g2_fill_2 FILLER_9_1334 ();
 sg13g2_decap_4 FILLER_9_1364 ();
 sg13g2_decap_8 FILLER_9_1396 ();
 sg13g2_decap_4 FILLER_9_1411 ();
 sg13g2_decap_8 FILLER_9_1420 ();
 sg13g2_fill_2 FILLER_9_1441 ();
 sg13g2_fill_1 FILLER_9_1443 ();
 sg13g2_decap_8 FILLER_9_1455 ();
 sg13g2_fill_1 FILLER_9_1462 ();
 sg13g2_fill_1 FILLER_9_1495 ();
 sg13g2_decap_8 FILLER_9_1520 ();
 sg13g2_fill_2 FILLER_9_1531 ();
 sg13g2_fill_2 FILLER_9_1546 ();
 sg13g2_fill_1 FILLER_9_1548 ();
 sg13g2_fill_1 FILLER_9_1562 ();
 sg13g2_decap_8 FILLER_9_1571 ();
 sg13g2_decap_8 FILLER_9_1578 ();
 sg13g2_fill_2 FILLER_9_1585 ();
 sg13g2_fill_1 FILLER_9_1587 ();
 sg13g2_decap_4 FILLER_9_1626 ();
 sg13g2_fill_2 FILLER_9_1647 ();
 sg13g2_fill_2 FILLER_9_1662 ();
 sg13g2_fill_1 FILLER_9_1664 ();
 sg13g2_fill_2 FILLER_9_1678 ();
 sg13g2_decap_4 FILLER_9_1686 ();
 sg13g2_fill_2 FILLER_9_1708 ();
 sg13g2_decap_8 FILLER_9_1714 ();
 sg13g2_fill_2 FILLER_9_1721 ();
 sg13g2_decap_8 FILLER_9_1751 ();
 sg13g2_decap_8 FILLER_9_1758 ();
 sg13g2_fill_2 FILLER_9_1765 ();
 sg13g2_fill_2 FILLER_9_1771 ();
 sg13g2_fill_1 FILLER_9_1781 ();
 sg13g2_fill_1 FILLER_9_1798 ();
 sg13g2_decap_4 FILLER_9_1824 ();
 sg13g2_fill_1 FILLER_9_1828 ();
 sg13g2_decap_4 FILLER_9_1839 ();
 sg13g2_fill_2 FILLER_9_1843 ();
 sg13g2_decap_4 FILLER_9_1866 ();
 sg13g2_fill_2 FILLER_9_1870 ();
 sg13g2_fill_2 FILLER_9_1884 ();
 sg13g2_fill_1 FILLER_9_1894 ();
 sg13g2_decap_8 FILLER_9_1904 ();
 sg13g2_fill_1 FILLER_9_1911 ();
 sg13g2_decap_8 FILLER_9_1920 ();
 sg13g2_decap_4 FILLER_9_1927 ();
 sg13g2_fill_2 FILLER_9_1931 ();
 sg13g2_decap_4 FILLER_9_1942 ();
 sg13g2_decap_8 FILLER_9_1964 ();
 sg13g2_fill_2 FILLER_9_1971 ();
 sg13g2_fill_1 FILLER_9_1973 ();
 sg13g2_decap_8 FILLER_9_1989 ();
 sg13g2_fill_1 FILLER_9_1996 ();
 sg13g2_decap_4 FILLER_9_2011 ();
 sg13g2_fill_2 FILLER_9_2015 ();
 sg13g2_decap_4 FILLER_9_2024 ();
 sg13g2_fill_1 FILLER_9_2028 ();
 sg13g2_fill_1 FILLER_9_2037 ();
 sg13g2_fill_1 FILLER_9_2055 ();
 sg13g2_fill_2 FILLER_9_2072 ();
 sg13g2_fill_1 FILLER_9_2074 ();
 sg13g2_decap_8 FILLER_9_2089 ();
 sg13g2_decap_8 FILLER_9_2096 ();
 sg13g2_fill_1 FILLER_9_2103 ();
 sg13g2_decap_8 FILLER_9_2111 ();
 sg13g2_fill_1 FILLER_9_2118 ();
 sg13g2_fill_2 FILLER_9_2125 ();
 sg13g2_decap_4 FILLER_9_2145 ();
 sg13g2_fill_2 FILLER_9_2149 ();
 sg13g2_decap_8 FILLER_9_2179 ();
 sg13g2_decap_4 FILLER_9_2186 ();
 sg13g2_fill_1 FILLER_9_2209 ();
 sg13g2_fill_2 FILLER_9_2225 ();
 sg13g2_fill_1 FILLER_9_2227 ();
 sg13g2_fill_2 FILLER_9_2247 ();
 sg13g2_fill_2 FILLER_9_2259 ();
 sg13g2_fill_2 FILLER_9_2265 ();
 sg13g2_fill_1 FILLER_9_2267 ();
 sg13g2_fill_2 FILLER_9_2289 ();
 sg13g2_fill_1 FILLER_9_2291 ();
 sg13g2_decap_4 FILLER_9_2312 ();
 sg13g2_fill_2 FILLER_9_2316 ();
 sg13g2_fill_2 FILLER_9_2336 ();
 sg13g2_fill_2 FILLER_9_2356 ();
 sg13g2_fill_2 FILLER_9_2368 ();
 sg13g2_decap_4 FILLER_9_2395 ();
 sg13g2_fill_1 FILLER_9_2399 ();
 sg13g2_decap_8 FILLER_9_2413 ();
 sg13g2_decap_8 FILLER_9_2420 ();
 sg13g2_fill_2 FILLER_9_2427 ();
 sg13g2_decap_4 FILLER_9_2438 ();
 sg13g2_fill_1 FILLER_9_2442 ();
 sg13g2_fill_2 FILLER_9_2469 ();
 sg13g2_fill_2 FILLER_9_2493 ();
 sg13g2_fill_1 FILLER_9_2495 ();
 sg13g2_fill_2 FILLER_9_2508 ();
 sg13g2_fill_1 FILLER_9_2510 ();
 sg13g2_decap_8 FILLER_9_2570 ();
 sg13g2_fill_2 FILLER_9_2587 ();
 sg13g2_fill_1 FILLER_9_2589 ();
 sg13g2_decap_8 FILLER_9_2599 ();
 sg13g2_fill_1 FILLER_9_2610 ();
 sg13g2_fill_1 FILLER_9_2615 ();
 sg13g2_fill_2 FILLER_9_2625 ();
 sg13g2_fill_1 FILLER_9_2627 ();
 sg13g2_decap_4 FILLER_9_2642 ();
 sg13g2_fill_2 FILLER_9_2646 ();
 sg13g2_fill_1 FILLER_9_2668 ();
 sg13g2_fill_1 FILLER_9_2702 ();
 sg13g2_fill_1 FILLER_9_2716 ();
 sg13g2_fill_1 FILLER_9_2730 ();
 sg13g2_fill_2 FILLER_9_2739 ();
 sg13g2_fill_1 FILLER_9_2741 ();
 sg13g2_fill_2 FILLER_9_2763 ();
 sg13g2_fill_1 FILLER_9_2765 ();
 sg13g2_decap_8 FILLER_9_2783 ();
 sg13g2_fill_2 FILLER_9_2790 ();
 sg13g2_fill_2 FILLER_9_2797 ();
 sg13g2_fill_2 FILLER_9_2809 ();
 sg13g2_fill_2 FILLER_9_2825 ();
 sg13g2_fill_1 FILLER_9_2827 ();
 sg13g2_fill_2 FILLER_9_2833 ();
 sg13g2_fill_1 FILLER_9_2835 ();
 sg13g2_fill_2 FILLER_9_2846 ();
 sg13g2_fill_1 FILLER_9_2848 ();
 sg13g2_fill_1 FILLER_9_2865 ();
 sg13g2_fill_2 FILLER_9_2887 ();
 sg13g2_fill_1 FILLER_9_2889 ();
 sg13g2_fill_1 FILLER_9_2923 ();
 sg13g2_decap_8 FILLER_9_2938 ();
 sg13g2_decap_8 FILLER_9_2945 ();
 sg13g2_decap_8 FILLER_9_2960 ();
 sg13g2_decap_4 FILLER_9_2967 ();
 sg13g2_fill_2 FILLER_9_2971 ();
 sg13g2_decap_4 FILLER_9_2981 ();
 sg13g2_fill_2 FILLER_9_2985 ();
 sg13g2_fill_1 FILLER_9_2992 ();
 sg13g2_decap_8 FILLER_9_3001 ();
 sg13g2_fill_2 FILLER_9_3008 ();
 sg13g2_fill_1 FILLER_9_3017 ();
 sg13g2_decap_4 FILLER_9_3026 ();
 sg13g2_fill_2 FILLER_9_3030 ();
 sg13g2_decap_8 FILLER_9_3045 ();
 sg13g2_fill_2 FILLER_9_3052 ();
 sg13g2_fill_1 FILLER_9_3054 ();
 sg13g2_fill_1 FILLER_9_3066 ();
 sg13g2_fill_2 FILLER_9_3088 ();
 sg13g2_fill_1 FILLER_9_3090 ();
 sg13g2_decap_8 FILLER_9_3096 ();
 sg13g2_decap_8 FILLER_9_3115 ();
 sg13g2_decap_4 FILLER_9_3138 ();
 sg13g2_fill_1 FILLER_9_3142 ();
 sg13g2_fill_1 FILLER_9_3148 ();
 sg13g2_fill_2 FILLER_9_3154 ();
 sg13g2_fill_1 FILLER_9_3160 ();
 sg13g2_decap_8 FILLER_9_3169 ();
 sg13g2_decap_4 FILLER_9_3176 ();
 sg13g2_decap_4 FILLER_9_3202 ();
 sg13g2_fill_1 FILLER_9_3206 ();
 sg13g2_fill_2 FILLER_9_3236 ();
 sg13g2_decap_4 FILLER_9_3270 ();
 sg13g2_fill_1 FILLER_9_3274 ();
 sg13g2_decap_4 FILLER_9_3279 ();
 sg13g2_fill_2 FILLER_9_3283 ();
 sg13g2_decap_4 FILLER_9_3292 ();
 sg13g2_fill_2 FILLER_9_3296 ();
 sg13g2_decap_4 FILLER_9_3311 ();
 sg13g2_fill_2 FILLER_9_3333 ();
 sg13g2_decap_8 FILLER_9_3340 ();
 sg13g2_fill_2 FILLER_9_3347 ();
 sg13g2_fill_1 FILLER_9_3355 ();
 sg13g2_fill_2 FILLER_9_3373 ();
 sg13g2_fill_1 FILLER_9_3375 ();
 sg13g2_decap_8 FILLER_9_3383 ();
 sg13g2_decap_8 FILLER_9_3390 ();
 sg13g2_fill_2 FILLER_9_3412 ();
 sg13g2_fill_1 FILLER_9_3429 ();
 sg13g2_fill_2 FILLER_9_3442 ();
 sg13g2_fill_1 FILLER_9_3444 ();
 sg13g2_decap_8 FILLER_9_3450 ();
 sg13g2_fill_1 FILLER_9_3457 ();
 sg13g2_fill_2 FILLER_9_3467 ();
 sg13g2_fill_1 FILLER_9_3469 ();
 sg13g2_decap_8 FILLER_9_3483 ();
 sg13g2_decap_8 FILLER_9_3490 ();
 sg13g2_fill_1 FILLER_9_3497 ();
 sg13g2_decap_8 FILLER_9_3533 ();
 sg13g2_decap_8 FILLER_9_3540 ();
 sg13g2_decap_8 FILLER_9_3547 ();
 sg13g2_decap_8 FILLER_9_3554 ();
 sg13g2_decap_8 FILLER_9_3561 ();
 sg13g2_decap_8 FILLER_9_3568 ();
 sg13g2_decap_4 FILLER_9_3575 ();
 sg13g2_fill_1 FILLER_9_3579 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_120 ();
 sg13g2_decap_4 FILLER_10_127 ();
 sg13g2_fill_1 FILLER_10_131 ();
 sg13g2_fill_1 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_146 ();
 sg13g2_decap_4 FILLER_10_162 ();
 sg13g2_fill_2 FILLER_10_183 ();
 sg13g2_fill_1 FILLER_10_185 ();
 sg13g2_decap_8 FILLER_10_199 ();
 sg13g2_fill_1 FILLER_10_206 ();
 sg13g2_decap_8 FILLER_10_230 ();
 sg13g2_fill_2 FILLER_10_237 ();
 sg13g2_fill_1 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_fill_2 FILLER_10_266 ();
 sg13g2_fill_2 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_326 ();
 sg13g2_decap_4 FILLER_10_341 ();
 sg13g2_fill_2 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_4 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_fill_2 FILLER_10_395 ();
 sg13g2_decap_4 FILLER_10_402 ();
 sg13g2_fill_2 FILLER_10_410 ();
 sg13g2_fill_1 FILLER_10_412 ();
 sg13g2_decap_4 FILLER_10_419 ();
 sg13g2_fill_1 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_4 FILLER_10_448 ();
 sg13g2_fill_1 FILLER_10_452 ();
 sg13g2_fill_2 FILLER_10_490 ();
 sg13g2_decap_4 FILLER_10_496 ();
 sg13g2_fill_1 FILLER_10_500 ();
 sg13g2_fill_2 FILLER_10_522 ();
 sg13g2_fill_2 FILLER_10_532 ();
 sg13g2_fill_1 FILLER_10_534 ();
 sg13g2_fill_1 FILLER_10_551 ();
 sg13g2_fill_2 FILLER_10_569 ();
 sg13g2_fill_1 FILLER_10_589 ();
 sg13g2_fill_2 FILLER_10_618 ();
 sg13g2_fill_1 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_643 ();
 sg13g2_fill_1 FILLER_10_650 ();
 sg13g2_fill_2 FILLER_10_677 ();
 sg13g2_decap_4 FILLER_10_702 ();
 sg13g2_fill_2 FILLER_10_706 ();
 sg13g2_decap_4 FILLER_10_718 ();
 sg13g2_fill_2 FILLER_10_722 ();
 sg13g2_decap_4 FILLER_10_737 ();
 sg13g2_decap_8 FILLER_10_745 ();
 sg13g2_decap_4 FILLER_10_752 ();
 sg13g2_fill_2 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_771 ();
 sg13g2_decap_4 FILLER_10_778 ();
 sg13g2_fill_1 FILLER_10_782 ();
 sg13g2_fill_2 FILLER_10_793 ();
 sg13g2_fill_2 FILLER_10_815 ();
 sg13g2_fill_2 FILLER_10_827 ();
 sg13g2_fill_1 FILLER_10_829 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_fill_2 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_910 ();
 sg13g2_decap_4 FILLER_10_917 ();
 sg13g2_fill_2 FILLER_10_947 ();
 sg13g2_fill_2 FILLER_10_954 ();
 sg13g2_fill_1 FILLER_10_956 ();
 sg13g2_decap_8 FILLER_10_967 ();
 sg13g2_fill_1 FILLER_10_974 ();
 sg13g2_fill_2 FILLER_10_990 ();
 sg13g2_fill_1 FILLER_10_992 ();
 sg13g2_decap_4 FILLER_10_1016 ();
 sg13g2_fill_1 FILLER_10_1024 ();
 sg13g2_fill_2 FILLER_10_1029 ();
 sg13g2_fill_2 FILLER_10_1053 ();
 sg13g2_fill_1 FILLER_10_1055 ();
 sg13g2_decap_4 FILLER_10_1082 ();
 sg13g2_fill_1 FILLER_10_1086 ();
 sg13g2_fill_2 FILLER_10_1091 ();
 sg13g2_decap_4 FILLER_10_1106 ();
 sg13g2_fill_1 FILLER_10_1110 ();
 sg13g2_fill_2 FILLER_10_1124 ();
 sg13g2_fill_1 FILLER_10_1126 ();
 sg13g2_fill_2 FILLER_10_1136 ();
 sg13g2_fill_2 FILLER_10_1161 ();
 sg13g2_fill_1 FILLER_10_1163 ();
 sg13g2_fill_2 FILLER_10_1169 ();
 sg13g2_fill_1 FILLER_10_1171 ();
 sg13g2_decap_8 FILLER_10_1187 ();
 sg13g2_decap_8 FILLER_10_1194 ();
 sg13g2_decap_8 FILLER_10_1201 ();
 sg13g2_decap_4 FILLER_10_1208 ();
 sg13g2_fill_2 FILLER_10_1212 ();
 sg13g2_decap_4 FILLER_10_1227 ();
 sg13g2_fill_1 FILLER_10_1249 ();
 sg13g2_fill_1 FILLER_10_1255 ();
 sg13g2_decap_4 FILLER_10_1261 ();
 sg13g2_decap_8 FILLER_10_1273 ();
 sg13g2_decap_4 FILLER_10_1280 ();
 sg13g2_fill_2 FILLER_10_1284 ();
 sg13g2_decap_8 FILLER_10_1301 ();
 sg13g2_fill_2 FILLER_10_1308 ();
 sg13g2_decap_8 FILLER_10_1319 ();
 sg13g2_fill_2 FILLER_10_1326 ();
 sg13g2_fill_1 FILLER_10_1328 ();
 sg13g2_fill_1 FILLER_10_1342 ();
 sg13g2_decap_8 FILLER_10_1356 ();
 sg13g2_decap_8 FILLER_10_1363 ();
 sg13g2_decap_4 FILLER_10_1370 ();
 sg13g2_fill_2 FILLER_10_1374 ();
 sg13g2_fill_1 FILLER_10_1381 ();
 sg13g2_decap_4 FILLER_10_1387 ();
 sg13g2_fill_2 FILLER_10_1396 ();
 sg13g2_fill_1 FILLER_10_1411 ();
 sg13g2_decap_8 FILLER_10_1416 ();
 sg13g2_decap_8 FILLER_10_1423 ();
 sg13g2_decap_8 FILLER_10_1430 ();
 sg13g2_decap_8 FILLER_10_1463 ();
 sg13g2_fill_1 FILLER_10_1470 ();
 sg13g2_fill_2 FILLER_10_1491 ();
 sg13g2_fill_2 FILLER_10_1502 ();
 sg13g2_fill_1 FILLER_10_1512 ();
 sg13g2_decap_8 FILLER_10_1526 ();
 sg13g2_fill_1 FILLER_10_1553 ();
 sg13g2_fill_1 FILLER_10_1574 ();
 sg13g2_fill_2 FILLER_10_1579 ();
 sg13g2_fill_2 FILLER_10_1594 ();
 sg13g2_decap_8 FILLER_10_1614 ();
 sg13g2_decap_8 FILLER_10_1621 ();
 sg13g2_fill_2 FILLER_10_1628 ();
 sg13g2_fill_1 FILLER_10_1630 ();
 sg13g2_fill_2 FILLER_10_1639 ();
 sg13g2_decap_8 FILLER_10_1662 ();
 sg13g2_decap_4 FILLER_10_1669 ();
 sg13g2_fill_1 FILLER_10_1673 ();
 sg13g2_fill_2 FILLER_10_1690 ();
 sg13g2_fill_2 FILLER_10_1697 ();
 sg13g2_fill_1 FILLER_10_1699 ();
 sg13g2_decap_8 FILLER_10_1727 ();
 sg13g2_decap_8 FILLER_10_1741 ();
 sg13g2_fill_2 FILLER_10_1748 ();
 sg13g2_fill_1 FILLER_10_1750 ();
 sg13g2_fill_2 FILLER_10_1762 ();
 sg13g2_fill_1 FILLER_10_1764 ();
 sg13g2_decap_8 FILLER_10_1785 ();
 sg13g2_decap_8 FILLER_10_1792 ();
 sg13g2_decap_8 FILLER_10_1799 ();
 sg13g2_decap_4 FILLER_10_1833 ();
 sg13g2_decap_8 FILLER_10_1845 ();
 sg13g2_fill_1 FILLER_10_1852 ();
 sg13g2_decap_8 FILLER_10_1869 ();
 sg13g2_decap_8 FILLER_10_1880 ();
 sg13g2_fill_2 FILLER_10_1906 ();
 sg13g2_fill_1 FILLER_10_1916 ();
 sg13g2_fill_2 FILLER_10_1930 ();
 sg13g2_fill_1 FILLER_10_1932 ();
 sg13g2_fill_2 FILLER_10_1942 ();
 sg13g2_fill_1 FILLER_10_1944 ();
 sg13g2_fill_2 FILLER_10_1962 ();
 sg13g2_fill_1 FILLER_10_1964 ();
 sg13g2_decap_8 FILLER_10_2017 ();
 sg13g2_decap_8 FILLER_10_2024 ();
 sg13g2_decap_8 FILLER_10_2040 ();
 sg13g2_decap_4 FILLER_10_2047 ();
 sg13g2_fill_1 FILLER_10_2056 ();
 sg13g2_fill_2 FILLER_10_2061 ();
 sg13g2_fill_1 FILLER_10_2063 ();
 sg13g2_fill_1 FILLER_10_2084 ();
 sg13g2_decap_8 FILLER_10_2113 ();
 sg13g2_decap_4 FILLER_10_2120 ();
 sg13g2_decap_8 FILLER_10_2137 ();
 sg13g2_decap_8 FILLER_10_2144 ();
 sg13g2_decap_4 FILLER_10_2151 ();
 sg13g2_fill_1 FILLER_10_2155 ();
 sg13g2_decap_4 FILLER_10_2160 ();
 sg13g2_decap_8 FILLER_10_2174 ();
 sg13g2_decap_4 FILLER_10_2181 ();
 sg13g2_fill_2 FILLER_10_2198 ();
 sg13g2_decap_4 FILLER_10_2239 ();
 sg13g2_fill_1 FILLER_10_2253 ();
 sg13g2_fill_1 FILLER_10_2269 ();
 sg13g2_decap_8 FILLER_10_2288 ();
 sg13g2_fill_1 FILLER_10_2311 ();
 sg13g2_fill_2 FILLER_10_2329 ();
 sg13g2_fill_1 FILLER_10_2331 ();
 sg13g2_fill_2 FILLER_10_2345 ();
 sg13g2_fill_2 FILLER_10_2350 ();
 sg13g2_decap_8 FILLER_10_2356 ();
 sg13g2_fill_2 FILLER_10_2363 ();
 sg13g2_fill_2 FILLER_10_2388 ();
 sg13g2_fill_1 FILLER_10_2390 ();
 sg13g2_fill_2 FILLER_10_2397 ();
 sg13g2_fill_1 FILLER_10_2399 ();
 sg13g2_decap_4 FILLER_10_2408 ();
 sg13g2_fill_1 FILLER_10_2412 ();
 sg13g2_decap_8 FILLER_10_2427 ();
 sg13g2_fill_2 FILLER_10_2434 ();
 sg13g2_decap_8 FILLER_10_2444 ();
 sg13g2_decap_4 FILLER_10_2451 ();
 sg13g2_fill_1 FILLER_10_2455 ();
 sg13g2_fill_2 FILLER_10_2475 ();
 sg13g2_fill_2 FILLER_10_2502 ();
 sg13g2_decap_4 FILLER_10_2524 ();
 sg13g2_fill_2 FILLER_10_2533 ();
 sg13g2_decap_4 FILLER_10_2545 ();
 sg13g2_fill_1 FILLER_10_2549 ();
 sg13g2_decap_8 FILLER_10_2561 ();
 sg13g2_fill_2 FILLER_10_2568 ();
 sg13g2_fill_1 FILLER_10_2590 ();
 sg13g2_decap_8 FILLER_10_2600 ();
 sg13g2_fill_2 FILLER_10_2607 ();
 sg13g2_fill_1 FILLER_10_2623 ();
 sg13g2_fill_1 FILLER_10_2628 ();
 sg13g2_decap_8 FILLER_10_2634 ();
 sg13g2_fill_1 FILLER_10_2641 ();
 sg13g2_fill_1 FILLER_10_2655 ();
 sg13g2_fill_1 FILLER_10_2661 ();
 sg13g2_decap_4 FILLER_10_2704 ();
 sg13g2_decap_4 FILLER_10_2738 ();
 sg13g2_fill_2 FILLER_10_2742 ();
 sg13g2_fill_2 FILLER_10_2758 ();
 sg13g2_fill_1 FILLER_10_2760 ();
 sg13g2_fill_2 FILLER_10_2781 ();
 sg13g2_fill_2 FILLER_10_2833 ();
 sg13g2_fill_1 FILLER_10_2835 ();
 sg13g2_fill_2 FILLER_10_2841 ();
 sg13g2_fill_1 FILLER_10_2843 ();
 sg13g2_fill_2 FILLER_10_2849 ();
 sg13g2_fill_1 FILLER_10_2851 ();
 sg13g2_fill_2 FILLER_10_2860 ();
 sg13g2_fill_2 FILLER_10_2872 ();
 sg13g2_fill_1 FILLER_10_2874 ();
 sg13g2_decap_8 FILLER_10_2888 ();
 sg13g2_decap_8 FILLER_10_2913 ();
 sg13g2_fill_2 FILLER_10_2920 ();
 sg13g2_fill_1 FILLER_10_2922 ();
 sg13g2_fill_2 FILLER_10_2936 ();
 sg13g2_fill_1 FILLER_10_2938 ();
 sg13g2_fill_2 FILLER_10_2943 ();
 sg13g2_fill_1 FILLER_10_2965 ();
 sg13g2_decap_8 FILLER_10_2971 ();
 sg13g2_decap_4 FILLER_10_2978 ();
 sg13g2_fill_1 FILLER_10_2982 ();
 sg13g2_decap_4 FILLER_10_3002 ();
 sg13g2_decap_4 FILLER_10_3049 ();
 sg13g2_fill_2 FILLER_10_3053 ();
 sg13g2_decap_8 FILLER_10_3071 ();
 sg13g2_fill_2 FILLER_10_3078 ();
 sg13g2_fill_1 FILLER_10_3080 ();
 sg13g2_fill_2 FILLER_10_3091 ();
 sg13g2_decap_8 FILLER_10_3122 ();
 sg13g2_fill_2 FILLER_10_3129 ();
 sg13g2_fill_1 FILLER_10_3131 ();
 sg13g2_fill_2 FILLER_10_3141 ();
 sg13g2_fill_1 FILLER_10_3143 ();
 sg13g2_fill_2 FILLER_10_3152 ();
 sg13g2_decap_4 FILLER_10_3172 ();
 sg13g2_fill_2 FILLER_10_3181 ();
 sg13g2_fill_1 FILLER_10_3183 ();
 sg13g2_fill_2 FILLER_10_3189 ();
 sg13g2_fill_2 FILLER_10_3209 ();
 sg13g2_decap_4 FILLER_10_3219 ();
 sg13g2_fill_2 FILLER_10_3231 ();
 sg13g2_fill_1 FILLER_10_3233 ();
 sg13g2_fill_2 FILLER_10_3238 ();
 sg13g2_fill_1 FILLER_10_3240 ();
 sg13g2_fill_1 FILLER_10_3263 ();
 sg13g2_decap_8 FILLER_10_3305 ();
 sg13g2_fill_1 FILLER_10_3317 ();
 sg13g2_decap_8 FILLER_10_3330 ();
 sg13g2_decap_8 FILLER_10_3354 ();
 sg13g2_fill_2 FILLER_10_3361 ();
 sg13g2_fill_2 FILLER_10_3368 ();
 sg13g2_decap_8 FILLER_10_3380 ();
 sg13g2_decap_4 FILLER_10_3400 ();
 sg13g2_decap_8 FILLER_10_3422 ();
 sg13g2_fill_2 FILLER_10_3429 ();
 sg13g2_fill_2 FILLER_10_3454 ();
 sg13g2_fill_1 FILLER_10_3456 ();
 sg13g2_decap_4 FILLER_10_3481 ();
 sg13g2_fill_2 FILLER_10_3485 ();
 sg13g2_decap_4 FILLER_10_3492 ();
 sg13g2_fill_2 FILLER_10_3496 ();
 sg13g2_fill_1 FILLER_10_3507 ();
 sg13g2_decap_8 FILLER_10_3517 ();
 sg13g2_decap_4 FILLER_10_3524 ();
 sg13g2_decap_8 FILLER_10_3537 ();
 sg13g2_decap_8 FILLER_10_3544 ();
 sg13g2_decap_8 FILLER_10_3551 ();
 sg13g2_decap_8 FILLER_10_3558 ();
 sg13g2_decap_8 FILLER_10_3565 ();
 sg13g2_decap_8 FILLER_10_3572 ();
 sg13g2_fill_1 FILLER_10_3579 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_fill_2 FILLER_11_86 ();
 sg13g2_fill_2 FILLER_11_96 ();
 sg13g2_fill_1 FILLER_11_98 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_146 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_4 FILLER_11_177 ();
 sg13g2_decap_4 FILLER_11_186 ();
 sg13g2_fill_1 FILLER_11_195 ();
 sg13g2_fill_2 FILLER_11_200 ();
 sg13g2_fill_2 FILLER_11_215 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_fill_2 FILLER_11_254 ();
 sg13g2_decap_8 FILLER_11_260 ();
 sg13g2_fill_2 FILLER_11_267 ();
 sg13g2_decap_4 FILLER_11_277 ();
 sg13g2_fill_2 FILLER_11_281 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_fill_2 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_4 FILLER_11_345 ();
 sg13g2_fill_2 FILLER_11_349 ();
 sg13g2_fill_2 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_4 FILLER_11_396 ();
 sg13g2_fill_1 FILLER_11_400 ();
 sg13g2_fill_1 FILLER_11_446 ();
 sg13g2_fill_2 FILLER_11_452 ();
 sg13g2_fill_1 FILLER_11_454 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_fill_1 FILLER_11_466 ();
 sg13g2_fill_1 FILLER_11_471 ();
 sg13g2_decap_4 FILLER_11_481 ();
 sg13g2_fill_2 FILLER_11_485 ();
 sg13g2_decap_8 FILLER_11_515 ();
 sg13g2_fill_1 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_536 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_fill_1 FILLER_11_581 ();
 sg13g2_fill_2 FILLER_11_591 ();
 sg13g2_fill_1 FILLER_11_593 ();
 sg13g2_fill_2 FILLER_11_615 ();
 sg13g2_fill_1 FILLER_11_617 ();
 sg13g2_fill_2 FILLER_11_640 ();
 sg13g2_fill_1 FILLER_11_642 ();
 sg13g2_fill_1 FILLER_11_675 ();
 sg13g2_fill_2 FILLER_11_681 ();
 sg13g2_decap_8 FILLER_11_691 ();
 sg13g2_fill_2 FILLER_11_698 ();
 sg13g2_fill_1 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_724 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_fill_1 FILLER_11_756 ();
 sg13g2_fill_2 FILLER_11_794 ();
 sg13g2_decap_4 FILLER_11_821 ();
 sg13g2_fill_1 FILLER_11_848 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_decap_4 FILLER_11_861 ();
 sg13g2_fill_2 FILLER_11_881 ();
 sg13g2_fill_2 FILLER_11_909 ();
 sg13g2_fill_2 FILLER_11_933 ();
 sg13g2_fill_1 FILLER_11_935 ();
 sg13g2_decap_4 FILLER_11_948 ();
 sg13g2_decap_4 FILLER_11_976 ();
 sg13g2_fill_2 FILLER_11_980 ();
 sg13g2_fill_2 FILLER_11_1020 ();
 sg13g2_fill_2 FILLER_11_1042 ();
 sg13g2_decap_4 FILLER_11_1056 ();
 sg13g2_fill_1 FILLER_11_1060 ();
 sg13g2_decap_8 FILLER_11_1077 ();
 sg13g2_fill_2 FILLER_11_1084 ();
 sg13g2_fill_1 FILLER_11_1086 ();
 sg13g2_fill_2 FILLER_11_1113 ();
 sg13g2_fill_1 FILLER_11_1115 ();
 sg13g2_decap_8 FILLER_11_1126 ();
 sg13g2_fill_1 FILLER_11_1133 ();
 sg13g2_fill_2 FILLER_11_1158 ();
 sg13g2_fill_1 FILLER_11_1160 ();
 sg13g2_decap_4 FILLER_11_1198 ();
 sg13g2_fill_1 FILLER_11_1202 ();
 sg13g2_fill_2 FILLER_11_1227 ();
 sg13g2_fill_1 FILLER_11_1229 ();
 sg13g2_fill_2 FILLER_11_1245 ();
 sg13g2_decap_4 FILLER_11_1275 ();
 sg13g2_fill_2 FILLER_11_1279 ();
 sg13g2_decap_8 FILLER_11_1306 ();
 sg13g2_decap_8 FILLER_11_1313 ();
 sg13g2_decap_4 FILLER_11_1320 ();
 sg13g2_decap_8 FILLER_11_1337 ();
 sg13g2_fill_1 FILLER_11_1344 ();
 sg13g2_decap_4 FILLER_11_1354 ();
 sg13g2_fill_2 FILLER_11_1358 ();
 sg13g2_fill_2 FILLER_11_1395 ();
 sg13g2_fill_1 FILLER_11_1397 ();
 sg13g2_decap_4 FILLER_11_1435 ();
 sg13g2_fill_2 FILLER_11_1439 ();
 sg13g2_decap_8 FILLER_11_1459 ();
 sg13g2_fill_2 FILLER_11_1466 ();
 sg13g2_decap_4 FILLER_11_1472 ();
 sg13g2_fill_1 FILLER_11_1476 ();
 sg13g2_decap_4 FILLER_11_1508 ();
 sg13g2_decap_8 FILLER_11_1520 ();
 sg13g2_fill_2 FILLER_11_1544 ();
 sg13g2_fill_2 FILLER_11_1554 ();
 sg13g2_fill_2 FILLER_11_1565 ();
 sg13g2_fill_2 FILLER_11_1585 ();
 sg13g2_fill_1 FILLER_11_1587 ();
 sg13g2_decap_8 FILLER_11_1596 ();
 sg13g2_fill_2 FILLER_11_1603 ();
 sg13g2_fill_2 FILLER_11_1613 ();
 sg13g2_decap_4 FILLER_11_1646 ();
 sg13g2_fill_2 FILLER_11_1663 ();
 sg13g2_decap_8 FILLER_11_1678 ();
 sg13g2_fill_2 FILLER_11_1691 ();
 sg13g2_fill_1 FILLER_11_1693 ();
 sg13g2_fill_1 FILLER_11_1714 ();
 sg13g2_fill_2 FILLER_11_1725 ();
 sg13g2_fill_1 FILLER_11_1759 ();
 sg13g2_fill_2 FILLER_11_1791 ();
 sg13g2_fill_1 FILLER_11_1793 ();
 sg13g2_fill_2 FILLER_11_1799 ();
 sg13g2_decap_8 FILLER_11_1824 ();
 sg13g2_decap_8 FILLER_11_1831 ();
 sg13g2_decap_4 FILLER_11_1838 ();
 sg13g2_fill_1 FILLER_11_1842 ();
 sg13g2_decap_8 FILLER_11_1856 ();
 sg13g2_decap_4 FILLER_11_1863 ();
 sg13g2_decap_8 FILLER_11_1884 ();
 sg13g2_decap_8 FILLER_11_1904 ();
 sg13g2_fill_1 FILLER_11_1911 ();
 sg13g2_fill_1 FILLER_11_1917 ();
 sg13g2_decap_8 FILLER_11_1925 ();
 sg13g2_fill_1 FILLER_11_1932 ();
 sg13g2_decap_8 FILLER_11_1962 ();
 sg13g2_fill_2 FILLER_11_1969 ();
 sg13g2_decap_8 FILLER_11_1983 ();
 sg13g2_decap_8 FILLER_11_1990 ();
 sg13g2_fill_2 FILLER_11_1997 ();
 sg13g2_fill_1 FILLER_11_1999 ();
 sg13g2_fill_1 FILLER_11_2028 ();
 sg13g2_fill_2 FILLER_11_2049 ();
 sg13g2_fill_2 FILLER_11_2068 ();
 sg13g2_fill_1 FILLER_11_2070 ();
 sg13g2_fill_2 FILLER_11_2080 ();
 sg13g2_fill_2 FILLER_11_2100 ();
 sg13g2_fill_1 FILLER_11_2102 ();
 sg13g2_fill_2 FILLER_11_2116 ();
 sg13g2_fill_1 FILLER_11_2146 ();
 sg13g2_decap_4 FILLER_11_2181 ();
 sg13g2_fill_2 FILLER_11_2195 ();
 sg13g2_fill_1 FILLER_11_2197 ();
 sg13g2_decap_8 FILLER_11_2210 ();
 sg13g2_decap_4 FILLER_11_2235 ();
 sg13g2_fill_2 FILLER_11_2239 ();
 sg13g2_fill_1 FILLER_11_2249 ();
 sg13g2_decap_8 FILLER_11_2283 ();
 sg13g2_decap_4 FILLER_11_2290 ();
 sg13g2_fill_2 FILLER_11_2294 ();
 sg13g2_fill_2 FILLER_11_2304 ();
 sg13g2_fill_1 FILLER_11_2306 ();
 sg13g2_fill_1 FILLER_11_2320 ();
 sg13g2_fill_2 FILLER_11_2343 ();
 sg13g2_decap_8 FILLER_11_2354 ();
 sg13g2_decap_8 FILLER_11_2361 ();
 sg13g2_decap_4 FILLER_11_2368 ();
 sg13g2_fill_2 FILLER_11_2389 ();
 sg13g2_decap_8 FILLER_11_2406 ();
 sg13g2_decap_4 FILLER_11_2441 ();
 sg13g2_fill_1 FILLER_11_2445 ();
 sg13g2_fill_2 FILLER_11_2471 ();
 sg13g2_decap_8 FILLER_11_2487 ();
 sg13g2_decap_8 FILLER_11_2494 ();
 sg13g2_fill_1 FILLER_11_2501 ();
 sg13g2_fill_2 FILLER_11_2516 ();
 sg13g2_fill_1 FILLER_11_2518 ();
 sg13g2_fill_2 FILLER_11_2558 ();
 sg13g2_fill_1 FILLER_11_2560 ();
 sg13g2_fill_1 FILLER_11_2569 ();
 sg13g2_decap_8 FILLER_11_2583 ();
 sg13g2_fill_2 FILLER_11_2610 ();
 sg13g2_fill_1 FILLER_11_2612 ();
 sg13g2_fill_1 FILLER_11_2618 ();
 sg13g2_fill_2 FILLER_11_2651 ();
 sg13g2_fill_2 FILLER_11_2658 ();
 sg13g2_fill_1 FILLER_11_2666 ();
 sg13g2_decap_8 FILLER_11_2688 ();
 sg13g2_fill_2 FILLER_11_2695 ();
 sg13g2_decap_8 FILLER_11_2706 ();
 sg13g2_decap_4 FILLER_11_2713 ();
 sg13g2_fill_2 FILLER_11_2717 ();
 sg13g2_decap_4 FILLER_11_2729 ();
 sg13g2_fill_1 FILLER_11_2733 ();
 sg13g2_fill_2 FILLER_11_2738 ();
 sg13g2_decap_4 FILLER_11_2758 ();
 sg13g2_fill_1 FILLER_11_2762 ();
 sg13g2_decap_8 FILLER_11_2781 ();
 sg13g2_fill_2 FILLER_11_2788 ();
 sg13g2_fill_2 FILLER_11_2807 ();
 sg13g2_fill_1 FILLER_11_2814 ();
 sg13g2_fill_1 FILLER_11_2823 ();
 sg13g2_fill_1 FILLER_11_2832 ();
 sg13g2_decap_8 FILLER_11_2838 ();
 sg13g2_decap_8 FILLER_11_2845 ();
 sg13g2_fill_2 FILLER_11_2852 ();
 sg13g2_fill_1 FILLER_11_2858 ();
 sg13g2_fill_1 FILLER_11_2863 ();
 sg13g2_decap_8 FILLER_11_2890 ();
 sg13g2_fill_1 FILLER_11_2897 ();
 sg13g2_decap_4 FILLER_11_2903 ();
 sg13g2_fill_1 FILLER_11_2907 ();
 sg13g2_decap_8 FILLER_11_2913 ();
 sg13g2_fill_2 FILLER_11_2920 ();
 sg13g2_decap_4 FILLER_11_2932 ();
 sg13g2_decap_8 FILLER_11_2945 ();
 sg13g2_fill_2 FILLER_11_2952 ();
 sg13g2_fill_2 FILLER_11_2959 ();
 sg13g2_fill_1 FILLER_11_2961 ();
 sg13g2_decap_4 FILLER_11_2974 ();
 sg13g2_fill_1 FILLER_11_2984 ();
 sg13g2_decap_8 FILLER_11_2994 ();
 sg13g2_fill_2 FILLER_11_3001 ();
 sg13g2_fill_1 FILLER_11_3003 ();
 sg13g2_fill_2 FILLER_11_3027 ();
 sg13g2_fill_2 FILLER_11_3047 ();
 sg13g2_fill_1 FILLER_11_3049 ();
 sg13g2_decap_4 FILLER_11_3063 ();
 sg13g2_fill_1 FILLER_11_3067 ();
 sg13g2_fill_2 FILLER_11_3072 ();
 sg13g2_fill_1 FILLER_11_3094 ();
 sg13g2_decap_4 FILLER_11_3103 ();
 sg13g2_fill_1 FILLER_11_3110 ();
 sg13g2_decap_8 FILLER_11_3121 ();
 sg13g2_decap_4 FILLER_11_3128 ();
 sg13g2_fill_2 FILLER_11_3132 ();
 sg13g2_decap_8 FILLER_11_3150 ();
 sg13g2_fill_1 FILLER_11_3157 ();
 sg13g2_decap_8 FILLER_11_3175 ();
 sg13g2_fill_2 FILLER_11_3182 ();
 sg13g2_fill_1 FILLER_11_3184 ();
 sg13g2_decap_8 FILLER_11_3206 ();
 sg13g2_fill_1 FILLER_11_3213 ();
 sg13g2_fill_2 FILLER_11_3239 ();
 sg13g2_fill_1 FILLER_11_3241 ();
 sg13g2_decap_8 FILLER_11_3270 ();
 sg13g2_decap_4 FILLER_11_3277 ();
 sg13g2_fill_1 FILLER_11_3281 ();
 sg13g2_decap_4 FILLER_11_3313 ();
 sg13g2_fill_2 FILLER_11_3330 ();
 sg13g2_decap_8 FILLER_11_3349 ();
 sg13g2_fill_2 FILLER_11_3356 ();
 sg13g2_fill_1 FILLER_11_3358 ();
 sg13g2_decap_4 FILLER_11_3379 ();
 sg13g2_fill_2 FILLER_11_3383 ();
 sg13g2_decap_8 FILLER_11_3390 ();
 sg13g2_fill_1 FILLER_11_3397 ();
 sg13g2_decap_8 FILLER_11_3420 ();
 sg13g2_fill_1 FILLER_11_3427 ();
 sg13g2_decap_8 FILLER_11_3436 ();
 sg13g2_decap_8 FILLER_11_3446 ();
 sg13g2_decap_8 FILLER_11_3453 ();
 sg13g2_decap_4 FILLER_11_3460 ();
 sg13g2_fill_2 FILLER_11_3464 ();
 sg13g2_fill_2 FILLER_11_3471 ();
 sg13g2_decap_4 FILLER_11_3485 ();
 sg13g2_decap_4 FILLER_11_3508 ();
 sg13g2_decap_8 FILLER_11_3542 ();
 sg13g2_decap_8 FILLER_11_3549 ();
 sg13g2_decap_8 FILLER_11_3556 ();
 sg13g2_decap_8 FILLER_11_3563 ();
 sg13g2_decap_8 FILLER_11_3570 ();
 sg13g2_fill_2 FILLER_11_3577 ();
 sg13g2_fill_1 FILLER_11_3579 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_fill_1 FILLER_12_63 ();
 sg13g2_decap_4 FILLER_12_76 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_fill_2 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_117 ();
 sg13g2_decap_4 FILLER_12_124 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_decap_8 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_160 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_fill_2 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_205 ();
 sg13g2_decap_4 FILLER_12_212 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_decap_4 FILLER_12_279 ();
 sg13g2_fill_2 FILLER_12_283 ();
 sg13g2_fill_1 FILLER_12_289 ();
 sg13g2_decap_4 FILLER_12_303 ();
 sg13g2_fill_2 FILLER_12_376 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_2 FILLER_12_402 ();
 sg13g2_fill_1 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_432 ();
 sg13g2_decap_8 FILLER_12_439 ();
 sg13g2_decap_4 FILLER_12_478 ();
 sg13g2_decap_4 FILLER_12_496 ();
 sg13g2_fill_2 FILLER_12_500 ();
 sg13g2_decap_8 FILLER_12_505 ();
 sg13g2_decap_8 FILLER_12_512 ();
 sg13g2_fill_2 FILLER_12_541 ();
 sg13g2_fill_1 FILLER_12_543 ();
 sg13g2_decap_8 FILLER_12_548 ();
 sg13g2_decap_8 FILLER_12_555 ();
 sg13g2_fill_2 FILLER_12_562 ();
 sg13g2_fill_1 FILLER_12_585 ();
 sg13g2_fill_2 FILLER_12_594 ();
 sg13g2_fill_2 FILLER_12_605 ();
 sg13g2_decap_4 FILLER_12_612 ();
 sg13g2_fill_2 FILLER_12_624 ();
 sg13g2_fill_1 FILLER_12_626 ();
 sg13g2_decap_8 FILLER_12_635 ();
 sg13g2_decap_4 FILLER_12_642 ();
 sg13g2_fill_2 FILLER_12_657 ();
 sg13g2_fill_1 FILLER_12_659 ();
 sg13g2_fill_2 FILLER_12_670 ();
 sg13g2_fill_1 FILLER_12_695 ();
 sg13g2_fill_2 FILLER_12_726 ();
 sg13g2_fill_1 FILLER_12_728 ();
 sg13g2_fill_2 FILLER_12_745 ();
 sg13g2_decap_8 FILLER_12_752 ();
 sg13g2_decap_4 FILLER_12_776 ();
 sg13g2_fill_1 FILLER_12_780 ();
 sg13g2_decap_8 FILLER_12_792 ();
 sg13g2_decap_8 FILLER_12_799 ();
 sg13g2_fill_2 FILLER_12_806 ();
 sg13g2_fill_2 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_4 FILLER_12_826 ();
 sg13g2_fill_1 FILLER_12_830 ();
 sg13g2_fill_2 FILLER_12_857 ();
 sg13g2_fill_1 FILLER_12_859 ();
 sg13g2_decap_8 FILLER_12_885 ();
 sg13g2_decap_4 FILLER_12_913 ();
 sg13g2_fill_2 FILLER_12_917 ();
 sg13g2_decap_8 FILLER_12_928 ();
 sg13g2_decap_4 FILLER_12_935 ();
 sg13g2_decap_4 FILLER_12_952 ();
 sg13g2_fill_2 FILLER_12_956 ();
 sg13g2_decap_8 FILLER_12_972 ();
 sg13g2_decap_8 FILLER_12_979 ();
 sg13g2_decap_4 FILLER_12_986 ();
 sg13g2_decap_4 FILLER_12_994 ();
 sg13g2_fill_1 FILLER_12_998 ();
 sg13g2_decap_8 FILLER_12_1018 ();
 sg13g2_fill_1 FILLER_12_1025 ();
 sg13g2_fill_2 FILLER_12_1047 ();
 sg13g2_fill_1 FILLER_12_1049 ();
 sg13g2_decap_8 FILLER_12_1055 ();
 sg13g2_decap_8 FILLER_12_1079 ();
 sg13g2_decap_8 FILLER_12_1086 ();
 sg13g2_decap_4 FILLER_12_1101 ();
 sg13g2_fill_2 FILLER_12_1109 ();
 sg13g2_fill_1 FILLER_12_1111 ();
 sg13g2_decap_4 FILLER_12_1116 ();
 sg13g2_decap_4 FILLER_12_1134 ();
 sg13g2_fill_2 FILLER_12_1138 ();
 sg13g2_decap_8 FILLER_12_1144 ();
 sg13g2_decap_8 FILLER_12_1156 ();
 sg13g2_decap_8 FILLER_12_1163 ();
 sg13g2_fill_1 FILLER_12_1170 ();
 sg13g2_decap_4 FILLER_12_1176 ();
 sg13g2_fill_2 FILLER_12_1180 ();
 sg13g2_decap_8 FILLER_12_1226 ();
 sg13g2_fill_1 FILLER_12_1233 ();
 sg13g2_decap_8 FILLER_12_1242 ();
 sg13g2_decap_8 FILLER_12_1249 ();
 sg13g2_fill_1 FILLER_12_1256 ();
 sg13g2_decap_8 FILLER_12_1262 ();
 sg13g2_decap_8 FILLER_12_1269 ();
 sg13g2_decap_4 FILLER_12_1276 ();
 sg13g2_fill_2 FILLER_12_1280 ();
 sg13g2_fill_1 FILLER_12_1291 ();
 sg13g2_decap_8 FILLER_12_1311 ();
 sg13g2_decap_8 FILLER_12_1336 ();
 sg13g2_decap_8 FILLER_12_1343 ();
 sg13g2_fill_1 FILLER_12_1369 ();
 sg13g2_decap_4 FILLER_12_1375 ();
 sg13g2_fill_2 FILLER_12_1384 ();
 sg13g2_fill_1 FILLER_12_1386 ();
 sg13g2_fill_1 FILLER_12_1395 ();
 sg13g2_fill_2 FILLER_12_1441 ();
 sg13g2_decap_4 FILLER_12_1499 ();
 sg13g2_decap_4 FILLER_12_1522 ();
 sg13g2_fill_1 FILLER_12_1526 ();
 sg13g2_fill_2 FILLER_12_1548 ();
 sg13g2_fill_1 FILLER_12_1550 ();
 sg13g2_decap_8 FILLER_12_1574 ();
 sg13g2_fill_2 FILLER_12_1594 ();
 sg13g2_decap_8 FILLER_12_1601 ();
 sg13g2_fill_2 FILLER_12_1624 ();
 sg13g2_fill_1 FILLER_12_1626 ();
 sg13g2_fill_2 FILLER_12_1635 ();
 sg13g2_fill_1 FILLER_12_1637 ();
 sg13g2_decap_4 FILLER_12_1650 ();
 sg13g2_fill_1 FILLER_12_1662 ();
 sg13g2_fill_2 FILLER_12_1675 ();
 sg13g2_decap_4 FILLER_12_1691 ();
 sg13g2_fill_1 FILLER_12_1700 ();
 sg13g2_fill_1 FILLER_12_1715 ();
 sg13g2_fill_2 FILLER_12_1753 ();
 sg13g2_fill_2 FILLER_12_1776 ();
 sg13g2_fill_1 FILLER_12_1778 ();
 sg13g2_fill_2 FILLER_12_1805 ();
 sg13g2_decap_8 FILLER_12_1833 ();
 sg13g2_decap_4 FILLER_12_1840 ();
 sg13g2_fill_2 FILLER_12_1861 ();
 sg13g2_fill_1 FILLER_12_1863 ();
 sg13g2_decap_8 FILLER_12_1880 ();
 sg13g2_fill_1 FILLER_12_1887 ();
 sg13g2_decap_4 FILLER_12_1916 ();
 sg13g2_fill_2 FILLER_12_1920 ();
 sg13g2_fill_1 FILLER_12_1944 ();
 sg13g2_fill_2 FILLER_12_1950 ();
 sg13g2_decap_4 FILLER_12_1961 ();
 sg13g2_decap_8 FILLER_12_1987 ();
 sg13g2_fill_1 FILLER_12_1994 ();
 sg13g2_fill_2 FILLER_12_2025 ();
 sg13g2_fill_1 FILLER_12_2027 ();
 sg13g2_fill_2 FILLER_12_2050 ();
 sg13g2_fill_1 FILLER_12_2052 ();
 sg13g2_decap_4 FILLER_12_2074 ();
 sg13g2_decap_4 FILLER_12_2081 ();
 sg13g2_fill_2 FILLER_12_2100 ();
 sg13g2_fill_1 FILLER_12_2102 ();
 sg13g2_decap_8 FILLER_12_2140 ();
 sg13g2_decap_8 FILLER_12_2147 ();
 sg13g2_decap_4 FILLER_12_2154 ();
 sg13g2_fill_2 FILLER_12_2158 ();
 sg13g2_fill_2 FILLER_12_2181 ();
 sg13g2_fill_1 FILLER_12_2183 ();
 sg13g2_fill_1 FILLER_12_2257 ();
 sg13g2_fill_1 FILLER_12_2270 ();
 sg13g2_decap_8 FILLER_12_2308 ();
 sg13g2_decap_8 FILLER_12_2315 ();
 sg13g2_fill_2 FILLER_12_2322 ();
 sg13g2_fill_1 FILLER_12_2324 ();
 sg13g2_decap_4 FILLER_12_2375 ();
 sg13g2_fill_2 FILLER_12_2379 ();
 sg13g2_decap_8 FILLER_12_2385 ();
 sg13g2_fill_2 FILLER_12_2392 ();
 sg13g2_fill_1 FILLER_12_2394 ();
 sg13g2_decap_4 FILLER_12_2398 ();
 sg13g2_fill_1 FILLER_12_2402 ();
 sg13g2_fill_2 FILLER_12_2407 ();
 sg13g2_decap_8 FILLER_12_2431 ();
 sg13g2_decap_4 FILLER_12_2438 ();
 sg13g2_decap_4 FILLER_12_2446 ();
 sg13g2_fill_1 FILLER_12_2450 ();
 sg13g2_decap_4 FILLER_12_2464 ();
 sg13g2_decap_8 FILLER_12_2490 ();
 sg13g2_decap_4 FILLER_12_2497 ();
 sg13g2_fill_2 FILLER_12_2513 ();
 sg13g2_fill_2 FILLER_12_2527 ();
 sg13g2_decap_8 FILLER_12_2561 ();
 sg13g2_decap_8 FILLER_12_2568 ();
 sg13g2_decap_4 FILLER_12_2575 ();
 sg13g2_fill_1 FILLER_12_2579 ();
 sg13g2_fill_1 FILLER_12_2585 ();
 sg13g2_decap_8 FILLER_12_2592 ();
 sg13g2_fill_2 FILLER_12_2599 ();
 sg13g2_fill_1 FILLER_12_2601 ();
 sg13g2_fill_1 FILLER_12_2606 ();
 sg13g2_decap_8 FILLER_12_2634 ();
 sg13g2_decap_4 FILLER_12_2645 ();
 sg13g2_fill_1 FILLER_12_2653 ();
 sg13g2_decap_8 FILLER_12_2685 ();
 sg13g2_decap_8 FILLER_12_2709 ();
 sg13g2_decap_4 FILLER_12_2716 ();
 sg13g2_fill_2 FILLER_12_2724 ();
 sg13g2_fill_1 FILLER_12_2726 ();
 sg13g2_decap_8 FILLER_12_2745 ();
 sg13g2_decap_8 FILLER_12_2752 ();
 sg13g2_fill_2 FILLER_12_2763 ();
 sg13g2_fill_1 FILLER_12_2793 ();
 sg13g2_decap_8 FILLER_12_2820 ();
 sg13g2_fill_2 FILLER_12_2827 ();
 sg13g2_fill_1 FILLER_12_2829 ();
 sg13g2_decap_4 FILLER_12_2839 ();
 sg13g2_fill_1 FILLER_12_2843 ();
 sg13g2_fill_2 FILLER_12_2853 ();
 sg13g2_decap_8 FILLER_12_2860 ();
 sg13g2_fill_1 FILLER_12_2867 ();
 sg13g2_fill_2 FILLER_12_2900 ();
 sg13g2_decap_4 FILLER_12_2907 ();
 sg13g2_decap_4 FILLER_12_2928 ();
 sg13g2_decap_8 FILLER_12_2950 ();
 sg13g2_decap_8 FILLER_12_2957 ();
 sg13g2_fill_2 FILLER_12_2978 ();
 sg13g2_fill_1 FILLER_12_2980 ();
 sg13g2_fill_2 FILLER_12_3032 ();
 sg13g2_fill_1 FILLER_12_3034 ();
 sg13g2_decap_8 FILLER_12_3048 ();
 sg13g2_decap_4 FILLER_12_3055 ();
 sg13g2_fill_2 FILLER_12_3065 ();
 sg13g2_fill_1 FILLER_12_3071 ();
 sg13g2_decap_4 FILLER_12_3078 ();
 sg13g2_fill_2 FILLER_12_3086 ();
 sg13g2_fill_2 FILLER_12_3092 ();
 sg13g2_decap_8 FILLER_12_3116 ();
 sg13g2_fill_2 FILLER_12_3123 ();
 sg13g2_decap_8 FILLER_12_3148 ();
 sg13g2_fill_2 FILLER_12_3155 ();
 sg13g2_fill_2 FILLER_12_3161 ();
 sg13g2_fill_1 FILLER_12_3163 ();
 sg13g2_decap_4 FILLER_12_3186 ();
 sg13g2_decap_4 FILLER_12_3203 ();
 sg13g2_fill_2 FILLER_12_3230 ();
 sg13g2_fill_1 FILLER_12_3232 ();
 sg13g2_fill_1 FILLER_12_3239 ();
 sg13g2_fill_2 FILLER_12_3257 ();
 sg13g2_fill_1 FILLER_12_3259 ();
 sg13g2_fill_2 FILLER_12_3312 ();
 sg13g2_fill_1 FILLER_12_3334 ();
 sg13g2_decap_8 FILLER_12_3339 ();
 sg13g2_fill_2 FILLER_12_3346 ();
 sg13g2_decap_4 FILLER_12_3353 ();
 sg13g2_fill_2 FILLER_12_3357 ();
 sg13g2_fill_2 FILLER_12_3372 ();
 sg13g2_decap_4 FILLER_12_3393 ();
 sg13g2_fill_1 FILLER_12_3397 ();
 sg13g2_decap_8 FILLER_12_3418 ();
 sg13g2_decap_4 FILLER_12_3425 ();
 sg13g2_fill_1 FILLER_12_3470 ();
 sg13g2_decap_4 FILLER_12_3496 ();
 sg13g2_fill_1 FILLER_12_3500 ();
 sg13g2_decap_4 FILLER_12_3511 ();
 sg13g2_fill_1 FILLER_12_3515 ();
 sg13g2_decap_8 FILLER_12_3558 ();
 sg13g2_decap_8 FILLER_12_3565 ();
 sg13g2_decap_8 FILLER_12_3572 ();
 sg13g2_fill_1 FILLER_12_3579 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_130 ();
 sg13g2_decap_4 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_180 ();
 sg13g2_fill_1 FILLER_13_208 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_fill_2 FILLER_13_265 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_fill_1 FILLER_13_310 ();
 sg13g2_fill_1 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_4 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_fill_1 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_fill_2 FILLER_13_398 ();
 sg13g2_fill_2 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_459 ();
 sg13g2_decap_8 FILLER_13_466 ();
 sg13g2_decap_4 FILLER_13_473 ();
 sg13g2_fill_2 FILLER_13_477 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_fill_2 FILLER_13_530 ();
 sg13g2_decap_4 FILLER_13_536 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_fill_2 FILLER_13_560 ();
 sg13g2_fill_2 FILLER_13_575 ();
 sg13g2_fill_1 FILLER_13_577 ();
 sg13g2_fill_2 FILLER_13_583 ();
 sg13g2_fill_1 FILLER_13_585 ();
 sg13g2_fill_1 FILLER_13_590 ();
 sg13g2_fill_1 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_601 ();
 sg13g2_fill_2 FILLER_13_616 ();
 sg13g2_decap_4 FILLER_13_644 ();
 sg13g2_fill_1 FILLER_13_648 ();
 sg13g2_fill_2 FILLER_13_665 ();
 sg13g2_decap_4 FILLER_13_699 ();
 sg13g2_fill_1 FILLER_13_703 ();
 sg13g2_fill_1 FILLER_13_716 ();
 sg13g2_fill_1 FILLER_13_739 ();
 sg13g2_decap_4 FILLER_13_759 ();
 sg13g2_fill_2 FILLER_13_763 ();
 sg13g2_decap_4 FILLER_13_769 ();
 sg13g2_fill_2 FILLER_13_773 ();
 sg13g2_fill_1 FILLER_13_802 ();
 sg13g2_fill_2 FILLER_13_813 ();
 sg13g2_fill_1 FILLER_13_815 ();
 sg13g2_decap_8 FILLER_13_859 ();
 sg13g2_fill_2 FILLER_13_866 ();
 sg13g2_decap_8 FILLER_13_880 ();
 sg13g2_fill_1 FILLER_13_887 ();
 sg13g2_fill_1 FILLER_13_893 ();
 sg13g2_decap_4 FILLER_13_917 ();
 sg13g2_fill_2 FILLER_13_921 ();
 sg13g2_decap_4 FILLER_13_927 ();
 sg13g2_fill_2 FILLER_13_931 ();
 sg13g2_fill_2 FILLER_13_944 ();
 sg13g2_fill_2 FILLER_13_954 ();
 sg13g2_fill_2 FILLER_13_969 ();
 sg13g2_decap_4 FILLER_13_1021 ();
 sg13g2_fill_2 FILLER_13_1025 ();
 sg13g2_fill_2 FILLER_13_1054 ();
 sg13g2_decap_8 FILLER_13_1085 ();
 sg13g2_decap_8 FILLER_13_1142 ();
 sg13g2_fill_2 FILLER_13_1149 ();
 sg13g2_fill_1 FILLER_13_1151 ();
 sg13g2_decap_8 FILLER_13_1185 ();
 sg13g2_fill_2 FILLER_13_1196 ();
 sg13g2_fill_1 FILLER_13_1198 ();
 sg13g2_fill_1 FILLER_13_1239 ();
 sg13g2_decap_4 FILLER_13_1269 ();
 sg13g2_fill_1 FILLER_13_1273 ();
 sg13g2_fill_2 FILLER_13_1294 ();
 sg13g2_fill_2 FILLER_13_1301 ();
 sg13g2_fill_2 FILLER_13_1320 ();
 sg13g2_decap_8 FILLER_13_1350 ();
 sg13g2_fill_1 FILLER_13_1357 ();
 sg13g2_fill_1 FILLER_13_1375 ();
 sg13g2_fill_2 FILLER_13_1381 ();
 sg13g2_fill_1 FILLER_13_1383 ();
 sg13g2_decap_8 FILLER_13_1403 ();
 sg13g2_decap_4 FILLER_13_1410 ();
 sg13g2_fill_1 FILLER_13_1432 ();
 sg13g2_fill_1 FILLER_13_1442 ();
 sg13g2_fill_2 FILLER_13_1454 ();
 sg13g2_fill_2 FILLER_13_1495 ();
 sg13g2_fill_2 FILLER_13_1508 ();
 sg13g2_decap_8 FILLER_13_1530 ();
 sg13g2_decap_8 FILLER_13_1537 ();
 sg13g2_fill_2 FILLER_13_1544 ();
 sg13g2_fill_1 FILLER_13_1558 ();
 sg13g2_decap_8 FILLER_13_1567 ();
 sg13g2_decap_8 FILLER_13_1574 ();
 sg13g2_decap_4 FILLER_13_1581 ();
 sg13g2_fill_2 FILLER_13_1585 ();
 sg13g2_decap_8 FILLER_13_1619 ();
 sg13g2_decap_8 FILLER_13_1626 ();
 sg13g2_fill_2 FILLER_13_1633 ();
 sg13g2_fill_1 FILLER_13_1635 ();
 sg13g2_decap_8 FILLER_13_1642 ();
 sg13g2_fill_1 FILLER_13_1649 ();
 sg13g2_fill_1 FILLER_13_1668 ();
 sg13g2_fill_2 FILLER_13_1685 ();
 sg13g2_decap_4 FILLER_13_1704 ();
 sg13g2_fill_1 FILLER_13_1708 ();
 sg13g2_decap_4 FILLER_13_1714 ();
 sg13g2_decap_8 FILLER_13_1735 ();
 sg13g2_decap_8 FILLER_13_1742 ();
 sg13g2_fill_1 FILLER_13_1749 ();
 sg13g2_fill_1 FILLER_13_1780 ();
 sg13g2_fill_1 FILLER_13_1794 ();
 sg13g2_decap_8 FILLER_13_1807 ();
 sg13g2_decap_8 FILLER_13_1819 ();
 sg13g2_fill_2 FILLER_13_1826 ();
 sg13g2_decap_8 FILLER_13_1838 ();
 sg13g2_fill_2 FILLER_13_1845 ();
 sg13g2_fill_1 FILLER_13_1847 ();
 sg13g2_decap_4 FILLER_13_1858 ();
 sg13g2_fill_1 FILLER_13_1862 ();
 sg13g2_fill_2 FILLER_13_1868 ();
 sg13g2_fill_1 FILLER_13_1870 ();
 sg13g2_fill_2 FILLER_13_1875 ();
 sg13g2_fill_2 FILLER_13_1886 ();
 sg13g2_fill_1 FILLER_13_1888 ();
 sg13g2_decap_8 FILLER_13_1907 ();
 sg13g2_decap_4 FILLER_13_1914 ();
 sg13g2_fill_1 FILLER_13_1930 ();
 sg13g2_decap_8 FILLER_13_1956 ();
 sg13g2_fill_1 FILLER_13_1963 ();
 sg13g2_decap_8 FILLER_13_1989 ();
 sg13g2_decap_8 FILLER_13_1996 ();
 sg13g2_fill_2 FILLER_13_2012 ();
 sg13g2_fill_1 FILLER_13_2014 ();
 sg13g2_fill_2 FILLER_13_2024 ();
 sg13g2_decap_8 FILLER_13_2038 ();
 sg13g2_decap_4 FILLER_13_2045 ();
 sg13g2_fill_1 FILLER_13_2049 ();
 sg13g2_decap_4 FILLER_13_2069 ();
 sg13g2_fill_2 FILLER_13_2073 ();
 sg13g2_fill_2 FILLER_13_2085 ();
 sg13g2_decap_8 FILLER_13_2095 ();
 sg13g2_fill_2 FILLER_13_2102 ();
 sg13g2_fill_1 FILLER_13_2104 ();
 sg13g2_fill_2 FILLER_13_2130 ();
 sg13g2_fill_1 FILLER_13_2132 ();
 sg13g2_decap_8 FILLER_13_2146 ();
 sg13g2_decap_4 FILLER_13_2153 ();
 sg13g2_fill_1 FILLER_13_2157 ();
 sg13g2_decap_8 FILLER_13_2175 ();
 sg13g2_decap_4 FILLER_13_2198 ();
 sg13g2_fill_1 FILLER_13_2202 ();
 sg13g2_decap_4 FILLER_13_2207 ();
 sg13g2_fill_2 FILLER_13_2260 ();
 sg13g2_decap_8 FILLER_13_2295 ();
 sg13g2_decap_8 FILLER_13_2302 ();
 sg13g2_decap_8 FILLER_13_2309 ();
 sg13g2_fill_2 FILLER_13_2316 ();
 sg13g2_decap_8 FILLER_13_2322 ();
 sg13g2_fill_1 FILLER_13_2329 ();
 sg13g2_fill_2 FILLER_13_2338 ();
 sg13g2_fill_1 FILLER_13_2340 ();
 sg13g2_fill_1 FILLER_13_2359 ();
 sg13g2_decap_8 FILLER_13_2392 ();
 sg13g2_decap_4 FILLER_13_2399 ();
 sg13g2_decap_8 FILLER_13_2407 ();
 sg13g2_fill_2 FILLER_13_2414 ();
 sg13g2_fill_1 FILLER_13_2416 ();
 sg13g2_fill_2 FILLER_13_2455 ();
 sg13g2_fill_1 FILLER_13_2457 ();
 sg13g2_fill_2 FILLER_13_2471 ();
 sg13g2_fill_1 FILLER_13_2473 ();
 sg13g2_fill_2 FILLER_13_2477 ();
 sg13g2_fill_1 FILLER_13_2479 ();
 sg13g2_fill_1 FILLER_13_2489 ();
 sg13g2_fill_2 FILLER_13_2512 ();
 sg13g2_fill_1 FILLER_13_2514 ();
 sg13g2_fill_2 FILLER_13_2532 ();
 sg13g2_decap_8 FILLER_13_2561 ();
 sg13g2_decap_8 FILLER_13_2568 ();
 sg13g2_fill_1 FILLER_13_2575 ();
 sg13g2_decap_8 FILLER_13_2593 ();
 sg13g2_decap_8 FILLER_13_2600 ();
 sg13g2_decap_4 FILLER_13_2607 ();
 sg13g2_fill_1 FILLER_13_2611 ();
 sg13g2_fill_1 FILLER_13_2640 ();
 sg13g2_fill_2 FILLER_13_2666 ();
 sg13g2_fill_2 FILLER_13_2680 ();
 sg13g2_fill_2 FILLER_13_2728 ();
 sg13g2_fill_1 FILLER_13_2730 ();
 sg13g2_fill_2 FILLER_13_2759 ();
 sg13g2_fill_1 FILLER_13_2761 ();
 sg13g2_decap_8 FILLER_13_2786 ();
 sg13g2_decap_4 FILLER_13_2793 ();
 sg13g2_fill_2 FILLER_13_2797 ();
 sg13g2_fill_2 FILLER_13_2827 ();
 sg13g2_fill_1 FILLER_13_2829 ();
 sg13g2_decap_4 FILLER_13_2883 ();
 sg13g2_fill_2 FILLER_13_2887 ();
 sg13g2_fill_2 FILLER_13_2975 ();
 sg13g2_decap_8 FILLER_13_3009 ();
 sg13g2_decap_8 FILLER_13_3021 ();
 sg13g2_decap_4 FILLER_13_3028 ();
 sg13g2_fill_2 FILLER_13_3032 ();
 sg13g2_fill_2 FILLER_13_3062 ();
 sg13g2_fill_2 FILLER_13_3072 ();
 sg13g2_decap_8 FILLER_13_3082 ();
 sg13g2_fill_2 FILLER_13_3089 ();
 sg13g2_fill_1 FILLER_13_3091 ();
 sg13g2_fill_1 FILLER_13_3096 ();
 sg13g2_decap_4 FILLER_13_3124 ();
 sg13g2_fill_2 FILLER_13_3128 ();
 sg13g2_decap_8 FILLER_13_3162 ();
 sg13g2_fill_2 FILLER_13_3169 ();
 sg13g2_fill_1 FILLER_13_3171 ();
 sg13g2_decap_8 FILLER_13_3204 ();
 sg13g2_decap_4 FILLER_13_3211 ();
 sg13g2_decap_8 FILLER_13_3252 ();
 sg13g2_fill_2 FILLER_13_3259 ();
 sg13g2_fill_1 FILLER_13_3265 ();
 sg13g2_fill_2 FILLER_13_3270 ();
 sg13g2_fill_1 FILLER_13_3272 ();
 sg13g2_fill_1 FILLER_13_3296 ();
 sg13g2_decap_8 FILLER_13_3305 ();
 sg13g2_fill_2 FILLER_13_3327 ();
 sg13g2_fill_1 FILLER_13_3343 ();
 sg13g2_fill_2 FILLER_13_3359 ();
 sg13g2_fill_1 FILLER_13_3361 ();
 sg13g2_decap_8 FILLER_13_3370 ();
 sg13g2_fill_2 FILLER_13_3377 ();
 sg13g2_fill_1 FILLER_13_3379 ();
 sg13g2_fill_1 FILLER_13_3388 ();
 sg13g2_fill_2 FILLER_13_3393 ();
 sg13g2_fill_1 FILLER_13_3395 ();
 sg13g2_decap_4 FILLER_13_3405 ();
 sg13g2_fill_2 FILLER_13_3420 ();
 sg13g2_fill_1 FILLER_13_3427 ();
 sg13g2_decap_4 FILLER_13_3441 ();
 sg13g2_fill_1 FILLER_13_3445 ();
 sg13g2_decap_8 FILLER_13_3451 ();
 sg13g2_decap_8 FILLER_13_3458 ();
 sg13g2_fill_2 FILLER_13_3480 ();
 sg13g2_fill_1 FILLER_13_3482 ();
 sg13g2_decap_4 FILLER_13_3500 ();
 sg13g2_fill_2 FILLER_13_3512 ();
 sg13g2_fill_1 FILLER_13_3514 ();
 sg13g2_fill_1 FILLER_13_3529 ();
 sg13g2_decap_8 FILLER_13_3543 ();
 sg13g2_decap_8 FILLER_13_3550 ();
 sg13g2_decap_8 FILLER_13_3557 ();
 sg13g2_decap_8 FILLER_13_3564 ();
 sg13g2_decap_8 FILLER_13_3571 ();
 sg13g2_fill_2 FILLER_13_3578 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_4 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_89 ();
 sg13g2_decap_8 FILLER_14_96 ();
 sg13g2_decap_8 FILLER_14_114 ();
 sg13g2_decap_4 FILLER_14_121 ();
 sg13g2_fill_2 FILLER_14_125 ();
 sg13g2_fill_2 FILLER_14_139 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_4 FILLER_14_175 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_fill_2 FILLER_14_189 ();
 sg13g2_decap_4 FILLER_14_196 ();
 sg13g2_fill_1 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_220 ();
 sg13g2_decap_4 FILLER_14_267 ();
 sg13g2_fill_2 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_4 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_365 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_fill_1 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_1 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_422 ();
 sg13g2_fill_2 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_14_444 ();
 sg13g2_fill_2 FILLER_14_451 ();
 sg13g2_fill_1 FILLER_14_453 ();
 sg13g2_decap_4 FILLER_14_485 ();
 sg13g2_decap_8 FILLER_14_493 ();
 sg13g2_decap_4 FILLER_14_500 ();
 sg13g2_fill_1 FILLER_14_504 ();
 sg13g2_fill_1 FILLER_14_559 ();
 sg13g2_decap_4 FILLER_14_581 ();
 sg13g2_fill_2 FILLER_14_604 ();
 sg13g2_decap_4 FILLER_14_612 ();
 sg13g2_fill_2 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_fill_1 FILLER_14_651 ();
 sg13g2_fill_1 FILLER_14_665 ();
 sg13g2_decap_4 FILLER_14_685 ();
 sg13g2_fill_1 FILLER_14_697 ();
 sg13g2_fill_2 FILLER_14_716 ();
 sg13g2_decap_4 FILLER_14_726 ();
 sg13g2_fill_1 FILLER_14_730 ();
 sg13g2_decap_8 FILLER_14_747 ();
 sg13g2_decap_4 FILLER_14_754 ();
 sg13g2_fill_2 FILLER_14_770 ();
 sg13g2_fill_1 FILLER_14_772 ();
 sg13g2_fill_2 FILLER_14_795 ();
 sg13g2_fill_1 FILLER_14_797 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_fill_1 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_823 ();
 sg13g2_decap_4 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_860 ();
 sg13g2_fill_2 FILLER_14_867 ();
 sg13g2_fill_1 FILLER_14_869 ();
 sg13g2_decap_8 FILLER_14_879 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_decap_8 FILLER_14_915 ();
 sg13g2_fill_2 FILLER_14_940 ();
 sg13g2_decap_8 FILLER_14_960 ();
 sg13g2_decap_4 FILLER_14_967 ();
 sg13g2_decap_4 FILLER_14_993 ();
 sg13g2_fill_1 FILLER_14_997 ();
 sg13g2_fill_2 FILLER_14_1037 ();
 sg13g2_decap_4 FILLER_14_1065 ();
 sg13g2_fill_1 FILLER_14_1069 ();
 sg13g2_fill_1 FILLER_14_1098 ();
 sg13g2_decap_8 FILLER_14_1112 ();
 sg13g2_fill_2 FILLER_14_1128 ();
 sg13g2_fill_1 FILLER_14_1158 ();
 sg13g2_decap_8 FILLER_14_1163 ();
 sg13g2_decap_8 FILLER_14_1196 ();
 sg13g2_decap_8 FILLER_14_1203 ();
 sg13g2_fill_2 FILLER_14_1210 ();
 sg13g2_decap_8 FILLER_14_1220 ();
 sg13g2_fill_1 FILLER_14_1236 ();
 sg13g2_fill_1 FILLER_14_1245 ();
 sg13g2_decap_8 FILLER_14_1262 ();
 sg13g2_decap_4 FILLER_14_1269 ();
 sg13g2_fill_1 FILLER_14_1273 ();
 sg13g2_fill_2 FILLER_14_1302 ();
 sg13g2_fill_1 FILLER_14_1304 ();
 sg13g2_decap_8 FILLER_14_1337 ();
 sg13g2_decap_8 FILLER_14_1344 ();
 sg13g2_fill_1 FILLER_14_1366 ();
 sg13g2_fill_1 FILLER_14_1377 ();
 sg13g2_fill_2 FILLER_14_1385 ();
 sg13g2_fill_1 FILLER_14_1387 ();
 sg13g2_decap_8 FILLER_14_1403 ();
 sg13g2_fill_2 FILLER_14_1410 ();
 sg13g2_fill_1 FILLER_14_1435 ();
 sg13g2_fill_2 FILLER_14_1448 ();
 sg13g2_fill_1 FILLER_14_1450 ();
 sg13g2_fill_2 FILLER_14_1502 ();
 sg13g2_fill_1 FILLER_14_1516 ();
 sg13g2_decap_8 FILLER_14_1521 ();
 sg13g2_decap_8 FILLER_14_1528 ();
 sg13g2_decap_4 FILLER_14_1535 ();
 sg13g2_fill_1 FILLER_14_1539 ();
 sg13g2_fill_2 FILLER_14_1553 ();
 sg13g2_decap_8 FILLER_14_1573 ();
 sg13g2_fill_2 FILLER_14_1580 ();
 sg13g2_fill_1 FILLER_14_1582 ();
 sg13g2_fill_1 FILLER_14_1587 ();
 sg13g2_decap_4 FILLER_14_1605 ();
 sg13g2_fill_2 FILLER_14_1609 ();
 sg13g2_decap_4 FILLER_14_1624 ();
 sg13g2_fill_2 FILLER_14_1628 ();
 sg13g2_decap_8 FILLER_14_1641 ();
 sg13g2_decap_8 FILLER_14_1648 ();
 sg13g2_fill_2 FILLER_14_1655 ();
 sg13g2_fill_2 FILLER_14_1685 ();
 sg13g2_fill_1 FILLER_14_1687 ();
 sg13g2_fill_1 FILLER_14_1697 ();
 sg13g2_decap_8 FILLER_14_1702 ();
 sg13g2_decap_4 FILLER_14_1709 ();
 sg13g2_fill_1 FILLER_14_1713 ();
 sg13g2_decap_8 FILLER_14_1750 ();
 sg13g2_fill_2 FILLER_14_1757 ();
 sg13g2_decap_4 FILLER_14_1772 ();
 sg13g2_fill_2 FILLER_14_1776 ();
 sg13g2_fill_2 FILLER_14_1791 ();
 sg13g2_fill_1 FILLER_14_1793 ();
 sg13g2_decap_8 FILLER_14_1802 ();
 sg13g2_decap_4 FILLER_14_1809 ();
 sg13g2_fill_2 FILLER_14_1813 ();
 sg13g2_decap_4 FILLER_14_1827 ();
 sg13g2_fill_2 FILLER_14_1847 ();
 sg13g2_decap_4 FILLER_14_1854 ();
 sg13g2_fill_2 FILLER_14_1875 ();
 sg13g2_fill_1 FILLER_14_1877 ();
 sg13g2_fill_2 FILLER_14_1887 ();
 sg13g2_fill_1 FILLER_14_1889 ();
 sg13g2_decap_8 FILLER_14_1911 ();
 sg13g2_decap_4 FILLER_14_1918 ();
 sg13g2_fill_1 FILLER_14_1922 ();
 sg13g2_fill_2 FILLER_14_1936 ();
 sg13g2_fill_1 FILLER_14_1938 ();
 sg13g2_fill_2 FILLER_14_1953 ();
 sg13g2_decap_8 FILLER_14_1959 ();
 sg13g2_fill_1 FILLER_14_1966 ();
 sg13g2_decap_4 FILLER_14_1984 ();
 sg13g2_fill_2 FILLER_14_1988 ();
 sg13g2_decap_8 FILLER_14_2045 ();
 sg13g2_decap_4 FILLER_14_2052 ();
 sg13g2_fill_1 FILLER_14_2056 ();
 sg13g2_decap_4 FILLER_14_2073 ();
 sg13g2_fill_2 FILLER_14_2077 ();
 sg13g2_decap_8 FILLER_14_2087 ();
 sg13g2_decap_8 FILLER_14_2099 ();
 sg13g2_decap_4 FILLER_14_2106 ();
 sg13g2_fill_1 FILLER_14_2110 ();
 sg13g2_fill_2 FILLER_14_2125 ();
 sg13g2_fill_1 FILLER_14_2127 ();
 sg13g2_fill_1 FILLER_14_2133 ();
 sg13g2_decap_8 FILLER_14_2147 ();
 sg13g2_fill_2 FILLER_14_2154 ();
 sg13g2_fill_1 FILLER_14_2156 ();
 sg13g2_decap_4 FILLER_14_2167 ();
 sg13g2_fill_1 FILLER_14_2171 ();
 sg13g2_fill_2 FILLER_14_2176 ();
 sg13g2_fill_1 FILLER_14_2185 ();
 sg13g2_decap_8 FILLER_14_2202 ();
 sg13g2_decap_4 FILLER_14_2209 ();
 sg13g2_decap_8 FILLER_14_2229 ();
 sg13g2_decap_8 FILLER_14_2236 ();
 sg13g2_fill_1 FILLER_14_2252 ();
 sg13g2_fill_2 FILLER_14_2257 ();
 sg13g2_fill_1 FILLER_14_2259 ();
 sg13g2_fill_2 FILLER_14_2263 ();
 sg13g2_fill_2 FILLER_14_2296 ();
 sg13g2_fill_1 FILLER_14_2298 ();
 sg13g2_fill_1 FILLER_14_2312 ();
 sg13g2_fill_1 FILLER_14_2379 ();
 sg13g2_fill_2 FILLER_14_2419 ();
 sg13g2_fill_1 FILLER_14_2421 ();
 sg13g2_fill_2 FILLER_14_2439 ();
 sg13g2_fill_1 FILLER_14_2441 ();
 sg13g2_fill_2 FILLER_14_2455 ();
 sg13g2_fill_2 FILLER_14_2485 ();
 sg13g2_fill_2 FILLER_14_2496 ();
 sg13g2_decap_8 FILLER_14_2532 ();
 sg13g2_decap_4 FILLER_14_2539 ();
 sg13g2_fill_2 FILLER_14_2579 ();
 sg13g2_decap_4 FILLER_14_2609 ();
 sg13g2_fill_2 FILLER_14_2613 ();
 sg13g2_decap_8 FILLER_14_2620 ();
 sg13g2_decap_4 FILLER_14_2627 ();
 sg13g2_fill_2 FILLER_14_2631 ();
 sg13g2_decap_4 FILLER_14_2642 ();
 sg13g2_fill_1 FILLER_14_2646 ();
 sg13g2_decap_8 FILLER_14_2655 ();
 sg13g2_decap_8 FILLER_14_2662 ();
 sg13g2_decap_8 FILLER_14_2677 ();
 sg13g2_decap_4 FILLER_14_2710 ();
 sg13g2_decap_8 FILLER_14_2735 ();
 sg13g2_fill_2 FILLER_14_2742 ();
 sg13g2_fill_2 FILLER_14_2770 ();
 sg13g2_fill_1 FILLER_14_2772 ();
 sg13g2_fill_2 FILLER_14_2795 ();
 sg13g2_fill_1 FILLER_14_2797 ();
 sg13g2_decap_4 FILLER_14_2803 ();
 sg13g2_decap_8 FILLER_14_2811 ();
 sg13g2_decap_8 FILLER_14_2818 ();
 sg13g2_decap_8 FILLER_14_2825 ();
 sg13g2_decap_4 FILLER_14_2832 ();
 sg13g2_fill_2 FILLER_14_2836 ();
 sg13g2_decap_4 FILLER_14_2851 ();
 sg13g2_fill_2 FILLER_14_2864 ();
 sg13g2_fill_2 FILLER_14_2887 ();
 sg13g2_fill_1 FILLER_14_2889 ();
 sg13g2_fill_2 FILLER_14_2902 ();
 sg13g2_fill_1 FILLER_14_2904 ();
 sg13g2_fill_2 FILLER_14_2913 ();
 sg13g2_fill_1 FILLER_14_2915 ();
 sg13g2_fill_2 FILLER_14_2942 ();
 sg13g2_fill_1 FILLER_14_2944 ();
 sg13g2_decap_8 FILLER_14_2988 ();
 sg13g2_decap_8 FILLER_14_2995 ();
 sg13g2_decap_4 FILLER_14_3002 ();
 sg13g2_fill_2 FILLER_14_3026 ();
 sg13g2_decap_8 FILLER_14_3031 ();
 sg13g2_decap_8 FILLER_14_3038 ();
 sg13g2_decap_8 FILLER_14_3045 ();
 sg13g2_decap_8 FILLER_14_3052 ();
 sg13g2_fill_2 FILLER_14_3059 ();
 sg13g2_decap_8 FILLER_14_3087 ();
 sg13g2_fill_1 FILLER_14_3094 ();
 sg13g2_decap_4 FILLER_14_3100 ();
 sg13g2_fill_2 FILLER_14_3104 ();
 sg13g2_decap_4 FILLER_14_3116 ();
 sg13g2_fill_2 FILLER_14_3120 ();
 sg13g2_fill_2 FILLER_14_3143 ();
 sg13g2_fill_2 FILLER_14_3187 ();
 sg13g2_fill_1 FILLER_14_3189 ();
 sg13g2_fill_1 FILLER_14_3203 ();
 sg13g2_decap_8 FILLER_14_3234 ();
 sg13g2_fill_2 FILLER_14_3241 ();
 sg13g2_fill_1 FILLER_14_3243 ();
 sg13g2_fill_1 FILLER_14_3292 ();
 sg13g2_decap_4 FILLER_14_3301 ();
 sg13g2_fill_1 FILLER_14_3313 ();
 sg13g2_fill_1 FILLER_14_3322 ();
 sg13g2_decap_8 FILLER_14_3327 ();
 sg13g2_decap_8 FILLER_14_3334 ();
 sg13g2_fill_2 FILLER_14_3341 ();
 sg13g2_fill_1 FILLER_14_3343 ();
 sg13g2_decap_8 FILLER_14_3371 ();
 sg13g2_decap_4 FILLER_14_3412 ();
 sg13g2_fill_1 FILLER_14_3426 ();
 sg13g2_decap_8 FILLER_14_3431 ();
 sg13g2_fill_1 FILLER_14_3447 ();
 sg13g2_fill_2 FILLER_14_3453 ();
 sg13g2_fill_2 FILLER_14_3487 ();
 sg13g2_fill_1 FILLER_14_3489 ();
 sg13g2_decap_8 FILLER_14_3503 ();
 sg13g2_fill_2 FILLER_14_3510 ();
 sg13g2_fill_2 FILLER_14_3529 ();
 sg13g2_decap_8 FILLER_14_3559 ();
 sg13g2_decap_8 FILLER_14_3566 ();
 sg13g2_decap_8 FILLER_14_3573 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_49 ();
 sg13g2_decap_4 FILLER_15_75 ();
 sg13g2_fill_1 FILLER_15_79 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_4 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_120 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_171 ();
 sg13g2_decap_8 FILLER_15_180 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_decap_4 FILLER_15_207 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_222 ();
 sg13g2_fill_1 FILLER_15_224 ();
 sg13g2_decap_4 FILLER_15_230 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_257 ();
 sg13g2_fill_2 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_292 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_decap_4 FILLER_15_320 ();
 sg13g2_fill_2 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_4 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_1 FILLER_15_366 ();
 sg13g2_fill_2 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_15_379 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_1 FILLER_15_415 ();
 sg13g2_decap_4 FILLER_15_435 ();
 sg13g2_fill_1 FILLER_15_439 ();
 sg13g2_fill_2 FILLER_15_446 ();
 sg13g2_fill_1 FILLER_15_448 ();
 sg13g2_fill_1 FILLER_15_463 ();
 sg13g2_decap_4 FILLER_15_492 ();
 sg13g2_decap_4 FILLER_15_504 ();
 sg13g2_fill_2 FILLER_15_513 ();
 sg13g2_decap_8 FILLER_15_528 ();
 sg13g2_fill_2 FILLER_15_535 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_decap_4 FILLER_15_564 ();
 sg13g2_fill_1 FILLER_15_568 ();
 sg13g2_fill_2 FILLER_15_573 ();
 sg13g2_decap_4 FILLER_15_583 ();
 sg13g2_fill_2 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_601 ();
 sg13g2_fill_2 FILLER_15_608 ();
 sg13g2_fill_2 FILLER_15_622 ();
 sg13g2_fill_1 FILLER_15_624 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_fill_1 FILLER_15_651 ();
 sg13g2_decap_4 FILLER_15_665 ();
 sg13g2_decap_4 FILLER_15_672 ();
 sg13g2_fill_1 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_694 ();
 sg13g2_fill_1 FILLER_15_701 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_4 FILLER_15_732 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_fill_1 FILLER_15_753 ();
 sg13g2_fill_2 FILLER_15_768 ();
 sg13g2_fill_1 FILLER_15_770 ();
 sg13g2_decap_4 FILLER_15_784 ();
 sg13g2_fill_2 FILLER_15_788 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_fill_1 FILLER_15_809 ();
 sg13g2_fill_2 FILLER_15_843 ();
 sg13g2_fill_1 FILLER_15_845 ();
 sg13g2_fill_2 FILLER_15_874 ();
 sg13g2_fill_1 FILLER_15_876 ();
 sg13g2_decap_8 FILLER_15_890 ();
 sg13g2_decap_4 FILLER_15_897 ();
 sg13g2_fill_1 FILLER_15_901 ();
 sg13g2_fill_1 FILLER_15_930 ();
 sg13g2_fill_2 FILLER_15_962 ();
 sg13g2_fill_1 FILLER_15_968 ();
 sg13g2_decap_8 FILLER_15_992 ();
 sg13g2_decap_4 FILLER_15_999 ();
 sg13g2_fill_2 FILLER_15_1008 ();
 sg13g2_decap_4 FILLER_15_1018 ();
 sg13g2_decap_8 FILLER_15_1027 ();
 sg13g2_decap_8 FILLER_15_1034 ();
 sg13g2_fill_2 FILLER_15_1041 ();
 sg13g2_fill_1 FILLER_15_1043 ();
 sg13g2_decap_8 FILLER_15_1072 ();
 sg13g2_decap_4 FILLER_15_1079 ();
 sg13g2_fill_2 FILLER_15_1095 ();
 sg13g2_fill_1 FILLER_15_1097 ();
 sg13g2_decap_8 FILLER_15_1130 ();
 sg13g2_decap_8 FILLER_15_1137 ();
 sg13g2_fill_2 FILLER_15_1144 ();
 sg13g2_decap_4 FILLER_15_1156 ();
 sg13g2_fill_1 FILLER_15_1160 ();
 sg13g2_decap_4 FILLER_15_1178 ();
 sg13g2_fill_1 FILLER_15_1210 ();
 sg13g2_fill_2 FILLER_15_1252 ();
 sg13g2_fill_1 FILLER_15_1254 ();
 sg13g2_decap_8 FILLER_15_1268 ();
 sg13g2_decap_4 FILLER_15_1275 ();
 sg13g2_fill_1 FILLER_15_1283 ();
 sg13g2_decap_8 FILLER_15_1316 ();
 sg13g2_decap_8 FILLER_15_1323 ();
 sg13g2_decap_8 FILLER_15_1334 ();
 sg13g2_fill_2 FILLER_15_1341 ();
 sg13g2_fill_2 FILLER_15_1369 ();
 sg13g2_decap_4 FILLER_15_1390 ();
 sg13g2_fill_2 FILLER_15_1394 ();
 sg13g2_decap_8 FILLER_15_1404 ();
 sg13g2_fill_1 FILLER_15_1429 ();
 sg13g2_decap_4 FILLER_15_1443 ();
 sg13g2_fill_2 FILLER_15_1451 ();
 sg13g2_fill_1 FILLER_15_1453 ();
 sg13g2_decap_8 FILLER_15_1462 ();
 sg13g2_decap_4 FILLER_15_1469 ();
 sg13g2_fill_2 FILLER_15_1488 ();
 sg13g2_fill_1 FILLER_15_1490 ();
 sg13g2_fill_2 FILLER_15_1523 ();
 sg13g2_decap_8 FILLER_15_1547 ();
 sg13g2_fill_2 FILLER_15_1554 ();
 sg13g2_fill_1 FILLER_15_1556 ();
 sg13g2_fill_2 FILLER_15_1593 ();
 sg13g2_fill_1 FILLER_15_1595 ();
 sg13g2_fill_1 FILLER_15_1604 ();
 sg13g2_fill_2 FILLER_15_1611 ();
 sg13g2_fill_1 FILLER_15_1613 ();
 sg13g2_decap_8 FILLER_15_1658 ();
 sg13g2_decap_4 FILLER_15_1665 ();
 sg13g2_fill_1 FILLER_15_1669 ();
 sg13g2_fill_2 FILLER_15_1674 ();
 sg13g2_fill_2 FILLER_15_1684 ();
 sg13g2_fill_2 FILLER_15_1692 ();
 sg13g2_decap_8 FILLER_15_1707 ();
 sg13g2_fill_2 FILLER_15_1714 ();
 sg13g2_fill_2 FILLER_15_1719 ();
 sg13g2_fill_1 FILLER_15_1721 ();
 sg13g2_decap_8 FILLER_15_1731 ();
 sg13g2_decap_8 FILLER_15_1738 ();
 sg13g2_decap_8 FILLER_15_1751 ();
 sg13g2_decap_8 FILLER_15_1758 ();
 sg13g2_fill_2 FILLER_15_1765 ();
 sg13g2_fill_1 FILLER_15_1767 ();
 sg13g2_fill_1 FILLER_15_1794 ();
 sg13g2_decap_4 FILLER_15_1817 ();
 sg13g2_fill_1 FILLER_15_1821 ();
 sg13g2_decap_8 FILLER_15_1858 ();
 sg13g2_fill_1 FILLER_15_1865 ();
 sg13g2_decap_4 FILLER_15_1875 ();
 sg13g2_fill_1 FILLER_15_1879 ();
 sg13g2_fill_2 FILLER_15_1896 ();
 sg13g2_fill_2 FILLER_15_1903 ();
 sg13g2_fill_1 FILLER_15_1905 ();
 sg13g2_decap_8 FILLER_15_1919 ();
 sg13g2_decap_8 FILLER_15_1926 ();
 sg13g2_fill_1 FILLER_15_1933 ();
 sg13g2_fill_1 FILLER_15_1939 ();
 sg13g2_fill_1 FILLER_15_1947 ();
 sg13g2_fill_1 FILLER_15_1968 ();
 sg13g2_fill_2 FILLER_15_1974 ();
 sg13g2_decap_8 FILLER_15_1981 ();
 sg13g2_decap_8 FILLER_15_1988 ();
 sg13g2_fill_2 FILLER_15_2017 ();
 sg13g2_fill_1 FILLER_15_2019 ();
 sg13g2_fill_2 FILLER_15_2047 ();
 sg13g2_fill_1 FILLER_15_2049 ();
 sg13g2_decap_8 FILLER_15_2075 ();
 sg13g2_decap_4 FILLER_15_2082 ();
 sg13g2_decap_4 FILLER_15_2112 ();
 sg13g2_fill_1 FILLER_15_2116 ();
 sg13g2_decap_4 FILLER_15_2132 ();
 sg13g2_fill_2 FILLER_15_2145 ();
 sg13g2_fill_2 FILLER_15_2152 ();
 sg13g2_fill_1 FILLER_15_2154 ();
 sg13g2_decap_8 FILLER_15_2199 ();
 sg13g2_decap_8 FILLER_15_2206 ();
 sg13g2_fill_2 FILLER_15_2213 ();
 sg13g2_decap_4 FILLER_15_2238 ();
 sg13g2_decap_8 FILLER_15_2258 ();
 sg13g2_decap_4 FILLER_15_2278 ();
 sg13g2_decap_4 FILLER_15_2326 ();
 sg13g2_fill_1 FILLER_15_2330 ();
 sg13g2_decap_4 FILLER_15_2336 ();
 sg13g2_fill_1 FILLER_15_2340 ();
 sg13g2_fill_1 FILLER_15_2348 ();
 sg13g2_decap_8 FILLER_15_2354 ();
 sg13g2_decap_8 FILLER_15_2361 ();
 sg13g2_fill_2 FILLER_15_2368 ();
 sg13g2_fill_1 FILLER_15_2370 ();
 sg13g2_decap_4 FILLER_15_2400 ();
 sg13g2_fill_2 FILLER_15_2408 ();
 sg13g2_decap_4 FILLER_15_2436 ();
 sg13g2_decap_8 FILLER_15_2456 ();
 sg13g2_fill_1 FILLER_15_2463 ();
 sg13g2_decap_8 FILLER_15_2502 ();
 sg13g2_fill_1 FILLER_15_2509 ();
 sg13g2_decap_4 FILLER_15_2520 ();
 sg13g2_decap_4 FILLER_15_2541 ();
 sg13g2_fill_1 FILLER_15_2545 ();
 sg13g2_fill_1 FILLER_15_2554 ();
 sg13g2_decap_8 FILLER_15_2560 ();
 sg13g2_decap_8 FILLER_15_2567 ();
 sg13g2_decap_8 FILLER_15_2574 ();
 sg13g2_fill_2 FILLER_15_2589 ();
 sg13g2_fill_1 FILLER_15_2591 ();
 sg13g2_decap_4 FILLER_15_2625 ();
 sg13g2_decap_8 FILLER_15_2646 ();
 sg13g2_fill_2 FILLER_15_2653 ();
 sg13g2_fill_2 FILLER_15_2694 ();
 sg13g2_fill_1 FILLER_15_2696 ();
 sg13g2_fill_2 FILLER_15_2706 ();
 sg13g2_fill_1 FILLER_15_2708 ();
 sg13g2_decap_4 FILLER_15_2727 ();
 sg13g2_fill_1 FILLER_15_2731 ();
 sg13g2_fill_1 FILLER_15_2763 ();
 sg13g2_fill_1 FILLER_15_2773 ();
 sg13g2_decap_8 FILLER_15_2784 ();
 sg13g2_fill_1 FILLER_15_2791 ();
 sg13g2_decap_8 FILLER_15_2832 ();
 sg13g2_decap_8 FILLER_15_2852 ();
 sg13g2_decap_4 FILLER_15_2859 ();
 sg13g2_fill_1 FILLER_15_2868 ();
 sg13g2_decap_8 FILLER_15_2879 ();
 sg13g2_decap_8 FILLER_15_2886 ();
 sg13g2_fill_1 FILLER_15_2893 ();
 sg13g2_decap_4 FILLER_15_2898 ();
 sg13g2_fill_1 FILLER_15_2902 ();
 sg13g2_decap_8 FILLER_15_2931 ();
 sg13g2_fill_2 FILLER_15_2938 ();
 sg13g2_fill_1 FILLER_15_2940 ();
 sg13g2_decap_8 FILLER_15_2954 ();
 sg13g2_decap_8 FILLER_15_2961 ();
 sg13g2_fill_1 FILLER_15_2968 ();
 sg13g2_decap_8 FILLER_15_2974 ();
 sg13g2_decap_8 FILLER_15_2981 ();
 sg13g2_fill_2 FILLER_15_2988 ();
 sg13g2_fill_1 FILLER_15_2990 ();
 sg13g2_fill_1 FILLER_15_3004 ();
 sg13g2_fill_1 FILLER_15_3019 ();
 sg13g2_fill_1 FILLER_15_3029 ();
 sg13g2_fill_2 FILLER_15_3035 ();
 sg13g2_fill_1 FILLER_15_3037 ();
 sg13g2_fill_2 FILLER_15_3048 ();
 sg13g2_decap_4 FILLER_15_3054 ();
 sg13g2_fill_1 FILLER_15_3058 ();
 sg13g2_fill_1 FILLER_15_3071 ();
 sg13g2_fill_2 FILLER_15_3080 ();
 sg13g2_fill_1 FILLER_15_3082 ();
 sg13g2_fill_2 FILLER_15_3089 ();
 sg13g2_fill_1 FILLER_15_3091 ();
 sg13g2_fill_2 FILLER_15_3100 ();
 sg13g2_fill_2 FILLER_15_3122 ();
 sg13g2_fill_1 FILLER_15_3124 ();
 sg13g2_decap_4 FILLER_15_3141 ();
 sg13g2_decap_4 FILLER_15_3167 ();
 sg13g2_fill_2 FILLER_15_3171 ();
 sg13g2_decap_8 FILLER_15_3189 ();
 sg13g2_decap_8 FILLER_15_3196 ();
 sg13g2_fill_2 FILLER_15_3203 ();
 sg13g2_fill_1 FILLER_15_3205 ();
 sg13g2_fill_1 FILLER_15_3224 ();
 sg13g2_fill_1 FILLER_15_3229 ();
 sg13g2_decap_8 FILLER_15_3238 ();
 sg13g2_decap_8 FILLER_15_3245 ();
 sg13g2_decap_8 FILLER_15_3252 ();
 sg13g2_decap_8 FILLER_15_3259 ();
 sg13g2_decap_4 FILLER_15_3266 ();
 sg13g2_fill_2 FILLER_15_3270 ();
 sg13g2_decap_4 FILLER_15_3298 ();
 sg13g2_fill_1 FILLER_15_3302 ();
 sg13g2_decap_4 FILLER_15_3326 ();
 sg13g2_decap_4 FILLER_15_3335 ();
 sg13g2_fill_1 FILLER_15_3339 ();
 sg13g2_fill_2 FILLER_15_3345 ();
 sg13g2_decap_8 FILLER_15_3362 ();
 sg13g2_decap_4 FILLER_15_3369 ();
 sg13g2_decap_8 FILLER_15_3402 ();
 sg13g2_fill_2 FILLER_15_3455 ();
 sg13g2_decap_8 FILLER_15_3480 ();
 sg13g2_fill_2 FILLER_15_3487 ();
 sg13g2_fill_1 FILLER_15_3489 ();
 sg13g2_decap_8 FILLER_15_3510 ();
 sg13g2_fill_1 FILLER_15_3517 ();
 sg13g2_fill_1 FILLER_15_3525 ();
 sg13g2_fill_1 FILLER_15_3535 ();
 sg13g2_decap_8 FILLER_15_3540 ();
 sg13g2_decap_8 FILLER_15_3547 ();
 sg13g2_decap_8 FILLER_15_3554 ();
 sg13g2_decap_8 FILLER_15_3561 ();
 sg13g2_decap_8 FILLER_15_3568 ();
 sg13g2_decap_4 FILLER_15_3575 ();
 sg13g2_fill_1 FILLER_15_3579 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_23 ();
 sg13g2_fill_1 FILLER_16_52 ();
 sg13g2_fill_2 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_96 ();
 sg13g2_decap_8 FILLER_16_103 ();
 sg13g2_fill_2 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_145 ();
 sg13g2_fill_2 FILLER_16_169 ();
 sg13g2_decap_4 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_decap_4 FILLER_16_232 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_decap_8 FILLER_16_257 ();
 sg13g2_fill_2 FILLER_16_273 ();
 sg13g2_fill_1 FILLER_16_275 ();
 sg13g2_fill_2 FILLER_16_292 ();
 sg13g2_fill_2 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_fill_1 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_347 ();
 sg13g2_decap_4 FILLER_16_359 ();
 sg13g2_fill_2 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_4 FILLER_16_377 ();
 sg13g2_decap_4 FILLER_16_394 ();
 sg13g2_fill_2 FILLER_16_398 ();
 sg13g2_fill_2 FILLER_16_429 ();
 sg13g2_fill_2 FILLER_16_448 ();
 sg13g2_fill_2 FILLER_16_455 ();
 sg13g2_fill_1 FILLER_16_457 ();
 sg13g2_fill_2 FILLER_16_475 ();
 sg13g2_fill_1 FILLER_16_482 ();
 sg13g2_fill_1 FILLER_16_491 ();
 sg13g2_decap_4 FILLER_16_499 ();
 sg13g2_decap_4 FILLER_16_530 ();
 sg13g2_decap_8 FILLER_16_554 ();
 sg13g2_decap_8 FILLER_16_561 ();
 sg13g2_decap_8 FILLER_16_568 ();
 sg13g2_fill_2 FILLER_16_588 ();
 sg13g2_fill_1 FILLER_16_590 ();
 sg13g2_decap_4 FILLER_16_604 ();
 sg13g2_decap_8 FILLER_16_612 ();
 sg13g2_decap_8 FILLER_16_619 ();
 sg13g2_fill_2 FILLER_16_626 ();
 sg13g2_decap_8 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_685 ();
 sg13g2_fill_2 FILLER_16_692 ();
 sg13g2_fill_1 FILLER_16_756 ();
 sg13g2_decap_4 FILLER_16_807 ();
 sg13g2_fill_1 FILLER_16_824 ();
 sg13g2_decap_8 FILLER_16_841 ();
 sg13g2_fill_2 FILLER_16_848 ();
 sg13g2_decap_8 FILLER_16_912 ();
 sg13g2_fill_2 FILLER_16_919 ();
 sg13g2_decap_4 FILLER_16_934 ();
 sg13g2_fill_1 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_943 ();
 sg13g2_decap_4 FILLER_16_950 ();
 sg13g2_fill_1 FILLER_16_954 ();
 sg13g2_fill_2 FILLER_16_967 ();
 sg13g2_fill_1 FILLER_16_969 ();
 sg13g2_fill_1 FILLER_16_1014 ();
 sg13g2_fill_1 FILLER_16_1023 ();
 sg13g2_fill_2 FILLER_16_1032 ();
 sg13g2_fill_2 FILLER_16_1063 ();
 sg13g2_fill_1 FILLER_16_1078 ();
 sg13g2_decap_8 FILLER_16_1100 ();
 sg13g2_fill_2 FILLER_16_1112 ();
 sg13g2_fill_1 FILLER_16_1114 ();
 sg13g2_fill_2 FILLER_16_1140 ();
 sg13g2_fill_1 FILLER_16_1142 ();
 sg13g2_fill_2 FILLER_16_1163 ();
 sg13g2_fill_1 FILLER_16_1165 ();
 sg13g2_decap_8 FILLER_16_1194 ();
 sg13g2_fill_2 FILLER_16_1201 ();
 sg13g2_fill_1 FILLER_16_1215 ();
 sg13g2_decap_8 FILLER_16_1242 ();
 sg13g2_decap_4 FILLER_16_1277 ();
 sg13g2_decap_8 FILLER_16_1310 ();
 sg13g2_decap_4 FILLER_16_1317 ();
 sg13g2_fill_1 FILLER_16_1321 ();
 sg13g2_fill_2 FILLER_16_1353 ();
 sg13g2_decap_4 FILLER_16_1368 ();
 sg13g2_decap_8 FILLER_16_1376 ();
 sg13g2_decap_4 FILLER_16_1383 ();
 sg13g2_decap_8 FILLER_16_1391 ();
 sg13g2_decap_4 FILLER_16_1407 ();
 sg13g2_fill_1 FILLER_16_1411 ();
 sg13g2_decap_4 FILLER_16_1416 ();
 sg13g2_fill_1 FILLER_16_1420 ();
 sg13g2_decap_8 FILLER_16_1425 ();
 sg13g2_fill_1 FILLER_16_1432 ();
 sg13g2_fill_2 FILLER_16_1484 ();
 sg13g2_fill_1 FILLER_16_1486 ();
 sg13g2_decap_8 FILLER_16_1516 ();
 sg13g2_fill_2 FILLER_16_1523 ();
 sg13g2_fill_1 FILLER_16_1525 ();
 sg13g2_fill_2 FILLER_16_1558 ();
 sg13g2_fill_1 FILLER_16_1573 ();
 sg13g2_decap_4 FILLER_16_1592 ();
 sg13g2_decap_8 FILLER_16_1612 ();
 sg13g2_fill_1 FILLER_16_1619 ();
 sg13g2_fill_2 FILLER_16_1623 ();
 sg13g2_fill_1 FILLER_16_1625 ();
 sg13g2_fill_2 FILLER_16_1643 ();
 sg13g2_decap_4 FILLER_16_1667 ();
 sg13g2_fill_1 FILLER_16_1671 ();
 sg13g2_fill_2 FILLER_16_1689 ();
 sg13g2_fill_1 FILLER_16_1691 ();
 sg13g2_fill_2 FILLER_16_1720 ();
 sg13g2_fill_1 FILLER_16_1722 ();
 sg13g2_decap_4 FILLER_16_1731 ();
 sg13g2_decap_8 FILLER_16_1770 ();
 sg13g2_fill_2 FILLER_16_1777 ();
 sg13g2_fill_1 FILLER_16_1779 ();
 sg13g2_fill_2 FILLER_16_1791 ();
 sg13g2_fill_1 FILLER_16_1793 ();
 sg13g2_decap_8 FILLER_16_1808 ();
 sg13g2_decap_8 FILLER_16_1815 ();
 sg13g2_decap_8 FILLER_16_1860 ();
 sg13g2_fill_2 FILLER_16_1905 ();
 sg13g2_fill_1 FILLER_16_1907 ();
 sg13g2_decap_8 FILLER_16_1913 ();
 sg13g2_decap_4 FILLER_16_1920 ();
 sg13g2_fill_1 FILLER_16_1924 ();
 sg13g2_decap_8 FILLER_16_1945 ();
 sg13g2_decap_8 FILLER_16_1952 ();
 sg13g2_decap_4 FILLER_16_1985 ();
 sg13g2_fill_2 FILLER_16_1998 ();
 sg13g2_fill_1 FILLER_16_2000 ();
 sg13g2_decap_8 FILLER_16_2029 ();
 sg13g2_fill_2 FILLER_16_2036 ();
 sg13g2_decap_8 FILLER_16_2043 ();
 sg13g2_decap_8 FILLER_16_2050 ();
 sg13g2_fill_2 FILLER_16_2068 ();
 sg13g2_decap_8 FILLER_16_2074 ();
 sg13g2_decap_8 FILLER_16_2081 ();
 sg13g2_fill_1 FILLER_16_2088 ();
 sg13g2_fill_1 FILLER_16_2107 ();
 sg13g2_fill_2 FILLER_16_2111 ();
 sg13g2_decap_4 FILLER_16_2130 ();
 sg13g2_fill_2 FILLER_16_2134 ();
 sg13g2_decap_8 FILLER_16_2171 ();
 sg13g2_fill_2 FILLER_16_2178 ();
 sg13g2_fill_1 FILLER_16_2180 ();
 sg13g2_fill_1 FILLER_16_2185 ();
 sg13g2_fill_1 FILLER_16_2204 ();
 sg13g2_fill_1 FILLER_16_2213 ();
 sg13g2_decap_4 FILLER_16_2242 ();
 sg13g2_fill_1 FILLER_16_2246 ();
 sg13g2_fill_2 FILLER_16_2260 ();
 sg13g2_decap_8 FILLER_16_2291 ();
 sg13g2_decap_8 FILLER_16_2298 ();
 sg13g2_decap_8 FILLER_16_2305 ();
 sg13g2_fill_1 FILLER_16_2312 ();
 sg13g2_fill_1 FILLER_16_2326 ();
 sg13g2_fill_1 FILLER_16_2340 ();
 sg13g2_decap_4 FILLER_16_2362 ();
 sg13g2_fill_1 FILLER_16_2366 ();
 sg13g2_decap_4 FILLER_16_2380 ();
 sg13g2_fill_2 FILLER_16_2384 ();
 sg13g2_fill_1 FILLER_16_2407 ();
 sg13g2_fill_2 FILLER_16_2413 ();
 sg13g2_fill_1 FILLER_16_2415 ();
 sg13g2_fill_2 FILLER_16_2429 ();
 sg13g2_decap_4 FILLER_16_2459 ();
 sg13g2_fill_2 FILLER_16_2489 ();
 sg13g2_fill_1 FILLER_16_2491 ();
 sg13g2_fill_2 FILLER_16_2523 ();
 sg13g2_fill_1 FILLER_16_2525 ();
 sg13g2_decap_8 FILLER_16_2568 ();
 sg13g2_fill_2 FILLER_16_2575 ();
 sg13g2_fill_2 FILLER_16_2586 ();
 sg13g2_fill_1 FILLER_16_2588 ();
 sg13g2_fill_2 FILLER_16_2598 ();
 sg13g2_decap_4 FILLER_16_2619 ();
 sg13g2_fill_2 FILLER_16_2623 ();
 sg13g2_decap_8 FILLER_16_2649 ();
 sg13g2_decap_4 FILLER_16_2656 ();
 sg13g2_fill_1 FILLER_16_2660 ();
 sg13g2_decap_8 FILLER_16_2670 ();
 sg13g2_decap_8 FILLER_16_2677 ();
 sg13g2_fill_1 FILLER_16_2684 ();
 sg13g2_decap_8 FILLER_16_2715 ();
 sg13g2_decap_8 FILLER_16_2722 ();
 sg13g2_fill_2 FILLER_16_2729 ();
 sg13g2_fill_1 FILLER_16_2739 ();
 sg13g2_decap_8 FILLER_16_2760 ();
 sg13g2_fill_2 FILLER_16_2767 ();
 sg13g2_decap_4 FILLER_16_2785 ();
 sg13g2_decap_4 FILLER_16_2793 ();
 sg13g2_fill_1 FILLER_16_2797 ();
 sg13g2_decap_8 FILLER_16_2802 ();
 sg13g2_fill_2 FILLER_16_2809 ();
 sg13g2_fill_1 FILLER_16_2811 ();
 sg13g2_decap_4 FILLER_16_2855 ();
 sg13g2_fill_2 FILLER_16_2859 ();
 sg13g2_decap_4 FILLER_16_2887 ();
 sg13g2_decap_8 FILLER_16_2903 ();
 sg13g2_decap_8 FILLER_16_2910 ();
 sg13g2_decap_8 FILLER_16_2922 ();
 sg13g2_fill_2 FILLER_16_2929 ();
 sg13g2_fill_1 FILLER_16_2944 ();
 sg13g2_decap_4 FILLER_16_2958 ();
 sg13g2_decap_4 FILLER_16_2966 ();
 sg13g2_fill_2 FILLER_16_2970 ();
 sg13g2_decap_4 FILLER_16_2977 ();
 sg13g2_decap_8 FILLER_16_2994 ();
 sg13g2_decap_8 FILLER_16_3001 ();
 sg13g2_decap_8 FILLER_16_3008 ();
 sg13g2_decap_8 FILLER_16_3023 ();
 sg13g2_fill_2 FILLER_16_3030 ();
 sg13g2_fill_1 FILLER_16_3037 ();
 sg13g2_decap_8 FILLER_16_3043 ();
 sg13g2_fill_2 FILLER_16_3050 ();
 sg13g2_decap_8 FILLER_16_3063 ();
 sg13g2_decap_8 FILLER_16_3070 ();
 sg13g2_fill_1 FILLER_16_3077 ();
 sg13g2_fill_2 FILLER_16_3084 ();
 sg13g2_decap_4 FILLER_16_3091 ();
 sg13g2_fill_1 FILLER_16_3095 ();
 sg13g2_fill_2 FILLER_16_3101 ();
 sg13g2_decap_8 FILLER_16_3107 ();
 sg13g2_fill_2 FILLER_16_3114 ();
 sg13g2_fill_1 FILLER_16_3116 ();
 sg13g2_decap_8 FILLER_16_3135 ();
 sg13g2_fill_1 FILLER_16_3142 ();
 sg13g2_fill_2 FILLER_16_3153 ();
 sg13g2_decap_8 FILLER_16_3160 ();
 sg13g2_decap_4 FILLER_16_3192 ();
 sg13g2_fill_1 FILLER_16_3196 ();
 sg13g2_fill_2 FILLER_16_3206 ();
 sg13g2_fill_1 FILLER_16_3221 ();
 sg13g2_fill_2 FILLER_16_3238 ();
 sg13g2_decap_8 FILLER_16_3260 ();
 sg13g2_fill_1 FILLER_16_3267 ();
 sg13g2_fill_2 FILLER_16_3281 ();
 sg13g2_decap_8 FILLER_16_3300 ();
 sg13g2_decap_4 FILLER_16_3307 ();
 sg13g2_fill_2 FILLER_16_3324 ();
 sg13g2_fill_2 FILLER_16_3339 ();
 sg13g2_fill_2 FILLER_16_3349 ();
 sg13g2_decap_4 FILLER_16_3371 ();
 sg13g2_fill_1 FILLER_16_3375 ();
 sg13g2_decap_4 FILLER_16_3379 ();
 sg13g2_fill_1 FILLER_16_3383 ();
 sg13g2_decap_8 FILLER_16_3425 ();
 sg13g2_fill_1 FILLER_16_3432 ();
 sg13g2_fill_1 FILLER_16_3443 ();
 sg13g2_decap_4 FILLER_16_3452 ();
 sg13g2_fill_2 FILLER_16_3456 ();
 sg13g2_fill_1 FILLER_16_3481 ();
 sg13g2_decap_8 FILLER_16_3510 ();
 sg13g2_decap_8 FILLER_16_3554 ();
 sg13g2_decap_8 FILLER_16_3561 ();
 sg13g2_decap_8 FILLER_16_3568 ();
 sg13g2_decap_4 FILLER_16_3575 ();
 sg13g2_fill_1 FILLER_16_3579 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_33 ();
 sg13g2_decap_8 FILLER_17_40 ();
 sg13g2_decap_4 FILLER_17_47 ();
 sg13g2_fill_2 FILLER_17_58 ();
 sg13g2_fill_1 FILLER_17_60 ();
 sg13g2_decap_8 FILLER_17_86 ();
 sg13g2_decap_8 FILLER_17_97 ();
 sg13g2_decap_4 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_decap_4 FILLER_17_143 ();
 sg13g2_decap_4 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_decap_8 FILLER_17_171 ();
 sg13g2_decap_8 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_4 FILLER_17_214 ();
 sg13g2_fill_2 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_256 ();
 sg13g2_fill_1 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_270 ();
 sg13g2_fill_2 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_285 ();
 sg13g2_decap_4 FILLER_17_298 ();
 sg13g2_decap_4 FILLER_17_320 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_fill_2 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_4 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_fill_1 FILLER_17_383 ();
 sg13g2_fill_1 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_449 ();
 sg13g2_fill_2 FILLER_17_456 ();
 sg13g2_decap_4 FILLER_17_491 ();
 sg13g2_fill_1 FILLER_17_504 ();
 sg13g2_decap_4 FILLER_17_567 ();
 sg13g2_fill_2 FILLER_17_599 ();
 sg13g2_fill_1 FILLER_17_601 ();
 sg13g2_fill_1 FILLER_17_618 ();
 sg13g2_fill_1 FILLER_17_632 ();
 sg13g2_decap_8 FILLER_17_646 ();
 sg13g2_fill_2 FILLER_17_653 ();
 sg13g2_decap_4 FILLER_17_662 ();
 sg13g2_fill_2 FILLER_17_666 ();
 sg13g2_decap_8 FILLER_17_681 ();
 sg13g2_decap_8 FILLER_17_719 ();
 sg13g2_decap_8 FILLER_17_726 ();
 sg13g2_fill_2 FILLER_17_733 ();
 sg13g2_fill_2 FILLER_17_753 ();
 sg13g2_fill_1 FILLER_17_755 ();
 sg13g2_fill_2 FILLER_17_760 ();
 sg13g2_fill_2 FILLER_17_766 ();
 sg13g2_decap_8 FILLER_17_781 ();
 sg13g2_decap_4 FILLER_17_788 ();
 sg13g2_fill_2 FILLER_17_792 ();
 sg13g2_fill_1 FILLER_17_827 ();
 sg13g2_decap_4 FILLER_17_895 ();
 sg13g2_fill_1 FILLER_17_915 ();
 sg13g2_fill_2 FILLER_17_938 ();
 sg13g2_decap_4 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_964 ();
 sg13g2_decap_4 FILLER_17_971 ();
 sg13g2_fill_1 FILLER_17_975 ();
 sg13g2_decap_4 FILLER_17_984 ();
 sg13g2_fill_2 FILLER_17_988 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_4 FILLER_17_1008 ();
 sg13g2_fill_2 FILLER_17_1012 ();
 sg13g2_fill_2 FILLER_17_1023 ();
 sg13g2_decap_4 FILLER_17_1038 ();
 sg13g2_fill_2 FILLER_17_1042 ();
 sg13g2_decap_8 FILLER_17_1067 ();
 sg13g2_decap_8 FILLER_17_1074 ();
 sg13g2_fill_2 FILLER_17_1081 ();
 sg13g2_fill_2 FILLER_17_1088 ();
 sg13g2_decap_4 FILLER_17_1100 ();
 sg13g2_fill_1 FILLER_17_1109 ();
 sg13g2_fill_2 FILLER_17_1115 ();
 sg13g2_decap_4 FILLER_17_1121 ();
 sg13g2_decap_8 FILLER_17_1133 ();
 sg13g2_decap_4 FILLER_17_1140 ();
 sg13g2_decap_8 FILLER_17_1164 ();
 sg13g2_fill_1 FILLER_17_1171 ();
 sg13g2_decap_8 FILLER_17_1176 ();
 sg13g2_decap_4 FILLER_17_1183 ();
 sg13g2_fill_2 FILLER_17_1187 ();
 sg13g2_decap_4 FILLER_17_1194 ();
 sg13g2_fill_2 FILLER_17_1198 ();
 sg13g2_decap_8 FILLER_17_1210 ();
 sg13g2_decap_8 FILLER_17_1217 ();
 sg13g2_decap_8 FILLER_17_1224 ();
 sg13g2_fill_2 FILLER_17_1235 ();
 sg13g2_decap_4 FILLER_17_1276 ();
 sg13g2_fill_2 FILLER_17_1280 ();
 sg13g2_fill_2 FILLER_17_1303 ();
 sg13g2_fill_2 FILLER_17_1326 ();
 sg13g2_decap_8 FILLER_17_1334 ();
 sg13g2_decap_8 FILLER_17_1341 ();
 sg13g2_decap_4 FILLER_17_1348 ();
 sg13g2_fill_2 FILLER_17_1352 ();
 sg13g2_decap_4 FILLER_17_1430 ();
 sg13g2_fill_2 FILLER_17_1443 ();
 sg13g2_decap_4 FILLER_17_1473 ();
 sg13g2_fill_2 FILLER_17_1490 ();
 sg13g2_fill_1 FILLER_17_1506 ();
 sg13g2_fill_2 FILLER_17_1535 ();
 sg13g2_decap_4 FILLER_17_1555 ();
 sg13g2_decap_4 FILLER_17_1621 ();
 sg13g2_decap_4 FILLER_17_1681 ();
 sg13g2_decap_8 FILLER_17_1693 ();
 sg13g2_decap_8 FILLER_17_1707 ();
 sg13g2_fill_2 FILLER_17_1714 ();
 sg13g2_decap_4 FILLER_17_1754 ();
 sg13g2_fill_1 FILLER_17_1758 ();
 sg13g2_decap_4 FILLER_17_1783 ();
 sg13g2_fill_1 FILLER_17_1792 ();
 sg13g2_fill_2 FILLER_17_1825 ();
 sg13g2_decap_8 FILLER_17_1830 ();
 sg13g2_fill_1 FILLER_17_1837 ();
 sg13g2_decap_8 FILLER_17_1859 ();
 sg13g2_fill_2 FILLER_17_1871 ();
 sg13g2_fill_1 FILLER_17_1883 ();
 sg13g2_decap_8 FILLER_17_1894 ();
 sg13g2_decap_8 FILLER_17_1901 ();
 sg13g2_decap_8 FILLER_17_1908 ();
 sg13g2_fill_1 FILLER_17_1915 ();
 sg13g2_fill_2 FILLER_17_1944 ();
 sg13g2_fill_1 FILLER_17_1968 ();
 sg13g2_fill_2 FILLER_17_1977 ();
 sg13g2_fill_1 FILLER_17_1979 ();
 sg13g2_decap_8 FILLER_17_1988 ();
 sg13g2_decap_4 FILLER_17_1995 ();
 sg13g2_fill_2 FILLER_17_2003 ();
 sg13g2_fill_1 FILLER_17_2013 ();
 sg13g2_fill_2 FILLER_17_2019 ();
 sg13g2_fill_1 FILLER_17_2021 ();
 sg13g2_fill_2 FILLER_17_2027 ();
 sg13g2_fill_1 FILLER_17_2029 ();
 sg13g2_fill_2 FILLER_17_2064 ();
 sg13g2_decap_4 FILLER_17_2079 ();
 sg13g2_fill_1 FILLER_17_2083 ();
 sg13g2_fill_1 FILLER_17_2096 ();
 sg13g2_decap_8 FILLER_17_2107 ();
 sg13g2_decap_4 FILLER_17_2114 ();
 sg13g2_fill_1 FILLER_17_2118 ();
 sg13g2_fill_2 FILLER_17_2124 ();
 sg13g2_fill_1 FILLER_17_2126 ();
 sg13g2_decap_8 FILLER_17_2132 ();
 sg13g2_decap_8 FILLER_17_2139 ();
 sg13g2_fill_1 FILLER_17_2146 ();
 sg13g2_fill_1 FILLER_17_2155 ();
 sg13g2_decap_4 FILLER_17_2165 ();
 sg13g2_fill_2 FILLER_17_2182 ();
 sg13g2_decap_8 FILLER_17_2199 ();
 sg13g2_decap_4 FILLER_17_2206 ();
 sg13g2_fill_2 FILLER_17_2220 ();
 sg13g2_fill_1 FILLER_17_2222 ();
 sg13g2_decap_8 FILLER_17_2241 ();
 sg13g2_decap_4 FILLER_17_2248 ();
 sg13g2_fill_1 FILLER_17_2252 ();
 sg13g2_decap_8 FILLER_17_2278 ();
 sg13g2_fill_1 FILLER_17_2285 ();
 sg13g2_fill_1 FILLER_17_2291 ();
 sg13g2_decap_4 FILLER_17_2333 ();
 sg13g2_fill_1 FILLER_17_2337 ();
 sg13g2_fill_2 FILLER_17_2353 ();
 sg13g2_fill_1 FILLER_17_2355 ();
 sg13g2_decap_4 FILLER_17_2361 ();
 sg13g2_fill_1 FILLER_17_2365 ();
 sg13g2_decap_4 FILLER_17_2383 ();
 sg13g2_fill_1 FILLER_17_2387 ();
 sg13g2_fill_1 FILLER_17_2396 ();
 sg13g2_fill_2 FILLER_17_2402 ();
 sg13g2_fill_1 FILLER_17_2404 ();
 sg13g2_decap_4 FILLER_17_2433 ();
 sg13g2_decap_8 FILLER_17_2452 ();
 sg13g2_decap_8 FILLER_17_2459 ();
 sg13g2_fill_1 FILLER_17_2466 ();
 sg13g2_fill_2 FILLER_17_2498 ();
 sg13g2_fill_2 FILLER_17_2505 ();
 sg13g2_fill_1 FILLER_17_2507 ();
 sg13g2_fill_2 FILLER_17_2525 ();
 sg13g2_decap_8 FILLER_17_2542 ();
 sg13g2_decap_4 FILLER_17_2549 ();
 sg13g2_fill_2 FILLER_17_2553 ();
 sg13g2_decap_8 FILLER_17_2567 ();
 sg13g2_fill_1 FILLER_17_2574 ();
 sg13g2_fill_1 FILLER_17_2588 ();
 sg13g2_decap_8 FILLER_17_2600 ();
 sg13g2_decap_8 FILLER_17_2607 ();
 sg13g2_decap_4 FILLER_17_2640 ();
 sg13g2_fill_2 FILLER_17_2644 ();
 sg13g2_fill_2 FILLER_17_2651 ();
 sg13g2_fill_1 FILLER_17_2653 ();
 sg13g2_fill_1 FILLER_17_2679 ();
 sg13g2_fill_1 FILLER_17_2696 ();
 sg13g2_fill_1 FILLER_17_2710 ();
 sg13g2_fill_2 FILLER_17_2731 ();
 sg13g2_fill_1 FILLER_17_2733 ();
 sg13g2_decap_4 FILLER_17_2739 ();
 sg13g2_decap_4 FILLER_17_2755 ();
 sg13g2_fill_2 FILLER_17_2759 ();
 sg13g2_fill_2 FILLER_17_2790 ();
 sg13g2_fill_1 FILLER_17_2792 ();
 sg13g2_decap_8 FILLER_17_2810 ();
 sg13g2_decap_4 FILLER_17_2817 ();
 sg13g2_fill_1 FILLER_17_2821 ();
 sg13g2_decap_8 FILLER_17_2827 ();
 sg13g2_fill_2 FILLER_17_2834 ();
 sg13g2_fill_2 FILLER_17_2850 ();
 sg13g2_fill_1 FILLER_17_2852 ();
 sg13g2_fill_1 FILLER_17_2861 ();
 sg13g2_decap_8 FILLER_17_2883 ();
 sg13g2_fill_2 FILLER_17_2890 ();
 sg13g2_fill_1 FILLER_17_2892 ();
 sg13g2_decap_8 FILLER_17_2911 ();
 sg13g2_fill_2 FILLER_17_2933 ();
 sg13g2_fill_1 FILLER_17_2943 ();
 sg13g2_decap_8 FILLER_17_2976 ();
 sg13g2_decap_4 FILLER_17_3004 ();
 sg13g2_fill_2 FILLER_17_3012 ();
 sg13g2_decap_4 FILLER_17_3031 ();
 sg13g2_fill_2 FILLER_17_3035 ();
 sg13g2_decap_4 FILLER_17_3059 ();
 sg13g2_fill_2 FILLER_17_3063 ();
 sg13g2_decap_8 FILLER_17_3079 ();
 sg13g2_fill_1 FILLER_17_3086 ();
 sg13g2_decap_4 FILLER_17_3102 ();
 sg13g2_fill_2 FILLER_17_3106 ();
 sg13g2_fill_1 FILLER_17_3121 ();
 sg13g2_decap_8 FILLER_17_3135 ();
 sg13g2_fill_2 FILLER_17_3142 ();
 sg13g2_fill_1 FILLER_17_3165 ();
 sg13g2_fill_2 FILLER_17_3185 ();
 sg13g2_decap_4 FILLER_17_3205 ();
 sg13g2_fill_2 FILLER_17_3209 ();
 sg13g2_fill_1 FILLER_17_3224 ();
 sg13g2_decap_4 FILLER_17_3239 ();
 sg13g2_fill_1 FILLER_17_3256 ();
 sg13g2_decap_8 FILLER_17_3276 ();
 sg13g2_fill_1 FILLER_17_3283 ();
 sg13g2_decap_4 FILLER_17_3297 ();
 sg13g2_fill_2 FILLER_17_3301 ();
 sg13g2_fill_1 FILLER_17_3323 ();
 sg13g2_decap_8 FILLER_17_3329 ();
 sg13g2_fill_2 FILLER_17_3336 ();
 sg13g2_fill_1 FILLER_17_3338 ();
 sg13g2_decap_4 FILLER_17_3343 ();
 sg13g2_fill_2 FILLER_17_3347 ();
 sg13g2_decap_8 FILLER_17_3353 ();
 sg13g2_fill_1 FILLER_17_3360 ();
 sg13g2_fill_1 FILLER_17_3366 ();
 sg13g2_decap_8 FILLER_17_3375 ();
 sg13g2_decap_4 FILLER_17_3382 ();
 sg13g2_fill_2 FILLER_17_3399 ();
 sg13g2_fill_1 FILLER_17_3401 ();
 sg13g2_decap_4 FILLER_17_3448 ();
 sg13g2_decap_8 FILLER_17_3457 ();
 sg13g2_fill_2 FILLER_17_3499 ();
 sg13g2_fill_2 FILLER_17_3505 ();
 sg13g2_decap_8 FILLER_17_3539 ();
 sg13g2_decap_8 FILLER_17_3546 ();
 sg13g2_decap_8 FILLER_17_3553 ();
 sg13g2_decap_8 FILLER_17_3560 ();
 sg13g2_decap_8 FILLER_17_3567 ();
 sg13g2_decap_4 FILLER_17_3574 ();
 sg13g2_fill_2 FILLER_17_3578 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_54 ();
 sg13g2_decap_4 FILLER_18_61 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_fill_2 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_fill_1 FILLER_18_142 ();
 sg13g2_decap_4 FILLER_18_173 ();
 sg13g2_fill_2 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_197 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_decap_4 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_286 ();
 sg13g2_decap_4 FILLER_18_293 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_decap_4 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_fill_2 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_fill_2 FILLER_18_399 ();
 sg13g2_fill_1 FILLER_18_405 ();
 sg13g2_fill_2 FILLER_18_419 ();
 sg13g2_fill_1 FILLER_18_421 ();
 sg13g2_decap_4 FILLER_18_426 ();
 sg13g2_fill_2 FILLER_18_430 ();
 sg13g2_fill_1 FILLER_18_473 ();
 sg13g2_decap_8 FILLER_18_527 ();
 sg13g2_fill_2 FILLER_18_543 ();
 sg13g2_fill_1 FILLER_18_545 ();
 sg13g2_fill_1 FILLER_18_551 ();
 sg13g2_fill_2 FILLER_18_573 ();
 sg13g2_fill_1 FILLER_18_575 ();
 sg13g2_fill_2 FILLER_18_580 ();
 sg13g2_fill_2 FILLER_18_596 ();
 sg13g2_fill_1 FILLER_18_598 ();
 sg13g2_decap_8 FILLER_18_620 ();
 sg13g2_decap_4 FILLER_18_627 ();
 sg13g2_fill_1 FILLER_18_659 ();
 sg13g2_decap_4 FILLER_18_693 ();
 sg13g2_fill_1 FILLER_18_697 ();
 sg13g2_fill_2 FILLER_18_701 ();
 sg13g2_decap_4 FILLER_18_764 ();
 sg13g2_fill_1 FILLER_18_768 ();
 sg13g2_fill_2 FILLER_18_782 ();
 sg13g2_decap_4 FILLER_18_819 ();
 sg13g2_fill_1 FILLER_18_823 ();
 sg13g2_decap_4 FILLER_18_828 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_fill_2 FILLER_18_850 ();
 sg13g2_fill_1 FILLER_18_852 ();
 sg13g2_fill_1 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_901 ();
 sg13g2_fill_2 FILLER_18_908 ();
 sg13g2_fill_1 FILLER_18_910 ();
 sg13g2_fill_2 FILLER_18_915 ();
 sg13g2_fill_1 FILLER_18_917 ();
 sg13g2_decap_4 FILLER_18_946 ();
 sg13g2_fill_1 FILLER_18_950 ();
 sg13g2_fill_1 FILLER_18_969 ();
 sg13g2_fill_2 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1011 ();
 sg13g2_fill_1 FILLER_18_1052 ();
 sg13g2_fill_1 FILLER_18_1061 ();
 sg13g2_decap_8 FILLER_18_1075 ();
 sg13g2_fill_2 FILLER_18_1082 ();
 sg13g2_fill_2 FILLER_18_1141 ();
 sg13g2_decap_4 FILLER_18_1173 ();
 sg13g2_fill_1 FILLER_18_1177 ();
 sg13g2_fill_2 FILLER_18_1194 ();
 sg13g2_fill_1 FILLER_18_1196 ();
 sg13g2_fill_1 FILLER_18_1216 ();
 sg13g2_fill_1 FILLER_18_1234 ();
 sg13g2_fill_1 FILLER_18_1240 ();
 sg13g2_fill_2 FILLER_18_1255 ();
 sg13g2_fill_1 FILLER_18_1294 ();
 sg13g2_fill_2 FILLER_18_1305 ();
 sg13g2_decap_8 FILLER_18_1312 ();
 sg13g2_fill_1 FILLER_18_1339 ();
 sg13g2_decap_8 FILLER_18_1344 ();
 sg13g2_decap_8 FILLER_18_1351 ();
 sg13g2_decap_4 FILLER_18_1358 ();
 sg13g2_fill_1 FILLER_18_1362 ();
 sg13g2_decap_4 FILLER_18_1373 ();
 sg13g2_decap_8 FILLER_18_1383 ();
 sg13g2_decap_4 FILLER_18_1390 ();
 sg13g2_fill_2 FILLER_18_1394 ();
 sg13g2_fill_1 FILLER_18_1413 ();
 sg13g2_fill_2 FILLER_18_1470 ();
 sg13g2_fill_1 FILLER_18_1472 ();
 sg13g2_decap_4 FILLER_18_1477 ();
 sg13g2_fill_1 FILLER_18_1481 ();
 sg13g2_fill_2 FILLER_18_1491 ();
 sg13g2_decap_8 FILLER_18_1526 ();
 sg13g2_decap_8 FILLER_18_1537 ();
 sg13g2_decap_8 FILLER_18_1544 ();
 sg13g2_decap_8 FILLER_18_1551 ();
 sg13g2_decap_4 FILLER_18_1558 ();
 sg13g2_decap_8 FILLER_18_1568 ();
 sg13g2_fill_2 FILLER_18_1575 ();
 sg13g2_fill_1 FILLER_18_1577 ();
 sg13g2_decap_8 FILLER_18_1582 ();
 sg13g2_decap_8 FILLER_18_1589 ();
 sg13g2_decap_8 FILLER_18_1596 ();
 sg13g2_fill_2 FILLER_18_1603 ();
 sg13g2_fill_1 FILLER_18_1605 ();
 sg13g2_fill_2 FILLER_18_1610 ();
 sg13g2_decap_8 FILLER_18_1617 ();
 sg13g2_decap_8 FILLER_18_1624 ();
 sg13g2_decap_4 FILLER_18_1631 ();
 sg13g2_fill_1 FILLER_18_1635 ();
 sg13g2_decap_8 FILLER_18_1647 ();
 sg13g2_decap_8 FILLER_18_1654 ();
 sg13g2_fill_1 FILLER_18_1661 ();
 sg13g2_fill_1 FILLER_18_1674 ();
 sg13g2_decap_4 FILLER_18_1680 ();
 sg13g2_fill_2 FILLER_18_1684 ();
 sg13g2_decap_8 FILLER_18_1712 ();
 sg13g2_decap_4 FILLER_18_1719 ();
 sg13g2_fill_2 FILLER_18_1723 ();
 sg13g2_decap_4 FILLER_18_1734 ();
 sg13g2_fill_1 FILLER_18_1738 ();
 sg13g2_fill_1 FILLER_18_1778 ();
 sg13g2_fill_1 FILLER_18_1801 ();
 sg13g2_decap_8 FILLER_18_1806 ();
 sg13g2_decap_8 FILLER_18_1813 ();
 sg13g2_decap_8 FILLER_18_1833 ();
 sg13g2_decap_4 FILLER_18_1840 ();
 sg13g2_fill_1 FILLER_18_1848 ();
 sg13g2_decap_8 FILLER_18_1852 ();
 sg13g2_fill_2 FILLER_18_1859 ();
 sg13g2_fill_1 FILLER_18_1861 ();
 sg13g2_fill_2 FILLER_18_1883 ();
 sg13g2_fill_1 FILLER_18_1892 ();
 sg13g2_fill_2 FILLER_18_1898 ();
 sg13g2_fill_1 FILLER_18_1900 ();
 sg13g2_fill_2 FILLER_18_1939 ();
 sg13g2_fill_1 FILLER_18_1941 ();
 sg13g2_decap_8 FILLER_18_1956 ();
 sg13g2_fill_1 FILLER_18_1963 ();
 sg13g2_decap_8 FILLER_18_1985 ();
 sg13g2_fill_2 FILLER_18_1992 ();
 sg13g2_fill_2 FILLER_18_2006 ();
 sg13g2_fill_1 FILLER_18_2008 ();
 sg13g2_fill_2 FILLER_18_2022 ();
 sg13g2_decap_4 FILLER_18_2064 ();
 sg13g2_fill_1 FILLER_18_2068 ();
 sg13g2_decap_8 FILLER_18_2110 ();
 sg13g2_decap_8 FILLER_18_2137 ();
 sg13g2_decap_4 FILLER_18_2144 ();
 sg13g2_fill_1 FILLER_18_2148 ();
 sg13g2_fill_2 FILLER_18_2177 ();
 sg13g2_fill_1 FILLER_18_2179 ();
 sg13g2_decap_4 FILLER_18_2224 ();
 sg13g2_fill_2 FILLER_18_2228 ();
 sg13g2_decap_8 FILLER_18_2235 ();
 sg13g2_fill_1 FILLER_18_2242 ();
 sg13g2_fill_2 FILLER_18_2256 ();
 sg13g2_fill_1 FILLER_18_2258 ();
 sg13g2_decap_8 FILLER_18_2264 ();
 sg13g2_decap_4 FILLER_18_2271 ();
 sg13g2_fill_2 FILLER_18_2275 ();
 sg13g2_fill_1 FILLER_18_2303 ();
 sg13g2_decap_8 FILLER_18_2331 ();
 sg13g2_fill_1 FILLER_18_2338 ();
 sg13g2_decap_8 FILLER_18_2364 ();
 sg13g2_fill_2 FILLER_18_2371 ();
 sg13g2_decap_8 FILLER_18_2383 ();
 sg13g2_decap_4 FILLER_18_2390 ();
 sg13g2_fill_1 FILLER_18_2394 ();
 sg13g2_fill_1 FILLER_18_2405 ();
 sg13g2_decap_8 FILLER_18_2424 ();
 sg13g2_fill_2 FILLER_18_2431 ();
 sg13g2_decap_8 FILLER_18_2456 ();
 sg13g2_fill_2 FILLER_18_2510 ();
 sg13g2_fill_1 FILLER_18_2512 ();
 sg13g2_decap_8 FILLER_18_2518 ();
 sg13g2_decap_8 FILLER_18_2525 ();
 sg13g2_fill_2 FILLER_18_2537 ();
 sg13g2_fill_1 FILLER_18_2539 ();
 sg13g2_fill_1 FILLER_18_2544 ();
 sg13g2_fill_1 FILLER_18_2549 ();
 sg13g2_decap_8 FILLER_18_2569 ();
 sg13g2_decap_8 FILLER_18_2576 ();
 sg13g2_decap_4 FILLER_18_2583 ();
 sg13g2_fill_1 FILLER_18_2587 ();
 sg13g2_fill_1 FILLER_18_2592 ();
 sg13g2_decap_4 FILLER_18_2610 ();
 sg13g2_decap_8 FILLER_18_2621 ();
 sg13g2_decap_8 FILLER_18_2628 ();
 sg13g2_fill_2 FILLER_18_2635 ();
 sg13g2_fill_2 FILLER_18_2655 ();
 sg13g2_fill_1 FILLER_18_2657 ();
 sg13g2_decap_8 FILLER_18_2671 ();
 sg13g2_decap_8 FILLER_18_2678 ();
 sg13g2_fill_1 FILLER_18_2689 ();
 sg13g2_decap_4 FILLER_18_2695 ();
 sg13g2_fill_2 FILLER_18_2723 ();
 sg13g2_fill_1 FILLER_18_2725 ();
 sg13g2_decap_8 FILLER_18_2749 ();
 sg13g2_fill_1 FILLER_18_2756 ();
 sg13g2_fill_2 FILLER_18_2766 ();
 sg13g2_fill_1 FILLER_18_2768 ();
 sg13g2_fill_2 FILLER_18_2774 ();
 sg13g2_fill_1 FILLER_18_2776 ();
 sg13g2_fill_2 FILLER_18_2811 ();
 sg13g2_fill_2 FILLER_18_2821 ();
 sg13g2_fill_1 FILLER_18_2876 ();
 sg13g2_decap_8 FILLER_18_2881 ();
 sg13g2_decap_4 FILLER_18_2888 ();
 sg13g2_fill_1 FILLER_18_2892 ();
 sg13g2_decap_4 FILLER_18_2935 ();
 sg13g2_fill_2 FILLER_18_2939 ();
 sg13g2_fill_2 FILLER_18_2950 ();
 sg13g2_fill_1 FILLER_18_2952 ();
 sg13g2_decap_8 FILLER_18_2965 ();
 sg13g2_decap_8 FILLER_18_2972 ();
 sg13g2_fill_1 FILLER_18_2979 ();
 sg13g2_decap_4 FILLER_18_3000 ();
 sg13g2_fill_1 FILLER_18_3015 ();
 sg13g2_fill_2 FILLER_18_3032 ();
 sg13g2_fill_2 FILLER_18_3052 ();
 sg13g2_fill_2 FILLER_18_3075 ();
 sg13g2_fill_1 FILLER_18_3077 ();
 sg13g2_fill_2 FILLER_18_3090 ();
 sg13g2_decap_4 FILLER_18_3110 ();
 sg13g2_fill_2 FILLER_18_3114 ();
 sg13g2_decap_8 FILLER_18_3123 ();
 sg13g2_decap_8 FILLER_18_3130 ();
 sg13g2_fill_2 FILLER_18_3137 ();
 sg13g2_fill_1 FILLER_18_3139 ();
 sg13g2_decap_8 FILLER_18_3161 ();
 sg13g2_fill_1 FILLER_18_3168 ();
 sg13g2_fill_1 FILLER_18_3174 ();
 sg13g2_fill_2 FILLER_18_3183 ();
 sg13g2_fill_1 FILLER_18_3185 ();
 sg13g2_fill_1 FILLER_18_3194 ();
 sg13g2_fill_1 FILLER_18_3203 ();
 sg13g2_decap_8 FILLER_18_3208 ();
 sg13g2_fill_2 FILLER_18_3215 ();
 sg13g2_fill_1 FILLER_18_3217 ();
 sg13g2_fill_1 FILLER_18_3267 ();
 sg13g2_fill_2 FILLER_18_3276 ();
 sg13g2_fill_1 FILLER_18_3278 ();
 sg13g2_fill_1 FILLER_18_3323 ();
 sg13g2_decap_8 FILLER_18_3332 ();
 sg13g2_decap_8 FILLER_18_3353 ();
 sg13g2_fill_1 FILLER_18_3360 ();
 sg13g2_fill_1 FILLER_18_3365 ();
 sg13g2_decap_8 FILLER_18_3371 ();
 sg13g2_decap_8 FILLER_18_3378 ();
 sg13g2_decap_8 FILLER_18_3389 ();
 sg13g2_decap_8 FILLER_18_3409 ();
 sg13g2_decap_4 FILLER_18_3416 ();
 sg13g2_decap_4 FILLER_18_3424 ();
 sg13g2_fill_2 FILLER_18_3428 ();
 sg13g2_decap_8 FILLER_18_3443 ();
 sg13g2_fill_2 FILLER_18_3476 ();
 sg13g2_fill_1 FILLER_18_3478 ();
 sg13g2_fill_1 FILLER_18_3497 ();
 sg13g2_fill_2 FILLER_18_3503 ();
 sg13g2_fill_1 FILLER_18_3505 ();
 sg13g2_fill_1 FILLER_18_3511 ();
 sg13g2_decap_8 FILLER_18_3516 ();
 sg13g2_decap_8 FILLER_18_3523 ();
 sg13g2_decap_8 FILLER_18_3530 ();
 sg13g2_decap_8 FILLER_18_3537 ();
 sg13g2_decap_8 FILLER_18_3544 ();
 sg13g2_decap_8 FILLER_18_3551 ();
 sg13g2_decap_8 FILLER_18_3558 ();
 sg13g2_decap_8 FILLER_18_3565 ();
 sg13g2_decap_8 FILLER_18_3572 ();
 sg13g2_fill_1 FILLER_18_3579 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_fill_1 FILLER_19_104 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_decap_4 FILLER_19_157 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_decap_4 FILLER_19_251 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_decap_4 FILLER_19_297 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_370 ();
 sg13g2_fill_2 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_1 FILLER_19_406 ();
 sg13g2_fill_2 FILLER_19_435 ();
 sg13g2_fill_1 FILLER_19_437 ();
 sg13g2_decap_4 FILLER_19_442 ();
 sg13g2_fill_2 FILLER_19_446 ();
 sg13g2_fill_2 FILLER_19_461 ();
 sg13g2_fill_1 FILLER_19_463 ();
 sg13g2_fill_1 FILLER_19_477 ();
 sg13g2_fill_1 FILLER_19_533 ();
 sg13g2_fill_2 FILLER_19_547 ();
 sg13g2_fill_1 FILLER_19_549 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_fill_1 FILLER_19_574 ();
 sg13g2_fill_1 FILLER_19_603 ();
 sg13g2_decap_4 FILLER_19_648 ();
 sg13g2_decap_8 FILLER_19_681 ();
 sg13g2_fill_2 FILLER_19_696 ();
 sg13g2_fill_1 FILLER_19_698 ();
 sg13g2_fill_1 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_4 FILLER_19_749 ();
 sg13g2_decap_4 FILLER_19_766 ();
 sg13g2_fill_1 FILLER_19_770 ();
 sg13g2_fill_2 FILLER_19_781 ();
 sg13g2_fill_1 FILLER_19_783 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_decap_8 FILLER_19_809 ();
 sg13g2_fill_2 FILLER_19_844 ();
 sg13g2_decap_8 FILLER_19_865 ();
 sg13g2_fill_2 FILLER_19_872 ();
 sg13g2_fill_1 FILLER_19_874 ();
 sg13g2_fill_1 FILLER_19_879 ();
 sg13g2_decap_8 FILLER_19_893 ();
 sg13g2_fill_2 FILLER_19_900 ();
 sg13g2_fill_1 FILLER_19_902 ();
 sg13g2_fill_1 FILLER_19_922 ();
 sg13g2_decap_4 FILLER_19_927 ();
 sg13g2_decap_8 FILLER_19_943 ();
 sg13g2_decap_8 FILLER_19_950 ();
 sg13g2_decap_8 FILLER_19_957 ();
 sg13g2_decap_8 FILLER_19_964 ();
 sg13g2_decap_8 FILLER_19_971 ();
 sg13g2_decap_8 FILLER_19_978 ();
 sg13g2_decap_4 FILLER_19_985 ();
 sg13g2_decap_8 FILLER_19_998 ();
 sg13g2_decap_8 FILLER_19_1005 ();
 sg13g2_decap_8 FILLER_19_1012 ();
 sg13g2_decap_8 FILLER_19_1019 ();
 sg13g2_decap_8 FILLER_19_1039 ();
 sg13g2_fill_1 FILLER_19_1054 ();
 sg13g2_fill_2 FILLER_19_1070 ();
 sg13g2_fill_1 FILLER_19_1072 ();
 sg13g2_decap_8 FILLER_19_1077 ();
 sg13g2_decap_8 FILLER_19_1084 ();
 sg13g2_fill_2 FILLER_19_1091 ();
 sg13g2_fill_1 FILLER_19_1093 ();
 sg13g2_fill_2 FILLER_19_1099 ();
 sg13g2_fill_2 FILLER_19_1106 ();
 sg13g2_decap_8 FILLER_19_1116 ();
 sg13g2_fill_1 FILLER_19_1123 ();
 sg13g2_decap_8 FILLER_19_1129 ();
 sg13g2_decap_8 FILLER_19_1136 ();
 sg13g2_decap_8 FILLER_19_1143 ();
 sg13g2_decap_8 FILLER_19_1150 ();
 sg13g2_decap_8 FILLER_19_1157 ();
 sg13g2_fill_2 FILLER_19_1164 ();
 sg13g2_decap_8 FILLER_19_1212 ();
 sg13g2_decap_4 FILLER_19_1228 ();
 sg13g2_decap_4 FILLER_19_1250 ();
 sg13g2_fill_2 FILLER_19_1254 ();
 sg13g2_fill_2 FILLER_19_1260 ();
 sg13g2_decap_8 FILLER_19_1266 ();
 sg13g2_fill_2 FILLER_19_1273 ();
 sg13g2_fill_1 FILLER_19_1275 ();
 sg13g2_fill_2 FILLER_19_1289 ();
 sg13g2_fill_1 FILLER_19_1291 ();
 sg13g2_decap_4 FILLER_19_1319 ();
 sg13g2_fill_1 FILLER_19_1323 ();
 sg13g2_decap_4 FILLER_19_1355 ();
 sg13g2_fill_1 FILLER_19_1359 ();
 sg13g2_fill_2 FILLER_19_1393 ();
 sg13g2_fill_1 FILLER_19_1395 ();
 sg13g2_decap_8 FILLER_19_1430 ();
 sg13g2_decap_4 FILLER_19_1482 ();
 sg13g2_fill_2 FILLER_19_1486 ();
 sg13g2_decap_8 FILLER_19_1520 ();
 sg13g2_decap_4 FILLER_19_1527 ();
 sg13g2_fill_2 FILLER_19_1531 ();
 sg13g2_fill_2 FILLER_19_1541 ();
 sg13g2_fill_2 FILLER_19_1556 ();
 sg13g2_fill_1 FILLER_19_1558 ();
 sg13g2_decap_4 FILLER_19_1575 ();
 sg13g2_decap_4 FILLER_19_1599 ();
 sg13g2_fill_1 FILLER_19_1603 ();
 sg13g2_fill_1 FILLER_19_1608 ();
 sg13g2_fill_2 FILLER_19_1628 ();
 sg13g2_decap_4 FILLER_19_1653 ();
 sg13g2_fill_2 FILLER_19_1657 ();
 sg13g2_decap_8 FILLER_19_1680 ();
 sg13g2_fill_2 FILLER_19_1687 ();
 sg13g2_decap_4 FILLER_19_1694 ();
 sg13g2_fill_2 FILLER_19_1698 ();
 sg13g2_decap_4 FILLER_19_1715 ();
 sg13g2_fill_1 FILLER_19_1732 ();
 sg13g2_decap_8 FILLER_19_1738 ();
 sg13g2_fill_2 FILLER_19_1745 ();
 sg13g2_fill_1 FILLER_19_1747 ();
 sg13g2_fill_1 FILLER_19_1752 ();
 sg13g2_fill_1 FILLER_19_1774 ();
 sg13g2_fill_2 FILLER_19_1787 ();
 sg13g2_fill_1 FILLER_19_1789 ();
 sg13g2_fill_1 FILLER_19_1823 ();
 sg13g2_decap_8 FILLER_19_1852 ();
 sg13g2_decap_8 FILLER_19_1859 ();
 sg13g2_fill_1 FILLER_19_1866 ();
 sg13g2_fill_1 FILLER_19_1871 ();
 sg13g2_fill_2 FILLER_19_1877 ();
 sg13g2_fill_1 FILLER_19_1879 ();
 sg13g2_fill_1 FILLER_19_1892 ();
 sg13g2_decap_4 FILLER_19_1915 ();
 sg13g2_fill_1 FILLER_19_1926 ();
 sg13g2_fill_2 FILLER_19_1940 ();
 sg13g2_fill_1 FILLER_19_1942 ();
 sg13g2_fill_1 FILLER_19_1947 ();
 sg13g2_decap_8 FILLER_19_1952 ();
 sg13g2_decap_4 FILLER_19_1959 ();
 sg13g2_fill_2 FILLER_19_1963 ();
 sg13g2_decap_8 FILLER_19_1975 ();
 sg13g2_decap_8 FILLER_19_1999 ();
 sg13g2_decap_4 FILLER_19_2006 ();
 sg13g2_fill_1 FILLER_19_2010 ();
 sg13g2_decap_8 FILLER_19_2019 ();
 sg13g2_decap_4 FILLER_19_2026 ();
 sg13g2_decap_8 FILLER_19_2041 ();
 sg13g2_decap_4 FILLER_19_2048 ();
 sg13g2_decap_8 FILLER_19_2062 ();
 sg13g2_decap_4 FILLER_19_2069 ();
 sg13g2_fill_2 FILLER_19_2073 ();
 sg13g2_decap_8 FILLER_19_2079 ();
 sg13g2_fill_1 FILLER_19_2086 ();
 sg13g2_fill_1 FILLER_19_2100 ();
 sg13g2_decap_8 FILLER_19_2166 ();
 sg13g2_decap_8 FILLER_19_2173 ();
 sg13g2_decap_8 FILLER_19_2180 ();
 sg13g2_fill_2 FILLER_19_2190 ();
 sg13g2_decap_8 FILLER_19_2196 ();
 sg13g2_decap_8 FILLER_19_2203 ();
 sg13g2_decap_4 FILLER_19_2210 ();
 sg13g2_fill_2 FILLER_19_2214 ();
 sg13g2_decap_4 FILLER_19_2231 ();
 sg13g2_fill_2 FILLER_19_2235 ();
 sg13g2_decap_4 FILLER_19_2261 ();
 sg13g2_fill_2 FILLER_19_2265 ();
 sg13g2_fill_2 FILLER_19_2302 ();
 sg13g2_fill_1 FILLER_19_2304 ();
 sg13g2_decap_4 FILLER_19_2324 ();
 sg13g2_fill_1 FILLER_19_2328 ();
 sg13g2_fill_1 FILLER_19_2334 ();
 sg13g2_decap_4 FILLER_19_2339 ();
 sg13g2_fill_1 FILLER_19_2343 ();
 sg13g2_fill_2 FILLER_19_2352 ();
 sg13g2_decap_8 FILLER_19_2373 ();
 sg13g2_decap_8 FILLER_19_2390 ();
 sg13g2_fill_1 FILLER_19_2397 ();
 sg13g2_decap_8 FILLER_19_2403 ();
 sg13g2_decap_4 FILLER_19_2432 ();
 sg13g2_fill_2 FILLER_19_2436 ();
 sg13g2_decap_8 FILLER_19_2460 ();
 sg13g2_decap_4 FILLER_19_2467 ();
 sg13g2_fill_1 FILLER_19_2471 ();
 sg13g2_decap_4 FILLER_19_2503 ();
 sg13g2_fill_2 FILLER_19_2507 ();
 sg13g2_decap_4 FILLER_19_2527 ();
 sg13g2_fill_2 FILLER_19_2568 ();
 sg13g2_fill_2 FILLER_19_2611 ();
 sg13g2_fill_1 FILLER_19_2613 ();
 sg13g2_decap_4 FILLER_19_2642 ();
 sg13g2_fill_2 FILLER_19_2646 ();
 sg13g2_fill_1 FILLER_19_2664 ();
 sg13g2_decap_8 FILLER_19_2676 ();
 sg13g2_decap_8 FILLER_19_2683 ();
 sg13g2_fill_2 FILLER_19_2690 ();
 sg13g2_decap_8 FILLER_19_2696 ();
 sg13g2_fill_1 FILLER_19_2703 ();
 sg13g2_decap_8 FILLER_19_2721 ();
 sg13g2_decap_4 FILLER_19_2728 ();
 sg13g2_fill_1 FILLER_19_2732 ();
 sg13g2_fill_2 FILLER_19_2738 ();
 sg13g2_fill_1 FILLER_19_2740 ();
 sg13g2_decap_8 FILLER_19_2746 ();
 sg13g2_decap_4 FILLER_19_2753 ();
 sg13g2_fill_2 FILLER_19_2777 ();
 sg13g2_fill_1 FILLER_19_2779 ();
 sg13g2_fill_2 FILLER_19_2796 ();
 sg13g2_decap_8 FILLER_19_2803 ();
 sg13g2_fill_2 FILLER_19_2810 ();
 sg13g2_decap_4 FILLER_19_2838 ();
 sg13g2_fill_2 FILLER_19_2842 ();
 sg13g2_fill_2 FILLER_19_2849 ();
 sg13g2_fill_1 FILLER_19_2861 ();
 sg13g2_fill_2 FILLER_19_2880 ();
 sg13g2_fill_2 FILLER_19_2895 ();
 sg13g2_decap_8 FILLER_19_2914 ();
 sg13g2_fill_1 FILLER_19_2921 ();
 sg13g2_fill_2 FILLER_19_2930 ();
 sg13g2_fill_1 FILLER_19_2949 ();
 sg13g2_fill_2 FILLER_19_2954 ();
 sg13g2_fill_1 FILLER_19_2956 ();
 sg13g2_fill_1 FILLER_19_2962 ();
 sg13g2_decap_4 FILLER_19_2968 ();
 sg13g2_fill_2 FILLER_19_2972 ();
 sg13g2_decap_8 FILLER_19_2983 ();
 sg13g2_fill_1 FILLER_19_2995 ();
 sg13g2_decap_8 FILLER_19_3000 ();
 sg13g2_decap_4 FILLER_19_3007 ();
 sg13g2_decap_8 FILLER_19_3030 ();
 sg13g2_fill_2 FILLER_19_3037 ();
 sg13g2_fill_2 FILLER_19_3048 ();
 sg13g2_decap_8 FILLER_19_3054 ();
 sg13g2_fill_1 FILLER_19_3061 ();
 sg13g2_decap_4 FILLER_19_3083 ();
 sg13g2_decap_4 FILLER_19_3091 ();
 sg13g2_fill_1 FILLER_19_3095 ();
 sg13g2_decap_8 FILLER_19_3111 ();
 sg13g2_fill_1 FILLER_19_3118 ();
 sg13g2_fill_1 FILLER_19_3124 ();
 sg13g2_fill_1 FILLER_19_3130 ();
 sg13g2_decap_4 FILLER_19_3144 ();
 sg13g2_fill_1 FILLER_19_3148 ();
 sg13g2_decap_8 FILLER_19_3167 ();
 sg13g2_decap_4 FILLER_19_3174 ();
 sg13g2_fill_2 FILLER_19_3178 ();
 sg13g2_fill_1 FILLER_19_3192 ();
 sg13g2_decap_8 FILLER_19_3204 ();
 sg13g2_decap_8 FILLER_19_3211 ();
 sg13g2_fill_1 FILLER_19_3232 ();
 sg13g2_decap_4 FILLER_19_3246 ();
 sg13g2_fill_1 FILLER_19_3250 ();
 sg13g2_fill_2 FILLER_19_3260 ();
 sg13g2_fill_1 FILLER_19_3262 ();
 sg13g2_decap_4 FILLER_19_3274 ();
 sg13g2_fill_2 FILLER_19_3278 ();
 sg13g2_decap_4 FILLER_19_3298 ();
 sg13g2_fill_1 FILLER_19_3302 ();
 sg13g2_decap_4 FILLER_19_3323 ();
 sg13g2_fill_2 FILLER_19_3327 ();
 sg13g2_fill_1 FILLER_19_3338 ();
 sg13g2_fill_2 FILLER_19_3393 ();
 sg13g2_fill_1 FILLER_19_3395 ();
 sg13g2_decap_8 FILLER_19_3416 ();
 sg13g2_decap_8 FILLER_19_3423 ();
 sg13g2_decap_8 FILLER_19_3430 ();
 sg13g2_fill_1 FILLER_19_3437 ();
 sg13g2_decap_4 FILLER_19_3459 ();
 sg13g2_fill_2 FILLER_19_3463 ();
 sg13g2_fill_1 FILLER_19_3474 ();
 sg13g2_fill_2 FILLER_19_3480 ();
 sg13g2_fill_1 FILLER_19_3482 ();
 sg13g2_fill_1 FILLER_19_3491 ();
 sg13g2_fill_2 FILLER_19_3496 ();
 sg13g2_fill_1 FILLER_19_3498 ();
 sg13g2_decap_8 FILLER_19_3514 ();
 sg13g2_decap_8 FILLER_19_3521 ();
 sg13g2_decap_8 FILLER_19_3528 ();
 sg13g2_decap_8 FILLER_19_3535 ();
 sg13g2_decap_8 FILLER_19_3542 ();
 sg13g2_decap_8 FILLER_19_3549 ();
 sg13g2_decap_8 FILLER_19_3556 ();
 sg13g2_decap_8 FILLER_19_3563 ();
 sg13g2_decap_8 FILLER_19_3570 ();
 sg13g2_fill_2 FILLER_19_3577 ();
 sg13g2_fill_1 FILLER_19_3579 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_4 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_52 ();
 sg13g2_decap_4 FILLER_20_59 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_122 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_163 ();
 sg13g2_decap_8 FILLER_20_176 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_215 ();
 sg13g2_decap_4 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_decap_4 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_decap_8 FILLER_20_288 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_2 FILLER_20_318 ();
 sg13g2_fill_2 FILLER_20_329 ();
 sg13g2_fill_1 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_345 ();
 sg13g2_fill_2 FILLER_20_365 ();
 sg13g2_fill_2 FILLER_20_383 ();
 sg13g2_fill_2 FILLER_20_398 ();
 sg13g2_fill_1 FILLER_20_400 ();
 sg13g2_fill_1 FILLER_20_414 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_fill_1 FILLER_20_430 ();
 sg13g2_decap_8 FILLER_20_457 ();
 sg13g2_fill_2 FILLER_20_464 ();
 sg13g2_fill_1 FILLER_20_466 ();
 sg13g2_fill_1 FILLER_20_480 ();
 sg13g2_fill_2 FILLER_20_485 ();
 sg13g2_fill_1 FILLER_20_499 ();
 sg13g2_decap_4 FILLER_20_517 ();
 sg13g2_fill_1 FILLER_20_521 ();
 sg13g2_decap_4 FILLER_20_526 ();
 sg13g2_fill_1 FILLER_20_530 ();
 sg13g2_fill_2 FILLER_20_535 ();
 sg13g2_fill_2 FILLER_20_545 ();
 sg13g2_fill_2 FILLER_20_556 ();
 sg13g2_fill_1 FILLER_20_558 ();
 sg13g2_decap_8 FILLER_20_563 ();
 sg13g2_decap_4 FILLER_20_570 ();
 sg13g2_fill_1 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_604 ();
 sg13g2_decap_8 FILLER_20_611 ();
 sg13g2_fill_2 FILLER_20_657 ();
 sg13g2_fill_1 FILLER_20_659 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_fill_1 FILLER_20_679 ();
 sg13g2_fill_2 FILLER_20_693 ();
 sg13g2_fill_1 FILLER_20_695 ();
 sg13g2_decap_4 FILLER_20_717 ();
 sg13g2_fill_1 FILLER_20_729 ();
 sg13g2_decap_4 FILLER_20_738 ();
 sg13g2_fill_1 FILLER_20_747 ();
 sg13g2_fill_2 FILLER_20_761 ();
 sg13g2_fill_2 FILLER_20_783 ();
 sg13g2_fill_1 FILLER_20_785 ();
 sg13g2_fill_2 FILLER_20_797 ();
 sg13g2_fill_1 FILLER_20_799 ();
 sg13g2_fill_2 FILLER_20_817 ();
 sg13g2_decap_8 FILLER_20_837 ();
 sg13g2_decap_4 FILLER_20_844 ();
 sg13g2_decap_8 FILLER_20_867 ();
 sg13g2_fill_2 FILLER_20_895 ();
 sg13g2_fill_2 FILLER_20_910 ();
 sg13g2_fill_2 FILLER_20_922 ();
 sg13g2_fill_2 FILLER_20_954 ();
 sg13g2_fill_1 FILLER_20_956 ();
 sg13g2_fill_2 FILLER_20_971 ();
 sg13g2_decap_8 FILLER_20_986 ();
 sg13g2_decap_4 FILLER_20_1001 ();
 sg13g2_fill_1 FILLER_20_1023 ();
 sg13g2_decap_8 FILLER_20_1034 ();
 sg13g2_decap_4 FILLER_20_1041 ();
 sg13g2_fill_1 FILLER_20_1045 ();
 sg13g2_decap_8 FILLER_20_1054 ();
 sg13g2_fill_1 FILLER_20_1061 ();
 sg13g2_fill_1 FILLER_20_1088 ();
 sg13g2_decap_8 FILLER_20_1136 ();
 sg13g2_decap_4 FILLER_20_1159 ();
 sg13g2_fill_1 FILLER_20_1189 ();
 sg13g2_fill_2 FILLER_20_1195 ();
 sg13g2_fill_1 FILLER_20_1197 ();
 sg13g2_fill_2 FILLER_20_1206 ();
 sg13g2_fill_1 FILLER_20_1208 ();
 sg13g2_fill_2 FILLER_20_1225 ();
 sg13g2_decap_4 FILLER_20_1232 ();
 sg13g2_decap_4 FILLER_20_1241 ();
 sg13g2_fill_2 FILLER_20_1245 ();
 sg13g2_fill_2 FILLER_20_1251 ();
 sg13g2_decap_4 FILLER_20_1257 ();
 sg13g2_fill_1 FILLER_20_1261 ();
 sg13g2_decap_4 FILLER_20_1271 ();
 sg13g2_fill_1 FILLER_20_1303 ();
 sg13g2_decap_8 FILLER_20_1309 ();
 sg13g2_decap_4 FILLER_20_1316 ();
 sg13g2_fill_2 FILLER_20_1320 ();
 sg13g2_decap_4 FILLER_20_1343 ();
 sg13g2_fill_2 FILLER_20_1347 ();
 sg13g2_decap_8 FILLER_20_1358 ();
 sg13g2_fill_2 FILLER_20_1365 ();
 sg13g2_fill_1 FILLER_20_1367 ();
 sg13g2_fill_1 FILLER_20_1392 ();
 sg13g2_fill_1 FILLER_20_1398 ();
 sg13g2_fill_2 FILLER_20_1404 ();
 sg13g2_fill_1 FILLER_20_1406 ();
 sg13g2_decap_4 FILLER_20_1423 ();
 sg13g2_fill_2 FILLER_20_1431 ();
 sg13g2_decap_4 FILLER_20_1467 ();
 sg13g2_decap_8 FILLER_20_1484 ();
 sg13g2_fill_1 FILLER_20_1491 ();
 sg13g2_fill_1 FILLER_20_1505 ();
 sg13g2_decap_8 FILLER_20_1514 ();
 sg13g2_decap_4 FILLER_20_1521 ();
 sg13g2_fill_2 FILLER_20_1525 ();
 sg13g2_fill_1 FILLER_20_1548 ();
 sg13g2_fill_2 FILLER_20_1564 ();
 sg13g2_decap_4 FILLER_20_1574 ();
 sg13g2_fill_2 FILLER_20_1578 ();
 sg13g2_fill_2 FILLER_20_1587 ();
 sg13g2_fill_2 FILLER_20_1610 ();
 sg13g2_fill_2 FILLER_20_1624 ();
 sg13g2_fill_2 FILLER_20_1634 ();
 sg13g2_fill_1 FILLER_20_1636 ();
 sg13g2_decap_8 FILLER_20_1655 ();
 sg13g2_fill_2 FILLER_20_1662 ();
 sg13g2_decap_8 FILLER_20_1682 ();
 sg13g2_decap_8 FILLER_20_1689 ();
 sg13g2_fill_1 FILLER_20_1696 ();
 sg13g2_fill_1 FILLER_20_1705 ();
 sg13g2_decap_8 FILLER_20_1710 ();
 sg13g2_fill_2 FILLER_20_1717 ();
 sg13g2_fill_1 FILLER_20_1719 ();
 sg13g2_decap_4 FILLER_20_1740 ();
 sg13g2_fill_1 FILLER_20_1766 ();
 sg13g2_fill_2 FILLER_20_1772 ();
 sg13g2_fill_1 FILLER_20_1774 ();
 sg13g2_decap_8 FILLER_20_1780 ();
 sg13g2_fill_2 FILLER_20_1792 ();
 sg13g2_decap_8 FILLER_20_1799 ();
 sg13g2_decap_8 FILLER_20_1806 ();
 sg13g2_fill_2 FILLER_20_1818 ();
 sg13g2_decap_8 FILLER_20_1830 ();
 sg13g2_fill_2 FILLER_20_1837 ();
 sg13g2_decap_4 FILLER_20_1853 ();
 sg13g2_decap_8 FILLER_20_1875 ();
 sg13g2_decap_8 FILLER_20_1882 ();
 sg13g2_fill_2 FILLER_20_1889 ();
 sg13g2_fill_2 FILLER_20_1900 ();
 sg13g2_fill_2 FILLER_20_1924 ();
 sg13g2_fill_2 FILLER_20_1952 ();
 sg13g2_fill_1 FILLER_20_1985 ();
 sg13g2_decap_8 FILLER_20_2006 ();
 sg13g2_fill_1 FILLER_20_2013 ();
 sg13g2_fill_2 FILLER_20_2024 ();
 sg13g2_fill_1 FILLER_20_2039 ();
 sg13g2_fill_2 FILLER_20_2045 ();
 sg13g2_fill_2 FILLER_20_2060 ();
 sg13g2_decap_8 FILLER_20_2080 ();
 sg13g2_decap_4 FILLER_20_2091 ();
 sg13g2_fill_2 FILLER_20_2107 ();
 sg13g2_fill_2 FILLER_20_2124 ();
 sg13g2_decap_4 FILLER_20_2161 ();
 sg13g2_fill_1 FILLER_20_2170 ();
 sg13g2_decap_8 FILLER_20_2180 ();
 sg13g2_decap_4 FILLER_20_2187 ();
 sg13g2_fill_2 FILLER_20_2191 ();
 sg13g2_fill_2 FILLER_20_2198 ();
 sg13g2_decap_8 FILLER_20_2205 ();
 sg13g2_decap_8 FILLER_20_2212 ();
 sg13g2_decap_8 FILLER_20_2237 ();
 sg13g2_decap_4 FILLER_20_2244 ();
 sg13g2_fill_1 FILLER_20_2248 ();
 sg13g2_fill_2 FILLER_20_2270 ();
 sg13g2_fill_2 FILLER_20_2276 ();
 sg13g2_fill_1 FILLER_20_2291 ();
 sg13g2_decap_4 FILLER_20_2308 ();
 sg13g2_decap_8 FILLER_20_2318 ();
 sg13g2_fill_1 FILLER_20_2325 ();
 sg13g2_decap_8 FILLER_20_2355 ();
 sg13g2_fill_2 FILLER_20_2362 ();
 sg13g2_fill_1 FILLER_20_2364 ();
 sg13g2_fill_2 FILLER_20_2386 ();
 sg13g2_fill_2 FILLER_20_2392 ();
 sg13g2_fill_2 FILLER_20_2443 ();
 sg13g2_fill_1 FILLER_20_2445 ();
 sg13g2_fill_1 FILLER_20_2450 ();
 sg13g2_fill_2 FILLER_20_2461 ();
 sg13g2_fill_1 FILLER_20_2463 ();
 sg13g2_decap_4 FILLER_20_2467 ();
 sg13g2_decap_8 FILLER_20_2499 ();
 sg13g2_decap_8 FILLER_20_2506 ();
 sg13g2_decap_4 FILLER_20_2513 ();
 sg13g2_fill_1 FILLER_20_2522 ();
 sg13g2_decap_8 FILLER_20_2537 ();
 sg13g2_decap_4 FILLER_20_2544 ();
 sg13g2_fill_2 FILLER_20_2548 ();
 sg13g2_fill_2 FILLER_20_2553 ();
 sg13g2_fill_1 FILLER_20_2555 ();
 sg13g2_decap_8 FILLER_20_2569 ();
 sg13g2_decap_4 FILLER_20_2576 ();
 sg13g2_fill_2 FILLER_20_2593 ();
 sg13g2_fill_1 FILLER_20_2595 ();
 sg13g2_decap_8 FILLER_20_2604 ();
 sg13g2_decap_8 FILLER_20_2611 ();
 sg13g2_fill_1 FILLER_20_2618 ();
 sg13g2_decap_4 FILLER_20_2623 ();
 sg13g2_fill_2 FILLER_20_2627 ();
 sg13g2_decap_8 FILLER_20_2634 ();
 sg13g2_decap_8 FILLER_20_2641 ();
 sg13g2_fill_1 FILLER_20_2648 ();
 sg13g2_fill_2 FILLER_20_2685 ();
 sg13g2_decap_8 FILLER_20_2715 ();
 sg13g2_decap_4 FILLER_20_2722 ();
 sg13g2_decap_4 FILLER_20_2758 ();
 sg13g2_fill_1 FILLER_20_2762 ();
 sg13g2_decap_8 FILLER_20_2788 ();
 sg13g2_fill_1 FILLER_20_2795 ();
 sg13g2_fill_2 FILLER_20_2815 ();
 sg13g2_decap_4 FILLER_20_2840 ();
 sg13g2_fill_1 FILLER_20_2844 ();
 sg13g2_fill_2 FILLER_20_2863 ();
 sg13g2_fill_1 FILLER_20_2865 ();
 sg13g2_decap_8 FILLER_20_2886 ();
 sg13g2_decap_8 FILLER_20_2893 ();
 sg13g2_fill_1 FILLER_20_2908 ();
 sg13g2_fill_1 FILLER_20_2917 ();
 sg13g2_decap_8 FILLER_20_2931 ();
 sg13g2_fill_2 FILLER_20_2938 ();
 sg13g2_fill_1 FILLER_20_2949 ();
 sg13g2_decap_8 FILLER_20_3004 ();
 sg13g2_fill_1 FILLER_20_3011 ();
 sg13g2_fill_1 FILLER_20_3035 ();
 sg13g2_decap_8 FILLER_20_3058 ();
 sg13g2_decap_8 FILLER_20_3065 ();
 sg13g2_fill_1 FILLER_20_3086 ();
 sg13g2_fill_2 FILLER_20_3117 ();
 sg13g2_fill_2 FILLER_20_3145 ();
 sg13g2_fill_1 FILLER_20_3147 ();
 sg13g2_fill_1 FILLER_20_3166 ();
 sg13g2_decap_8 FILLER_20_3189 ();
 sg13g2_fill_1 FILLER_20_3216 ();
 sg13g2_fill_2 FILLER_20_3257 ();
 sg13g2_decap_8 FILLER_20_3281 ();
 sg13g2_decap_8 FILLER_20_3288 ();
 sg13g2_fill_2 FILLER_20_3295 ();
 sg13g2_fill_2 FILLER_20_3308 ();
 sg13g2_decap_8 FILLER_20_3328 ();
 sg13g2_fill_2 FILLER_20_3335 ();
 sg13g2_fill_1 FILLER_20_3337 ();
 sg13g2_decap_4 FILLER_20_3342 ();
 sg13g2_decap_8 FILLER_20_3367 ();
 sg13g2_decap_4 FILLER_20_3374 ();
 sg13g2_decap_8 FILLER_20_3390 ();
 sg13g2_decap_8 FILLER_20_3414 ();
 sg13g2_decap_8 FILLER_20_3421 ();
 sg13g2_fill_2 FILLER_20_3438 ();
 sg13g2_fill_2 FILLER_20_3462 ();
 sg13g2_fill_2 FILLER_20_3501 ();
 sg13g2_fill_1 FILLER_20_3503 ();
 sg13g2_decap_8 FILLER_20_3523 ();
 sg13g2_decap_8 FILLER_20_3530 ();
 sg13g2_decap_8 FILLER_20_3537 ();
 sg13g2_decap_8 FILLER_20_3544 ();
 sg13g2_decap_8 FILLER_20_3551 ();
 sg13g2_decap_8 FILLER_20_3558 ();
 sg13g2_decap_8 FILLER_20_3565 ();
 sg13g2_decap_8 FILLER_20_3572 ();
 sg13g2_fill_1 FILLER_20_3579 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_94 ();
 sg13g2_decap_4 FILLER_21_101 ();
 sg13g2_fill_2 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_164 ();
 sg13g2_fill_1 FILLER_21_178 ();
 sg13g2_decap_4 FILLER_21_189 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_fill_1 FILLER_21_215 ();
 sg13g2_decap_4 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_245 ();
 sg13g2_decap_4 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_299 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_21_353 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_375 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_fill_1 FILLER_21_409 ();
 sg13g2_fill_2 FILLER_21_436 ();
 sg13g2_fill_2 FILLER_21_451 ();
 sg13g2_fill_1 FILLER_21_453 ();
 sg13g2_fill_2 FILLER_21_467 ();
 sg13g2_decap_4 FILLER_21_482 ();
 sg13g2_fill_1 FILLER_21_486 ();
 sg13g2_fill_2 FILLER_21_503 ();
 sg13g2_fill_1 FILLER_21_505 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_4 FILLER_21_518 ();
 sg13g2_decap_4 FILLER_21_527 ();
 sg13g2_fill_2 FILLER_21_531 ();
 sg13g2_fill_2 FILLER_21_561 ();
 sg13g2_fill_2 FILLER_21_593 ();
 sg13g2_fill_2 FILLER_21_599 ();
 sg13g2_fill_1 FILLER_21_613 ();
 sg13g2_decap_4 FILLER_21_627 ();
 sg13g2_fill_1 FILLER_21_631 ();
 sg13g2_decap_4 FILLER_21_650 ();
 sg13g2_fill_2 FILLER_21_654 ();
 sg13g2_fill_2 FILLER_21_700 ();
 sg13g2_fill_2 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_744 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_fill_2 FILLER_21_770 ();
 sg13g2_fill_1 FILLER_21_772 ();
 sg13g2_fill_1 FILLER_21_783 ();
 sg13g2_decap_8 FILLER_21_797 ();
 sg13g2_fill_2 FILLER_21_822 ();
 sg13g2_fill_2 FILLER_21_828 ();
 sg13g2_fill_1 FILLER_21_830 ();
 sg13g2_decap_4 FILLER_21_836 ();
 sg13g2_fill_2 FILLER_21_840 ();
 sg13g2_fill_1 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_867 ();
 sg13g2_fill_2 FILLER_21_900 ();
 sg13g2_decap_8 FILLER_21_923 ();
 sg13g2_fill_2 FILLER_21_930 ();
 sg13g2_fill_2 FILLER_21_938 ();
 sg13g2_decap_4 FILLER_21_945 ();
 sg13g2_fill_1 FILLER_21_949 ();
 sg13g2_fill_2 FILLER_21_974 ();
 sg13g2_fill_1 FILLER_21_976 ();
 sg13g2_decap_4 FILLER_21_986 ();
 sg13g2_fill_1 FILLER_21_990 ();
 sg13g2_decap_8 FILLER_21_1052 ();
 sg13g2_fill_1 FILLER_21_1068 ();
 sg13g2_fill_1 FILLER_21_1078 ();
 sg13g2_fill_1 FILLER_21_1087 ();
 sg13g2_fill_1 FILLER_21_1115 ();
 sg13g2_fill_1 FILLER_21_1119 ();
 sg13g2_fill_2 FILLER_21_1161 ();
 sg13g2_fill_1 FILLER_21_1163 ();
 sg13g2_decap_8 FILLER_21_1168 ();
 sg13g2_decap_8 FILLER_21_1175 ();
 sg13g2_decap_4 FILLER_21_1182 ();
 sg13g2_decap_8 FILLER_21_1211 ();
 sg13g2_decap_4 FILLER_21_1218 ();
 sg13g2_fill_2 FILLER_21_1222 ();
 sg13g2_decap_4 FILLER_21_1275 ();
 sg13g2_fill_1 FILLER_21_1279 ();
 sg13g2_decap_8 FILLER_21_1309 ();
 sg13g2_fill_2 FILLER_21_1316 ();
 sg13g2_fill_1 FILLER_21_1318 ();
 sg13g2_fill_1 FILLER_21_1332 ();
 sg13g2_decap_4 FILLER_21_1342 ();
 sg13g2_fill_1 FILLER_21_1346 ();
 sg13g2_decap_4 FILLER_21_1365 ();
 sg13g2_decap_4 FILLER_21_1383 ();
 sg13g2_fill_2 FILLER_21_1387 ();
 sg13g2_decap_8 FILLER_21_1404 ();
 sg13g2_decap_8 FILLER_21_1411 ();
 sg13g2_fill_1 FILLER_21_1418 ();
 sg13g2_decap_8 FILLER_21_1428 ();
 sg13g2_decap_4 FILLER_21_1435 ();
 sg13g2_fill_1 FILLER_21_1439 ();
 sg13g2_decap_4 FILLER_21_1454 ();
 sg13g2_fill_1 FILLER_21_1458 ();
 sg13g2_fill_2 FILLER_21_1472 ();
 sg13g2_fill_1 FILLER_21_1474 ();
 sg13g2_fill_2 FILLER_21_1488 ();
 sg13g2_fill_1 FILLER_21_1490 ();
 sg13g2_decap_8 FILLER_21_1508 ();
 sg13g2_decap_8 FILLER_21_1515 ();
 sg13g2_fill_2 FILLER_21_1522 ();
 sg13g2_decap_8 FILLER_21_1545 ();
 sg13g2_decap_4 FILLER_21_1568 ();
 sg13g2_fill_2 FILLER_21_1572 ();
 sg13g2_fill_2 FILLER_21_1597 ();
 sg13g2_fill_1 FILLER_21_1599 ();
 sg13g2_decap_4 FILLER_21_1618 ();
 sg13g2_fill_2 FILLER_21_1622 ();
 sg13g2_decap_8 FILLER_21_1642 ();
 sg13g2_fill_1 FILLER_21_1649 ();
 sg13g2_decap_8 FILLER_21_1655 ();
 sg13g2_fill_1 FILLER_21_1662 ();
 sg13g2_fill_2 FILLER_21_1681 ();
 sg13g2_fill_2 FILLER_21_1707 ();
 sg13g2_decap_4 FILLER_21_1737 ();
 sg13g2_fill_2 FILLER_21_1741 ();
 sg13g2_decap_4 FILLER_21_1752 ();
 sg13g2_fill_2 FILLER_21_1761 ();
 sg13g2_fill_1 FILLER_21_1776 ();
 sg13g2_fill_2 FILLER_21_1785 ();
 sg13g2_fill_2 FILLER_21_1799 ();
 sg13g2_fill_1 FILLER_21_1801 ();
 sg13g2_fill_2 FILLER_21_1812 ();
 sg13g2_fill_1 FILLER_21_1824 ();
 sg13g2_fill_2 FILLER_21_1838 ();
 sg13g2_fill_1 FILLER_21_1840 ();
 sg13g2_decap_4 FILLER_21_1869 ();
 sg13g2_decap_8 FILLER_21_1931 ();
 sg13g2_decap_4 FILLER_21_1938 ();
 sg13g2_fill_2 FILLER_21_1952 ();
 sg13g2_fill_2 FILLER_21_1980 ();
 sg13g2_fill_1 FILLER_21_1982 ();
 sg13g2_decap_4 FILLER_21_2013 ();
 sg13g2_fill_1 FILLER_21_2017 ();
 sg13g2_decap_4 FILLER_21_2050 ();
 sg13g2_fill_2 FILLER_21_2054 ();
 sg13g2_fill_1 FILLER_21_2081 ();
 sg13g2_fill_1 FILLER_21_2087 ();
 sg13g2_decap_8 FILLER_21_2123 ();
 sg13g2_fill_1 FILLER_21_2143 ();
 sg13g2_fill_1 FILLER_21_2169 ();
 sg13g2_fill_2 FILLER_21_2178 ();
 sg13g2_fill_2 FILLER_21_2214 ();
 sg13g2_fill_1 FILLER_21_2216 ();
 sg13g2_fill_1 FILLER_21_2246 ();
 sg13g2_decap_4 FILLER_21_2266 ();
 sg13g2_decap_8 FILLER_21_2278 ();
 sg13g2_decap_4 FILLER_21_2285 ();
 sg13g2_fill_1 FILLER_21_2289 ();
 sg13g2_fill_2 FILLER_21_2318 ();
 sg13g2_decap_4 FILLER_21_2333 ();
 sg13g2_fill_2 FILLER_21_2337 ();
 sg13g2_decap_8 FILLER_21_2359 ();
 sg13g2_decap_8 FILLER_21_2406 ();
 sg13g2_decap_4 FILLER_21_2413 ();
 sg13g2_fill_1 FILLER_21_2417 ();
 sg13g2_decap_8 FILLER_21_2430 ();
 sg13g2_fill_1 FILLER_21_2437 ();
 sg13g2_decap_8 FILLER_21_2463 ();
 sg13g2_decap_4 FILLER_21_2470 ();
 sg13g2_fill_1 FILLER_21_2474 ();
 sg13g2_decap_8 FILLER_21_2484 ();
 sg13g2_decap_8 FILLER_21_2491 ();
 sg13g2_fill_1 FILLER_21_2498 ();
 sg13g2_fill_2 FILLER_21_2523 ();
 sg13g2_decap_4 FILLER_21_2538 ();
 sg13g2_fill_2 FILLER_21_2542 ();
 sg13g2_decap_8 FILLER_21_2568 ();
 sg13g2_fill_2 FILLER_21_2575 ();
 sg13g2_decap_8 FILLER_21_2593 ();
 sg13g2_fill_2 FILLER_21_2610 ();
 sg13g2_fill_2 FILLER_21_2616 ();
 sg13g2_fill_2 FILLER_21_2634 ();
 sg13g2_fill_2 FILLER_21_2645 ();
 sg13g2_decap_8 FILLER_21_2665 ();
 sg13g2_fill_1 FILLER_21_2672 ();
 sg13g2_fill_1 FILLER_21_2691 ();
 sg13g2_decap_4 FILLER_21_2695 ();
 sg13g2_decap_8 FILLER_21_2718 ();
 sg13g2_fill_1 FILLER_21_2733 ();
 sg13g2_fill_2 FILLER_21_2746 ();
 sg13g2_decap_4 FILLER_21_2761 ();
 sg13g2_fill_1 FILLER_21_2765 ();
 sg13g2_fill_1 FILLER_21_2776 ();
 sg13g2_decap_4 FILLER_21_2781 ();
 sg13g2_fill_2 FILLER_21_2785 ();
 sg13g2_decap_8 FILLER_21_2798 ();
 sg13g2_fill_1 FILLER_21_2805 ();
 sg13g2_decap_4 FILLER_21_2811 ();
 sg13g2_fill_1 FILLER_21_2815 ();
 sg13g2_decap_8 FILLER_21_2820 ();
 sg13g2_decap_8 FILLER_21_2827 ();
 sg13g2_decap_8 FILLER_21_2834 ();
 sg13g2_fill_2 FILLER_21_2841 ();
 sg13g2_fill_1 FILLER_21_2843 ();
 sg13g2_decap_8 FILLER_21_2857 ();
 sg13g2_decap_4 FILLER_21_2869 ();
 sg13g2_fill_1 FILLER_21_2873 ();
 sg13g2_decap_4 FILLER_21_2886 ();
 sg13g2_fill_2 FILLER_21_2890 ();
 sg13g2_decap_4 FILLER_21_2905 ();
 sg13g2_decap_8 FILLER_21_2914 ();
 sg13g2_fill_1 FILLER_21_2921 ();
 sg13g2_fill_1 FILLER_21_2927 ();
 sg13g2_decap_8 FILLER_21_2938 ();
 sg13g2_decap_8 FILLER_21_2945 ();
 sg13g2_fill_2 FILLER_21_2952 ();
 sg13g2_fill_1 FILLER_21_2954 ();
 sg13g2_fill_2 FILLER_21_2964 ();
 sg13g2_fill_1 FILLER_21_2966 ();
 sg13g2_fill_2 FILLER_21_2971 ();
 sg13g2_decap_8 FILLER_21_2987 ();
 sg13g2_decap_4 FILLER_21_2994 ();
 sg13g2_decap_8 FILLER_21_3011 ();
 sg13g2_fill_2 FILLER_21_3027 ();
 sg13g2_fill_1 FILLER_21_3029 ();
 sg13g2_decap_4 FILLER_21_3034 ();
 sg13g2_decap_4 FILLER_21_3056 ();
 sg13g2_fill_2 FILLER_21_3060 ();
 sg13g2_fill_2 FILLER_21_3067 ();
 sg13g2_decap_8 FILLER_21_3073 ();
 sg13g2_decap_8 FILLER_21_3080 ();
 sg13g2_decap_8 FILLER_21_3087 ();
 sg13g2_decap_8 FILLER_21_3094 ();
 sg13g2_decap_8 FILLER_21_3101 ();
 sg13g2_decap_4 FILLER_21_3108 ();
 sg13g2_fill_2 FILLER_21_3112 ();
 sg13g2_fill_2 FILLER_21_3131 ();
 sg13g2_fill_1 FILLER_21_3133 ();
 sg13g2_decap_4 FILLER_21_3138 ();
 sg13g2_fill_2 FILLER_21_3142 ();
 sg13g2_fill_1 FILLER_21_3157 ();
 sg13g2_decap_8 FILLER_21_3163 ();
 sg13g2_decap_4 FILLER_21_3188 ();
 sg13g2_fill_1 FILLER_21_3192 ();
 sg13g2_fill_2 FILLER_21_3201 ();
 sg13g2_fill_1 FILLER_21_3203 ();
 sg13g2_decap_8 FILLER_21_3213 ();
 sg13g2_decap_8 FILLER_21_3220 ();
 sg13g2_decap_4 FILLER_21_3227 ();
 sg13g2_decap_8 FILLER_21_3240 ();
 sg13g2_decap_8 FILLER_21_3247 ();
 sg13g2_fill_2 FILLER_21_3254 ();
 sg13g2_fill_2 FILLER_21_3269 ();
 sg13g2_fill_2 FILLER_21_3302 ();
 sg13g2_fill_1 FILLER_21_3304 ();
 sg13g2_decap_8 FILLER_21_3309 ();
 sg13g2_decap_4 FILLER_21_3316 ();
 sg13g2_decap_4 FILLER_21_3325 ();
 sg13g2_fill_1 FILLER_21_3329 ();
 sg13g2_fill_2 FILLER_21_3361 ();
 sg13g2_fill_2 FILLER_21_3372 ();
 sg13g2_fill_1 FILLER_21_3386 ();
 sg13g2_decap_4 FILLER_21_3391 ();
 sg13g2_fill_2 FILLER_21_3395 ();
 sg13g2_decap_8 FILLER_21_3419 ();
 sg13g2_fill_1 FILLER_21_3426 ();
 sg13g2_decap_4 FILLER_21_3432 ();
 sg13g2_fill_1 FILLER_21_3436 ();
 sg13g2_decap_8 FILLER_21_3441 ();
 sg13g2_decap_4 FILLER_21_3448 ();
 sg13g2_fill_2 FILLER_21_3452 ();
 sg13g2_decap_4 FILLER_21_3458 ();
 sg13g2_decap_8 FILLER_21_3466 ();
 sg13g2_decap_8 FILLER_21_3473 ();
 sg13g2_fill_2 FILLER_21_3480 ();
 sg13g2_fill_1 FILLER_21_3482 ();
 sg13g2_fill_1 FILLER_21_3488 ();
 sg13g2_decap_4 FILLER_21_3493 ();
 sg13g2_fill_1 FILLER_21_3497 ();
 sg13g2_decap_8 FILLER_21_3515 ();
 sg13g2_decap_8 FILLER_21_3522 ();
 sg13g2_decap_8 FILLER_21_3529 ();
 sg13g2_decap_8 FILLER_21_3536 ();
 sg13g2_decap_8 FILLER_21_3543 ();
 sg13g2_decap_8 FILLER_21_3550 ();
 sg13g2_decap_8 FILLER_21_3557 ();
 sg13g2_decap_8 FILLER_21_3564 ();
 sg13g2_decap_8 FILLER_21_3571 ();
 sg13g2_fill_2 FILLER_21_3578 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_46 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_decap_4 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_decap_8 FILLER_22_136 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_169 ();
 sg13g2_decap_8 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_183 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_decap_4 FILLER_22_202 ();
 sg13g2_fill_1 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_decap_8 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_fill_2 FILLER_22_253 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_decap_4 FILLER_22_274 ();
 sg13g2_fill_2 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_292 ();
 sg13g2_decap_4 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_decap_4 FILLER_22_327 ();
 sg13g2_decap_4 FILLER_22_357 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_decap_4 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_4 FILLER_22_402 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_decap_4 FILLER_22_429 ();
 sg13g2_fill_2 FILLER_22_438 ();
 sg13g2_decap_4 FILLER_22_501 ();
 sg13g2_fill_1 FILLER_22_505 ();
 sg13g2_fill_1 FILLER_22_558 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_4 FILLER_22_595 ();
 sg13g2_fill_1 FILLER_22_599 ();
 sg13g2_fill_2 FILLER_22_613 ();
 sg13g2_fill_1 FILLER_22_615 ();
 sg13g2_fill_2 FILLER_22_625 ();
 sg13g2_fill_1 FILLER_22_627 ();
 sg13g2_fill_2 FILLER_22_641 ();
 sg13g2_fill_1 FILLER_22_643 ();
 sg13g2_fill_2 FILLER_22_696 ();
 sg13g2_decap_8 FILLER_22_715 ();
 sg13g2_decap_4 FILLER_22_722 ();
 sg13g2_fill_2 FILLER_22_729 ();
 sg13g2_fill_1 FILLER_22_731 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_fill_1 FILLER_22_769 ();
 sg13g2_decap_8 FILLER_22_775 ();
 sg13g2_decap_4 FILLER_22_782 ();
 sg13g2_fill_1 FILLER_22_786 ();
 sg13g2_fill_1 FILLER_22_800 ();
 sg13g2_fill_2 FILLER_22_806 ();
 sg13g2_decap_4 FILLER_22_817 ();
 sg13g2_fill_1 FILLER_22_821 ();
 sg13g2_fill_2 FILLER_22_831 ();
 sg13g2_fill_1 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_839 ();
 sg13g2_fill_2 FILLER_22_846 ();
 sg13g2_fill_1 FILLER_22_848 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_893 ();
 sg13g2_fill_1 FILLER_22_900 ();
 sg13g2_fill_1 FILLER_22_919 ();
 sg13g2_decap_8 FILLER_22_923 ();
 sg13g2_decap_8 FILLER_22_930 ();
 sg13g2_decap_4 FILLER_22_950 ();
 sg13g2_fill_2 FILLER_22_954 ();
 sg13g2_fill_2 FILLER_22_964 ();
 sg13g2_fill_2 FILLER_22_978 ();
 sg13g2_decap_4 FILLER_22_987 ();
 sg13g2_fill_2 FILLER_22_991 ();
 sg13g2_fill_2 FILLER_22_1009 ();
 sg13g2_fill_1 FILLER_22_1011 ();
 sg13g2_decap_4 FILLER_22_1020 ();
 sg13g2_fill_2 FILLER_22_1024 ();
 sg13g2_fill_2 FILLER_22_1031 ();
 sg13g2_fill_1 FILLER_22_1037 ();
 sg13g2_decap_8 FILLER_22_1043 ();
 sg13g2_fill_1 FILLER_22_1050 ();
 sg13g2_decap_8 FILLER_22_1055 ();
 sg13g2_decap_4 FILLER_22_1062 ();
 sg13g2_fill_2 FILLER_22_1066 ();
 sg13g2_decap_8 FILLER_22_1086 ();
 sg13g2_decap_8 FILLER_22_1106 ();
 sg13g2_decap_8 FILLER_22_1117 ();
 sg13g2_decap_4 FILLER_22_1124 ();
 sg13g2_fill_1 FILLER_22_1128 ();
 sg13g2_decap_8 FILLER_22_1133 ();
 sg13g2_decap_4 FILLER_22_1140 ();
 sg13g2_fill_2 FILLER_22_1144 ();
 sg13g2_fill_2 FILLER_22_1156 ();
 sg13g2_fill_1 FILLER_22_1158 ();
 sg13g2_fill_2 FILLER_22_1164 ();
 sg13g2_decap_8 FILLER_22_1171 ();
 sg13g2_fill_2 FILLER_22_1178 ();
 sg13g2_decap_8 FILLER_22_1193 ();
 sg13g2_fill_1 FILLER_22_1200 ();
 sg13g2_decap_8 FILLER_22_1239 ();
 sg13g2_decap_8 FILLER_22_1246 ();
 sg13g2_decap_8 FILLER_22_1253 ();
 sg13g2_fill_2 FILLER_22_1260 ();
 sg13g2_fill_1 FILLER_22_1275 ();
 sg13g2_fill_2 FILLER_22_1313 ();
 sg13g2_decap_4 FILLER_22_1328 ();
 sg13g2_fill_2 FILLER_22_1332 ();
 sg13g2_decap_8 FILLER_22_1349 ();
 sg13g2_fill_2 FILLER_22_1356 ();
 sg13g2_fill_1 FILLER_22_1358 ();
 sg13g2_fill_1 FILLER_22_1363 ();
 sg13g2_decap_8 FILLER_22_1369 ();
 sg13g2_decap_8 FILLER_22_1376 ();
 sg13g2_fill_2 FILLER_22_1383 ();
 sg13g2_decap_4 FILLER_22_1397 ();
 sg13g2_decap_4 FILLER_22_1415 ();
 sg13g2_decap_8 FILLER_22_1423 ();
 sg13g2_fill_2 FILLER_22_1430 ();
 sg13g2_fill_1 FILLER_22_1432 ();
 sg13g2_fill_2 FILLER_22_1446 ();
 sg13g2_fill_2 FILLER_22_1453 ();
 sg13g2_decap_4 FILLER_22_1509 ();
 sg13g2_fill_2 FILLER_22_1513 ();
 sg13g2_fill_2 FILLER_22_1599 ();
 sg13g2_fill_2 FILLER_22_1611 ();
 sg13g2_fill_1 FILLER_22_1613 ();
 sg13g2_decap_8 FILLER_22_1618 ();
 sg13g2_decap_8 FILLER_22_1625 ();
 sg13g2_fill_2 FILLER_22_1632 ();
 sg13g2_fill_1 FILLER_22_1634 ();
 sg13g2_decap_8 FILLER_22_1658 ();
 sg13g2_decap_8 FILLER_22_1665 ();
 sg13g2_fill_2 FILLER_22_1672 ();
 sg13g2_fill_1 FILLER_22_1674 ();
 sg13g2_decap_4 FILLER_22_1680 ();
 sg13g2_decap_8 FILLER_22_1710 ();
 sg13g2_fill_1 FILLER_22_1717 ();
 sg13g2_decap_8 FILLER_22_1728 ();
 sg13g2_decap_8 FILLER_22_1750 ();
 sg13g2_decap_8 FILLER_22_1757 ();
 sg13g2_decap_8 FILLER_22_1764 ();
 sg13g2_fill_2 FILLER_22_1771 ();
 sg13g2_decap_8 FILLER_22_1788 ();
 sg13g2_fill_1 FILLER_22_1795 ();
 sg13g2_fill_2 FILLER_22_1800 ();
 sg13g2_decap_8 FILLER_22_1807 ();
 sg13g2_decap_4 FILLER_22_1814 ();
 sg13g2_fill_2 FILLER_22_1832 ();
 sg13g2_fill_1 FILLER_22_1834 ();
 sg13g2_fill_1 FILLER_22_1860 ();
 sg13g2_decap_4 FILLER_22_1874 ();
 sg13g2_fill_1 FILLER_22_1913 ();
 sg13g2_decap_8 FILLER_22_1976 ();
 sg13g2_decap_4 FILLER_22_1983 ();
 sg13g2_fill_2 FILLER_22_1992 ();
 sg13g2_decap_8 FILLER_22_2020 ();
 sg13g2_decap_4 FILLER_22_2031 ();
 sg13g2_fill_1 FILLER_22_2049 ();
 sg13g2_decap_4 FILLER_22_2055 ();
 sg13g2_fill_2 FILLER_22_2064 ();
 sg13g2_decap_4 FILLER_22_2081 ();
 sg13g2_fill_1 FILLER_22_2101 ();
 sg13g2_fill_2 FILLER_22_2116 ();
 sg13g2_fill_1 FILLER_22_2118 ();
 sg13g2_decap_8 FILLER_22_2132 ();
 sg13g2_fill_2 FILLER_22_2152 ();
 sg13g2_fill_2 FILLER_22_2164 ();
 sg13g2_fill_1 FILLER_22_2166 ();
 sg13g2_decap_8 FILLER_22_2174 ();
 sg13g2_decap_8 FILLER_22_2181 ();
 sg13g2_fill_1 FILLER_22_2188 ();
 sg13g2_fill_2 FILLER_22_2194 ();
 sg13g2_decap_8 FILLER_22_2205 ();
 sg13g2_decap_8 FILLER_22_2212 ();
 sg13g2_fill_1 FILLER_22_2239 ();
 sg13g2_decap_4 FILLER_22_2289 ();
 sg13g2_fill_2 FILLER_22_2293 ();
 sg13g2_decap_8 FILLER_22_2299 ();
 sg13g2_decap_8 FILLER_22_2306 ();
 sg13g2_decap_4 FILLER_22_2313 ();
 sg13g2_fill_1 FILLER_22_2317 ();
 sg13g2_fill_2 FILLER_22_2335 ();
 sg13g2_fill_1 FILLER_22_2337 ();
 sg13g2_fill_2 FILLER_22_2343 ();
 sg13g2_fill_2 FILLER_22_2352 ();
 sg13g2_decap_4 FILLER_22_2367 ();
 sg13g2_fill_1 FILLER_22_2371 ();
 sg13g2_fill_1 FILLER_22_2402 ();
 sg13g2_fill_2 FILLER_22_2416 ();
 sg13g2_fill_1 FILLER_22_2418 ();
 sg13g2_fill_2 FILLER_22_2441 ();
 sg13g2_fill_2 FILLER_22_2465 ();
 sg13g2_decap_8 FILLER_22_2487 ();
 sg13g2_decap_8 FILLER_22_2494 ();
 sg13g2_decap_8 FILLER_22_2501 ();
 sg13g2_decap_4 FILLER_22_2518 ();
 sg13g2_decap_8 FILLER_22_2533 ();
 sg13g2_decap_4 FILLER_22_2540 ();
 sg13g2_fill_2 FILLER_22_2544 ();
 sg13g2_fill_1 FILLER_22_2552 ();
 sg13g2_fill_1 FILLER_22_2558 ();
 sg13g2_decap_8 FILLER_22_2563 ();
 sg13g2_decap_8 FILLER_22_2570 ();
 sg13g2_fill_2 FILLER_22_2601 ();
 sg13g2_fill_2 FILLER_22_2613 ();
 sg13g2_fill_1 FILLER_22_2615 ();
 sg13g2_fill_2 FILLER_22_2622 ();
 sg13g2_fill_1 FILLER_22_2624 ();
 sg13g2_fill_2 FILLER_22_2644 ();
 sg13g2_decap_4 FILLER_22_2656 ();
 sg13g2_fill_1 FILLER_22_2660 ();
 sg13g2_fill_2 FILLER_22_2691 ();
 sg13g2_fill_1 FILLER_22_2693 ();
 sg13g2_fill_1 FILLER_22_2707 ();
 sg13g2_fill_2 FILLER_22_2750 ();
 sg13g2_decap_8 FILLER_22_2757 ();
 sg13g2_decap_8 FILLER_22_2764 ();
 sg13g2_fill_2 FILLER_22_2775 ();
 sg13g2_fill_1 FILLER_22_2777 ();
 sg13g2_decap_4 FILLER_22_2839 ();
 sg13g2_fill_2 FILLER_22_2856 ();
 sg13g2_decap_8 FILLER_22_2866 ();
 sg13g2_fill_1 FILLER_22_2883 ();
 sg13g2_decap_8 FILLER_22_2889 ();
 sg13g2_fill_1 FILLER_22_2896 ();
 sg13g2_fill_2 FILLER_22_2918 ();
 sg13g2_decap_4 FILLER_22_2929 ();
 sg13g2_decap_4 FILLER_22_2945 ();
 sg13g2_decap_8 FILLER_22_2989 ();
 sg13g2_decap_8 FILLER_22_2996 ();
 sg13g2_fill_1 FILLER_22_3003 ();
 sg13g2_fill_2 FILLER_22_3012 ();
 sg13g2_fill_1 FILLER_22_3014 ();
 sg13g2_decap_8 FILLER_22_3041 ();
 sg13g2_decap_8 FILLER_22_3048 ();
 sg13g2_fill_2 FILLER_22_3109 ();
 sg13g2_decap_4 FILLER_22_3132 ();
 sg13g2_fill_1 FILLER_22_3136 ();
 sg13g2_decap_4 FILLER_22_3158 ();
 sg13g2_fill_2 FILLER_22_3166 ();
 sg13g2_fill_1 FILLER_22_3168 ();
 sg13g2_decap_4 FILLER_22_3182 ();
 sg13g2_fill_2 FILLER_22_3186 ();
 sg13g2_decap_8 FILLER_22_3214 ();
 sg13g2_decap_8 FILLER_22_3241 ();
 sg13g2_decap_8 FILLER_22_3248 ();
 sg13g2_decap_4 FILLER_22_3255 ();
 sg13g2_decap_4 FILLER_22_3275 ();
 sg13g2_fill_2 FILLER_22_3279 ();
 sg13g2_fill_2 FILLER_22_3285 ();
 sg13g2_decap_8 FILLER_22_3292 ();
 sg13g2_fill_1 FILLER_22_3299 ();
 sg13g2_decap_8 FILLER_22_3334 ();
 sg13g2_decap_8 FILLER_22_3341 ();
 sg13g2_fill_2 FILLER_22_3357 ();
 sg13g2_fill_1 FILLER_22_3359 ();
 sg13g2_fill_2 FILLER_22_3373 ();
 sg13g2_fill_1 FILLER_22_3375 ();
 sg13g2_decap_4 FILLER_22_3424 ();
 sg13g2_decap_8 FILLER_22_3476 ();
 sg13g2_fill_1 FILLER_22_3483 ();
 sg13g2_decap_8 FILLER_22_3509 ();
 sg13g2_decap_8 FILLER_22_3516 ();
 sg13g2_decap_8 FILLER_22_3523 ();
 sg13g2_decap_8 FILLER_22_3530 ();
 sg13g2_decap_8 FILLER_22_3537 ();
 sg13g2_decap_8 FILLER_22_3544 ();
 sg13g2_decap_8 FILLER_22_3551 ();
 sg13g2_decap_8 FILLER_22_3558 ();
 sg13g2_decap_8 FILLER_22_3565 ();
 sg13g2_decap_8 FILLER_22_3572 ();
 sg13g2_fill_1 FILLER_22_3579 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_111 ();
 sg13g2_decap_4 FILLER_23_139 ();
 sg13g2_fill_2 FILLER_23_143 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_159 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_decap_4 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_253 ();
 sg13g2_decap_4 FILLER_23_264 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_389 ();
 sg13g2_decap_4 FILLER_23_402 ();
 sg13g2_fill_1 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_23_449 ();
 sg13g2_fill_1 FILLER_23_456 ();
 sg13g2_fill_1 FILLER_23_480 ();
 sg13g2_fill_2 FILLER_23_489 ();
 sg13g2_fill_2 FILLER_23_495 ();
 sg13g2_fill_2 FILLER_23_521 ();
 sg13g2_fill_2 FILLER_23_536 ();
 sg13g2_fill_1 FILLER_23_538 ();
 sg13g2_fill_2 FILLER_23_588 ();
 sg13g2_fill_1 FILLER_23_590 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_fill_2 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_fill_2 FILLER_23_623 ();
 sg13g2_fill_2 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_fill_2 FILLER_23_686 ();
 sg13g2_decap_4 FILLER_23_699 ();
 sg13g2_decap_8 FILLER_23_741 ();
 sg13g2_decap_4 FILLER_23_748 ();
 sg13g2_fill_2 FILLER_23_752 ();
 sg13g2_decap_8 FILLER_23_782 ();
 sg13g2_decap_4 FILLER_23_789 ();
 sg13g2_fill_2 FILLER_23_798 ();
 sg13g2_fill_1 FILLER_23_800 ();
 sg13g2_decap_4 FILLER_23_819 ();
 sg13g2_fill_2 FILLER_23_823 ();
 sg13g2_fill_1 FILLER_23_836 ();
 sg13g2_decap_8 FILLER_23_842 ();
 sg13g2_decap_8 FILLER_23_849 ();
 sg13g2_decap_8 FILLER_23_856 ();
 sg13g2_fill_2 FILLER_23_891 ();
 sg13g2_fill_1 FILLER_23_893 ();
 sg13g2_decap_4 FILLER_23_921 ();
 sg13g2_fill_1 FILLER_23_925 ();
 sg13g2_decap_8 FILLER_23_954 ();
 sg13g2_fill_2 FILLER_23_989 ();
 sg13g2_fill_1 FILLER_23_991 ();
 sg13g2_fill_2 FILLER_23_1002 ();
 sg13g2_decap_8 FILLER_23_1009 ();
 sg13g2_fill_2 FILLER_23_1016 ();
 sg13g2_fill_1 FILLER_23_1027 ();
 sg13g2_fill_2 FILLER_23_1038 ();
 sg13g2_decap_8 FILLER_23_1053 ();
 sg13g2_fill_1 FILLER_23_1060 ();
 sg13g2_fill_2 FILLER_23_1065 ();
 sg13g2_decap_4 FILLER_23_1080 ();
 sg13g2_decap_8 FILLER_23_1117 ();
 sg13g2_decap_4 FILLER_23_1124 ();
 sg13g2_fill_2 FILLER_23_1128 ();
 sg13g2_decap_8 FILLER_23_1152 ();
 sg13g2_decap_4 FILLER_23_1159 ();
 sg13g2_decap_4 FILLER_23_1176 ();
 sg13g2_decap_8 FILLER_23_1197 ();
 sg13g2_decap_4 FILLER_23_1204 ();
 sg13g2_fill_1 FILLER_23_1208 ();
 sg13g2_decap_4 FILLER_23_1234 ();
 sg13g2_fill_2 FILLER_23_1289 ();
 sg13g2_fill_1 FILLER_23_1291 ();
 sg13g2_fill_2 FILLER_23_1310 ();
 sg13g2_fill_2 FILLER_23_1316 ();
 sg13g2_fill_1 FILLER_23_1318 ();
 sg13g2_fill_1 FILLER_23_1332 ();
 sg13g2_fill_2 FILLER_23_1412 ();
 sg13g2_fill_2 FILLER_23_1442 ();
 sg13g2_decap_4 FILLER_23_1452 ();
 sg13g2_fill_1 FILLER_23_1460 ();
 sg13g2_decap_8 FILLER_23_1487 ();
 sg13g2_decap_8 FILLER_23_1494 ();
 sg13g2_fill_2 FILLER_23_1501 ();
 sg13g2_fill_1 FILLER_23_1503 ();
 sg13g2_decap_8 FILLER_23_1517 ();
 sg13g2_fill_2 FILLER_23_1538 ();
 sg13g2_fill_1 FILLER_23_1540 ();
 sg13g2_decap_4 FILLER_23_1546 ();
 sg13g2_decap_8 FILLER_23_1564 ();
 sg13g2_fill_1 FILLER_23_1571 ();
 sg13g2_fill_2 FILLER_23_1585 ();
 sg13g2_fill_1 FILLER_23_1587 ();
 sg13g2_fill_1 FILLER_23_1601 ();
 sg13g2_fill_2 FILLER_23_1630 ();
 sg13g2_fill_2 FILLER_23_1640 ();
 sg13g2_decap_4 FILLER_23_1656 ();
 sg13g2_fill_2 FILLER_23_1660 ();
 sg13g2_fill_2 FILLER_23_1674 ();
 sg13g2_fill_1 FILLER_23_1676 ();
 sg13g2_decap_8 FILLER_23_1683 ();
 sg13g2_decap_8 FILLER_23_1716 ();
 sg13g2_decap_4 FILLER_23_1723 ();
 sg13g2_fill_2 FILLER_23_1727 ();
 sg13g2_decap_8 FILLER_23_1736 ();
 sg13g2_decap_4 FILLER_23_1743 ();
 sg13g2_fill_2 FILLER_23_1752 ();
 sg13g2_fill_2 FILLER_23_1772 ();
 sg13g2_fill_2 FILLER_23_1781 ();
 sg13g2_fill_1 FILLER_23_1783 ();
 sg13g2_decap_8 FILLER_23_1790 ();
 sg13g2_decap_4 FILLER_23_1797 ();
 sg13g2_decap_4 FILLER_23_1819 ();
 sg13g2_fill_2 FILLER_23_1823 ();
 sg13g2_decap_4 FILLER_23_1851 ();
 sg13g2_fill_2 FILLER_23_1855 ();
 sg13g2_fill_2 FILLER_23_1861 ();
 sg13g2_fill_1 FILLER_23_1863 ();
 sg13g2_decap_4 FILLER_23_1913 ();
 sg13g2_fill_1 FILLER_23_1917 ();
 sg13g2_fill_2 FILLER_23_1944 ();
 sg13g2_decap_8 FILLER_23_1962 ();
 sg13g2_decap_4 FILLER_23_1969 ();
 sg13g2_fill_2 FILLER_23_1973 ();
 sg13g2_decap_8 FILLER_23_2012 ();
 sg13g2_decap_8 FILLER_23_2019 ();
 sg13g2_fill_1 FILLER_23_2026 ();
 sg13g2_decap_4 FILLER_23_2069 ();
 sg13g2_fill_2 FILLER_23_2073 ();
 sg13g2_decap_8 FILLER_23_2097 ();
 sg13g2_fill_2 FILLER_23_2104 ();
 sg13g2_fill_1 FILLER_23_2106 ();
 sg13g2_fill_1 FILLER_23_2119 ();
 sg13g2_decap_8 FILLER_23_2128 ();
 sg13g2_fill_2 FILLER_23_2135 ();
 sg13g2_fill_1 FILLER_23_2165 ();
 sg13g2_decap_4 FILLER_23_2182 ();
 sg13g2_fill_2 FILLER_23_2186 ();
 sg13g2_decap_4 FILLER_23_2209 ();
 sg13g2_decap_8 FILLER_23_2239 ();
 sg13g2_fill_2 FILLER_23_2246 ();
 sg13g2_fill_2 FILLER_23_2258 ();
 sg13g2_decap_8 FILLER_23_2265 ();
 sg13g2_fill_2 FILLER_23_2272 ();
 sg13g2_fill_1 FILLER_23_2274 ();
 sg13g2_decap_8 FILLER_23_2285 ();
 sg13g2_fill_2 FILLER_23_2292 ();
 sg13g2_fill_1 FILLER_23_2294 ();
 sg13g2_fill_2 FILLER_23_2313 ();
 sg13g2_decap_8 FILLER_23_2321 ();
 sg13g2_decap_8 FILLER_23_2335 ();
 sg13g2_fill_2 FILLER_23_2342 ();
 sg13g2_decap_4 FILLER_23_2347 ();
 sg13g2_decap_4 FILLER_23_2369 ();
 sg13g2_fill_1 FILLER_23_2388 ();
 sg13g2_fill_2 FILLER_23_2398 ();
 sg13g2_fill_1 FILLER_23_2400 ();
 sg13g2_fill_1 FILLER_23_2406 ();
 sg13g2_decap_8 FILLER_23_2417 ();
 sg13g2_fill_2 FILLER_23_2451 ();
 sg13g2_fill_1 FILLER_23_2453 ();
 sg13g2_fill_1 FILLER_23_2461 ();
 sg13g2_decap_4 FILLER_23_2465 ();
 sg13g2_fill_1 FILLER_23_2469 ();
 sg13g2_decap_4 FILLER_23_2474 ();
 sg13g2_fill_2 FILLER_23_2478 ();
 sg13g2_fill_2 FILLER_23_2520 ();
 sg13g2_fill_1 FILLER_23_2522 ();
 sg13g2_decap_4 FILLER_23_2574 ();
 sg13g2_fill_2 FILLER_23_2578 ();
 sg13g2_fill_2 FILLER_23_2589 ();
 sg13g2_decap_4 FILLER_23_2596 ();
 sg13g2_fill_2 FILLER_23_2600 ();
 sg13g2_fill_1 FILLER_23_2620 ();
 sg13g2_fill_2 FILLER_23_2628 ();
 sg13g2_decap_4 FILLER_23_2638 ();
 sg13g2_decap_8 FILLER_23_2660 ();
 sg13g2_fill_2 FILLER_23_2667 ();
 sg13g2_decap_8 FILLER_23_2690 ();
 sg13g2_fill_2 FILLER_23_2697 ();
 sg13g2_fill_1 FILLER_23_2699 ();
 sg13g2_fill_1 FILLER_23_2715 ();
 sg13g2_decap_4 FILLER_23_2732 ();
 sg13g2_fill_2 FILLER_23_2748 ();
 sg13g2_fill_2 FILLER_23_2764 ();
 sg13g2_decap_4 FILLER_23_2774 ();
 sg13g2_decap_8 FILLER_23_2786 ();
 sg13g2_fill_1 FILLER_23_2793 ();
 sg13g2_decap_8 FILLER_23_2798 ();
 sg13g2_fill_2 FILLER_23_2805 ();
 sg13g2_fill_1 FILLER_23_2810 ();
 sg13g2_decap_8 FILLER_23_2819 ();
 sg13g2_fill_2 FILLER_23_2826 ();
 sg13g2_fill_1 FILLER_23_2828 ();
 sg13g2_decap_8 FILLER_23_2842 ();
 sg13g2_fill_2 FILLER_23_2849 ();
 sg13g2_fill_1 FILLER_23_2851 ();
 sg13g2_fill_2 FILLER_23_2872 ();
 sg13g2_fill_1 FILLER_23_2874 ();
 sg13g2_decap_8 FILLER_23_2883 ();
 sg13g2_fill_2 FILLER_23_2890 ();
 sg13g2_fill_1 FILLER_23_2892 ();
 sg13g2_fill_2 FILLER_23_2906 ();
 sg13g2_fill_2 FILLER_23_2926 ();
 sg13g2_fill_1 FILLER_23_2928 ();
 sg13g2_fill_1 FILLER_23_2945 ();
 sg13g2_fill_1 FILLER_23_2959 ();
 sg13g2_fill_2 FILLER_23_2964 ();
 sg13g2_decap_4 FILLER_23_2998 ();
 sg13g2_fill_1 FILLER_23_3002 ();
 sg13g2_fill_2 FILLER_23_3015 ();
 sg13g2_fill_1 FILLER_23_3017 ();
 sg13g2_fill_1 FILLER_23_3035 ();
 sg13g2_decap_8 FILLER_23_3047 ();
 sg13g2_decap_8 FILLER_23_3054 ();
 sg13g2_decap_8 FILLER_23_3079 ();
 sg13g2_fill_1 FILLER_23_3086 ();
 sg13g2_fill_2 FILLER_23_3107 ();
 sg13g2_decap_8 FILLER_23_3132 ();
 sg13g2_fill_2 FILLER_23_3139 ();
 sg13g2_fill_2 FILLER_23_3154 ();
 sg13g2_decap_8 FILLER_23_3179 ();
 sg13g2_decap_4 FILLER_23_3186 ();
 sg13g2_fill_1 FILLER_23_3190 ();
 sg13g2_decap_4 FILLER_23_3209 ();
 sg13g2_fill_1 FILLER_23_3253 ();
 sg13g2_fill_2 FILLER_23_3272 ();
 sg13g2_decap_8 FILLER_23_3299 ();
 sg13g2_fill_2 FILLER_23_3306 ();
 sg13g2_decap_8 FILLER_23_3363 ();
 sg13g2_decap_8 FILLER_23_3370 ();
 sg13g2_decap_8 FILLER_23_3377 ();
 sg13g2_fill_2 FILLER_23_3384 ();
 sg13g2_decap_4 FILLER_23_3396 ();
 sg13g2_fill_2 FILLER_23_3400 ();
 sg13g2_decap_4 FILLER_23_3426 ();
 sg13g2_fill_1 FILLER_23_3430 ();
 sg13g2_fill_1 FILLER_23_3443 ();
 sg13g2_decap_8 FILLER_23_3454 ();
 sg13g2_decap_4 FILLER_23_3461 ();
 sg13g2_decap_8 FILLER_23_3478 ();
 sg13g2_fill_2 FILLER_23_3485 ();
 sg13g2_fill_1 FILLER_23_3487 ();
 sg13g2_decap_8 FILLER_23_3503 ();
 sg13g2_decap_8 FILLER_23_3510 ();
 sg13g2_decap_8 FILLER_23_3517 ();
 sg13g2_decap_8 FILLER_23_3524 ();
 sg13g2_decap_8 FILLER_23_3531 ();
 sg13g2_decap_8 FILLER_23_3538 ();
 sg13g2_decap_8 FILLER_23_3545 ();
 sg13g2_decap_8 FILLER_23_3552 ();
 sg13g2_decap_8 FILLER_23_3559 ();
 sg13g2_decap_8 FILLER_23_3566 ();
 sg13g2_decap_8 FILLER_23_3573 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_51 ();
 sg13g2_decap_4 FILLER_24_58 ();
 sg13g2_fill_2 FILLER_24_62 ();
 sg13g2_decap_4 FILLER_24_81 ();
 sg13g2_decap_4 FILLER_24_90 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_decap_4 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_120 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_fill_2 FILLER_24_150 ();
 sg13g2_decap_4 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_decap_4 FILLER_24_203 ();
 sg13g2_decap_4 FILLER_24_218 ();
 sg13g2_decap_4 FILLER_24_226 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_decap_4 FILLER_24_379 ();
 sg13g2_fill_1 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_1 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_24_421 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_fill_1 FILLER_24_430 ();
 sg13g2_fill_2 FILLER_24_444 ();
 sg13g2_decap_8 FILLER_24_451 ();
 sg13g2_decap_8 FILLER_24_458 ();
 sg13g2_fill_1 FILLER_24_465 ();
 sg13g2_decap_8 FILLER_24_480 ();
 sg13g2_decap_4 FILLER_24_487 ();
 sg13g2_fill_2 FILLER_24_491 ();
 sg13g2_decap_8 FILLER_24_507 ();
 sg13g2_decap_8 FILLER_24_514 ();
 sg13g2_decap_8 FILLER_24_521 ();
 sg13g2_decap_4 FILLER_24_528 ();
 sg13g2_decap_4 FILLER_24_538 ();
 sg13g2_fill_2 FILLER_24_542 ();
 sg13g2_decap_4 FILLER_24_548 ();
 sg13g2_fill_2 FILLER_24_557 ();
 sg13g2_decap_8 FILLER_24_562 ();
 sg13g2_decap_8 FILLER_24_569 ();
 sg13g2_decap_8 FILLER_24_576 ();
 sg13g2_fill_2 FILLER_24_583 ();
 sg13g2_fill_2 FILLER_24_620 ();
 sg13g2_fill_1 FILLER_24_644 ();
 sg13g2_decap_4 FILLER_24_677 ();
 sg13g2_decap_8 FILLER_24_713 ();
 sg13g2_decap_8 FILLER_24_720 ();
 sg13g2_decap_4 FILLER_24_727 ();
 sg13g2_decap_8 FILLER_24_748 ();
 sg13g2_fill_1 FILLER_24_755 ();
 sg13g2_fill_2 FILLER_24_763 ();
 sg13g2_fill_1 FILLER_24_765 ();
 sg13g2_decap_8 FILLER_24_781 ();
 sg13g2_fill_1 FILLER_24_788 ();
 sg13g2_decap_4 FILLER_24_801 ();
 sg13g2_fill_2 FILLER_24_805 ();
 sg13g2_decap_4 FILLER_24_825 ();
 sg13g2_fill_1 FILLER_24_829 ();
 sg13g2_decap_4 FILLER_24_850 ();
 sg13g2_decap_8 FILLER_24_867 ();
 sg13g2_fill_2 FILLER_24_874 ();
 sg13g2_fill_1 FILLER_24_876 ();
 sg13g2_decap_8 FILLER_24_886 ();
 sg13g2_decap_8 FILLER_24_893 ();
 sg13g2_fill_2 FILLER_24_900 ();
 sg13g2_fill_1 FILLER_24_902 ();
 sg13g2_decap_8 FILLER_24_923 ();
 sg13g2_fill_2 FILLER_24_930 ();
 sg13g2_decap_8 FILLER_24_936 ();
 sg13g2_decap_8 FILLER_24_943 ();
 sg13g2_fill_2 FILLER_24_950 ();
 sg13g2_fill_1 FILLER_24_952 ();
 sg13g2_fill_2 FILLER_24_968 ();
 sg13g2_decap_4 FILLER_24_975 ();
 sg13g2_fill_2 FILLER_24_986 ();
 sg13g2_fill_1 FILLER_24_988 ();
 sg13g2_decap_4 FILLER_24_993 ();
 sg13g2_fill_1 FILLER_24_997 ();
 sg13g2_fill_1 FILLER_24_1002 ();
 sg13g2_decap_8 FILLER_24_1008 ();
 sg13g2_fill_2 FILLER_24_1033 ();
 sg13g2_decap_4 FILLER_24_1039 ();
 sg13g2_fill_1 FILLER_24_1043 ();
 sg13g2_decap_4 FILLER_24_1078 ();
 sg13g2_fill_2 FILLER_24_1086 ();
 sg13g2_decap_8 FILLER_24_1098 ();
 sg13g2_fill_2 FILLER_24_1105 ();
 sg13g2_fill_2 FILLER_24_1124 ();
 sg13g2_fill_1 FILLER_24_1126 ();
 sg13g2_fill_1 FILLER_24_1144 ();
 sg13g2_fill_1 FILLER_24_1152 ();
 sg13g2_decap_4 FILLER_24_1159 ();
 sg13g2_decap_8 FILLER_24_1202 ();
 sg13g2_decap_4 FILLER_24_1209 ();
 sg13g2_fill_1 FILLER_24_1213 ();
 sg13g2_decap_8 FILLER_24_1240 ();
 sg13g2_decap_4 FILLER_24_1263 ();
 sg13g2_fill_2 FILLER_24_1276 ();
 sg13g2_fill_2 FILLER_24_1303 ();
 sg13g2_fill_1 FILLER_24_1305 ();
 sg13g2_decap_8 FILLER_24_1332 ();
 sg13g2_fill_1 FILLER_24_1339 ();
 sg13g2_decap_8 FILLER_24_1352 ();
 sg13g2_decap_4 FILLER_24_1359 ();
 sg13g2_fill_1 FILLER_24_1363 ();
 sg13g2_fill_2 FILLER_24_1386 ();
 sg13g2_fill_1 FILLER_24_1388 ();
 sg13g2_decap_4 FILLER_24_1393 ();
 sg13g2_fill_1 FILLER_24_1397 ();
 sg13g2_decap_8 FILLER_24_1403 ();
 sg13g2_decap_8 FILLER_24_1410 ();
 sg13g2_fill_1 FILLER_24_1417 ();
 sg13g2_decap_8 FILLER_24_1431 ();
 sg13g2_fill_1 FILLER_24_1438 ();
 sg13g2_decap_4 FILLER_24_1443 ();
 sg13g2_decap_8 FILLER_24_1452 ();
 sg13g2_fill_2 FILLER_24_1459 ();
 sg13g2_fill_1 FILLER_24_1461 ();
 sg13g2_fill_2 FILLER_24_1471 ();
 sg13g2_fill_1 FILLER_24_1473 ();
 sg13g2_fill_2 FILLER_24_1530 ();
 sg13g2_decap_8 FILLER_24_1550 ();
 sg13g2_fill_2 FILLER_24_1557 ();
 sg13g2_fill_2 FILLER_24_1569 ();
 sg13g2_decap_8 FILLER_24_1584 ();
 sg13g2_fill_1 FILLER_24_1591 ();
 sg13g2_fill_2 FILLER_24_1605 ();
 sg13g2_decap_4 FILLER_24_1611 ();
 sg13g2_fill_2 FILLER_24_1615 ();
 sg13g2_fill_2 FILLER_24_1634 ();
 sg13g2_fill_2 FILLER_24_1655 ();
 sg13g2_fill_1 FILLER_24_1657 ();
 sg13g2_decap_8 FILLER_24_1678 ();
 sg13g2_decap_4 FILLER_24_1685 ();
 sg13g2_fill_1 FILLER_24_1689 ();
 sg13g2_fill_2 FILLER_24_1722 ();
 sg13g2_fill_1 FILLER_24_1745 ();
 sg13g2_decap_8 FILLER_24_1758 ();
 sg13g2_decap_4 FILLER_24_1765 ();
 sg13g2_decap_8 FILLER_24_1797 ();
 sg13g2_fill_2 FILLER_24_1804 ();
 sg13g2_decap_4 FILLER_24_1824 ();
 sg13g2_fill_2 FILLER_24_1828 ();
 sg13g2_fill_1 FILLER_24_1849 ();
 sg13g2_decap_8 FILLER_24_1858 ();
 sg13g2_decap_4 FILLER_24_1865 ();
 sg13g2_fill_2 FILLER_24_1869 ();
 sg13g2_decap_4 FILLER_24_1878 ();
 sg13g2_fill_2 FILLER_24_1882 ();
 sg13g2_fill_2 FILLER_24_1893 ();
 sg13g2_fill_1 FILLER_24_1895 ();
 sg13g2_decap_8 FILLER_24_1924 ();
 sg13g2_decap_4 FILLER_24_1949 ();
 sg13g2_fill_1 FILLER_24_1953 ();
 sg13g2_fill_2 FILLER_24_1957 ();
 sg13g2_fill_2 FILLER_24_1968 ();
 sg13g2_fill_1 FILLER_24_1970 ();
 sg13g2_fill_2 FILLER_24_2016 ();
 sg13g2_fill_1 FILLER_24_2028 ();
 sg13g2_fill_2 FILLER_24_2050 ();
 sg13g2_decap_4 FILLER_24_2060 ();
 sg13g2_fill_2 FILLER_24_2064 ();
 sg13g2_fill_2 FILLER_24_2075 ();
 sg13g2_fill_1 FILLER_24_2077 ();
 sg13g2_fill_1 FILLER_24_2084 ();
 sg13g2_decap_4 FILLER_24_2091 ();
 sg13g2_fill_2 FILLER_24_2095 ();
 sg13g2_decap_4 FILLER_24_2102 ();
 sg13g2_decap_8 FILLER_24_2125 ();
 sg13g2_decap_4 FILLER_24_2132 ();
 sg13g2_fill_2 FILLER_24_2136 ();
 sg13g2_decap_8 FILLER_24_2148 ();
 sg13g2_fill_2 FILLER_24_2155 ();
 sg13g2_fill_1 FILLER_24_2157 ();
 sg13g2_decap_8 FILLER_24_2179 ();
 sg13g2_decap_4 FILLER_24_2186 ();
 sg13g2_decap_8 FILLER_24_2203 ();
 sg13g2_decap_8 FILLER_24_2210 ();
 sg13g2_fill_2 FILLER_24_2217 ();
 sg13g2_decap_8 FILLER_24_2236 ();
 sg13g2_decap_8 FILLER_24_2250 ();
 sg13g2_decap_4 FILLER_24_2257 ();
 sg13g2_fill_2 FILLER_24_2261 ();
 sg13g2_decap_4 FILLER_24_2266 ();
 sg13g2_fill_2 FILLER_24_2270 ();
 sg13g2_fill_2 FILLER_24_2278 ();
 sg13g2_decap_4 FILLER_24_2285 ();
 sg13g2_decap_4 FILLER_24_2306 ();
 sg13g2_fill_2 FILLER_24_2310 ();
 sg13g2_fill_1 FILLER_24_2328 ();
 sg13g2_decap_8 FILLER_24_2333 ();
 sg13g2_decap_8 FILLER_24_2340 ();
 sg13g2_decap_8 FILLER_24_2347 ();
 sg13g2_fill_2 FILLER_24_2354 ();
 sg13g2_fill_2 FILLER_24_2369 ();
 sg13g2_fill_2 FILLER_24_2387 ();
 sg13g2_fill_1 FILLER_24_2389 ();
 sg13g2_decap_4 FILLER_24_2399 ();
 sg13g2_fill_2 FILLER_24_2403 ();
 sg13g2_decap_8 FILLER_24_2423 ();
 sg13g2_decap_4 FILLER_24_2430 ();
 sg13g2_fill_1 FILLER_24_2434 ();
 sg13g2_decap_4 FILLER_24_2448 ();
 sg13g2_decap_8 FILLER_24_2460 ();
 sg13g2_decap_8 FILLER_24_2467 ();
 sg13g2_decap_4 FILLER_24_2474 ();
 sg13g2_fill_2 FILLER_24_2489 ();
 sg13g2_fill_1 FILLER_24_2491 ();
 sg13g2_decap_8 FILLER_24_2496 ();
 sg13g2_fill_2 FILLER_24_2503 ();
 sg13g2_decap_4 FILLER_24_2514 ();
 sg13g2_fill_1 FILLER_24_2518 ();
 sg13g2_decap_8 FILLER_24_2530 ();
 sg13g2_decap_4 FILLER_24_2537 ();
 sg13g2_fill_1 FILLER_24_2541 ();
 sg13g2_decap_8 FILLER_24_2559 ();
 sg13g2_decap_8 FILLER_24_2566 ();
 sg13g2_fill_2 FILLER_24_2573 ();
 sg13g2_fill_2 FILLER_24_2592 ();
 sg13g2_decap_8 FILLER_24_2631 ();
 sg13g2_fill_2 FILLER_24_2638 ();
 sg13g2_fill_1 FILLER_24_2640 ();
 sg13g2_decap_4 FILLER_24_2655 ();
 sg13g2_fill_2 FILLER_24_2687 ();
 sg13g2_fill_1 FILLER_24_2689 ();
 sg13g2_decap_8 FILLER_24_2698 ();
 sg13g2_fill_1 FILLER_24_2705 ();
 sg13g2_fill_1 FILLER_24_2716 ();
 sg13g2_decap_4 FILLER_24_2726 ();
 sg13g2_fill_1 FILLER_24_2730 ();
 sg13g2_decap_8 FILLER_24_2735 ();
 sg13g2_decap_8 FILLER_24_2742 ();
 sg13g2_decap_8 FILLER_24_2749 ();
 sg13g2_decap_4 FILLER_24_2756 ();
 sg13g2_fill_1 FILLER_24_2760 ();
 sg13g2_fill_1 FILLER_24_2798 ();
 sg13g2_fill_1 FILLER_24_2811 ();
 sg13g2_fill_2 FILLER_24_2827 ();
 sg13g2_fill_2 FILLER_24_2851 ();
 sg13g2_fill_2 FILLER_24_2869 ();
 sg13g2_fill_1 FILLER_24_2871 ();
 sg13g2_fill_2 FILLER_24_2889 ();
 sg13g2_fill_1 FILLER_24_2914 ();
 sg13g2_decap_4 FILLER_24_2920 ();
 sg13g2_fill_2 FILLER_24_2948 ();
 sg13g2_fill_1 FILLER_24_2950 ();
 sg13g2_decap_8 FILLER_24_2993 ();
 sg13g2_decap_8 FILLER_24_3000 ();
 sg13g2_fill_1 FILLER_24_3015 ();
 sg13g2_fill_2 FILLER_24_3022 ();
 sg13g2_fill_1 FILLER_24_3024 ();
 sg13g2_fill_2 FILLER_24_3042 ();
 sg13g2_fill_1 FILLER_24_3044 ();
 sg13g2_fill_2 FILLER_24_3056 ();
 sg13g2_fill_2 FILLER_24_3063 ();
 sg13g2_fill_2 FILLER_24_3085 ();
 sg13g2_fill_1 FILLER_24_3087 ();
 sg13g2_decap_4 FILLER_24_3105 ();
 sg13g2_fill_2 FILLER_24_3109 ();
 sg13g2_fill_2 FILLER_24_3128 ();
 sg13g2_fill_2 FILLER_24_3164 ();
 sg13g2_fill_1 FILLER_24_3166 ();
 sg13g2_decap_4 FILLER_24_3187 ();
 sg13g2_decap_8 FILLER_24_3211 ();
 sg13g2_decap_4 FILLER_24_3218 ();
 sg13g2_decap_4 FILLER_24_3256 ();
 sg13g2_fill_1 FILLER_24_3260 ();
 sg13g2_fill_2 FILLER_24_3265 ();
 sg13g2_decap_8 FILLER_24_3272 ();
 sg13g2_fill_2 FILLER_24_3279 ();
 sg13g2_fill_1 FILLER_24_3281 ();
 sg13g2_decap_8 FILLER_24_3290 ();
 sg13g2_fill_1 FILLER_24_3297 ();
 sg13g2_fill_1 FILLER_24_3305 ();
 sg13g2_decap_8 FILLER_24_3310 ();
 sg13g2_decap_8 FILLER_24_3317 ();
 sg13g2_decap_4 FILLER_24_3331 ();
 sg13g2_fill_1 FILLER_24_3335 ();
 sg13g2_fill_2 FILLER_24_3358 ();
 sg13g2_fill_1 FILLER_24_3360 ();
 sg13g2_decap_4 FILLER_24_3374 ();
 sg13g2_fill_2 FILLER_24_3378 ();
 sg13g2_decap_8 FILLER_24_3399 ();
 sg13g2_decap_4 FILLER_24_3406 ();
 sg13g2_fill_2 FILLER_24_3410 ();
 sg13g2_fill_1 FILLER_24_3417 ();
 sg13g2_decap_8 FILLER_24_3428 ();
 sg13g2_fill_1 FILLER_24_3435 ();
 sg13g2_fill_1 FILLER_24_3455 ();
 sg13g2_fill_1 FILLER_24_3469 ();
 sg13g2_decap_8 FILLER_24_3486 ();
 sg13g2_fill_1 FILLER_24_3498 ();
 sg13g2_fill_1 FILLER_24_3502 ();
 sg13g2_decap_8 FILLER_24_3507 ();
 sg13g2_decap_8 FILLER_24_3514 ();
 sg13g2_decap_8 FILLER_24_3521 ();
 sg13g2_decap_8 FILLER_24_3528 ();
 sg13g2_decap_8 FILLER_24_3535 ();
 sg13g2_decap_8 FILLER_24_3542 ();
 sg13g2_decap_8 FILLER_24_3549 ();
 sg13g2_decap_8 FILLER_24_3556 ();
 sg13g2_decap_8 FILLER_24_3563 ();
 sg13g2_decap_8 FILLER_24_3570 ();
 sg13g2_fill_2 FILLER_24_3577 ();
 sg13g2_fill_1 FILLER_24_3579 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_decap_8 FILLER_25_104 ();
 sg13g2_decap_4 FILLER_25_111 ();
 sg13g2_decap_8 FILLER_25_120 ();
 sg13g2_decap_4 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_135 ();
 sg13g2_decap_4 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_153 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_177 ();
 sg13g2_decap_8 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_decap_4 FILLER_25_209 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_271 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_354 ();
 sg13g2_decap_4 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_decap_4 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_403 ();
 sg13g2_decap_4 FILLER_25_415 ();
 sg13g2_fill_2 FILLER_25_419 ();
 sg13g2_decap_8 FILLER_25_426 ();
 sg13g2_fill_1 FILLER_25_433 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_fill_1 FILLER_25_462 ();
 sg13g2_fill_2 FILLER_25_483 ();
 sg13g2_fill_1 FILLER_25_485 ();
 sg13g2_decap_4 FILLER_25_504 ();
 sg13g2_decap_4 FILLER_25_525 ();
 sg13g2_fill_1 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_fill_2 FILLER_25_560 ();
 sg13g2_fill_1 FILLER_25_562 ();
 sg13g2_decap_4 FILLER_25_584 ();
 sg13g2_fill_1 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_600 ();
 sg13g2_decap_8 FILLER_25_607 ();
 sg13g2_decap_8 FILLER_25_614 ();
 sg13g2_decap_4 FILLER_25_621 ();
 sg13g2_decap_4 FILLER_25_633 ();
 sg13g2_fill_1 FILLER_25_642 ();
 sg13g2_decap_8 FILLER_25_673 ();
 sg13g2_fill_2 FILLER_25_680 ();
 sg13g2_fill_1 FILLER_25_682 ();
 sg13g2_fill_2 FILLER_25_691 ();
 sg13g2_decap_4 FILLER_25_719 ();
 sg13g2_fill_2 FILLER_25_723 ();
 sg13g2_decap_4 FILLER_25_756 ();
 sg13g2_fill_1 FILLER_25_760 ();
 sg13g2_fill_2 FILLER_25_767 ();
 sg13g2_fill_1 FILLER_25_769 ();
 sg13g2_fill_2 FILLER_25_777 ();
 sg13g2_decap_4 FILLER_25_784 ();
 sg13g2_fill_1 FILLER_25_788 ();
 sg13g2_decap_4 FILLER_25_797 ();
 sg13g2_decap_8 FILLER_25_818 ();
 sg13g2_fill_2 FILLER_25_825 ();
 sg13g2_decap_4 FILLER_25_848 ();
 sg13g2_fill_2 FILLER_25_884 ();
 sg13g2_fill_1 FILLER_25_886 ();
 sg13g2_fill_2 FILLER_25_891 ();
 sg13g2_decap_4 FILLER_25_904 ();
 sg13g2_decap_4 FILLER_25_966 ();
 sg13g2_fill_2 FILLER_25_970 ();
 sg13g2_fill_2 FILLER_25_999 ();
 sg13g2_fill_1 FILLER_25_1001 ();
 sg13g2_fill_1 FILLER_25_1015 ();
 sg13g2_fill_2 FILLER_25_1037 ();
 sg13g2_fill_1 FILLER_25_1039 ();
 sg13g2_fill_1 FILLER_25_1058 ();
 sg13g2_fill_2 FILLER_25_1063 ();
 sg13g2_decap_8 FILLER_25_1091 ();
 sg13g2_decap_4 FILLER_25_1125 ();
 sg13g2_fill_2 FILLER_25_1142 ();
 sg13g2_fill_1 FILLER_25_1144 ();
 sg13g2_fill_2 FILLER_25_1153 ();
 sg13g2_fill_1 FILLER_25_1162 ();
 sg13g2_decap_8 FILLER_25_1176 ();
 sg13g2_fill_1 FILLER_25_1183 ();
 sg13g2_fill_2 FILLER_25_1206 ();
 sg13g2_fill_1 FILLER_25_1226 ();
 sg13g2_fill_2 FILLER_25_1239 ();
 sg13g2_fill_1 FILLER_25_1241 ();
 sg13g2_fill_2 FILLER_25_1298 ();
 sg13g2_decap_4 FILLER_25_1305 ();
 sg13g2_fill_1 FILLER_25_1309 ();
 sg13g2_decap_4 FILLER_25_1314 ();
 sg13g2_decap_8 FILLER_25_1322 ();
 sg13g2_fill_2 FILLER_25_1329 ();
 sg13g2_fill_1 FILLER_25_1331 ();
 sg13g2_fill_2 FILLER_25_1356 ();
 sg13g2_decap_8 FILLER_25_1377 ();
 sg13g2_decap_4 FILLER_25_1384 ();
 sg13g2_fill_2 FILLER_25_1388 ();
 sg13g2_decap_4 FILLER_25_1402 ();
 sg13g2_decap_4 FILLER_25_1411 ();
 sg13g2_fill_1 FILLER_25_1441 ();
 sg13g2_decap_8 FILLER_25_1470 ();
 sg13g2_fill_2 FILLER_25_1477 ();
 sg13g2_fill_2 FILLER_25_1483 ();
 sg13g2_fill_1 FILLER_25_1485 ();
 sg13g2_decap_4 FILLER_25_1503 ();
 sg13g2_fill_1 FILLER_25_1507 ();
 sg13g2_fill_1 FILLER_25_1525 ();
 sg13g2_decap_8 FILLER_25_1538 ();
 sg13g2_decap_4 FILLER_25_1545 ();
 sg13g2_fill_2 FILLER_25_1574 ();
 sg13g2_fill_2 FILLER_25_1583 ();
 sg13g2_fill_2 FILLER_25_1590 ();
 sg13g2_decap_4 FILLER_25_1609 ();
 sg13g2_fill_1 FILLER_25_1613 ();
 sg13g2_decap_8 FILLER_25_1619 ();
 sg13g2_fill_2 FILLER_25_1631 ();
 sg13g2_fill_1 FILLER_25_1633 ();
 sg13g2_fill_2 FILLER_25_1640 ();
 sg13g2_fill_2 FILLER_25_1648 ();
 sg13g2_fill_1 FILLER_25_1650 ();
 sg13g2_fill_2 FILLER_25_1662 ();
 sg13g2_fill_1 FILLER_25_1664 ();
 sg13g2_decap_8 FILLER_25_1681 ();
 sg13g2_decap_8 FILLER_25_1688 ();
 sg13g2_decap_4 FILLER_25_1695 ();
 sg13g2_decap_8 FILLER_25_1703 ();
 sg13g2_fill_2 FILLER_25_1710 ();
 sg13g2_fill_1 FILLER_25_1712 ();
 sg13g2_fill_2 FILLER_25_1726 ();
 sg13g2_fill_1 FILLER_25_1728 ();
 sg13g2_decap_8 FILLER_25_1734 ();
 sg13g2_fill_1 FILLER_25_1762 ();
 sg13g2_fill_2 FILLER_25_1778 ();
 sg13g2_decap_8 FILLER_25_1785 ();
 sg13g2_decap_4 FILLER_25_1792 ();
 sg13g2_fill_1 FILLER_25_1796 ();
 sg13g2_fill_1 FILLER_25_1818 ();
 sg13g2_decap_8 FILLER_25_1823 ();
 sg13g2_decap_4 FILLER_25_1835 ();
 sg13g2_fill_1 FILLER_25_1839 ();
 sg13g2_fill_1 FILLER_25_1844 ();
 sg13g2_decap_4 FILLER_25_1855 ();
 sg13g2_decap_8 FILLER_25_1888 ();
 sg13g2_decap_4 FILLER_25_1895 ();
 sg13g2_fill_1 FILLER_25_1899 ();
 sg13g2_decap_8 FILLER_25_1909 ();
 sg13g2_decap_4 FILLER_25_1916 ();
 sg13g2_fill_2 FILLER_25_1933 ();
 sg13g2_fill_1 FILLER_25_1935 ();
 sg13g2_fill_2 FILLER_25_1976 ();
 sg13g2_fill_2 FILLER_25_2000 ();
 sg13g2_fill_2 FILLER_25_2019 ();
 sg13g2_fill_1 FILLER_25_2034 ();
 sg13g2_decap_8 FILLER_25_2039 ();
 sg13g2_decap_4 FILLER_25_2046 ();
 sg13g2_decap_8 FILLER_25_2065 ();
 sg13g2_decap_4 FILLER_25_2072 ();
 sg13g2_fill_1 FILLER_25_2076 ();
 sg13g2_decap_4 FILLER_25_2126 ();
 sg13g2_fill_1 FILLER_25_2130 ();
 sg13g2_decap_4 FILLER_25_2138 ();
 sg13g2_fill_1 FILLER_25_2142 ();
 sg13g2_decap_4 FILLER_25_2180 ();
 sg13g2_decap_4 FILLER_25_2302 ();
 sg13g2_fill_2 FILLER_25_2306 ();
 sg13g2_decap_4 FILLER_25_2351 ();
 sg13g2_fill_1 FILLER_25_2355 ();
 sg13g2_fill_1 FILLER_25_2369 ();
 sg13g2_decap_4 FILLER_25_2396 ();
 sg13g2_fill_2 FILLER_25_2400 ();
 sg13g2_fill_2 FILLER_25_2429 ();
 sg13g2_fill_1 FILLER_25_2431 ();
 sg13g2_fill_1 FILLER_25_2445 ();
 sg13g2_decap_4 FILLER_25_2481 ();
 sg13g2_fill_2 FILLER_25_2517 ();
 sg13g2_fill_1 FILLER_25_2519 ();
 sg13g2_fill_1 FILLER_25_2553 ();
 sg13g2_decap_8 FILLER_25_2561 ();
 sg13g2_decap_8 FILLER_25_2568 ();
 sg13g2_fill_2 FILLER_25_2575 ();
 sg13g2_fill_1 FILLER_25_2577 ();
 sg13g2_decap_8 FILLER_25_2588 ();
 sg13g2_fill_2 FILLER_25_2595 ();
 sg13g2_fill_2 FILLER_25_2605 ();
 sg13g2_decap_4 FILLER_25_2615 ();
 sg13g2_decap_8 FILLER_25_2631 ();
 sg13g2_fill_2 FILLER_25_2638 ();
 sg13g2_fill_1 FILLER_25_2640 ();
 sg13g2_decap_4 FILLER_25_2661 ();
 sg13g2_decap_8 FILLER_25_2681 ();
 sg13g2_decap_8 FILLER_25_2688 ();
 sg13g2_fill_2 FILLER_25_2695 ();
 sg13g2_decap_8 FILLER_25_2704 ();
 sg13g2_decap_8 FILLER_25_2711 ();
 sg13g2_decap_4 FILLER_25_2718 ();
 sg13g2_fill_2 FILLER_25_2722 ();
 sg13g2_fill_2 FILLER_25_2737 ();
 sg13g2_fill_1 FILLER_25_2739 ();
 sg13g2_decap_8 FILLER_25_2744 ();
 sg13g2_fill_2 FILLER_25_2751 ();
 sg13g2_fill_2 FILLER_25_2757 ();
 sg13g2_fill_1 FILLER_25_2759 ();
 sg13g2_fill_2 FILLER_25_2786 ();
 sg13g2_fill_1 FILLER_25_2788 ();
 sg13g2_fill_2 FILLER_25_2807 ();
 sg13g2_fill_1 FILLER_25_2809 ();
 sg13g2_decap_4 FILLER_25_2818 ();
 sg13g2_fill_1 FILLER_25_2822 ();
 sg13g2_decap_4 FILLER_25_2830 ();
 sg13g2_fill_1 FILLER_25_2834 ();
 sg13g2_decap_4 FILLER_25_2843 ();
 sg13g2_decap_4 FILLER_25_2875 ();
 sg13g2_fill_1 FILLER_25_2879 ();
 sg13g2_fill_1 FILLER_25_2884 ();
 sg13g2_decap_8 FILLER_25_2913 ();
 sg13g2_decap_8 FILLER_25_2920 ();
 sg13g2_fill_1 FILLER_25_2927 ();
 sg13g2_decap_4 FILLER_25_2944 ();
 sg13g2_decap_4 FILLER_25_2965 ();
 sg13g2_decap_8 FILLER_25_3004 ();
 sg13g2_fill_2 FILLER_25_3011 ();
 sg13g2_fill_1 FILLER_25_3049 ();
 sg13g2_fill_1 FILLER_25_3074 ();
 sg13g2_decap_8 FILLER_25_3104 ();
 sg13g2_decap_8 FILLER_25_3111 ();
 sg13g2_fill_1 FILLER_25_3118 ();
 sg13g2_decap_8 FILLER_25_3123 ();
 sg13g2_decap_8 FILLER_25_3159 ();
 sg13g2_fill_2 FILLER_25_3166 ();
 sg13g2_decap_8 FILLER_25_3183 ();
 sg13g2_decap_8 FILLER_25_3190 ();
 sg13g2_fill_2 FILLER_25_3197 ();
 sg13g2_decap_8 FILLER_25_3207 ();
 sg13g2_decap_8 FILLER_25_3214 ();
 sg13g2_fill_2 FILLER_25_3221 ();
 sg13g2_fill_1 FILLER_25_3223 ();
 sg13g2_fill_2 FILLER_25_3233 ();
 sg13g2_fill_1 FILLER_25_3235 ();
 sg13g2_decap_8 FILLER_25_3251 ();
 sg13g2_decap_4 FILLER_25_3258 ();
 sg13g2_fill_2 FILLER_25_3262 ();
 sg13g2_fill_2 FILLER_25_3270 ();
 sg13g2_fill_1 FILLER_25_3300 ();
 sg13g2_fill_1 FILLER_25_3329 ();
 sg13g2_decap_4 FILLER_25_3335 ();
 sg13g2_fill_1 FILLER_25_3339 ();
 sg13g2_decap_8 FILLER_25_3400 ();
 sg13g2_decap_4 FILLER_25_3407 ();
 sg13g2_fill_1 FILLER_25_3411 ();
 sg13g2_decap_8 FILLER_25_3432 ();
 sg13g2_decap_8 FILLER_25_3439 ();
 sg13g2_fill_1 FILLER_25_3450 ();
 sg13g2_decap_4 FILLER_25_3456 ();
 sg13g2_fill_2 FILLER_25_3460 ();
 sg13g2_fill_2 FILLER_25_3480 ();
 sg13g2_fill_2 FILLER_25_3489 ();
 sg13g2_fill_1 FILLER_25_3497 ();
 sg13g2_decap_8 FILLER_25_3526 ();
 sg13g2_decap_8 FILLER_25_3533 ();
 sg13g2_decap_8 FILLER_25_3540 ();
 sg13g2_decap_8 FILLER_25_3547 ();
 sg13g2_decap_8 FILLER_25_3554 ();
 sg13g2_decap_8 FILLER_25_3561 ();
 sg13g2_decap_8 FILLER_25_3568 ();
 sg13g2_decap_4 FILLER_25_3575 ();
 sg13g2_fill_1 FILLER_25_3579 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_49 ();
 sg13g2_decap_4 FILLER_26_87 ();
 sg13g2_decap_8 FILLER_26_96 ();
 sg13g2_decap_8 FILLER_26_103 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_135 ();
 sg13g2_fill_2 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_decap_8 FILLER_26_233 ();
 sg13g2_decap_4 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_4 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_2 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_344 ();
 sg13g2_fill_2 FILLER_26_374 ();
 sg13g2_fill_1 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_402 ();
 sg13g2_fill_2 FILLER_26_431 ();
 sg13g2_decap_4 FILLER_26_436 ();
 sg13g2_fill_1 FILLER_26_440 ();
 sg13g2_fill_2 FILLER_26_454 ();
 sg13g2_fill_1 FILLER_26_456 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_fill_2 FILLER_26_476 ();
 sg13g2_fill_1 FILLER_26_550 ();
 sg13g2_fill_2 FILLER_26_556 ();
 sg13g2_fill_2 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_617 ();
 sg13g2_decap_4 FILLER_26_624 ();
 sg13g2_fill_2 FILLER_26_628 ();
 sg13g2_decap_4 FILLER_26_643 ();
 sg13g2_decap_4 FILLER_26_673 ();
 sg13g2_decap_8 FILLER_26_689 ();
 sg13g2_decap_8 FILLER_26_696 ();
 sg13g2_decap_4 FILLER_26_703 ();
 sg13g2_fill_2 FILLER_26_707 ();
 sg13g2_decap_4 FILLER_26_722 ();
 sg13g2_fill_1 FILLER_26_726 ();
 sg13g2_fill_2 FILLER_26_730 ();
 sg13g2_fill_1 FILLER_26_732 ();
 sg13g2_decap_8 FILLER_26_750 ();
 sg13g2_fill_2 FILLER_26_757 ();
 sg13g2_fill_2 FILLER_26_782 ();
 sg13g2_fill_1 FILLER_26_792 ();
 sg13g2_decap_8 FILLER_26_797 ();
 sg13g2_decap_8 FILLER_26_804 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_4 FILLER_26_852 ();
 sg13g2_decap_4 FILLER_26_868 ();
 sg13g2_fill_1 FILLER_26_872 ();
 sg13g2_decap_8 FILLER_26_904 ();
 sg13g2_fill_2 FILLER_26_928 ();
 sg13g2_fill_1 FILLER_26_930 ();
 sg13g2_decap_8 FILLER_26_936 ();
 sg13g2_decap_4 FILLER_26_943 ();
 sg13g2_fill_2 FILLER_26_947 ();
 sg13g2_fill_2 FILLER_26_963 ();
 sg13g2_fill_2 FILLER_26_973 ();
 sg13g2_decap_8 FILLER_26_983 ();
 sg13g2_decap_8 FILLER_26_990 ();
 sg13g2_fill_2 FILLER_26_1002 ();
 sg13g2_fill_1 FILLER_26_1004 ();
 sg13g2_fill_2 FILLER_26_1009 ();
 sg13g2_fill_1 FILLER_26_1011 ();
 sg13g2_fill_2 FILLER_26_1025 ();
 sg13g2_decap_8 FILLER_26_1041 ();
 sg13g2_fill_1 FILLER_26_1048 ();
 sg13g2_decap_4 FILLER_26_1052 ();
 sg13g2_fill_1 FILLER_26_1056 ();
 sg13g2_decap_4 FILLER_26_1067 ();
 sg13g2_fill_1 FILLER_26_1071 ();
 sg13g2_decap_8 FILLER_26_1084 ();
 sg13g2_decap_8 FILLER_26_1091 ();
 sg13g2_decap_4 FILLER_26_1130 ();
 sg13g2_fill_2 FILLER_26_1134 ();
 sg13g2_decap_8 FILLER_26_1144 ();
 sg13g2_fill_2 FILLER_26_1151 ();
 sg13g2_fill_1 FILLER_26_1153 ();
 sg13g2_fill_1 FILLER_26_1159 ();
 sg13g2_decap_4 FILLER_26_1164 ();
 sg13g2_fill_2 FILLER_26_1181 ();
 sg13g2_fill_1 FILLER_26_1183 ();
 sg13g2_decap_8 FILLER_26_1209 ();
 sg13g2_fill_2 FILLER_26_1216 ();
 sg13g2_decap_8 FILLER_26_1231 ();
 sg13g2_fill_1 FILLER_26_1238 ();
 sg13g2_fill_1 FILLER_26_1252 ();
 sg13g2_decap_8 FILLER_26_1263 ();
 sg13g2_decap_8 FILLER_26_1270 ();
 sg13g2_decap_4 FILLER_26_1277 ();
 sg13g2_decap_8 FILLER_26_1297 ();
 sg13g2_decap_4 FILLER_26_1304 ();
 sg13g2_fill_1 FILLER_26_1308 ();
 sg13g2_fill_2 FILLER_26_1319 ();
 sg13g2_fill_1 FILLER_26_1321 ();
 sg13g2_fill_2 FILLER_26_1349 ();
 sg13g2_fill_1 FILLER_26_1351 ();
 sg13g2_decap_4 FILLER_26_1357 ();
 sg13g2_fill_2 FILLER_26_1361 ();
 sg13g2_fill_2 FILLER_26_1368 ();
 sg13g2_decap_8 FILLER_26_1374 ();
 sg13g2_fill_2 FILLER_26_1381 ();
 sg13g2_fill_2 FILLER_26_1395 ();
 sg13g2_fill_1 FILLER_26_1397 ();
 sg13g2_fill_1 FILLER_26_1409 ();
 sg13g2_decap_8 FILLER_26_1414 ();
 sg13g2_fill_1 FILLER_26_1421 ();
 sg13g2_fill_2 FILLER_26_1427 ();
 sg13g2_fill_1 FILLER_26_1429 ();
 sg13g2_decap_8 FILLER_26_1445 ();
 sg13g2_decap_8 FILLER_26_1456 ();
 sg13g2_decap_8 FILLER_26_1463 ();
 sg13g2_fill_1 FILLER_26_1470 ();
 sg13g2_fill_2 FILLER_26_1475 ();
 sg13g2_fill_1 FILLER_26_1477 ();
 sg13g2_fill_2 FILLER_26_1519 ();
 sg13g2_fill_1 FILLER_26_1521 ();
 sg13g2_fill_2 FILLER_26_1554 ();
 sg13g2_fill_1 FILLER_26_1556 ();
 sg13g2_fill_2 FILLER_26_1562 ();
 sg13g2_fill_2 FILLER_26_1576 ();
 sg13g2_decap_8 FILLER_26_1583 ();
 sg13g2_decap_4 FILLER_26_1590 ();
 sg13g2_fill_2 FILLER_26_1594 ();
 sg13g2_decap_8 FILLER_26_1609 ();
 sg13g2_fill_1 FILLER_26_1616 ();
 sg13g2_decap_4 FILLER_26_1622 ();
 sg13g2_fill_1 FILLER_26_1626 ();
 sg13g2_fill_2 FILLER_26_1635 ();
 sg13g2_decap_8 FILLER_26_1650 ();
 sg13g2_fill_2 FILLER_26_1665 ();
 sg13g2_fill_1 FILLER_26_1679 ();
 sg13g2_decap_4 FILLER_26_1695 ();
 sg13g2_fill_2 FILLER_26_1699 ();
 sg13g2_decap_8 FILLER_26_1732 ();
 sg13g2_fill_2 FILLER_26_1766 ();
 sg13g2_fill_1 FILLER_26_1777 ();
 sg13g2_fill_1 FILLER_26_1801 ();
 sg13g2_fill_2 FILLER_26_1820 ();
 sg13g2_fill_1 FILLER_26_1822 ();
 sg13g2_decap_8 FILLER_26_1852 ();
 sg13g2_decap_8 FILLER_26_1859 ();
 sg13g2_decap_8 FILLER_26_1866 ();
 sg13g2_fill_2 FILLER_26_1886 ();
 sg13g2_fill_1 FILLER_26_1888 ();
 sg13g2_decap_4 FILLER_26_1910 ();
 sg13g2_fill_1 FILLER_26_1914 ();
 sg13g2_decap_4 FILLER_26_1957 ();
 sg13g2_fill_2 FILLER_26_1961 ();
 sg13g2_fill_2 FILLER_26_1998 ();
 sg13g2_fill_1 FILLER_26_2000 ();
 sg13g2_decap_8 FILLER_26_2013 ();
 sg13g2_decap_8 FILLER_26_2020 ();
 sg13g2_decap_4 FILLER_26_2043 ();
 sg13g2_fill_1 FILLER_26_2047 ();
 sg13g2_fill_2 FILLER_26_2075 ();
 sg13g2_decap_4 FILLER_26_2099 ();
 sg13g2_fill_2 FILLER_26_2103 ();
 sg13g2_decap_8 FILLER_26_2115 ();
 sg13g2_fill_2 FILLER_26_2122 ();
 sg13g2_fill_1 FILLER_26_2124 ();
 sg13g2_decap_4 FILLER_26_2153 ();
 sg13g2_fill_2 FILLER_26_2161 ();
 sg13g2_fill_2 FILLER_26_2167 ();
 sg13g2_fill_1 FILLER_26_2169 ();
 sg13g2_fill_2 FILLER_26_2179 ();
 sg13g2_fill_2 FILLER_26_2185 ();
 sg13g2_decap_4 FILLER_26_2200 ();
 sg13g2_fill_1 FILLER_26_2213 ();
 sg13g2_fill_2 FILLER_26_2218 ();
 sg13g2_fill_1 FILLER_26_2220 ();
 sg13g2_decap_8 FILLER_26_2225 ();
 sg13g2_decap_8 FILLER_26_2232 ();
 sg13g2_decap_4 FILLER_26_2239 ();
 sg13g2_fill_1 FILLER_26_2243 ();
 sg13g2_decap_8 FILLER_26_2252 ();
 sg13g2_decap_8 FILLER_26_2259 ();
 sg13g2_decap_8 FILLER_26_2266 ();
 sg13g2_fill_1 FILLER_26_2273 ();
 sg13g2_decap_8 FILLER_26_2308 ();
 sg13g2_fill_1 FILLER_26_2315 ();
 sg13g2_fill_1 FILLER_26_2328 ();
 sg13g2_decap_8 FILLER_26_2357 ();
 sg13g2_decap_8 FILLER_26_2364 ();
 sg13g2_decap_8 FILLER_26_2403 ();
 sg13g2_fill_2 FILLER_26_2410 ();
 sg13g2_fill_1 FILLER_26_2412 ();
 sg13g2_fill_1 FILLER_26_2430 ();
 sg13g2_decap_8 FILLER_26_2445 ();
 sg13g2_decap_4 FILLER_26_2452 ();
 sg13g2_fill_1 FILLER_26_2456 ();
 sg13g2_decap_4 FILLER_26_2466 ();
 sg13g2_decap_4 FILLER_26_2483 ();
 sg13g2_fill_1 FILLER_26_2504 ();
 sg13g2_fill_2 FILLER_26_2518 ();
 sg13g2_fill_1 FILLER_26_2520 ();
 sg13g2_decap_8 FILLER_26_2530 ();
 sg13g2_decap_8 FILLER_26_2537 ();
 sg13g2_fill_2 FILLER_26_2544 ();
 sg13g2_fill_1 FILLER_26_2546 ();
 sg13g2_fill_1 FILLER_26_2579 ();
 sg13g2_decap_4 FILLER_26_2585 ();
 sg13g2_decap_8 FILLER_26_2616 ();
 sg13g2_fill_2 FILLER_26_2623 ();
 sg13g2_fill_1 FILLER_26_2625 ();
 sg13g2_decap_4 FILLER_26_2654 ();
 sg13g2_fill_2 FILLER_26_2658 ();
 sg13g2_fill_2 FILLER_26_2689 ();
 sg13g2_fill_1 FILLER_26_2691 ();
 sg13g2_decap_8 FILLER_26_2720 ();
 sg13g2_decap_8 FILLER_26_2727 ();
 sg13g2_fill_1 FILLER_26_2734 ();
 sg13g2_fill_1 FILLER_26_2763 ();
 sg13g2_decap_8 FILLER_26_2781 ();
 sg13g2_fill_2 FILLER_26_2796 ();
 sg13g2_fill_1 FILLER_26_2798 ();
 sg13g2_decap_8 FILLER_26_2811 ();
 sg13g2_fill_2 FILLER_26_2818 ();
 sg13g2_fill_1 FILLER_26_2820 ();
 sg13g2_decap_4 FILLER_26_2849 ();
 sg13g2_decap_4 FILLER_26_2867 ();
 sg13g2_decap_8 FILLER_26_2884 ();
 sg13g2_decap_8 FILLER_26_2891 ();
 sg13g2_decap_4 FILLER_26_2898 ();
 sg13g2_decap_8 FILLER_26_2906 ();
 sg13g2_fill_1 FILLER_26_2913 ();
 sg13g2_decap_8 FILLER_26_2927 ();
 sg13g2_decap_8 FILLER_26_2934 ();
 sg13g2_decap_8 FILLER_26_2941 ();
 sg13g2_fill_1 FILLER_26_2948 ();
 sg13g2_fill_2 FILLER_26_2975 ();
 sg13g2_fill_2 FILLER_26_2989 ();
 sg13g2_fill_1 FILLER_26_2991 ();
 sg13g2_decap_8 FILLER_26_3004 ();
 sg13g2_decap_4 FILLER_26_3011 ();
 sg13g2_fill_2 FILLER_26_3015 ();
 sg13g2_decap_8 FILLER_26_3024 ();
 sg13g2_decap_8 FILLER_26_3031 ();
 sg13g2_decap_8 FILLER_26_3038 ();
 sg13g2_decap_8 FILLER_26_3045 ();
 sg13g2_fill_2 FILLER_26_3052 ();
 sg13g2_fill_1 FILLER_26_3054 ();
 sg13g2_decap_8 FILLER_26_3065 ();
 sg13g2_fill_2 FILLER_26_3072 ();
 sg13g2_fill_1 FILLER_26_3074 ();
 sg13g2_fill_2 FILLER_26_3088 ();
 sg13g2_fill_2 FILLER_26_3099 ();
 sg13g2_decap_8 FILLER_26_3108 ();
 sg13g2_decap_8 FILLER_26_3120 ();
 sg13g2_decap_8 FILLER_26_3134 ();
 sg13g2_decap_4 FILLER_26_3141 ();
 sg13g2_fill_2 FILLER_26_3145 ();
 sg13g2_decap_8 FILLER_26_3154 ();
 sg13g2_decap_8 FILLER_26_3161 ();
 sg13g2_decap_4 FILLER_26_3168 ();
 sg13g2_decap_8 FILLER_26_3210 ();
 sg13g2_decap_4 FILLER_26_3217 ();
 sg13g2_fill_2 FILLER_26_3256 ();
 sg13g2_decap_4 FILLER_26_3297 ();
 sg13g2_fill_1 FILLER_26_3301 ();
 sg13g2_fill_2 FILLER_26_3315 ();
 sg13g2_fill_1 FILLER_26_3317 ();
 sg13g2_decap_4 FILLER_26_3324 ();
 sg13g2_fill_1 FILLER_26_3328 ();
 sg13g2_fill_2 FILLER_26_3341 ();
 sg13g2_fill_2 FILLER_26_3374 ();
 sg13g2_fill_1 FILLER_26_3376 ();
 sg13g2_decap_8 FILLER_26_3386 ();
 sg13g2_decap_4 FILLER_26_3393 ();
 sg13g2_fill_1 FILLER_26_3397 ();
 sg13g2_decap_8 FILLER_26_3432 ();
 sg13g2_fill_1 FILLER_26_3439 ();
 sg13g2_fill_2 FILLER_26_3465 ();
 sg13g2_fill_1 FILLER_26_3467 ();
 sg13g2_decap_8 FILLER_26_3509 ();
 sg13g2_decap_8 FILLER_26_3516 ();
 sg13g2_decap_8 FILLER_26_3523 ();
 sg13g2_decap_8 FILLER_26_3530 ();
 sg13g2_decap_8 FILLER_26_3537 ();
 sg13g2_decap_8 FILLER_26_3544 ();
 sg13g2_decap_8 FILLER_26_3551 ();
 sg13g2_decap_8 FILLER_26_3558 ();
 sg13g2_decap_8 FILLER_26_3565 ();
 sg13g2_decap_8 FILLER_26_3572 ();
 sg13g2_fill_1 FILLER_26_3579 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_53 ();
 sg13g2_decap_4 FILLER_27_59 ();
 sg13g2_fill_2 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_143 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_decap_4 FILLER_27_199 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_215 ();
 sg13g2_fill_2 FILLER_27_245 ();
 sg13g2_fill_1 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_fill_2 FILLER_27_312 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_decap_4 FILLER_27_384 ();
 sg13g2_fill_2 FILLER_27_388 ();
 sg13g2_fill_1 FILLER_27_406 ();
 sg13g2_fill_2 FILLER_27_436 ();
 sg13g2_decap_8 FILLER_27_475 ();
 sg13g2_decap_8 FILLER_27_482 ();
 sg13g2_decap_8 FILLER_27_489 ();
 sg13g2_decap_8 FILLER_27_496 ();
 sg13g2_decap_8 FILLER_27_503 ();
 sg13g2_decap_4 FILLER_27_510 ();
 sg13g2_fill_1 FILLER_27_514 ();
 sg13g2_decap_8 FILLER_27_544 ();
 sg13g2_decap_4 FILLER_27_551 ();
 sg13g2_fill_2 FILLER_27_555 ();
 sg13g2_fill_2 FILLER_27_562 ();
 sg13g2_decap_4 FILLER_27_585 ();
 sg13g2_fill_2 FILLER_27_589 ();
 sg13g2_decap_8 FILLER_27_629 ();
 sg13g2_fill_2 FILLER_27_636 ();
 sg13g2_fill_1 FILLER_27_638 ();
 sg13g2_fill_1 FILLER_27_680 ();
 sg13g2_fill_2 FILLER_27_694 ();
 sg13g2_fill_1 FILLER_27_696 ();
 sg13g2_fill_2 FILLER_27_708 ();
 sg13g2_fill_1 FILLER_27_729 ();
 sg13g2_decap_8 FILLER_27_738 ();
 sg13g2_decap_4 FILLER_27_745 ();
 sg13g2_decap_8 FILLER_27_754 ();
 sg13g2_fill_1 FILLER_27_761 ();
 sg13g2_fill_2 FILLER_27_770 ();
 sg13g2_fill_2 FILLER_27_780 ();
 sg13g2_fill_1 FILLER_27_795 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_4 FILLER_27_819 ();
 sg13g2_fill_1 FILLER_27_826 ();
 sg13g2_fill_2 FILLER_27_831 ();
 sg13g2_decap_8 FILLER_27_837 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_4 FILLER_27_851 ();
 sg13g2_decap_8 FILLER_27_904 ();
 sg13g2_decap_8 FILLER_27_911 ();
 sg13g2_fill_2 FILLER_27_918 ();
 sg13g2_fill_1 FILLER_27_920 ();
 sg13g2_decap_8 FILLER_27_944 ();
 sg13g2_decap_8 FILLER_27_951 ();
 sg13g2_decap_4 FILLER_27_958 ();
 sg13g2_fill_1 FILLER_27_962 ();
 sg13g2_decap_4 FILLER_27_967 ();
 sg13g2_fill_1 FILLER_27_976 ();
 sg13g2_decap_8 FILLER_27_981 ();
 sg13g2_fill_1 FILLER_27_988 ();
 sg13g2_decap_8 FILLER_27_992 ();
 sg13g2_decap_8 FILLER_27_1027 ();
 sg13g2_fill_2 FILLER_27_1034 ();
 sg13g2_decap_8 FILLER_27_1041 ();
 sg13g2_decap_4 FILLER_27_1048 ();
 sg13g2_fill_2 FILLER_27_1063 ();
 sg13g2_decap_8 FILLER_27_1069 ();
 sg13g2_fill_2 FILLER_27_1076 ();
 sg13g2_fill_1 FILLER_27_1078 ();
 sg13g2_fill_2 FILLER_27_1105 ();
 sg13g2_decap_8 FILLER_27_1111 ();
 sg13g2_decap_4 FILLER_27_1118 ();
 sg13g2_fill_1 FILLER_27_1122 ();
 sg13g2_decap_8 FILLER_27_1156 ();
 sg13g2_fill_2 FILLER_27_1163 ();
 sg13g2_fill_1 FILLER_27_1165 ();
 sg13g2_decap_8 FILLER_27_1220 ();
 sg13g2_decap_4 FILLER_27_1227 ();
 sg13g2_fill_2 FILLER_27_1231 ();
 sg13g2_fill_1 FILLER_27_1240 ();
 sg13g2_decap_8 FILLER_27_1245 ();
 sg13g2_fill_2 FILLER_27_1252 ();
 sg13g2_fill_1 FILLER_27_1254 ();
 sg13g2_decap_8 FILLER_27_1259 ();
 sg13g2_fill_1 FILLER_27_1266 ();
 sg13g2_fill_2 FILLER_27_1280 ();
 sg13g2_fill_1 FILLER_27_1282 ();
 sg13g2_decap_8 FILLER_27_1297 ();
 sg13g2_decap_8 FILLER_27_1304 ();
 sg13g2_decap_8 FILLER_27_1319 ();
 sg13g2_decap_4 FILLER_27_1326 ();
 sg13g2_fill_2 FILLER_27_1330 ();
 sg13g2_decap_4 FILLER_27_1353 ();
 sg13g2_fill_2 FILLER_27_1357 ();
 sg13g2_decap_4 FILLER_27_1379 ();
 sg13g2_fill_2 FILLER_27_1383 ();
 sg13g2_fill_1 FILLER_27_1411 ();
 sg13g2_decap_8 FILLER_27_1420 ();
 sg13g2_decap_8 FILLER_27_1427 ();
 sg13g2_decap_8 FILLER_27_1439 ();
 sg13g2_decap_8 FILLER_27_1446 ();
 sg13g2_decap_4 FILLER_27_1453 ();
 sg13g2_fill_1 FILLER_27_1457 ();
 sg13g2_fill_2 FILLER_27_1507 ();
 sg13g2_fill_1 FILLER_27_1509 ();
 sg13g2_fill_2 FILLER_27_1523 ();
 sg13g2_fill_1 FILLER_27_1525 ();
 sg13g2_decap_8 FILLER_27_1552 ();
 sg13g2_fill_1 FILLER_27_1559 ();
 sg13g2_fill_1 FILLER_27_1581 ();
 sg13g2_fill_2 FILLER_27_1587 ();
 sg13g2_decap_4 FILLER_27_1612 ();
 sg13g2_fill_1 FILLER_27_1616 ();
 sg13g2_decap_8 FILLER_27_1621 ();
 sg13g2_decap_4 FILLER_27_1628 ();
 sg13g2_fill_2 FILLER_27_1632 ();
 sg13g2_decap_8 FILLER_27_1661 ();
 sg13g2_fill_2 FILLER_27_1668 ();
 sg13g2_fill_1 FILLER_27_1670 ();
 sg13g2_decap_8 FILLER_27_1699 ();
 sg13g2_fill_1 FILLER_27_1722 ();
 sg13g2_decap_8 FILLER_27_1737 ();
 sg13g2_fill_2 FILLER_27_1744 ();
 sg13g2_fill_1 FILLER_27_1765 ();
 sg13g2_decap_8 FILLER_27_1770 ();
 sg13g2_decap_8 FILLER_27_1777 ();
 sg13g2_decap_8 FILLER_27_1784 ();
 sg13g2_decap_8 FILLER_27_1791 ();
 sg13g2_fill_2 FILLER_27_1810 ();
 sg13g2_fill_1 FILLER_27_1828 ();
 sg13g2_decap_4 FILLER_27_1838 ();
 sg13g2_fill_2 FILLER_27_1846 ();
 sg13g2_fill_1 FILLER_27_1848 ();
 sg13g2_decap_8 FILLER_27_1857 ();
 sg13g2_fill_1 FILLER_27_1864 ();
 sg13g2_fill_2 FILLER_27_1870 ();
 sg13g2_fill_2 FILLER_27_1884 ();
 sg13g2_fill_1 FILLER_27_1886 ();
 sg13g2_decap_8 FILLER_27_1900 ();
 sg13g2_decap_8 FILLER_27_1907 ();
 sg13g2_fill_2 FILLER_27_1914 ();
 sg13g2_fill_1 FILLER_27_1916 ();
 sg13g2_decap_4 FILLER_27_1935 ();
 sg13g2_fill_2 FILLER_27_1939 ();
 sg13g2_decap_8 FILLER_27_1958 ();
 sg13g2_decap_4 FILLER_27_1965 ();
 sg13g2_fill_2 FILLER_27_1969 ();
 sg13g2_fill_1 FILLER_27_1975 ();
 sg13g2_decap_8 FILLER_27_1997 ();
 sg13g2_decap_4 FILLER_27_2022 ();
 sg13g2_fill_1 FILLER_27_2026 ();
 sg13g2_decap_8 FILLER_27_2038 ();
 sg13g2_decap_8 FILLER_27_2045 ();
 sg13g2_decap_4 FILLER_27_2052 ();
 sg13g2_fill_1 FILLER_27_2056 ();
 sg13g2_decap_8 FILLER_27_2070 ();
 sg13g2_decap_4 FILLER_27_2077 ();
 sg13g2_fill_1 FILLER_27_2081 ();
 sg13g2_decap_8 FILLER_27_2087 ();
 sg13g2_fill_2 FILLER_27_2094 ();
 sg13g2_fill_1 FILLER_27_2096 ();
 sg13g2_decap_4 FILLER_27_2109 ();
 sg13g2_decap_8 FILLER_27_2121 ();
 sg13g2_fill_2 FILLER_27_2128 ();
 sg13g2_decap_8 FILLER_27_2134 ();
 sg13g2_decap_4 FILLER_27_2141 ();
 sg13g2_fill_1 FILLER_27_2145 ();
 sg13g2_fill_2 FILLER_27_2154 ();
 sg13g2_fill_1 FILLER_27_2156 ();
 sg13g2_fill_1 FILLER_27_2163 ();
 sg13g2_fill_2 FILLER_27_2170 ();
 sg13g2_fill_1 FILLER_27_2172 ();
 sg13g2_fill_1 FILLER_27_2182 ();
 sg13g2_fill_2 FILLER_27_2209 ();
 sg13g2_fill_1 FILLER_27_2262 ();
 sg13g2_fill_2 FILLER_27_2285 ();
 sg13g2_fill_2 FILLER_27_2295 ();
 sg13g2_fill_1 FILLER_27_2297 ();
 sg13g2_decap_8 FILLER_27_2340 ();
 sg13g2_decap_4 FILLER_27_2347 ();
 sg13g2_fill_1 FILLER_27_2351 ();
 sg13g2_decap_4 FILLER_27_2367 ();
 sg13g2_fill_1 FILLER_27_2371 ();
 sg13g2_decap_4 FILLER_27_2385 ();
 sg13g2_decap_8 FILLER_27_2396 ();
 sg13g2_fill_2 FILLER_27_2403 ();
 sg13g2_fill_2 FILLER_27_2418 ();
 sg13g2_fill_1 FILLER_27_2448 ();
 sg13g2_fill_1 FILLER_27_2474 ();
 sg13g2_fill_2 FILLER_27_2516 ();
 sg13g2_fill_1 FILLER_27_2518 ();
 sg13g2_decap_8 FILLER_27_2536 ();
 sg13g2_decap_8 FILLER_27_2561 ();
 sg13g2_decap_4 FILLER_27_2568 ();
 sg13g2_fill_1 FILLER_27_2572 ();
 sg13g2_fill_1 FILLER_27_2596 ();
 sg13g2_fill_1 FILLER_27_2602 ();
 sg13g2_decap_8 FILLER_27_2613 ();
 sg13g2_decap_4 FILLER_27_2620 ();
 sg13g2_decap_8 FILLER_27_2641 ();
 sg13g2_decap_8 FILLER_27_2648 ();
 sg13g2_fill_2 FILLER_27_2681 ();
 sg13g2_fill_1 FILLER_27_2683 ();
 sg13g2_decap_4 FILLER_27_2693 ();
 sg13g2_fill_2 FILLER_27_2701 ();
 sg13g2_fill_1 FILLER_27_2703 ();
 sg13g2_fill_2 FILLER_27_2762 ();
 sg13g2_decap_8 FILLER_27_2779 ();
 sg13g2_fill_2 FILLER_27_2786 ();
 sg13g2_decap_8 FILLER_27_2816 ();
 sg13g2_fill_2 FILLER_27_2823 ();
 sg13g2_fill_1 FILLER_27_2825 ();
 sg13g2_decap_8 FILLER_27_2830 ();
 sg13g2_decap_8 FILLER_27_2837 ();
 sg13g2_decap_4 FILLER_27_2844 ();
 sg13g2_fill_2 FILLER_27_2848 ();
 sg13g2_decap_4 FILLER_27_2860 ();
 sg13g2_decap_4 FILLER_27_2908 ();
 sg13g2_decap_4 FILLER_27_2940 ();
 sg13g2_decap_4 FILLER_27_2951 ();
 sg13g2_fill_2 FILLER_27_2955 ();
 sg13g2_decap_4 FILLER_27_2983 ();
 sg13g2_fill_1 FILLER_27_3015 ();
 sg13g2_fill_1 FILLER_27_3057 ();
 sg13g2_fill_2 FILLER_27_3086 ();
 sg13g2_decap_4 FILLER_27_3120 ();
 sg13g2_fill_1 FILLER_27_3124 ();
 sg13g2_fill_2 FILLER_27_3185 ();
 sg13g2_decap_8 FILLER_27_3192 ();
 sg13g2_decap_8 FILLER_27_3227 ();
 sg13g2_decap_4 FILLER_27_3234 ();
 sg13g2_decap_8 FILLER_27_3243 ();
 sg13g2_fill_1 FILLER_27_3282 ();
 sg13g2_fill_1 FILLER_27_3288 ();
 sg13g2_fill_1 FILLER_27_3294 ();
 sg13g2_decap_8 FILLER_27_3300 ();
 sg13g2_decap_4 FILLER_27_3307 ();
 sg13g2_fill_2 FILLER_27_3360 ();
 sg13g2_fill_1 FILLER_27_3362 ();
 sg13g2_fill_1 FILLER_27_3374 ();
 sg13g2_fill_1 FILLER_27_3386 ();
 sg13g2_decap_4 FILLER_27_3392 ();
 sg13g2_fill_1 FILLER_27_3396 ();
 sg13g2_decap_8 FILLER_27_3402 ();
 sg13g2_fill_2 FILLER_27_3409 ();
 sg13g2_fill_1 FILLER_27_3411 ();
 sg13g2_fill_1 FILLER_27_3433 ();
 sg13g2_decap_8 FILLER_27_3460 ();
 sg13g2_decap_8 FILLER_27_3467 ();
 sg13g2_decap_8 FILLER_27_3474 ();
 sg13g2_decap_4 FILLER_27_3481 ();
 sg13g2_fill_1 FILLER_27_3485 ();
 sg13g2_decap_4 FILLER_27_3490 ();
 sg13g2_decap_8 FILLER_27_3498 ();
 sg13g2_decap_8 FILLER_27_3505 ();
 sg13g2_decap_8 FILLER_27_3512 ();
 sg13g2_decap_8 FILLER_27_3519 ();
 sg13g2_decap_8 FILLER_27_3526 ();
 sg13g2_decap_8 FILLER_27_3533 ();
 sg13g2_decap_8 FILLER_27_3540 ();
 sg13g2_decap_8 FILLER_27_3547 ();
 sg13g2_decap_8 FILLER_27_3554 ();
 sg13g2_decap_8 FILLER_27_3561 ();
 sg13g2_decap_8 FILLER_27_3568 ();
 sg13g2_decap_4 FILLER_27_3575 ();
 sg13g2_fill_1 FILLER_27_3579 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_decap_4 FILLER_28_85 ();
 sg13g2_fill_2 FILLER_28_107 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_117 ();
 sg13g2_decap_8 FILLER_28_135 ();
 sg13g2_decap_8 FILLER_28_142 ();
 sg13g2_decap_8 FILLER_28_166 ();
 sg13g2_decap_4 FILLER_28_173 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_decap_4 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_237 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_decap_4 FILLER_28_278 ();
 sg13g2_decap_4 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_decap_4 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_decap_4 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_fill_2 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_28_409 ();
 sg13g2_decap_8 FILLER_28_423 ();
 sg13g2_decap_8 FILLER_28_430 ();
 sg13g2_decap_4 FILLER_28_437 ();
 sg13g2_decap_4 FILLER_28_466 ();
 sg13g2_fill_2 FILLER_28_505 ();
 sg13g2_fill_1 FILLER_28_507 ();
 sg13g2_fill_1 FILLER_28_524 ();
 sg13g2_fill_2 FILLER_28_530 ();
 sg13g2_fill_1 FILLER_28_532 ();
 sg13g2_fill_2 FILLER_28_545 ();
 sg13g2_fill_1 FILLER_28_547 ();
 sg13g2_decap_8 FILLER_28_552 ();
 sg13g2_fill_1 FILLER_28_572 ();
 sg13g2_decap_8 FILLER_28_593 ();
 sg13g2_fill_2 FILLER_28_613 ();
 sg13g2_fill_1 FILLER_28_615 ();
 sg13g2_decap_4 FILLER_28_646 ();
 sg13g2_fill_2 FILLER_28_650 ();
 sg13g2_fill_2 FILLER_28_670 ();
 sg13g2_fill_1 FILLER_28_672 ();
 sg13g2_decap_4 FILLER_28_720 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_decap_4 FILLER_28_741 ();
 sg13g2_fill_2 FILLER_28_758 ();
 sg13g2_fill_1 FILLER_28_760 ();
 sg13g2_decap_4 FILLER_28_856 ();
 sg13g2_fill_1 FILLER_28_860 ();
 sg13g2_fill_1 FILLER_28_891 ();
 sg13g2_decap_8 FILLER_28_946 ();
 sg13g2_fill_1 FILLER_28_957 ();
 sg13g2_fill_2 FILLER_28_1001 ();
 sg13g2_fill_1 FILLER_28_1055 ();
 sg13g2_fill_2 FILLER_28_1088 ();
 sg13g2_fill_1 FILLER_28_1090 ();
 sg13g2_decap_4 FILLER_28_1126 ();
 sg13g2_decap_8 FILLER_28_1166 ();
 sg13g2_decap_8 FILLER_28_1225 ();
 sg13g2_decap_4 FILLER_28_1232 ();
 sg13g2_decap_4 FILLER_28_1264 ();
 sg13g2_fill_2 FILLER_28_1281 ();
 sg13g2_decap_4 FILLER_28_1298 ();
 sg13g2_decap_8 FILLER_28_1320 ();
 sg13g2_decap_4 FILLER_28_1327 ();
 sg13g2_fill_2 FILLER_28_1331 ();
 sg13g2_fill_2 FILLER_28_1337 ();
 sg13g2_fill_2 FILLER_28_1349 ();
 sg13g2_decap_8 FILLER_28_1356 ();
 sg13g2_fill_2 FILLER_28_1363 ();
 sg13g2_fill_1 FILLER_28_1365 ();
 sg13g2_fill_2 FILLER_28_1446 ();
 sg13g2_fill_1 FILLER_28_1479 ();
 sg13g2_fill_1 FILLER_28_1506 ();
 sg13g2_decap_8 FILLER_28_1551 ();
 sg13g2_fill_2 FILLER_28_1558 ();
 sg13g2_fill_1 FILLER_28_1560 ();
 sg13g2_fill_1 FILLER_28_1578 ();
 sg13g2_decap_8 FILLER_28_1583 ();
 sg13g2_fill_1 FILLER_28_1590 ();
 sg13g2_decap_8 FILLER_28_1606 ();
 sg13g2_fill_1 FILLER_28_1619 ();
 sg13g2_decap_4 FILLER_28_1636 ();
 sg13g2_fill_2 FILLER_28_1640 ();
 sg13g2_fill_2 FILLER_28_1677 ();
 sg13g2_decap_8 FILLER_28_1697 ();
 sg13g2_decap_8 FILLER_28_1704 ();
 sg13g2_decap_8 FILLER_28_1711 ();
 sg13g2_fill_2 FILLER_28_1718 ();
 sg13g2_fill_1 FILLER_28_1720 ();
 sg13g2_decap_4 FILLER_28_1726 ();
 sg13g2_fill_1 FILLER_28_1730 ();
 sg13g2_decap_8 FILLER_28_1767 ();
 sg13g2_fill_2 FILLER_28_1778 ();
 sg13g2_decap_8 FILLER_28_1784 ();
 sg13g2_decap_8 FILLER_28_1791 ();
 sg13g2_decap_8 FILLER_28_1798 ();
 sg13g2_decap_4 FILLER_28_1805 ();
 sg13g2_decap_8 FILLER_28_1821 ();
 sg13g2_decap_8 FILLER_28_1828 ();
 sg13g2_decap_8 FILLER_28_1835 ();
 sg13g2_fill_2 FILLER_28_1863 ();
 sg13g2_decap_8 FILLER_28_1886 ();
 sg13g2_decap_8 FILLER_28_1893 ();
 sg13g2_decap_4 FILLER_28_1900 ();
 sg13g2_decap_4 FILLER_28_1933 ();
 sg13g2_fill_2 FILLER_28_1937 ();
 sg13g2_decap_4 FILLER_28_1952 ();
 sg13g2_fill_1 FILLER_28_1984 ();
 sg13g2_decap_4 FILLER_28_2002 ();
 sg13g2_fill_2 FILLER_28_2006 ();
 sg13g2_fill_1 FILLER_28_2013 ();
 sg13g2_fill_1 FILLER_28_2019 ();
 sg13g2_fill_2 FILLER_28_2024 ();
 sg13g2_fill_2 FILLER_28_2046 ();
 sg13g2_fill_1 FILLER_28_2048 ();
 sg13g2_fill_2 FILLER_28_2070 ();
 sg13g2_decap_4 FILLER_28_2096 ();
 sg13g2_fill_1 FILLER_28_2100 ();
 sg13g2_decap_4 FILLER_28_2130 ();
 sg13g2_fill_2 FILLER_28_2134 ();
 sg13g2_fill_2 FILLER_28_2152 ();
 sg13g2_fill_1 FILLER_28_2154 ();
 sg13g2_decap_4 FILLER_28_2180 ();
 sg13g2_decap_8 FILLER_28_2200 ();
 sg13g2_decap_4 FILLER_28_2207 ();
 sg13g2_fill_1 FILLER_28_2211 ();
 sg13g2_decap_8 FILLER_28_2233 ();
 sg13g2_fill_1 FILLER_28_2240 ();
 sg13g2_fill_1 FILLER_28_2258 ();
 sg13g2_decap_8 FILLER_28_2272 ();
 sg13g2_fill_1 FILLER_28_2279 ();
 sg13g2_decap_4 FILLER_28_2289 ();
 sg13g2_fill_2 FILLER_28_2293 ();
 sg13g2_decap_4 FILLER_28_2323 ();
 sg13g2_decap_8 FILLER_28_2369 ();
 sg13g2_decap_4 FILLER_28_2376 ();
 sg13g2_fill_2 FILLER_28_2380 ();
 sg13g2_fill_2 FILLER_28_2401 ();
 sg13g2_fill_1 FILLER_28_2403 ();
 sg13g2_decap_4 FILLER_28_2409 ();
 sg13g2_fill_1 FILLER_28_2413 ();
 sg13g2_decap_8 FILLER_28_2425 ();
 sg13g2_decap_8 FILLER_28_2432 ();
 sg13g2_decap_8 FILLER_28_2439 ();
 sg13g2_decap_8 FILLER_28_2446 ();
 sg13g2_decap_4 FILLER_28_2453 ();
 sg13g2_decap_4 FILLER_28_2465 ();
 sg13g2_fill_2 FILLER_28_2487 ();
 sg13g2_fill_1 FILLER_28_2489 ();
 sg13g2_fill_2 FILLER_28_2508 ();
 sg13g2_fill_1 FILLER_28_2510 ();
 sg13g2_fill_2 FILLER_28_2526 ();
 sg13g2_decap_4 FILLER_28_2538 ();
 sg13g2_fill_2 FILLER_28_2542 ();
 sg13g2_decap_8 FILLER_28_2558 ();
 sg13g2_decap_8 FILLER_28_2565 ();
 sg13g2_fill_1 FILLER_28_2581 ();
 sg13g2_fill_2 FILLER_28_2587 ();
 sg13g2_fill_1 FILLER_28_2589 ();
 sg13g2_decap_4 FILLER_28_2602 ();
 sg13g2_decap_4 FILLER_28_2618 ();
 sg13g2_fill_1 FILLER_28_2622 ();
 sg13g2_fill_2 FILLER_28_2636 ();
 sg13g2_decap_4 FILLER_28_2648 ();
 sg13g2_fill_1 FILLER_28_2652 ();
 sg13g2_fill_1 FILLER_28_2681 ();
 sg13g2_decap_4 FILLER_28_2692 ();
 sg13g2_fill_1 FILLER_28_2696 ();
 sg13g2_decap_4 FILLER_28_2727 ();
 sg13g2_decap_8 FILLER_28_2778 ();
 sg13g2_fill_2 FILLER_28_2785 ();
 sg13g2_fill_1 FILLER_28_2787 ();
 sg13g2_fill_2 FILLER_28_2799 ();
 sg13g2_fill_1 FILLER_28_2801 ();
 sg13g2_fill_1 FILLER_28_2815 ();
 sg13g2_fill_2 FILLER_28_2851 ();
 sg13g2_fill_1 FILLER_28_2853 ();
 sg13g2_decap_4 FILLER_28_2876 ();
 sg13g2_decap_8 FILLER_28_2890 ();
 sg13g2_decap_8 FILLER_28_2897 ();
 sg13g2_decap_4 FILLER_28_2914 ();
 sg13g2_fill_1 FILLER_28_2918 ();
 sg13g2_fill_1 FILLER_28_2924 ();
 sg13g2_decap_4 FILLER_28_2930 ();
 sg13g2_fill_1 FILLER_28_2934 ();
 sg13g2_decap_4 FILLER_28_2943 ();
 sg13g2_decap_8 FILLER_28_2960 ();
 sg13g2_decap_4 FILLER_28_2967 ();
 sg13g2_decap_8 FILLER_28_3000 ();
 sg13g2_fill_2 FILLER_28_3007 ();
 sg13g2_decap_8 FILLER_28_3014 ();
 sg13g2_decap_8 FILLER_28_3025 ();
 sg13g2_decap_8 FILLER_28_3032 ();
 sg13g2_decap_4 FILLER_28_3039 ();
 sg13g2_fill_2 FILLER_28_3056 ();
 sg13g2_decap_4 FILLER_28_3078 ();
 sg13g2_fill_1 FILLER_28_3082 ();
 sg13g2_fill_1 FILLER_28_3124 ();
 sg13g2_decap_8 FILLER_28_3142 ();
 sg13g2_fill_2 FILLER_28_3149 ();
 sg13g2_decap_8 FILLER_28_3155 ();
 sg13g2_decap_4 FILLER_28_3167 ();
 sg13g2_fill_1 FILLER_28_3171 ();
 sg13g2_fill_2 FILLER_28_3202 ();
 sg13g2_decap_8 FILLER_28_3208 ();
 sg13g2_fill_1 FILLER_28_3228 ();
 sg13g2_decap_8 FILLER_28_3251 ();
 sg13g2_fill_2 FILLER_28_3281 ();
 sg13g2_decap_8 FILLER_28_3316 ();
 sg13g2_decap_4 FILLER_28_3323 ();
 sg13g2_fill_2 FILLER_28_3327 ();
 sg13g2_fill_1 FILLER_28_3338 ();
 sg13g2_fill_2 FILLER_28_3348 ();
 sg13g2_fill_1 FILLER_28_3350 ();
 sg13g2_decap_4 FILLER_28_3371 ();
 sg13g2_fill_2 FILLER_28_3380 ();
 sg13g2_decap_8 FILLER_28_3390 ();
 sg13g2_decap_4 FILLER_28_3397 ();
 sg13g2_decap_4 FILLER_28_3406 ();
 sg13g2_fill_1 FILLER_28_3410 ();
 sg13g2_decap_8 FILLER_28_3414 ();
 sg13g2_fill_2 FILLER_28_3421 ();
 sg13g2_fill_1 FILLER_28_3423 ();
 sg13g2_decap_4 FILLER_28_3438 ();
 sg13g2_fill_1 FILLER_28_3442 ();
 sg13g2_fill_2 FILLER_28_3451 ();
 sg13g2_decap_4 FILLER_28_3484 ();
 sg13g2_fill_1 FILLER_28_3506 ();
 sg13g2_decap_8 FILLER_28_3516 ();
 sg13g2_decap_8 FILLER_28_3523 ();
 sg13g2_decap_8 FILLER_28_3530 ();
 sg13g2_decap_8 FILLER_28_3537 ();
 sg13g2_decap_8 FILLER_28_3544 ();
 sg13g2_decap_8 FILLER_28_3551 ();
 sg13g2_decap_8 FILLER_28_3558 ();
 sg13g2_decap_8 FILLER_28_3565 ();
 sg13g2_decap_8 FILLER_28_3572 ();
 sg13g2_fill_1 FILLER_28_3579 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_117 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_fill_2 FILLER_29_385 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_decap_4 FILLER_29_410 ();
 sg13g2_fill_1 FILLER_29_414 ();
 sg13g2_decap_4 FILLER_29_419 ();
 sg13g2_fill_2 FILLER_29_423 ();
 sg13g2_decap_4 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_29_446 ();
 sg13g2_decap_4 FILLER_29_452 ();
 sg13g2_fill_1 FILLER_29_456 ();
 sg13g2_fill_1 FILLER_29_475 ();
 sg13g2_decap_8 FILLER_29_493 ();
 sg13g2_decap_4 FILLER_29_518 ();
 sg13g2_fill_1 FILLER_29_522 ();
 sg13g2_decap_4 FILLER_29_528 ();
 sg13g2_fill_1 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_548 ();
 sg13g2_fill_1 FILLER_29_555 ();
 sg13g2_fill_2 FILLER_29_576 ();
 sg13g2_fill_1 FILLER_29_592 ();
 sg13g2_decap_8 FILLER_29_626 ();
 sg13g2_decap_4 FILLER_29_633 ();
 sg13g2_fill_1 FILLER_29_637 ();
 sg13g2_decap_4 FILLER_29_663 ();
 sg13g2_fill_2 FILLER_29_667 ();
 sg13g2_decap_8 FILLER_29_695 ();
 sg13g2_decap_4 FILLER_29_702 ();
 sg13g2_fill_2 FILLER_29_706 ();
 sg13g2_fill_2 FILLER_29_735 ();
 sg13g2_decap_4 FILLER_29_765 ();
 sg13g2_fill_2 FILLER_29_769 ();
 sg13g2_fill_2 FILLER_29_780 ();
 sg13g2_decap_8 FILLER_29_792 ();
 sg13g2_decap_4 FILLER_29_799 ();
 sg13g2_fill_2 FILLER_29_803 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_4 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_4 FILLER_29_842 ();
 sg13g2_fill_2 FILLER_29_846 ();
 sg13g2_fill_1 FILLER_29_891 ();
 sg13g2_fill_2 FILLER_29_904 ();
 sg13g2_decap_8 FILLER_29_966 ();
 sg13g2_decap_4 FILLER_29_973 ();
 sg13g2_fill_2 FILLER_29_977 ();
 sg13g2_fill_2 FILLER_29_984 ();
 sg13g2_fill_1 FILLER_29_986 ();
 sg13g2_decap_8 FILLER_29_1015 ();
 sg13g2_fill_2 FILLER_29_1022 ();
 sg13g2_decap_4 FILLER_29_1029 ();
 sg13g2_decap_4 FILLER_29_1037 ();
 sg13g2_fill_1 FILLER_29_1041 ();
 sg13g2_fill_1 FILLER_29_1055 ();
 sg13g2_decap_8 FILLER_29_1059 ();
 sg13g2_decap_8 FILLER_29_1066 ();
 sg13g2_fill_2 FILLER_29_1073 ();
 sg13g2_fill_1 FILLER_29_1075 ();
 sg13g2_fill_1 FILLER_29_1089 ();
 sg13g2_decap_8 FILLER_29_1113 ();
 sg13g2_decap_4 FILLER_29_1120 ();
 sg13g2_fill_1 FILLER_29_1169 ();
 sg13g2_fill_1 FILLER_29_1209 ();
 sg13g2_decap_8 FILLER_29_1234 ();
 sg13g2_decap_8 FILLER_29_1241 ();
 sg13g2_decap_4 FILLER_29_1258 ();
 sg13g2_decap_8 FILLER_29_1275 ();
 sg13g2_fill_2 FILLER_29_1282 ();
 sg13g2_fill_1 FILLER_29_1284 ();
 sg13g2_decap_4 FILLER_29_1302 ();
 sg13g2_fill_2 FILLER_29_1306 ();
 sg13g2_decap_4 FILLER_29_1325 ();
 sg13g2_fill_2 FILLER_29_1329 ();
 sg13g2_fill_2 FILLER_29_1343 ();
 sg13g2_fill_1 FILLER_29_1345 ();
 sg13g2_decap_8 FILLER_29_1366 ();
 sg13g2_decap_8 FILLER_29_1373 ();
 sg13g2_decap_8 FILLER_29_1380 ();
 sg13g2_fill_1 FILLER_29_1399 ();
 sg13g2_fill_1 FILLER_29_1424 ();
 sg13g2_decap_4 FILLER_29_1444 ();
 sg13g2_fill_2 FILLER_29_1448 ();
 sg13g2_fill_1 FILLER_29_1495 ();
 sg13g2_fill_2 FILLER_29_1519 ();
 sg13g2_fill_1 FILLER_29_1542 ();
 sg13g2_decap_4 FILLER_29_1548 ();
 sg13g2_decap_4 FILLER_29_1572 ();
 sg13g2_fill_2 FILLER_29_1576 ();
 sg13g2_decap_8 FILLER_29_1588 ();
 sg13g2_fill_1 FILLER_29_1595 ();
 sg13g2_fill_2 FILLER_29_1601 ();
 sg13g2_fill_1 FILLER_29_1603 ();
 sg13g2_fill_2 FILLER_29_1622 ();
 sg13g2_decap_4 FILLER_29_1648 ();
 sg13g2_fill_2 FILLER_29_1652 ();
 sg13g2_fill_2 FILLER_29_1658 ();
 sg13g2_fill_1 FILLER_29_1660 ();
 sg13g2_decap_4 FILLER_29_1666 ();
 sg13g2_fill_1 FILLER_29_1670 ();
 sg13g2_fill_2 FILLER_29_1676 ();
 sg13g2_fill_1 FILLER_29_1678 ();
 sg13g2_fill_1 FILLER_29_1691 ();
 sg13g2_fill_2 FILLER_29_1724 ();
 sg13g2_fill_1 FILLER_29_1726 ();
 sg13g2_decap_4 FILLER_29_1736 ();
 sg13g2_decap_8 FILLER_29_1744 ();
 sg13g2_fill_2 FILLER_29_1751 ();
 sg13g2_fill_1 FILLER_29_1753 ();
 sg13g2_fill_2 FILLER_29_1764 ();
 sg13g2_decap_4 FILLER_29_1771 ();
 sg13g2_fill_1 FILLER_29_1803 ();
 sg13g2_decap_8 FILLER_29_1840 ();
 sg13g2_fill_2 FILLER_29_1847 ();
 sg13g2_fill_1 FILLER_29_1849 ();
 sg13g2_decap_8 FILLER_29_1860 ();
 sg13g2_fill_2 FILLER_29_1867 ();
 sg13g2_decap_4 FILLER_29_1915 ();
 sg13g2_fill_1 FILLER_29_1919 ();
 sg13g2_decap_8 FILLER_29_1934 ();
 sg13g2_decap_4 FILLER_29_1941 ();
 sg13g2_fill_1 FILLER_29_1975 ();
 sg13g2_fill_2 FILLER_29_1990 ();
 sg13g2_fill_1 FILLER_29_1992 ();
 sg13g2_decap_8 FILLER_29_1998 ();
 sg13g2_fill_1 FILLER_29_2005 ();
 sg13g2_decap_4 FILLER_29_2018 ();
 sg13g2_fill_1 FILLER_29_2022 ();
 sg13g2_fill_1 FILLER_29_2028 ();
 sg13g2_fill_1 FILLER_29_2034 ();
 sg13g2_fill_1 FILLER_29_2045 ();
 sg13g2_decap_4 FILLER_29_2051 ();
 sg13g2_fill_1 FILLER_29_2055 ();
 sg13g2_decap_8 FILLER_29_2072 ();
 sg13g2_fill_2 FILLER_29_2079 ();
 sg13g2_decap_8 FILLER_29_2099 ();
 sg13g2_decap_4 FILLER_29_2106 ();
 sg13g2_fill_2 FILLER_29_2110 ();
 sg13g2_decap_8 FILLER_29_2123 ();
 sg13g2_decap_8 FILLER_29_2130 ();
 sg13g2_fill_2 FILLER_29_2150 ();
 sg13g2_fill_1 FILLER_29_2165 ();
 sg13g2_fill_2 FILLER_29_2177 ();
 sg13g2_fill_1 FILLER_29_2179 ();
 sg13g2_decap_8 FILLER_29_2203 ();
 sg13g2_decap_8 FILLER_29_2210 ();
 sg13g2_fill_2 FILLER_29_2217 ();
 sg13g2_decap_8 FILLER_29_2224 ();
 sg13g2_decap_4 FILLER_29_2231 ();
 sg13g2_fill_1 FILLER_29_2235 ();
 sg13g2_decap_8 FILLER_29_2252 ();
 sg13g2_fill_2 FILLER_29_2274 ();
 sg13g2_decap_4 FILLER_29_2312 ();
 sg13g2_fill_1 FILLER_29_2316 ();
 sg13g2_fill_1 FILLER_29_2358 ();
 sg13g2_decap_8 FILLER_29_2377 ();
 sg13g2_decap_4 FILLER_29_2392 ();
 sg13g2_fill_1 FILLER_29_2396 ();
 sg13g2_fill_2 FILLER_29_2405 ();
 sg13g2_fill_2 FILLER_29_2413 ();
 sg13g2_fill_1 FILLER_29_2420 ();
 sg13g2_fill_1 FILLER_29_2426 ();
 sg13g2_fill_2 FILLER_29_2447 ();
 sg13g2_fill_1 FILLER_29_2449 ();
 sg13g2_decap_8 FILLER_29_2482 ();
 sg13g2_decap_8 FILLER_29_2489 ();
 sg13g2_fill_2 FILLER_29_2496 ();
 sg13g2_fill_2 FILLER_29_2513 ();
 sg13g2_fill_1 FILLER_29_2515 ();
 sg13g2_decap_4 FILLER_29_2524 ();
 sg13g2_fill_2 FILLER_29_2546 ();
 sg13g2_fill_1 FILLER_29_2548 ();
 sg13g2_fill_1 FILLER_29_2562 ();
 sg13g2_decap_4 FILLER_29_2580 ();
 sg13g2_decap_8 FILLER_29_2596 ();
 sg13g2_fill_2 FILLER_29_2603 ();
 sg13g2_fill_1 FILLER_29_2605 ();
 sg13g2_fill_1 FILLER_29_2616 ();
 sg13g2_decap_8 FILLER_29_2626 ();
 sg13g2_fill_1 FILLER_29_2633 ();
 sg13g2_decap_4 FILLER_29_2660 ();
 sg13g2_fill_1 FILLER_29_2664 ();
 sg13g2_decap_8 FILLER_29_2687 ();
 sg13g2_decap_4 FILLER_29_2694 ();
 sg13g2_fill_1 FILLER_29_2712 ();
 sg13g2_fill_2 FILLER_29_2731 ();
 sg13g2_decap_8 FILLER_29_2737 ();
 sg13g2_fill_2 FILLER_29_2744 ();
 sg13g2_fill_2 FILLER_29_2754 ();
 sg13g2_fill_1 FILLER_29_2756 ();
 sg13g2_decap_4 FILLER_29_2762 ();
 sg13g2_decap_8 FILLER_29_2776 ();
 sg13g2_decap_8 FILLER_29_2783 ();
 sg13g2_fill_1 FILLER_29_2795 ();
 sg13g2_fill_2 FILLER_29_2826 ();
 sg13g2_decap_8 FILLER_29_2832 ();
 sg13g2_decap_8 FILLER_29_2839 ();
 sg13g2_fill_1 FILLER_29_2846 ();
 sg13g2_decap_8 FILLER_29_2861 ();
 sg13g2_fill_1 FILLER_29_2868 ();
 sg13g2_decap_4 FILLER_29_2890 ();
 sg13g2_fill_2 FILLER_29_2917 ();
 sg13g2_fill_1 FILLER_29_2919 ();
 sg13g2_decap_8 FILLER_29_2930 ();
 sg13g2_decap_4 FILLER_29_2937 ();
 sg13g2_fill_2 FILLER_29_2946 ();
 sg13g2_fill_1 FILLER_29_2953 ();
 sg13g2_decap_8 FILLER_29_2967 ();
 sg13g2_decap_4 FILLER_29_2974 ();
 sg13g2_fill_1 FILLER_29_2978 ();
 sg13g2_fill_2 FILLER_29_2985 ();
 sg13g2_fill_1 FILLER_29_2987 ();
 sg13g2_fill_2 FILLER_29_3003 ();
 sg13g2_fill_1 FILLER_29_3005 ();
 sg13g2_decap_8 FILLER_29_3027 ();
 sg13g2_decap_4 FILLER_29_3034 ();
 sg13g2_fill_2 FILLER_29_3038 ();
 sg13g2_decap_8 FILLER_29_3048 ();
 sg13g2_decap_8 FILLER_29_3055 ();
 sg13g2_decap_8 FILLER_29_3062 ();
 sg13g2_decap_4 FILLER_29_3069 ();
 sg13g2_fill_1 FILLER_29_3077 ();
 sg13g2_decap_8 FILLER_29_3091 ();
 sg13g2_fill_1 FILLER_29_3098 ();
 sg13g2_decap_4 FILLER_29_3110 ();
 sg13g2_fill_2 FILLER_29_3119 ();
 sg13g2_fill_1 FILLER_29_3121 ();
 sg13g2_decap_8 FILLER_29_3173 ();
 sg13g2_fill_2 FILLER_29_3180 ();
 sg13g2_decap_4 FILLER_29_3192 ();
 sg13g2_fill_2 FILLER_29_3196 ();
 sg13g2_fill_2 FILLER_29_3215 ();
 sg13g2_decap_4 FILLER_29_3229 ();
 sg13g2_fill_1 FILLER_29_3233 ();
 sg13g2_decap_4 FILLER_29_3241 ();
 sg13g2_fill_2 FILLER_29_3245 ();
 sg13g2_fill_1 FILLER_29_3252 ();
 sg13g2_fill_2 FILLER_29_3265 ();
 sg13g2_decap_8 FILLER_29_3277 ();
 sg13g2_decap_8 FILLER_29_3284 ();
 sg13g2_fill_1 FILLER_29_3305 ();
 sg13g2_fill_2 FILLER_29_3354 ();
 sg13g2_fill_1 FILLER_29_3356 ();
 sg13g2_fill_2 FILLER_29_3369 ();
 sg13g2_decap_4 FILLER_29_3398 ();
 sg13g2_fill_2 FILLER_29_3410 ();
 sg13g2_fill_2 FILLER_29_3420 ();
 sg13g2_decap_8 FILLER_29_3436 ();
 sg13g2_fill_2 FILLER_29_3456 ();
 sg13g2_decap_4 FILLER_29_3483 ();
 sg13g2_fill_2 FILLER_29_3487 ();
 sg13g2_decap_8 FILLER_29_3521 ();
 sg13g2_decap_8 FILLER_29_3528 ();
 sg13g2_decap_8 FILLER_29_3535 ();
 sg13g2_decap_8 FILLER_29_3542 ();
 sg13g2_decap_8 FILLER_29_3549 ();
 sg13g2_decap_8 FILLER_29_3556 ();
 sg13g2_decap_8 FILLER_29_3563 ();
 sg13g2_decap_8 FILLER_29_3570 ();
 sg13g2_fill_2 FILLER_29_3577 ();
 sg13g2_fill_1 FILLER_29_3579 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_decap_8 FILLER_30_73 ();
 sg13g2_decap_8 FILLER_30_80 ();
 sg13g2_decap_4 FILLER_30_87 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_decap_4 FILLER_30_155 ();
 sg13g2_fill_2 FILLER_30_159 ();
 sg13g2_decap_8 FILLER_30_185 ();
 sg13g2_decap_8 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_decap_4 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_234 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_decap_8 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_330 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_decap_4 FILLER_30_351 ();
 sg13g2_fill_2 FILLER_30_355 ();
 sg13g2_decap_4 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_401 ();
 sg13g2_fill_2 FILLER_30_414 ();
 sg13g2_fill_2 FILLER_30_430 ();
 sg13g2_fill_1 FILLER_30_432 ();
 sg13g2_fill_1 FILLER_30_438 ();
 sg13g2_fill_1 FILLER_30_444 ();
 sg13g2_fill_2 FILLER_30_453 ();
 sg13g2_decap_8 FILLER_30_467 ();
 sg13g2_decap_8 FILLER_30_474 ();
 sg13g2_decap_4 FILLER_30_481 ();
 sg13g2_fill_2 FILLER_30_499 ();
 sg13g2_fill_2 FILLER_30_509 ();
 sg13g2_fill_1 FILLER_30_511 ();
 sg13g2_fill_2 FILLER_30_524 ();
 sg13g2_fill_2 FILLER_30_546 ();
 sg13g2_fill_1 FILLER_30_548 ();
 sg13g2_decap_8 FILLER_30_573 ();
 sg13g2_decap_8 FILLER_30_580 ();
 sg13g2_fill_1 FILLER_30_587 ();
 sg13g2_decap_4 FILLER_30_605 ();
 sg13g2_fill_1 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_618 ();
 sg13g2_decap_4 FILLER_30_625 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_4 FILLER_30_644 ();
 sg13g2_fill_1 FILLER_30_648 ();
 sg13g2_decap_8 FILLER_30_654 ();
 sg13g2_decap_8 FILLER_30_661 ();
 sg13g2_decap_4 FILLER_30_668 ();
 sg13g2_decap_8 FILLER_30_692 ();
 sg13g2_decap_8 FILLER_30_699 ();
 sg13g2_decap_4 FILLER_30_706 ();
 sg13g2_fill_1 FILLER_30_731 ();
 sg13g2_fill_2 FILLER_30_741 ();
 sg13g2_fill_1 FILLER_30_751 ();
 sg13g2_decap_4 FILLER_30_794 ();
 sg13g2_decap_4 FILLER_30_818 ();
 sg13g2_fill_1 FILLER_30_822 ();
 sg13g2_fill_2 FILLER_30_844 ();
 sg13g2_fill_1 FILLER_30_846 ();
 sg13g2_decap_4 FILLER_30_858 ();
 sg13g2_decap_4 FILLER_30_866 ();
 sg13g2_fill_2 FILLER_30_870 ();
 sg13g2_decap_4 FILLER_30_946 ();
 sg13g2_fill_2 FILLER_30_966 ();
 sg13g2_fill_1 FILLER_30_968 ();
 sg13g2_fill_1 FILLER_30_992 ();
 sg13g2_decap_8 FILLER_30_997 ();
 sg13g2_decap_8 FILLER_30_1004 ();
 sg13g2_decap_4 FILLER_30_1011 ();
 sg13g2_decap_4 FILLER_30_1065 ();
 sg13g2_decap_8 FILLER_30_1097 ();
 sg13g2_fill_2 FILLER_30_1109 ();
 sg13g2_fill_1 FILLER_30_1111 ();
 sg13g2_decap_8 FILLER_30_1140 ();
 sg13g2_decap_8 FILLER_30_1147 ();
 sg13g2_fill_1 FILLER_30_1154 ();
 sg13g2_decap_8 FILLER_30_1171 ();
 sg13g2_decap_4 FILLER_30_1178 ();
 sg13g2_fill_2 FILLER_30_1182 ();
 sg13g2_fill_1 FILLER_30_1197 ();
 sg13g2_fill_1 FILLER_30_1216 ();
 sg13g2_decap_4 FILLER_30_1238 ();
 sg13g2_fill_2 FILLER_30_1275 ();
 sg13g2_decap_8 FILLER_30_1285 ();
 sg13g2_decap_4 FILLER_30_1292 ();
 sg13g2_fill_2 FILLER_30_1296 ();
 sg13g2_fill_1 FILLER_30_1304 ();
 sg13g2_fill_2 FILLER_30_1310 ();
 sg13g2_fill_2 FILLER_30_1329 ();
 sg13g2_fill_1 FILLER_30_1331 ();
 sg13g2_fill_1 FILLER_30_1360 ();
 sg13g2_decap_8 FILLER_30_1369 ();
 sg13g2_fill_1 FILLER_30_1376 ();
 sg13g2_fill_2 FILLER_30_1395 ();
 sg13g2_fill_2 FILLER_30_1405 ();
 sg13g2_decap_4 FILLER_30_1422 ();
 sg13g2_fill_2 FILLER_30_1426 ();
 sg13g2_fill_2 FILLER_30_1479 ();
 sg13g2_fill_1 FILLER_30_1520 ();
 sg13g2_fill_2 FILLER_30_1526 ();
 sg13g2_decap_4 FILLER_30_1546 ();
 sg13g2_fill_2 FILLER_30_1550 ();
 sg13g2_fill_1 FILLER_30_1565 ();
 sg13g2_decap_4 FILLER_30_1577 ();
 sg13g2_decap_8 FILLER_30_1586 ();
 sg13g2_decap_4 FILLER_30_1593 ();
 sg13g2_fill_2 FILLER_30_1603 ();
 sg13g2_fill_1 FILLER_30_1622 ();
 sg13g2_decap_4 FILLER_30_1628 ();
 sg13g2_fill_1 FILLER_30_1632 ();
 sg13g2_decap_8 FILLER_30_1650 ();
 sg13g2_decap_4 FILLER_30_1657 ();
 sg13g2_fill_1 FILLER_30_1661 ();
 sg13g2_fill_1 FILLER_30_1678 ();
 sg13g2_decap_8 FILLER_30_1692 ();
 sg13g2_fill_2 FILLER_30_1699 ();
 sg13g2_fill_1 FILLER_30_1701 ();
 sg13g2_decap_8 FILLER_30_1706 ();
 sg13g2_fill_2 FILLER_30_1713 ();
 sg13g2_fill_2 FILLER_30_1730 ();
 sg13g2_fill_2 FILLER_30_1741 ();
 sg13g2_fill_2 FILLER_30_1754 ();
 sg13g2_decap_8 FILLER_30_1776 ();
 sg13g2_decap_8 FILLER_30_1795 ();
 sg13g2_fill_2 FILLER_30_1802 ();
 sg13g2_fill_1 FILLER_30_1804 ();
 sg13g2_fill_2 FILLER_30_1837 ();
 sg13g2_fill_1 FILLER_30_1850 ();
 sg13g2_fill_2 FILLER_30_1864 ();
 sg13g2_decap_4 FILLER_30_1871 ();
 sg13g2_fill_1 FILLER_30_1893 ();
 sg13g2_fill_1 FILLER_30_1904 ();
 sg13g2_decap_8 FILLER_30_1910 ();
 sg13g2_decap_4 FILLER_30_1917 ();
 sg13g2_fill_1 FILLER_30_1925 ();
 sg13g2_decap_8 FILLER_30_1939 ();
 sg13g2_decap_8 FILLER_30_1946 ();
 sg13g2_decap_4 FILLER_30_1981 ();
 sg13g2_decap_8 FILLER_30_1989 ();
 sg13g2_decap_4 FILLER_30_1996 ();
 sg13g2_decap_8 FILLER_30_2014 ();
 sg13g2_decap_8 FILLER_30_2021 ();
 sg13g2_fill_2 FILLER_30_2028 ();
 sg13g2_fill_1 FILLER_30_2033 ();
 sg13g2_fill_2 FILLER_30_2047 ();
 sg13g2_decap_8 FILLER_30_2076 ();
 sg13g2_fill_2 FILLER_30_2083 ();
 sg13g2_fill_1 FILLER_30_2085 ();
 sg13g2_decap_8 FILLER_30_2094 ();
 sg13g2_decap_8 FILLER_30_2101 ();
 sg13g2_fill_2 FILLER_30_2108 ();
 sg13g2_decap_8 FILLER_30_2130 ();
 sg13g2_fill_2 FILLER_30_2137 ();
 sg13g2_fill_2 FILLER_30_2147 ();
 sg13g2_fill_1 FILLER_30_2149 ();
 sg13g2_fill_1 FILLER_30_2159 ();
 sg13g2_fill_2 FILLER_30_2179 ();
 sg13g2_fill_1 FILLER_30_2181 ();
 sg13g2_decap_4 FILLER_30_2207 ();
 sg13g2_fill_2 FILLER_30_2211 ();
 sg13g2_decap_8 FILLER_30_2234 ();
 sg13g2_fill_2 FILLER_30_2241 ();
 sg13g2_decap_8 FILLER_30_2248 ();
 sg13g2_decap_8 FILLER_30_2276 ();
 sg13g2_decap_4 FILLER_30_2283 ();
 sg13g2_decap_8 FILLER_30_2313 ();
 sg13g2_decap_4 FILLER_30_2320 ();
 sg13g2_fill_2 FILLER_30_2338 ();
 sg13g2_fill_2 FILLER_30_2358 ();
 sg13g2_fill_1 FILLER_30_2360 ();
 sg13g2_decap_4 FILLER_30_2372 ();
 sg13g2_fill_1 FILLER_30_2376 ();
 sg13g2_fill_2 FILLER_30_2399 ();
 sg13g2_fill_1 FILLER_30_2401 ();
 sg13g2_decap_8 FILLER_30_2427 ();
 sg13g2_decap_8 FILLER_30_2434 ();
 sg13g2_fill_2 FILLER_30_2441 ();
 sg13g2_fill_1 FILLER_30_2459 ();
 sg13g2_fill_2 FILLER_30_2465 ();
 sg13g2_decap_4 FILLER_30_2489 ();
 sg13g2_fill_2 FILLER_30_2521 ();
 sg13g2_fill_2 FILLER_30_2528 ();
 sg13g2_fill_1 FILLER_30_2530 ();
 sg13g2_fill_1 FILLER_30_2558 ();
 sg13g2_fill_2 FILLER_30_2569 ();
 sg13g2_fill_1 FILLER_30_2571 ();
 sg13g2_decap_4 FILLER_30_2576 ();
 sg13g2_decap_4 FILLER_30_2607 ();
 sg13g2_fill_1 FILLER_30_2626 ();
 sg13g2_fill_2 FILLER_30_2635 ();
 sg13g2_fill_1 FILLER_30_2637 ();
 sg13g2_decap_8 FILLER_30_2658 ();
 sg13g2_decap_4 FILLER_30_2693 ();
 sg13g2_fill_1 FILLER_30_2697 ();
 sg13g2_decap_4 FILLER_30_2707 ();
 sg13g2_fill_2 FILLER_30_2753 ();
 sg13g2_fill_2 FILLER_30_2782 ();
 sg13g2_fill_2 FILLER_30_2807 ();
 sg13g2_fill_1 FILLER_30_2809 ();
 sg13g2_decap_8 FILLER_30_2822 ();
 sg13g2_fill_2 FILLER_30_2829 ();
 sg13g2_decap_4 FILLER_30_2863 ();
 sg13g2_fill_1 FILLER_30_2867 ();
 sg13g2_decap_8 FILLER_30_2895 ();
 sg13g2_fill_2 FILLER_30_2902 ();
 sg13g2_decap_4 FILLER_30_2917 ();
 sg13g2_fill_1 FILLER_30_2921 ();
 sg13g2_decap_4 FILLER_30_2939 ();
 sg13g2_fill_1 FILLER_30_2943 ();
 sg13g2_decap_8 FILLER_30_2970 ();
 sg13g2_fill_2 FILLER_30_2977 ();
 sg13g2_fill_1 FILLER_30_2979 ();
 sg13g2_decap_4 FILLER_30_2988 ();
 sg13g2_fill_1 FILLER_30_3016 ();
 sg13g2_fill_1 FILLER_30_3033 ();
 sg13g2_fill_2 FILLER_30_3060 ();
 sg13g2_fill_2 FILLER_30_3066 ();
 sg13g2_fill_1 FILLER_30_3068 ();
 sg13g2_fill_1 FILLER_30_3108 ();
 sg13g2_fill_2 FILLER_30_3124 ();
 sg13g2_fill_1 FILLER_30_3126 ();
 sg13g2_decap_8 FILLER_30_3162 ();
 sg13g2_fill_1 FILLER_30_3169 ();
 sg13g2_decap_8 FILLER_30_3186 ();
 sg13g2_decap_4 FILLER_30_3193 ();
 sg13g2_fill_1 FILLER_30_3202 ();
 sg13g2_decap_8 FILLER_30_3221 ();
 sg13g2_fill_2 FILLER_30_3228 ();
 sg13g2_fill_1 FILLER_30_3230 ();
 sg13g2_fill_1 FILLER_30_3267 ();
 sg13g2_decap_8 FILLER_30_3281 ();
 sg13g2_fill_1 FILLER_30_3288 ();
 sg13g2_decap_8 FILLER_30_3309 ();
 sg13g2_fill_2 FILLER_30_3338 ();
 sg13g2_fill_2 FILLER_30_3344 ();
 sg13g2_fill_1 FILLER_30_3346 ();
 sg13g2_fill_2 FILLER_30_3355 ();
 sg13g2_fill_1 FILLER_30_3357 ();
 sg13g2_fill_1 FILLER_30_3366 ();
 sg13g2_decap_4 FILLER_30_3375 ();
 sg13g2_fill_1 FILLER_30_3379 ();
 sg13g2_decap_4 FILLER_30_3398 ();
 sg13g2_fill_1 FILLER_30_3409 ();
 sg13g2_fill_2 FILLER_30_3416 ();
 sg13g2_fill_1 FILLER_30_3426 ();
 sg13g2_decap_8 FILLER_30_3431 ();
 sg13g2_decap_8 FILLER_30_3438 ();
 sg13g2_fill_2 FILLER_30_3453 ();
 sg13g2_decap_4 FILLER_30_3485 ();
 sg13g2_decap_8 FILLER_30_3500 ();
 sg13g2_decap_8 FILLER_30_3507 ();
 sg13g2_decap_8 FILLER_30_3514 ();
 sg13g2_decap_8 FILLER_30_3521 ();
 sg13g2_decap_8 FILLER_30_3528 ();
 sg13g2_decap_8 FILLER_30_3535 ();
 sg13g2_decap_8 FILLER_30_3542 ();
 sg13g2_decap_8 FILLER_30_3549 ();
 sg13g2_decap_8 FILLER_30_3556 ();
 sg13g2_decap_8 FILLER_30_3563 ();
 sg13g2_decap_8 FILLER_30_3570 ();
 sg13g2_fill_2 FILLER_30_3577 ();
 sg13g2_fill_1 FILLER_30_3579 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_111 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_decap_8 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_2 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_236 ();
 sg13g2_fill_1 FILLER_31_243 ();
 sg13g2_decap_8 FILLER_31_249 ();
 sg13g2_fill_2 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_258 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_decap_4 FILLER_31_342 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_31_369 ();
 sg13g2_fill_2 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_445 ();
 sg13g2_fill_2 FILLER_31_452 ();
 sg13g2_fill_1 FILLER_31_454 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_4 FILLER_31_476 ();
 sg13g2_fill_1 FILLER_31_500 ();
 sg13g2_fill_1 FILLER_31_528 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_fill_2 FILLER_31_546 ();
 sg13g2_fill_2 FILLER_31_579 ();
 sg13g2_fill_1 FILLER_31_581 ();
 sg13g2_fill_1 FILLER_31_589 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_fill_2 FILLER_31_622 ();
 sg13g2_fill_2 FILLER_31_652 ();
 sg13g2_fill_1 FILLER_31_654 ();
 sg13g2_fill_2 FILLER_31_702 ();
 sg13g2_decap_8 FILLER_31_712 ();
 sg13g2_decap_4 FILLER_31_719 ();
 sg13g2_fill_1 FILLER_31_723 ();
 sg13g2_fill_1 FILLER_31_744 ();
 sg13g2_fill_1 FILLER_31_750 ();
 sg13g2_fill_1 FILLER_31_760 ();
 sg13g2_decap_8 FILLER_31_765 ();
 sg13g2_fill_1 FILLER_31_772 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_4 FILLER_31_798 ();
 sg13g2_fill_1 FILLER_31_811 ();
 sg13g2_fill_1 FILLER_31_824 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_fill_1 FILLER_31_849 ();
 sg13g2_decap_8 FILLER_31_865 ();
 sg13g2_fill_1 FILLER_31_884 ();
 sg13g2_decap_4 FILLER_31_898 ();
 sg13g2_fill_1 FILLER_31_902 ();
 sg13g2_decap_4 FILLER_31_919 ();
 sg13g2_fill_1 FILLER_31_944 ();
 sg13g2_decap_4 FILLER_31_954 ();
 sg13g2_fill_2 FILLER_31_963 ();
 sg13g2_fill_1 FILLER_31_965 ();
 sg13g2_decap_4 FILLER_31_970 ();
 sg13g2_fill_2 FILLER_31_974 ();
 sg13g2_decap_8 FILLER_31_981 ();
 sg13g2_decap_4 FILLER_31_988 ();
 sg13g2_fill_1 FILLER_31_992 ();
 sg13g2_decap_8 FILLER_31_1035 ();
 sg13g2_fill_2 FILLER_31_1042 ();
 sg13g2_fill_1 FILLER_31_1044 ();
 sg13g2_decap_4 FILLER_31_1070 ();
 sg13g2_fill_1 FILLER_31_1074 ();
 sg13g2_decap_8 FILLER_31_1087 ();
 sg13g2_fill_2 FILLER_31_1094 ();
 sg13g2_decap_4 FILLER_31_1104 ();
 sg13g2_fill_2 FILLER_31_1128 ();
 sg13g2_fill_2 FILLER_31_1142 ();
 sg13g2_fill_1 FILLER_31_1144 ();
 sg13g2_decap_4 FILLER_31_1148 ();
 sg13g2_fill_1 FILLER_31_1152 ();
 sg13g2_fill_2 FILLER_31_1181 ();
 sg13g2_fill_2 FILLER_31_1221 ();
 sg13g2_fill_1 FILLER_31_1223 ();
 sg13g2_decap_8 FILLER_31_1229 ();
 sg13g2_decap_4 FILLER_31_1236 ();
 sg13g2_decap_4 FILLER_31_1250 ();
 sg13g2_fill_1 FILLER_31_1254 ();
 sg13g2_decap_4 FILLER_31_1280 ();
 sg13g2_fill_2 FILLER_31_1289 ();
 sg13g2_fill_1 FILLER_31_1291 ();
 sg13g2_decap_4 FILLER_31_1305 ();
 sg13g2_fill_2 FILLER_31_1309 ();
 sg13g2_fill_2 FILLER_31_1319 ();
 sg13g2_fill_1 FILLER_31_1321 ();
 sg13g2_decap_4 FILLER_31_1328 ();
 sg13g2_fill_1 FILLER_31_1332 ();
 sg13g2_fill_2 FILLER_31_1337 ();
 sg13g2_decap_8 FILLER_31_1366 ();
 sg13g2_decap_8 FILLER_31_1373 ();
 sg13g2_fill_1 FILLER_31_1380 ();
 sg13g2_decap_8 FILLER_31_1395 ();
 sg13g2_fill_1 FILLER_31_1402 ();
 sg13g2_decap_4 FILLER_31_1407 ();
 sg13g2_fill_2 FILLER_31_1411 ();
 sg13g2_fill_2 FILLER_31_1425 ();
 sg13g2_fill_2 FILLER_31_1432 ();
 sg13g2_fill_1 FILLER_31_1434 ();
 sg13g2_fill_1 FILLER_31_1462 ();
 sg13g2_decap_8 FILLER_31_1480 ();
 sg13g2_fill_2 FILLER_31_1487 ();
 sg13g2_fill_1 FILLER_31_1489 ();
 sg13g2_fill_2 FILLER_31_1511 ();
 sg13g2_fill_1 FILLER_31_1513 ();
 sg13g2_fill_2 FILLER_31_1524 ();
 sg13g2_decap_4 FILLER_31_1541 ();
 sg13g2_fill_1 FILLER_31_1545 ();
 sg13g2_fill_1 FILLER_31_1571 ();
 sg13g2_fill_2 FILLER_31_1576 ();
 sg13g2_fill_1 FILLER_31_1586 ();
 sg13g2_decap_4 FILLER_31_1599 ();
 sg13g2_fill_1 FILLER_31_1611 ();
 sg13g2_fill_1 FILLER_31_1622 ();
 sg13g2_decap_8 FILLER_31_1633 ();
 sg13g2_decap_4 FILLER_31_1640 ();
 sg13g2_fill_1 FILLER_31_1644 ();
 sg13g2_fill_1 FILLER_31_1662 ();
 sg13g2_fill_2 FILLER_31_1672 ();
 sg13g2_fill_1 FILLER_31_1674 ();
 sg13g2_fill_2 FILLER_31_1685 ();
 sg13g2_decap_8 FILLER_31_1695 ();
 sg13g2_decap_4 FILLER_31_1702 ();
 sg13g2_fill_1 FILLER_31_1706 ();
 sg13g2_decap_8 FILLER_31_1735 ();
 sg13g2_decap_4 FILLER_31_1742 ();
 sg13g2_fill_2 FILLER_31_1746 ();
 sg13g2_decap_8 FILLER_31_1753 ();
 sg13g2_decap_8 FILLER_31_1760 ();
 sg13g2_fill_2 FILLER_31_1767 ();
 sg13g2_fill_1 FILLER_31_1769 ();
 sg13g2_fill_2 FILLER_31_1807 ();
 sg13g2_fill_1 FILLER_31_1837 ();
 sg13g2_fill_2 FILLER_31_1854 ();
 sg13g2_fill_1 FILLER_31_1856 ();
 sg13g2_decap_4 FILLER_31_1910 ();
 sg13g2_fill_2 FILLER_31_1914 ();
 sg13g2_decap_4 FILLER_31_1941 ();
 sg13g2_fill_1 FILLER_31_1945 ();
 sg13g2_fill_1 FILLER_31_1959 ();
 sg13g2_fill_2 FILLER_31_1971 ();
 sg13g2_decap_8 FILLER_31_1977 ();
 sg13g2_decap_8 FILLER_31_2027 ();
 sg13g2_decap_4 FILLER_31_2034 ();
 sg13g2_decap_8 FILLER_31_2053 ();
 sg13g2_fill_1 FILLER_31_2060 ();
 sg13g2_decap_4 FILLER_31_2077 ();
 sg13g2_decap_4 FILLER_31_2110 ();
 sg13g2_decap_8 FILLER_31_2123 ();
 sg13g2_decap_4 FILLER_31_2130 ();
 sg13g2_fill_2 FILLER_31_2134 ();
 sg13g2_decap_4 FILLER_31_2141 ();
 sg13g2_fill_1 FILLER_31_2145 ();
 sg13g2_fill_2 FILLER_31_2159 ();
 sg13g2_decap_8 FILLER_31_2170 ();
 sg13g2_decap_8 FILLER_31_2177 ();
 sg13g2_fill_2 FILLER_31_2184 ();
 sg13g2_fill_2 FILLER_31_2196 ();
 sg13g2_fill_1 FILLER_31_2198 ();
 sg13g2_fill_2 FILLER_31_2207 ();
 sg13g2_decap_4 FILLER_31_2213 ();
 sg13g2_fill_1 FILLER_31_2217 ();
 sg13g2_decap_4 FILLER_31_2279 ();
 sg13g2_fill_1 FILLER_31_2283 ();
 sg13g2_fill_1 FILLER_31_2318 ();
 sg13g2_fill_2 FILLER_31_2339 ();
 sg13g2_fill_1 FILLER_31_2341 ();
 sg13g2_fill_2 FILLER_31_2358 ();
 sg13g2_fill_1 FILLER_31_2360 ();
 sg13g2_decap_8 FILLER_31_2366 ();
 sg13g2_decap_8 FILLER_31_2373 ();
 sg13g2_fill_2 FILLER_31_2380 ();
 sg13g2_fill_2 FILLER_31_2392 ();
 sg13g2_fill_1 FILLER_31_2394 ();
 sg13g2_fill_2 FILLER_31_2423 ();
 sg13g2_decap_4 FILLER_31_2449 ();
 sg13g2_fill_1 FILLER_31_2453 ();
 sg13g2_fill_2 FILLER_31_2473 ();
 sg13g2_decap_8 FILLER_31_2487 ();
 sg13g2_fill_2 FILLER_31_2511 ();
 sg13g2_fill_2 FILLER_31_2521 ();
 sg13g2_fill_1 FILLER_31_2530 ();
 sg13g2_fill_2 FILLER_31_2549 ();
 sg13g2_fill_1 FILLER_31_2551 ();
 sg13g2_fill_2 FILLER_31_2557 ();
 sg13g2_fill_1 FILLER_31_2559 ();
 sg13g2_decap_4 FILLER_31_2570 ();
 sg13g2_fill_1 FILLER_31_2574 ();
 sg13g2_decap_8 FILLER_31_2594 ();
 sg13g2_decap_8 FILLER_31_2601 ();
 sg13g2_decap_8 FILLER_31_2621 ();
 sg13g2_fill_2 FILLER_31_2628 ();
 sg13g2_fill_1 FILLER_31_2630 ();
 sg13g2_decap_8 FILLER_31_2647 ();
 sg13g2_decap_4 FILLER_31_2654 ();
 sg13g2_fill_2 FILLER_31_2674 ();
 sg13g2_fill_2 FILLER_31_2681 ();
 sg13g2_decap_8 FILLER_31_2688 ();
 sg13g2_fill_2 FILLER_31_2695 ();
 sg13g2_fill_1 FILLER_31_2697 ();
 sg13g2_decap_8 FILLER_31_2717 ();
 sg13g2_fill_1 FILLER_31_2724 ();
 sg13g2_fill_2 FILLER_31_2729 ();
 sg13g2_decap_8 FILLER_31_2735 ();
 sg13g2_decap_4 FILLER_31_2742 ();
 sg13g2_fill_2 FILLER_31_2746 ();
 sg13g2_fill_1 FILLER_31_2752 ();
 sg13g2_decap_8 FILLER_31_2763 ();
 sg13g2_decap_4 FILLER_31_2770 ();
 sg13g2_fill_1 FILLER_31_2774 ();
 sg13g2_fill_1 FILLER_31_2789 ();
 sg13g2_fill_1 FILLER_31_2804 ();
 sg13g2_decap_4 FILLER_31_2827 ();
 sg13g2_fill_1 FILLER_31_2831 ();
 sg13g2_fill_1 FILLER_31_2835 ();
 sg13g2_fill_2 FILLER_31_2845 ();
 sg13g2_decap_4 FILLER_31_2864 ();
 sg13g2_fill_1 FILLER_31_2868 ();
 sg13g2_decap_4 FILLER_31_2875 ();
 sg13g2_fill_1 FILLER_31_2879 ();
 sg13g2_fill_2 FILLER_31_2894 ();
 sg13g2_fill_2 FILLER_31_2941 ();
 sg13g2_fill_1 FILLER_31_2953 ();
 sg13g2_fill_2 FILLER_31_2963 ();
 sg13g2_decap_8 FILLER_31_2975 ();
 sg13g2_decap_4 FILLER_31_2982 ();
 sg13g2_fill_1 FILLER_31_3024 ();
 sg13g2_fill_2 FILLER_31_3035 ();
 sg13g2_decap_8 FILLER_31_3050 ();
 sg13g2_fill_1 FILLER_31_3076 ();
 sg13g2_fill_2 FILLER_31_3082 ();
 sg13g2_fill_1 FILLER_31_3084 ();
 sg13g2_decap_8 FILLER_31_3090 ();
 sg13g2_decap_8 FILLER_31_3097 ();
 sg13g2_fill_2 FILLER_31_3104 ();
 sg13g2_fill_1 FILLER_31_3106 ();
 sg13g2_fill_2 FILLER_31_3112 ();
 sg13g2_fill_2 FILLER_31_3127 ();
 sg13g2_fill_1 FILLER_31_3129 ();
 sg13g2_decap_8 FILLER_31_3138 ();
 sg13g2_fill_1 FILLER_31_3145 ();
 sg13g2_fill_1 FILLER_31_3154 ();
 sg13g2_fill_2 FILLER_31_3173 ();
 sg13g2_fill_1 FILLER_31_3175 ();
 sg13g2_fill_2 FILLER_31_3197 ();
 sg13g2_fill_1 FILLER_31_3199 ();
 sg13g2_fill_1 FILLER_31_3221 ();
 sg13g2_decap_8 FILLER_31_3230 ();
 sg13g2_decap_8 FILLER_31_3237 ();
 sg13g2_fill_1 FILLER_31_3244 ();
 sg13g2_fill_2 FILLER_31_3250 ();
 sg13g2_fill_1 FILLER_31_3252 ();
 sg13g2_fill_1 FILLER_31_3261 ();
 sg13g2_decap_8 FILLER_31_3274 ();
 sg13g2_fill_1 FILLER_31_3294 ();
 sg13g2_decap_8 FILLER_31_3307 ();
 sg13g2_fill_2 FILLER_31_3364 ();
 sg13g2_fill_1 FILLER_31_3420 ();
 sg13g2_fill_1 FILLER_31_3470 ();
 sg13g2_fill_1 FILLER_31_3490 ();
 sg13g2_decap_8 FILLER_31_3519 ();
 sg13g2_decap_8 FILLER_31_3526 ();
 sg13g2_decap_8 FILLER_31_3533 ();
 sg13g2_decap_8 FILLER_31_3540 ();
 sg13g2_decap_8 FILLER_31_3547 ();
 sg13g2_decap_8 FILLER_31_3554 ();
 sg13g2_decap_8 FILLER_31_3561 ();
 sg13g2_decap_8 FILLER_31_3568 ();
 sg13g2_decap_4 FILLER_31_3575 ();
 sg13g2_fill_1 FILLER_31_3579 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_4 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_80 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_fill_2 FILLER_32_156 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_183 ();
 sg13g2_decap_4 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_decap_4 FILLER_32_287 ();
 sg13g2_fill_2 FILLER_32_302 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_decap_4 FILLER_32_388 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_32_414 ();
 sg13g2_fill_2 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_32_444 ();
 sg13g2_decap_4 FILLER_32_476 ();
 sg13g2_fill_2 FILLER_32_499 ();
 sg13g2_fill_1 FILLER_32_501 ();
 sg13g2_decap_4 FILLER_32_507 ();
 sg13g2_fill_1 FILLER_32_511 ();
 sg13g2_fill_1 FILLER_32_529 ();
 sg13g2_decap_8 FILLER_32_542 ();
 sg13g2_decap_8 FILLER_32_549 ();
 sg13g2_decap_8 FILLER_32_556 ();
 sg13g2_fill_2 FILLER_32_563 ();
 sg13g2_fill_1 FILLER_32_565 ();
 sg13g2_decap_4 FILLER_32_571 ();
 sg13g2_fill_2 FILLER_32_575 ();
 sg13g2_decap_8 FILLER_32_607 ();
 sg13g2_fill_1 FILLER_32_614 ();
 sg13g2_fill_1 FILLER_32_637 ();
 sg13g2_fill_1 FILLER_32_647 ();
 sg13g2_decap_4 FILLER_32_656 ();
 sg13g2_fill_2 FILLER_32_664 ();
 sg13g2_fill_1 FILLER_32_666 ();
 sg13g2_decap_8 FILLER_32_697 ();
 sg13g2_decap_4 FILLER_32_704 ();
 sg13g2_fill_1 FILLER_32_708 ();
 sg13g2_fill_2 FILLER_32_717 ();
 sg13g2_fill_2 FILLER_32_726 ();
 sg13g2_decap_8 FILLER_32_755 ();
 sg13g2_fill_2 FILLER_32_776 ();
 sg13g2_decap_4 FILLER_32_783 ();
 sg13g2_fill_2 FILLER_32_787 ();
 sg13g2_fill_1 FILLER_32_813 ();
 sg13g2_fill_1 FILLER_32_836 ();
 sg13g2_decap_4 FILLER_32_863 ();
 sg13g2_fill_1 FILLER_32_867 ();
 sg13g2_fill_1 FILLER_32_884 ();
 sg13g2_fill_2 FILLER_32_894 ();
 sg13g2_fill_1 FILLER_32_896 ();
 sg13g2_decap_8 FILLER_32_902 ();
 sg13g2_fill_1 FILLER_32_927 ();
 sg13g2_fill_1 FILLER_32_932 ();
 sg13g2_decap_4 FILLER_32_938 ();
 sg13g2_fill_2 FILLER_32_951 ();
 sg13g2_decap_4 FILLER_32_982 ();
 sg13g2_fill_2 FILLER_32_1007 ();
 sg13g2_fill_1 FILLER_32_1009 ();
 sg13g2_fill_2 FILLER_32_1025 ();
 sg13g2_fill_1 FILLER_32_1027 ();
 sg13g2_fill_2 FILLER_32_1090 ();
 sg13g2_fill_1 FILLER_32_1092 ();
 sg13g2_decap_4 FILLER_32_1121 ();
 sg13g2_fill_1 FILLER_32_1134 ();
 sg13g2_fill_1 FILLER_32_1167 ();
 sg13g2_fill_1 FILLER_32_1173 ();
 sg13g2_decap_4 FILLER_32_1183 ();
 sg13g2_fill_2 FILLER_32_1187 ();
 sg13g2_fill_2 FILLER_32_1196 ();
 sg13g2_decap_8 FILLER_32_1226 ();
 sg13g2_decap_8 FILLER_32_1233 ();
 sg13g2_fill_2 FILLER_32_1245 ();
 sg13g2_decap_4 FILLER_32_1256 ();
 sg13g2_fill_2 FILLER_32_1277 ();
 sg13g2_decap_4 FILLER_32_1301 ();
 sg13g2_fill_1 FILLER_32_1305 ();
 sg13g2_fill_2 FILLER_32_1319 ();
 sg13g2_fill_1 FILLER_32_1335 ();
 sg13g2_decap_4 FILLER_32_1341 ();
 sg13g2_decap_4 FILLER_32_1350 ();
 sg13g2_fill_2 FILLER_32_1354 ();
 sg13g2_fill_2 FILLER_32_1364 ();
 sg13g2_fill_1 FILLER_32_1366 ();
 sg13g2_fill_2 FILLER_32_1400 ();
 sg13g2_fill_1 FILLER_32_1402 ();
 sg13g2_decap_4 FILLER_32_1407 ();
 sg13g2_decap_8 FILLER_32_1419 ();
 sg13g2_decap_8 FILLER_32_1443 ();
 sg13g2_decap_8 FILLER_32_1450 ();
 sg13g2_decap_4 FILLER_32_1457 ();
 sg13g2_fill_2 FILLER_32_1461 ();
 sg13g2_decap_4 FILLER_32_1500 ();
 sg13g2_decap_4 FILLER_32_1513 ();
 sg13g2_decap_4 FILLER_32_1525 ();
 sg13g2_decap_8 FILLER_32_1534 ();
 sg13g2_fill_2 FILLER_32_1544 ();
 sg13g2_fill_2 FILLER_32_1550 ();
 sg13g2_fill_1 FILLER_32_1552 ();
 sg13g2_fill_1 FILLER_32_1564 ();
 sg13g2_decap_8 FILLER_32_1587 ();
 sg13g2_fill_1 FILLER_32_1594 ();
 sg13g2_decap_4 FILLER_32_1600 ();
 sg13g2_fill_2 FILLER_32_1604 ();
 sg13g2_decap_4 FILLER_32_1614 ();
 sg13g2_fill_2 FILLER_32_1628 ();
 sg13g2_fill_1 FILLER_32_1630 ();
 sg13g2_fill_1 FILLER_32_1640 ();
 sg13g2_fill_1 FILLER_32_1658 ();
 sg13g2_fill_2 FILLER_32_1672 ();
 sg13g2_fill_1 FILLER_32_1674 ();
 sg13g2_fill_2 FILLER_32_1682 ();
 sg13g2_decap_8 FILLER_32_1692 ();
 sg13g2_decap_8 FILLER_32_1699 ();
 sg13g2_fill_2 FILLER_32_1706 ();
 sg13g2_fill_1 FILLER_32_1708 ();
 sg13g2_decap_4 FILLER_32_1728 ();
 sg13g2_fill_1 FILLER_32_1759 ();
 sg13g2_decap_4 FILLER_32_1767 ();
 sg13g2_decap_8 FILLER_32_1778 ();
 sg13g2_decap_8 FILLER_32_1785 ();
 sg13g2_fill_2 FILLER_32_1792 ();
 sg13g2_fill_1 FILLER_32_1794 ();
 sg13g2_decap_8 FILLER_32_1809 ();
 sg13g2_decap_8 FILLER_32_1829 ();
 sg13g2_fill_1 FILLER_32_1836 ();
 sg13g2_decap_8 FILLER_32_1859 ();
 sg13g2_fill_2 FILLER_32_1866 ();
 sg13g2_decap_8 FILLER_32_1881 ();
 sg13g2_fill_2 FILLER_32_1888 ();
 sg13g2_decap_4 FILLER_32_1894 ();
 sg13g2_decap_4 FILLER_32_1926 ();
 sg13g2_fill_2 FILLER_32_1930 ();
 sg13g2_fill_2 FILLER_32_1960 ();
 sg13g2_fill_1 FILLER_32_1962 ();
 sg13g2_fill_2 FILLER_32_1972 ();
 sg13g2_decap_4 FILLER_32_1979 ();
 sg13g2_fill_2 FILLER_32_2008 ();
 sg13g2_fill_1 FILLER_32_2020 ();
 sg13g2_fill_2 FILLER_32_2025 ();
 sg13g2_fill_2 FILLER_32_2032 ();
 sg13g2_fill_1 FILLER_32_2034 ();
 sg13g2_fill_1 FILLER_32_2042 ();
 sg13g2_fill_2 FILLER_32_2055 ();
 sg13g2_fill_1 FILLER_32_2080 ();
 sg13g2_decap_8 FILLER_32_2101 ();
 sg13g2_decap_8 FILLER_32_2108 ();
 sg13g2_fill_1 FILLER_32_2115 ();
 sg13g2_fill_2 FILLER_32_2124 ();
 sg13g2_fill_1 FILLER_32_2126 ();
 sg13g2_fill_2 FILLER_32_2154 ();
 sg13g2_decap_8 FILLER_32_2164 ();
 sg13g2_decap_4 FILLER_32_2171 ();
 sg13g2_fill_2 FILLER_32_2183 ();
 sg13g2_decap_4 FILLER_32_2214 ();
 sg13g2_fill_1 FILLER_32_2231 ();
 sg13g2_fill_1 FILLER_32_2236 ();
 sg13g2_decap_4 FILLER_32_2242 ();
 sg13g2_fill_2 FILLER_32_2254 ();
 sg13g2_fill_1 FILLER_32_2256 ();
 sg13g2_decap_8 FILLER_32_2274 ();
 sg13g2_decap_8 FILLER_32_2281 ();
 sg13g2_fill_2 FILLER_32_2304 ();
 sg13g2_decap_8 FILLER_32_2310 ();
 sg13g2_decap_8 FILLER_32_2317 ();
 sg13g2_fill_2 FILLER_32_2324 ();
 sg13g2_fill_1 FILLER_32_2326 ();
 sg13g2_decap_8 FILLER_32_2337 ();
 sg13g2_decap_8 FILLER_32_2344 ();
 sg13g2_fill_2 FILLER_32_2351 ();
 sg13g2_fill_1 FILLER_32_2353 ();
 sg13g2_decap_4 FILLER_32_2374 ();
 sg13g2_fill_1 FILLER_32_2378 ();
 sg13g2_decap_4 FILLER_32_2393 ();
 sg13g2_decap_4 FILLER_32_2402 ();
 sg13g2_decap_8 FILLER_32_2414 ();
 sg13g2_decap_8 FILLER_32_2421 ();
 sg13g2_decap_8 FILLER_32_2443 ();
 sg13g2_decap_4 FILLER_32_2450 ();
 sg13g2_fill_1 FILLER_32_2454 ();
 sg13g2_fill_2 FILLER_32_2468 ();
 sg13g2_fill_1 FILLER_32_2470 ();
 sg13g2_fill_2 FILLER_32_2475 ();
 sg13g2_fill_1 FILLER_32_2477 ();
 sg13g2_decap_4 FILLER_32_2495 ();
 sg13g2_fill_2 FILLER_32_2499 ();
 sg13g2_decap_4 FILLER_32_2504 ();
 sg13g2_decap_4 FILLER_32_2540 ();
 sg13g2_fill_2 FILLER_32_2544 ();
 sg13g2_fill_2 FILLER_32_2551 ();
 sg13g2_decap_4 FILLER_32_2569 ();
 sg13g2_fill_2 FILLER_32_2573 ();
 sg13g2_decap_8 FILLER_32_2588 ();
 sg13g2_decap_8 FILLER_32_2595 ();
 sg13g2_fill_1 FILLER_32_2602 ();
 sg13g2_fill_1 FILLER_32_2619 ();
 sg13g2_decap_8 FILLER_32_2634 ();
 sg13g2_decap_8 FILLER_32_2641 ();
 sg13g2_decap_4 FILLER_32_2652 ();
 sg13g2_decap_8 FILLER_32_2689 ();
 sg13g2_fill_1 FILLER_32_2696 ();
 sg13g2_decap_4 FILLER_32_2709 ();
 sg13g2_decap_8 FILLER_32_2734 ();
 sg13g2_fill_2 FILLER_32_2749 ();
 sg13g2_fill_1 FILLER_32_2751 ();
 sg13g2_fill_1 FILLER_32_2771 ();
 sg13g2_decap_8 FILLER_32_2775 ();
 sg13g2_decap_4 FILLER_32_2790 ();
 sg13g2_fill_1 FILLER_32_2794 ();
 sg13g2_decap_8 FILLER_32_2821 ();
 sg13g2_fill_1 FILLER_32_2841 ();
 sg13g2_fill_2 FILLER_32_2859 ();
 sg13g2_fill_1 FILLER_32_2871 ();
 sg13g2_decap_8 FILLER_32_2877 ();
 sg13g2_fill_2 FILLER_32_2884 ();
 sg13g2_fill_2 FILLER_32_2891 ();
 sg13g2_fill_1 FILLER_32_2893 ();
 sg13g2_fill_2 FILLER_32_2897 ();
 sg13g2_decap_8 FILLER_32_2926 ();
 sg13g2_decap_4 FILLER_32_2933 ();
 sg13g2_fill_2 FILLER_32_2937 ();
 sg13g2_fill_1 FILLER_32_2959 ();
 sg13g2_decap_8 FILLER_32_2978 ();
 sg13g2_fill_1 FILLER_32_2997 ();
 sg13g2_fill_1 FILLER_32_3006 ();
 sg13g2_fill_2 FILLER_32_3022 ();
 sg13g2_fill_1 FILLER_32_3024 ();
 sg13g2_fill_1 FILLER_32_3030 ();
 sg13g2_decap_8 FILLER_32_3041 ();
 sg13g2_decap_8 FILLER_32_3053 ();
 sg13g2_fill_2 FILLER_32_3060 ();
 sg13g2_fill_1 FILLER_32_3062 ();
 sg13g2_fill_2 FILLER_32_3071 ();
 sg13g2_fill_1 FILLER_32_3073 ();
 sg13g2_fill_2 FILLER_32_3108 ();
 sg13g2_fill_1 FILLER_32_3139 ();
 sg13g2_fill_2 FILLER_32_3166 ();
 sg13g2_fill_1 FILLER_32_3168 ();
 sg13g2_fill_2 FILLER_32_3188 ();
 sg13g2_fill_1 FILLER_32_3194 ();
 sg13g2_fill_2 FILLER_32_3210 ();
 sg13g2_fill_1 FILLER_32_3212 ();
 sg13g2_decap_4 FILLER_32_3230 ();
 sg13g2_fill_1 FILLER_32_3241 ();
 sg13g2_fill_2 FILLER_32_3257 ();
 sg13g2_fill_1 FILLER_32_3259 ();
 sg13g2_fill_1 FILLER_32_3265 ();
 sg13g2_decap_8 FILLER_32_3306 ();
 sg13g2_decap_4 FILLER_32_3313 ();
 sg13g2_fill_1 FILLER_32_3317 ();
 sg13g2_decap_4 FILLER_32_3323 ();
 sg13g2_fill_1 FILLER_32_3327 ();
 sg13g2_decap_8 FILLER_32_3336 ();
 sg13g2_decap_8 FILLER_32_3343 ();
 sg13g2_fill_2 FILLER_32_3360 ();
 sg13g2_fill_1 FILLER_32_3362 ();
 sg13g2_fill_2 FILLER_32_3366 ();
 sg13g2_fill_1 FILLER_32_3372 ();
 sg13g2_decap_4 FILLER_32_3378 ();
 sg13g2_fill_1 FILLER_32_3382 ();
 sg13g2_decap_8 FILLER_32_3403 ();
 sg13g2_decap_8 FILLER_32_3410 ();
 sg13g2_decap_4 FILLER_32_3442 ();
 sg13g2_fill_1 FILLER_32_3446 ();
 sg13g2_decap_8 FILLER_32_3452 ();
 sg13g2_decap_4 FILLER_32_3459 ();
 sg13g2_decap_8 FILLER_32_3479 ();
 sg13g2_decap_8 FILLER_32_3486 ();
 sg13g2_decap_8 FILLER_32_3493 ();
 sg13g2_decap_8 FILLER_32_3500 ();
 sg13g2_decap_8 FILLER_32_3507 ();
 sg13g2_decap_8 FILLER_32_3514 ();
 sg13g2_decap_8 FILLER_32_3521 ();
 sg13g2_decap_8 FILLER_32_3528 ();
 sg13g2_decap_8 FILLER_32_3535 ();
 sg13g2_decap_8 FILLER_32_3542 ();
 sg13g2_decap_8 FILLER_32_3549 ();
 sg13g2_decap_8 FILLER_32_3556 ();
 sg13g2_decap_8 FILLER_32_3563 ();
 sg13g2_decap_8 FILLER_32_3570 ();
 sg13g2_fill_2 FILLER_32_3577 ();
 sg13g2_fill_1 FILLER_32_3579 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_117 ();
 sg13g2_decap_8 FILLER_33_124 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_163 ();
 sg13g2_fill_1 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_206 ();
 sg13g2_fill_1 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_decap_4 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_308 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_328 ();
 sg13g2_decap_8 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_fill_1 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_405 ();
 sg13g2_fill_1 FILLER_33_412 ();
 sg13g2_fill_2 FILLER_33_426 ();
 sg13g2_fill_1 FILLER_33_428 ();
 sg13g2_decap_8 FILLER_33_470 ();
 sg13g2_fill_2 FILLER_33_477 ();
 sg13g2_fill_2 FILLER_33_482 ();
 sg13g2_fill_1 FILLER_33_484 ();
 sg13g2_fill_2 FILLER_33_489 ();
 sg13g2_fill_1 FILLER_33_491 ();
 sg13g2_decap_8 FILLER_33_496 ();
 sg13g2_decap_8 FILLER_33_503 ();
 sg13g2_decap_4 FILLER_33_510 ();
 sg13g2_fill_1 FILLER_33_514 ();
 sg13g2_decap_4 FILLER_33_525 ();
 sg13g2_fill_1 FILLER_33_529 ();
 sg13g2_decap_8 FILLER_33_558 ();
 sg13g2_decap_8 FILLER_33_565 ();
 sg13g2_decap_8 FILLER_33_572 ();
 sg13g2_decap_4 FILLER_33_579 ();
 sg13g2_fill_2 FILLER_33_583 ();
 sg13g2_fill_2 FILLER_33_590 ();
 sg13g2_fill_1 FILLER_33_592 ();
 sg13g2_fill_1 FILLER_33_621 ();
 sg13g2_fill_1 FILLER_33_634 ();
 sg13g2_fill_1 FILLER_33_643 ();
 sg13g2_decap_8 FILLER_33_650 ();
 sg13g2_decap_8 FILLER_33_657 ();
 sg13g2_decap_4 FILLER_33_664 ();
 sg13g2_fill_1 FILLER_33_668 ();
 sg13g2_fill_1 FILLER_33_682 ();
 sg13g2_fill_1 FILLER_33_716 ();
 sg13g2_fill_2 FILLER_33_721 ();
 sg13g2_fill_1 FILLER_33_731 ();
 sg13g2_decap_4 FILLER_33_736 ();
 sg13g2_fill_1 FILLER_33_756 ();
 sg13g2_decap_4 FILLER_33_765 ();
 sg13g2_fill_2 FILLER_33_769 ();
 sg13g2_fill_2 FILLER_33_785 ();
 sg13g2_fill_1 FILLER_33_787 ();
 sg13g2_fill_2 FILLER_33_796 ();
 sg13g2_fill_2 FILLER_33_824 ();
 sg13g2_fill_2 FILLER_33_841 ();
 sg13g2_fill_1 FILLER_33_843 ();
 sg13g2_fill_2 FILLER_33_871 ();
 sg13g2_fill_1 FILLER_33_873 ();
 sg13g2_fill_2 FILLER_33_882 ();
 sg13g2_decap_8 FILLER_33_897 ();
 sg13g2_decap_8 FILLER_33_904 ();
 sg13g2_fill_1 FILLER_33_911 ();
 sg13g2_fill_2 FILLER_33_938 ();
 sg13g2_fill_2 FILLER_33_950 ();
 sg13g2_fill_1 FILLER_33_952 ();
 sg13g2_decap_8 FILLER_33_958 ();
 sg13g2_decap_4 FILLER_33_980 ();
 sg13g2_fill_2 FILLER_33_1001 ();
 sg13g2_fill_2 FILLER_33_1012 ();
 sg13g2_fill_1 FILLER_33_1014 ();
 sg13g2_decap_8 FILLER_33_1023 ();
 sg13g2_fill_2 FILLER_33_1030 ();
 sg13g2_fill_1 FILLER_33_1032 ();
 sg13g2_decap_4 FILLER_33_1036 ();
 sg13g2_decap_8 FILLER_33_1058 ();
 sg13g2_fill_1 FILLER_33_1065 ();
 sg13g2_decap_8 FILLER_33_1082 ();
 sg13g2_decap_4 FILLER_33_1089 ();
 sg13g2_fill_2 FILLER_33_1132 ();
 sg13g2_fill_2 FILLER_33_1139 ();
 sg13g2_fill_1 FILLER_33_1154 ();
 sg13g2_fill_2 FILLER_33_1164 ();
 sg13g2_fill_2 FILLER_33_1171 ();
 sg13g2_decap_8 FILLER_33_1177 ();
 sg13g2_fill_1 FILLER_33_1184 ();
 sg13g2_fill_2 FILLER_33_1221 ();
 sg13g2_fill_2 FILLER_33_1228 ();
 sg13g2_fill_1 FILLER_33_1230 ();
 sg13g2_fill_1 FILLER_33_1251 ();
 sg13g2_decap_8 FILLER_33_1274 ();
 sg13g2_fill_2 FILLER_33_1285 ();
 sg13g2_fill_1 FILLER_33_1287 ();
 sg13g2_fill_2 FILLER_33_1304 ();
 sg13g2_fill_1 FILLER_33_1306 ();
 sg13g2_fill_2 FILLER_33_1315 ();
 sg13g2_decap_8 FILLER_33_1322 ();
 sg13g2_decap_8 FILLER_33_1329 ();
 sg13g2_decap_4 FILLER_33_1336 ();
 sg13g2_fill_1 FILLER_33_1340 ();
 sg13g2_decap_8 FILLER_33_1358 ();
 sg13g2_decap_8 FILLER_33_1365 ();
 sg13g2_decap_8 FILLER_33_1372 ();
 sg13g2_decap_4 FILLER_33_1379 ();
 sg13g2_fill_2 FILLER_33_1389 ();
 sg13g2_fill_2 FILLER_33_1403 ();
 sg13g2_fill_1 FILLER_33_1405 ();
 sg13g2_fill_1 FILLER_33_1422 ();
 sg13g2_fill_2 FILLER_33_1428 ();
 sg13g2_fill_1 FILLER_33_1430 ();
 sg13g2_decap_8 FILLER_33_1444 ();
 sg13g2_fill_2 FILLER_33_1451 ();
 sg13g2_decap_8 FILLER_33_1483 ();
 sg13g2_fill_2 FILLER_33_1490 ();
 sg13g2_fill_1 FILLER_33_1492 ();
 sg13g2_decap_8 FILLER_33_1515 ();
 sg13g2_decap_4 FILLER_33_1522 ();
 sg13g2_decap_4 FILLER_33_1530 ();
 sg13g2_fill_1 FILLER_33_1534 ();
 sg13g2_fill_1 FILLER_33_1545 ();
 sg13g2_decap_4 FILLER_33_1554 ();
 sg13g2_fill_1 FILLER_33_1558 ();
 sg13g2_fill_1 FILLER_33_1564 ();
 sg13g2_decap_4 FILLER_33_1569 ();
 sg13g2_decap_8 FILLER_33_1581 ();
 sg13g2_fill_2 FILLER_33_1588 ();
 sg13g2_fill_2 FILLER_33_1624 ();
 sg13g2_decap_8 FILLER_33_1630 ();
 sg13g2_decap_8 FILLER_33_1637 ();
 sg13g2_fill_2 FILLER_33_1644 ();
 sg13g2_fill_1 FILLER_33_1646 ();
 sg13g2_decap_8 FILLER_33_1660 ();
 sg13g2_decap_4 FILLER_33_1667 ();
 sg13g2_fill_1 FILLER_33_1671 ();
 sg13g2_decap_8 FILLER_33_1693 ();
 sg13g2_decap_8 FILLER_33_1700 ();
 sg13g2_decap_4 FILLER_33_1707 ();
 sg13g2_fill_1 FILLER_33_1711 ();
 sg13g2_decap_8 FILLER_33_1734 ();
 sg13g2_fill_1 FILLER_33_1741 ();
 sg13g2_decap_4 FILLER_33_1778 ();
 sg13g2_decap_8 FILLER_33_1808 ();
 sg13g2_decap_8 FILLER_33_1829 ();
 sg13g2_fill_2 FILLER_33_1836 ();
 sg13g2_decap_8 FILLER_33_1856 ();
 sg13g2_fill_1 FILLER_33_1863 ();
 sg13g2_decap_4 FILLER_33_1886 ();
 sg13g2_fill_1 FILLER_33_1890 ();
 sg13g2_decap_8 FILLER_33_1917 ();
 sg13g2_fill_2 FILLER_33_1924 ();
 sg13g2_fill_1 FILLER_33_1926 ();
 sg13g2_fill_2 FILLER_33_1953 ();
 sg13g2_fill_1 FILLER_33_1983 ();
 sg13g2_fill_1 FILLER_33_2003 ();
 sg13g2_decap_8 FILLER_33_2017 ();
 sg13g2_decap_8 FILLER_33_2024 ();
 sg13g2_decap_8 FILLER_33_2031 ();
 sg13g2_fill_2 FILLER_33_2038 ();
 sg13g2_fill_2 FILLER_33_2057 ();
 sg13g2_fill_1 FILLER_33_2059 ();
 sg13g2_decap_4 FILLER_33_2078 ();
 sg13g2_fill_2 FILLER_33_2082 ();
 sg13g2_decap_4 FILLER_33_2087 ();
 sg13g2_decap_8 FILLER_33_2099 ();
 sg13g2_fill_2 FILLER_33_2106 ();
 sg13g2_fill_1 FILLER_33_2108 ();
 sg13g2_fill_2 FILLER_33_2144 ();
 sg13g2_fill_1 FILLER_33_2146 ();
 sg13g2_decap_8 FILLER_33_2155 ();
 sg13g2_fill_2 FILLER_33_2162 ();
 sg13g2_fill_1 FILLER_33_2164 ();
 sg13g2_decap_8 FILLER_33_2168 ();
 sg13g2_decap_4 FILLER_33_2175 ();
 sg13g2_fill_2 FILLER_33_2187 ();
 sg13g2_decap_4 FILLER_33_2194 ();
 sg13g2_fill_2 FILLER_33_2198 ();
 sg13g2_fill_2 FILLER_33_2211 ();
 sg13g2_decap_8 FILLER_33_2236 ();
 sg13g2_decap_8 FILLER_33_2243 ();
 sg13g2_fill_2 FILLER_33_2250 ();
 sg13g2_fill_1 FILLER_33_2252 ();
 sg13g2_decap_8 FILLER_33_2275 ();
 sg13g2_decap_8 FILLER_33_2282 ();
 sg13g2_fill_1 FILLER_33_2289 ();
 sg13g2_fill_1 FILLER_33_2322 ();
 sg13g2_fill_2 FILLER_33_2346 ();
 sg13g2_decap_8 FILLER_33_2375 ();
 sg13g2_fill_1 FILLER_33_2382 ();
 sg13g2_fill_2 FILLER_33_2393 ();
 sg13g2_fill_1 FILLER_33_2395 ();
 sg13g2_fill_2 FILLER_33_2413 ();
 sg13g2_fill_1 FILLER_33_2419 ();
 sg13g2_fill_1 FILLER_33_2430 ();
 sg13g2_decap_8 FILLER_33_2449 ();
 sg13g2_decap_4 FILLER_33_2456 ();
 sg13g2_decap_8 FILLER_33_2468 ();
 sg13g2_decap_8 FILLER_33_2475 ();
 sg13g2_fill_2 FILLER_33_2482 ();
 sg13g2_fill_1 FILLER_33_2484 ();
 sg13g2_decap_8 FILLER_33_2511 ();
 sg13g2_decap_8 FILLER_33_2518 ();
 sg13g2_fill_2 FILLER_33_2528 ();
 sg13g2_fill_2 FILLER_33_2538 ();
 sg13g2_fill_1 FILLER_33_2553 ();
 sg13g2_fill_2 FILLER_33_2579 ();
 sg13g2_fill_2 FILLER_33_2594 ();
 sg13g2_decap_4 FILLER_33_2619 ();
 sg13g2_decap_8 FILLER_33_2640 ();
 sg13g2_fill_2 FILLER_33_2647 ();
 sg13g2_fill_1 FILLER_33_2649 ();
 sg13g2_fill_1 FILLER_33_2668 ();
 sg13g2_fill_1 FILLER_33_2673 ();
 sg13g2_decap_4 FILLER_33_2687 ();
 sg13g2_fill_1 FILLER_33_2691 ();
 sg13g2_decap_8 FILLER_33_2730 ();
 sg13g2_fill_2 FILLER_33_2737 ();
 sg13g2_fill_1 FILLER_33_2739 ();
 sg13g2_decap_4 FILLER_33_2744 ();
 sg13g2_fill_1 FILLER_33_2761 ();
 sg13g2_fill_2 FILLER_33_2766 ();
 sg13g2_decap_8 FILLER_33_2810 ();
 sg13g2_decap_8 FILLER_33_2817 ();
 sg13g2_fill_1 FILLER_33_2836 ();
 sg13g2_fill_1 FILLER_33_2849 ();
 sg13g2_decap_8 FILLER_33_2860 ();
 sg13g2_fill_1 FILLER_33_2867 ();
 sg13g2_decap_8 FILLER_33_2872 ();
 sg13g2_fill_2 FILLER_33_2879 ();
 sg13g2_fill_2 FILLER_33_2886 ();
 sg13g2_fill_1 FILLER_33_2888 ();
 sg13g2_decap_4 FILLER_33_2907 ();
 sg13g2_fill_1 FILLER_33_2911 ();
 sg13g2_decap_8 FILLER_33_2938 ();
 sg13g2_fill_2 FILLER_33_2945 ();
 sg13g2_fill_1 FILLER_33_2947 ();
 sg13g2_decap_8 FILLER_33_2953 ();
 sg13g2_decap_4 FILLER_33_2960 ();
 sg13g2_fill_1 FILLER_33_2964 ();
 sg13g2_fill_1 FILLER_33_2982 ();
 sg13g2_fill_2 FILLER_33_3014 ();
 sg13g2_fill_2 FILLER_33_3023 ();
 sg13g2_fill_2 FILLER_33_3030 ();
 sg13g2_fill_1 FILLER_33_3032 ();
 sg13g2_fill_1 FILLER_33_3052 ();
 sg13g2_decap_8 FILLER_33_3063 ();
 sg13g2_fill_2 FILLER_33_3078 ();
 sg13g2_fill_1 FILLER_33_3080 ();
 sg13g2_decap_8 FILLER_33_3086 ();
 sg13g2_fill_2 FILLER_33_3102 ();
 sg13g2_fill_1 FILLER_33_3104 ();
 sg13g2_fill_2 FILLER_33_3140 ();
 sg13g2_fill_1 FILLER_33_3142 ();
 sg13g2_fill_2 FILLER_33_3160 ();
 sg13g2_decap_8 FILLER_33_3184 ();
 sg13g2_decap_4 FILLER_33_3191 ();
 sg13g2_decap_4 FILLER_33_3228 ();
 sg13g2_decap_4 FILLER_33_3236 ();
 sg13g2_fill_2 FILLER_33_3240 ();
 sg13g2_decap_8 FILLER_33_3251 ();
 sg13g2_fill_2 FILLER_33_3258 ();
 sg13g2_fill_1 FILLER_33_3260 ();
 sg13g2_fill_1 FILLER_33_3265 ();
 sg13g2_fill_2 FILLER_33_3275 ();
 sg13g2_fill_1 FILLER_33_3277 ();
 sg13g2_fill_1 FILLER_33_3281 ();
 sg13g2_decap_8 FILLER_33_3304 ();
 sg13g2_decap_4 FILLER_33_3311 ();
 sg13g2_decap_8 FILLER_33_3321 ();
 sg13g2_fill_2 FILLER_33_3328 ();
 sg13g2_decap_8 FILLER_33_3334 ();
 sg13g2_fill_2 FILLER_33_3341 ();
 sg13g2_fill_1 FILLER_33_3343 ();
 sg13g2_fill_2 FILLER_33_3381 ();
 sg13g2_fill_1 FILLER_33_3383 ();
 sg13g2_decap_4 FILLER_33_3400 ();
 sg13g2_fill_1 FILLER_33_3416 ();
 sg13g2_fill_2 FILLER_33_3486 ();
 sg13g2_fill_1 FILLER_33_3488 ();
 sg13g2_decap_8 FILLER_33_3502 ();
 sg13g2_decap_8 FILLER_33_3509 ();
 sg13g2_decap_8 FILLER_33_3516 ();
 sg13g2_decap_8 FILLER_33_3523 ();
 sg13g2_decap_8 FILLER_33_3530 ();
 sg13g2_decap_8 FILLER_33_3537 ();
 sg13g2_decap_8 FILLER_33_3544 ();
 sg13g2_decap_8 FILLER_33_3551 ();
 sg13g2_decap_8 FILLER_33_3558 ();
 sg13g2_decap_8 FILLER_33_3565 ();
 sg13g2_decap_8 FILLER_33_3572 ();
 sg13g2_fill_1 FILLER_33_3579 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_4 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_81 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_decap_8 FILLER_34_115 ();
 sg13g2_decap_8 FILLER_34_122 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_171 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_decap_4 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_264 ();
 sg13g2_decap_4 FILLER_34_292 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_378 ();
 sg13g2_decap_4 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_409 ();
 sg13g2_fill_2 FILLER_34_439 ();
 sg13g2_decap_8 FILLER_34_445 ();
 sg13g2_fill_1 FILLER_34_457 ();
 sg13g2_decap_4 FILLER_34_466 ();
 sg13g2_fill_2 FILLER_34_470 ();
 sg13g2_fill_2 FILLER_34_528 ();
 sg13g2_fill_1 FILLER_34_530 ();
 sg13g2_decap_8 FILLER_34_548 ();
 sg13g2_fill_2 FILLER_34_555 ();
 sg13g2_decap_8 FILLER_34_570 ();
 sg13g2_fill_2 FILLER_34_577 ();
 sg13g2_fill_1 FILLER_34_579 ();
 sg13g2_fill_2 FILLER_34_620 ();
 sg13g2_fill_2 FILLER_34_639 ();
 sg13g2_fill_1 FILLER_34_641 ();
 sg13g2_decap_8 FILLER_34_646 ();
 sg13g2_decap_8 FILLER_34_653 ();
 sg13g2_decap_4 FILLER_34_665 ();
 sg13g2_fill_2 FILLER_34_669 ();
 sg13g2_decap_8 FILLER_34_706 ();
 sg13g2_decap_8 FILLER_34_730 ();
 sg13g2_fill_1 FILLER_34_737 ();
 sg13g2_decap_8 FILLER_34_774 ();
 sg13g2_decap_8 FILLER_34_781 ();
 sg13g2_decap_4 FILLER_34_788 ();
 sg13g2_fill_2 FILLER_34_792 ();
 sg13g2_fill_2 FILLER_34_808 ();
 sg13g2_fill_1 FILLER_34_810 ();
 sg13g2_decap_8 FILLER_34_830 ();
 sg13g2_fill_2 FILLER_34_837 ();
 sg13g2_fill_1 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_866 ();
 sg13g2_decap_8 FILLER_34_873 ();
 sg13g2_decap_4 FILLER_34_880 ();
 sg13g2_fill_2 FILLER_34_917 ();
 sg13g2_decap_8 FILLER_34_923 ();
 sg13g2_decap_8 FILLER_34_930 ();
 sg13g2_decap_8 FILLER_34_937 ();
 sg13g2_decap_4 FILLER_34_944 ();
 sg13g2_fill_2 FILLER_34_964 ();
 sg13g2_fill_1 FILLER_34_970 ();
 sg13g2_decap_8 FILLER_34_976 ();
 sg13g2_decap_4 FILLER_34_983 ();
 sg13g2_fill_1 FILLER_34_1008 ();
 sg13g2_fill_1 FILLER_34_1035 ();
 sg13g2_decap_8 FILLER_34_1055 ();
 sg13g2_fill_2 FILLER_34_1062 ();
 sg13g2_fill_1 FILLER_34_1064 ();
 sg13g2_decap_4 FILLER_34_1082 ();
 sg13g2_fill_2 FILLER_34_1119 ();
 sg13g2_fill_2 FILLER_34_1138 ();
 sg13g2_fill_1 FILLER_34_1153 ();
 sg13g2_fill_1 FILLER_34_1167 ();
 sg13g2_decap_4 FILLER_34_1176 ();
 sg13g2_fill_1 FILLER_34_1180 ();
 sg13g2_decap_8 FILLER_34_1199 ();
 sg13g2_fill_2 FILLER_34_1206 ();
 sg13g2_fill_2 FILLER_34_1216 ();
 sg13g2_decap_8 FILLER_34_1226 ();
 sg13g2_decap_4 FILLER_34_1233 ();
 sg13g2_decap_8 FILLER_34_1266 ();
 sg13g2_decap_8 FILLER_34_1273 ();
 sg13g2_decap_4 FILLER_34_1285 ();
 sg13g2_fill_1 FILLER_34_1289 ();
 sg13g2_fill_1 FILLER_34_1299 ();
 sg13g2_decap_8 FILLER_34_1322 ();
 sg13g2_decap_8 FILLER_34_1329 ();
 sg13g2_fill_2 FILLER_34_1336 ();
 sg13g2_fill_2 FILLER_34_1347 ();
 sg13g2_decap_8 FILLER_34_1361 ();
 sg13g2_decap_8 FILLER_34_1409 ();
 sg13g2_decap_8 FILLER_34_1416 ();
 sg13g2_fill_2 FILLER_34_1423 ();
 sg13g2_fill_1 FILLER_34_1425 ();
 sg13g2_decap_4 FILLER_34_1459 ();
 sg13g2_fill_2 FILLER_34_1463 ();
 sg13g2_decap_8 FILLER_34_1483 ();
 sg13g2_fill_1 FILLER_34_1490 ();
 sg13g2_fill_1 FILLER_34_1519 ();
 sg13g2_fill_2 FILLER_34_1538 ();
 sg13g2_fill_1 FILLER_34_1540 ();
 sg13g2_decap_8 FILLER_34_1545 ();
 sg13g2_fill_2 FILLER_34_1552 ();
 sg13g2_fill_1 FILLER_34_1554 ();
 sg13g2_decap_4 FILLER_34_1562 ();
 sg13g2_decap_8 FILLER_34_1570 ();
 sg13g2_decap_8 FILLER_34_1577 ();
 sg13g2_fill_1 FILLER_34_1616 ();
 sg13g2_decap_8 FILLER_34_1634 ();
 sg13g2_fill_1 FILLER_34_1641 ();
 sg13g2_decap_8 FILLER_34_1651 ();
 sg13g2_fill_2 FILLER_34_1658 ();
 sg13g2_fill_1 FILLER_34_1660 ();
 sg13g2_decap_4 FILLER_34_1665 ();
 sg13g2_fill_1 FILLER_34_1669 ();
 sg13g2_decap_4 FILLER_34_1674 ();
 sg13g2_fill_2 FILLER_34_1691 ();
 sg13g2_fill_1 FILLER_34_1693 ();
 sg13g2_fill_1 FILLER_34_1719 ();
 sg13g2_fill_1 FILLER_34_1728 ();
 sg13g2_decap_4 FILLER_34_1737 ();
 sg13g2_fill_1 FILLER_34_1741 ();
 sg13g2_decap_8 FILLER_34_1750 ();
 sg13g2_fill_2 FILLER_34_1757 ();
 sg13g2_fill_2 FILLER_34_1782 ();
 sg13g2_decap_8 FILLER_34_1801 ();
 sg13g2_fill_1 FILLER_34_1808 ();
 sg13g2_fill_2 FILLER_34_1833 ();
 sg13g2_decap_8 FILLER_34_1840 ();
 sg13g2_decap_8 FILLER_34_1847 ();
 sg13g2_decap_8 FILLER_34_1854 ();
 sg13g2_fill_1 FILLER_34_1861 ();
 sg13g2_decap_4 FILLER_34_1884 ();
 sg13g2_fill_1 FILLER_34_1900 ();
 sg13g2_fill_2 FILLER_34_1927 ();
 sg13g2_fill_2 FILLER_34_1946 ();
 sg13g2_fill_1 FILLER_34_1948 ();
 sg13g2_decap_8 FILLER_34_1975 ();
 sg13g2_fill_2 FILLER_34_1982 ();
 sg13g2_fill_1 FILLER_34_1984 ();
 sg13g2_decap_4 FILLER_34_1988 ();
 sg13g2_fill_2 FILLER_34_2013 ();
 sg13g2_fill_1 FILLER_34_2015 ();
 sg13g2_decap_4 FILLER_34_2034 ();
 sg13g2_fill_1 FILLER_34_2038 ();
 sg13g2_fill_2 FILLER_34_2053 ();
 sg13g2_fill_1 FILLER_34_2055 ();
 sg13g2_fill_2 FILLER_34_2060 ();
 sg13g2_fill_1 FILLER_34_2067 ();
 sg13g2_fill_2 FILLER_34_2073 ();
 sg13g2_fill_1 FILLER_34_2075 ();
 sg13g2_fill_2 FILLER_34_2104 ();
 sg13g2_fill_1 FILLER_34_2106 ();
 sg13g2_fill_2 FILLER_34_2124 ();
 sg13g2_fill_1 FILLER_34_2139 ();
 sg13g2_fill_2 FILLER_34_2154 ();
 sg13g2_decap_4 FILLER_34_2192 ();
 sg13g2_fill_1 FILLER_34_2196 ();
 sg13g2_decap_8 FILLER_34_2205 ();
 sg13g2_fill_1 FILLER_34_2212 ();
 sg13g2_decap_8 FILLER_34_2227 ();
 sg13g2_fill_2 FILLER_34_2234 ();
 sg13g2_fill_2 FILLER_34_2276 ();
 sg13g2_fill_2 FILLER_34_2282 ();
 sg13g2_fill_1 FILLER_34_2284 ();
 sg13g2_fill_2 FILLER_34_2298 ();
 sg13g2_fill_2 FILLER_34_2326 ();
 sg13g2_fill_1 FILLER_34_2340 ();
 sg13g2_decap_8 FILLER_34_2344 ();
 sg13g2_fill_2 FILLER_34_2351 ();
 sg13g2_fill_2 FILLER_34_2372 ();
 sg13g2_fill_1 FILLER_34_2374 ();
 sg13g2_decap_8 FILLER_34_2388 ();
 sg13g2_fill_2 FILLER_34_2395 ();
 sg13g2_fill_1 FILLER_34_2401 ();
 sg13g2_decap_4 FILLER_34_2419 ();
 sg13g2_fill_1 FILLER_34_2423 ();
 sg13g2_fill_2 FILLER_34_2445 ();
 sg13g2_fill_1 FILLER_34_2447 ();
 sg13g2_decap_4 FILLER_34_2474 ();
 sg13g2_fill_1 FILLER_34_2478 ();
 sg13g2_fill_2 FILLER_34_2533 ();
 sg13g2_decap_4 FILLER_34_2544 ();
 sg13g2_fill_1 FILLER_34_2548 ();
 sg13g2_fill_1 FILLER_34_2558 ();
 sg13g2_decap_8 FILLER_34_2572 ();
 sg13g2_fill_1 FILLER_34_2579 ();
 sg13g2_fill_2 FILLER_34_2649 ();
 sg13g2_decap_8 FILLER_34_2679 ();
 sg13g2_decap_8 FILLER_34_2686 ();
 sg13g2_decap_4 FILLER_34_2693 ();
 sg13g2_fill_1 FILLER_34_2697 ();
 sg13g2_decap_8 FILLER_34_2741 ();
 sg13g2_fill_1 FILLER_34_2748 ();
 sg13g2_fill_1 FILLER_34_2774 ();
 sg13g2_decap_4 FILLER_34_2798 ();
 sg13g2_fill_2 FILLER_34_2802 ();
 sg13g2_fill_2 FILLER_34_2829 ();
 sg13g2_decap_4 FILLER_34_2840 ();
 sg13g2_fill_1 FILLER_34_2866 ();
 sg13g2_decap_4 FILLER_34_2902 ();
 sg13g2_fill_1 FILLER_34_2906 ();
 sg13g2_decap_4 FILLER_34_2957 ();
 sg13g2_fill_2 FILLER_34_2961 ();
 sg13g2_fill_2 FILLER_34_2981 ();
 sg13g2_decap_8 FILLER_34_3014 ();
 sg13g2_fill_2 FILLER_34_3031 ();
 sg13g2_fill_1 FILLER_34_3033 ();
 sg13g2_fill_1 FILLER_34_3039 ();
 sg13g2_fill_2 FILLER_34_3045 ();
 sg13g2_fill_1 FILLER_34_3047 ();
 sg13g2_decap_8 FILLER_34_3061 ();
 sg13g2_decap_4 FILLER_34_3068 ();
 sg13g2_fill_2 FILLER_34_3089 ();
 sg13g2_decap_8 FILLER_34_3108 ();
 sg13g2_decap_8 FILLER_34_3134 ();
 sg13g2_fill_2 FILLER_34_3141 ();
 sg13g2_fill_2 FILLER_34_3169 ();
 sg13g2_fill_1 FILLER_34_3171 ();
 sg13g2_decap_4 FILLER_34_3176 ();
 sg13g2_fill_1 FILLER_34_3180 ();
 sg13g2_fill_1 FILLER_34_3189 ();
 sg13g2_fill_2 FILLER_34_3201 ();
 sg13g2_decap_4 FILLER_34_3211 ();
 sg13g2_fill_2 FILLER_34_3220 ();
 sg13g2_fill_1 FILLER_34_3222 ();
 sg13g2_decap_8 FILLER_34_3240 ();
 sg13g2_decap_8 FILLER_34_3247 ();
 sg13g2_fill_1 FILLER_34_3266 ();
 sg13g2_fill_1 FILLER_34_3281 ();
 sg13g2_fill_2 FILLER_34_3323 ();
 sg13g2_fill_2 FILLER_34_3389 ();
 sg13g2_fill_1 FILLER_34_3391 ();
 sg13g2_decap_8 FILLER_34_3406 ();
 sg13g2_fill_1 FILLER_34_3426 ();
 sg13g2_decap_8 FILLER_34_3431 ();
 sg13g2_decap_8 FILLER_34_3438 ();
 sg13g2_decap_4 FILLER_34_3445 ();
 sg13g2_fill_2 FILLER_34_3449 ();
 sg13g2_fill_2 FILLER_34_3461 ();
 sg13g2_decap_8 FILLER_34_3467 ();
 sg13g2_decap_8 FILLER_34_3474 ();
 sg13g2_fill_2 FILLER_34_3481 ();
 sg13g2_fill_1 FILLER_34_3483 ();
 sg13g2_decap_8 FILLER_34_3497 ();
 sg13g2_decap_8 FILLER_34_3504 ();
 sg13g2_decap_8 FILLER_34_3511 ();
 sg13g2_decap_8 FILLER_34_3518 ();
 sg13g2_decap_8 FILLER_34_3525 ();
 sg13g2_decap_8 FILLER_34_3532 ();
 sg13g2_decap_8 FILLER_34_3539 ();
 sg13g2_decap_8 FILLER_34_3546 ();
 sg13g2_decap_8 FILLER_34_3553 ();
 sg13g2_decap_8 FILLER_34_3560 ();
 sg13g2_decap_8 FILLER_34_3567 ();
 sg13g2_decap_4 FILLER_34_3574 ();
 sg13g2_fill_2 FILLER_34_3578 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_4 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_226 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_241 ();
 sg13g2_decap_8 FILLER_35_248 ();
 sg13g2_decap_4 FILLER_35_255 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_271 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_decap_4 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_314 ();
 sg13g2_decap_4 FILLER_35_321 ();
 sg13g2_fill_2 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_343 ();
 sg13g2_decap_4 FILLER_35_348 ();
 sg13g2_decap_4 FILLER_35_380 ();
 sg13g2_fill_2 FILLER_35_425 ();
 sg13g2_fill_1 FILLER_35_427 ();
 sg13g2_decap_4 FILLER_35_474 ();
 sg13g2_fill_2 FILLER_35_483 ();
 sg13g2_decap_4 FILLER_35_510 ();
 sg13g2_fill_2 FILLER_35_514 ();
 sg13g2_decap_8 FILLER_35_549 ();
 sg13g2_decap_4 FILLER_35_556 ();
 sg13g2_decap_8 FILLER_35_572 ();
 sg13g2_fill_1 FILLER_35_587 ();
 sg13g2_decap_4 FILLER_35_592 ();
 sg13g2_fill_2 FILLER_35_641 ();
 sg13g2_fill_1 FILLER_35_643 ();
 sg13g2_fill_1 FILLER_35_680 ();
 sg13g2_fill_2 FILLER_35_717 ();
 sg13g2_fill_1 FILLER_35_719 ();
 sg13g2_decap_8 FILLER_35_725 ();
 sg13g2_fill_1 FILLER_35_760 ();
 sg13g2_fill_1 FILLER_35_766 ();
 sg13g2_decap_4 FILLER_35_780 ();
 sg13g2_fill_2 FILLER_35_784 ();
 sg13g2_decap_4 FILLER_35_798 ();
 sg13g2_fill_2 FILLER_35_820 ();
 sg13g2_fill_1 FILLER_35_822 ();
 sg13g2_decap_4 FILLER_35_827 ();
 sg13g2_fill_2 FILLER_35_831 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_fill_2 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_fill_2 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_35_880 ();
 sg13g2_decap_8 FILLER_35_887 ();
 sg13g2_decap_8 FILLER_35_898 ();
 sg13g2_fill_2 FILLER_35_905 ();
 sg13g2_fill_2 FILLER_35_923 ();
 sg13g2_decap_8 FILLER_35_943 ();
 sg13g2_fill_2 FILLER_35_950 ();
 sg13g2_fill_1 FILLER_35_952 ();
 sg13g2_fill_1 FILLER_35_957 ();
 sg13g2_fill_2 FILLER_35_968 ();
 sg13g2_decap_8 FILLER_35_978 ();
 sg13g2_fill_1 FILLER_35_985 ();
 sg13g2_fill_1 FILLER_35_1003 ();
 sg13g2_fill_1 FILLER_35_1021 ();
 sg13g2_fill_2 FILLER_35_1036 ();
 sg13g2_decap_4 FILLER_35_1060 ();
 sg13g2_fill_2 FILLER_35_1064 ();
 sg13g2_fill_2 FILLER_35_1098 ();
 sg13g2_fill_2 FILLER_35_1128 ();
 sg13g2_fill_1 FILLER_35_1143 ();
 sg13g2_fill_1 FILLER_35_1157 ();
 sg13g2_fill_2 FILLER_35_1165 ();
 sg13g2_decap_4 FILLER_35_1172 ();
 sg13g2_fill_2 FILLER_35_1176 ();
 sg13g2_decap_8 FILLER_35_1196 ();
 sg13g2_decap_8 FILLER_35_1203 ();
 sg13g2_fill_1 FILLER_35_1210 ();
 sg13g2_fill_2 FILLER_35_1219 ();
 sg13g2_fill_1 FILLER_35_1221 ();
 sg13g2_fill_2 FILLER_35_1226 ();
 sg13g2_fill_2 FILLER_35_1258 ();
 sg13g2_decap_8 FILLER_35_1268 ();
 sg13g2_decap_4 FILLER_35_1275 ();
 sg13g2_fill_2 FILLER_35_1279 ();
 sg13g2_fill_1 FILLER_35_1294 ();
 sg13g2_decap_4 FILLER_35_1330 ();
 sg13g2_fill_1 FILLER_35_1334 ();
 sg13g2_fill_2 FILLER_35_1344 ();
 sg13g2_decap_8 FILLER_35_1382 ();
 sg13g2_decap_8 FILLER_35_1402 ();
 sg13g2_fill_2 FILLER_35_1409 ();
 sg13g2_fill_2 FILLER_35_1416 ();
 sg13g2_fill_1 FILLER_35_1440 ();
 sg13g2_decap_8 FILLER_35_1454 ();
 sg13g2_decap_8 FILLER_35_1461 ();
 sg13g2_fill_2 FILLER_35_1494 ();
 sg13g2_fill_1 FILLER_35_1496 ();
 sg13g2_decap_4 FILLER_35_1518 ();
 sg13g2_fill_1 FILLER_35_1588 ();
 sg13g2_decap_8 FILLER_35_1607 ();
 sg13g2_fill_2 FILLER_35_1614 ();
 sg13g2_fill_1 FILLER_35_1616 ();
 sg13g2_fill_2 FILLER_35_1657 ();
 sg13g2_fill_1 FILLER_35_1659 ();
 sg13g2_decap_4 FILLER_35_1721 ();
 sg13g2_fill_1 FILLER_35_1725 ();
 sg13g2_decap_8 FILLER_35_1730 ();
 sg13g2_fill_2 FILLER_35_1737 ();
 sg13g2_fill_1 FILLER_35_1739 ();
 sg13g2_decap_8 FILLER_35_1744 ();
 sg13g2_fill_1 FILLER_35_1751 ();
 sg13g2_fill_1 FILLER_35_1769 ();
 sg13g2_decap_4 FILLER_35_1779 ();
 sg13g2_fill_2 FILLER_35_1783 ();
 sg13g2_decap_8 FILLER_35_1789 ();
 sg13g2_decap_8 FILLER_35_1796 ();
 sg13g2_fill_2 FILLER_35_1803 ();
 sg13g2_fill_1 FILLER_35_1805 ();
 sg13g2_fill_1 FILLER_35_1815 ();
 sg13g2_fill_2 FILLER_35_1868 ();
 sg13g2_decap_4 FILLER_35_1907 ();
 sg13g2_fill_1 FILLER_35_1911 ();
 sg13g2_fill_2 FILLER_35_1925 ();
 sg13g2_decap_8 FILLER_35_1942 ();
 sg13g2_fill_2 FILLER_35_1949 ();
 sg13g2_fill_1 FILLER_35_1951 ();
 sg13g2_decap_4 FILLER_35_1974 ();
 sg13g2_fill_2 FILLER_35_1978 ();
 sg13g2_decap_4 FILLER_35_2012 ();
 sg13g2_fill_2 FILLER_35_2016 ();
 sg13g2_fill_1 FILLER_35_2050 ();
 sg13g2_fill_2 FILLER_35_2054 ();
 sg13g2_fill_1 FILLER_35_2056 ();
 sg13g2_fill_2 FILLER_35_2079 ();
 sg13g2_decap_8 FILLER_35_2094 ();
 sg13g2_decap_4 FILLER_35_2101 ();
 sg13g2_fill_1 FILLER_35_2105 ();
 sg13g2_decap_8 FILLER_35_2178 ();
 sg13g2_decap_8 FILLER_35_2185 ();
 sg13g2_decap_4 FILLER_35_2192 ();
 sg13g2_fill_1 FILLER_35_2196 ();
 sg13g2_decap_8 FILLER_35_2201 ();
 sg13g2_fill_2 FILLER_35_2208 ();
 sg13g2_decap_4 FILLER_35_2247 ();
 sg13g2_fill_1 FILLER_35_2251 ();
 sg13g2_fill_2 FILLER_35_2298 ();
 sg13g2_fill_1 FILLER_35_2300 ();
 sg13g2_fill_1 FILLER_35_2310 ();
 sg13g2_fill_1 FILLER_35_2324 ();
 sg13g2_fill_1 FILLER_35_2335 ();
 sg13g2_fill_1 FILLER_35_2341 ();
 sg13g2_fill_1 FILLER_35_2360 ();
 sg13g2_fill_1 FILLER_35_2366 ();
 sg13g2_decap_4 FILLER_35_2393 ();
 sg13g2_fill_2 FILLER_35_2397 ();
 sg13g2_fill_2 FILLER_35_2404 ();
 sg13g2_decap_8 FILLER_35_2410 ();
 sg13g2_decap_8 FILLER_35_2417 ();
 sg13g2_decap_8 FILLER_35_2441 ();
 sg13g2_fill_2 FILLER_35_2448 ();
 sg13g2_fill_1 FILLER_35_2450 ();
 sg13g2_decap_4 FILLER_35_2484 ();
 sg13g2_fill_1 FILLER_35_2488 ();
 sg13g2_fill_2 FILLER_35_2502 ();
 sg13g2_fill_1 FILLER_35_2504 ();
 sg13g2_fill_1 FILLER_35_2512 ();
 sg13g2_fill_1 FILLER_35_2534 ();
 sg13g2_fill_2 FILLER_35_2568 ();
 sg13g2_fill_1 FILLER_35_2570 ();
 sg13g2_fill_1 FILLER_35_2584 ();
 sg13g2_fill_2 FILLER_35_2591 ();
 sg13g2_fill_1 FILLER_35_2593 ();
 sg13g2_decap_8 FILLER_35_2598 ();
 sg13g2_decap_4 FILLER_35_2605 ();
 sg13g2_fill_2 FILLER_35_2609 ();
 sg13g2_fill_2 FILLER_35_2618 ();
 sg13g2_decap_8 FILLER_35_2624 ();
 sg13g2_decap_4 FILLER_35_2631 ();
 sg13g2_fill_2 FILLER_35_2635 ();
 sg13g2_fill_1 FILLER_35_2655 ();
 sg13g2_decap_8 FILLER_35_2663 ();
 sg13g2_decap_4 FILLER_35_2670 ();
 sg13g2_fill_2 FILLER_35_2674 ();
 sg13g2_decap_4 FILLER_35_2704 ();
 sg13g2_decap_4 FILLER_35_2721 ();
 sg13g2_fill_1 FILLER_35_2725 ();
 sg13g2_fill_2 FILLER_35_2810 ();
 sg13g2_decap_4 FILLER_35_2826 ();
 sg13g2_fill_1 FILLER_35_2830 ();
 sg13g2_decap_8 FILLER_35_2839 ();
 sg13g2_decap_4 FILLER_35_2846 ();
 sg13g2_fill_1 FILLER_35_2850 ();
 sg13g2_decap_8 FILLER_35_2858 ();
 sg13g2_decap_8 FILLER_35_2865 ();
 sg13g2_decap_4 FILLER_35_2883 ();
 sg13g2_fill_1 FILLER_35_2887 ();
 sg13g2_decap_8 FILLER_35_2900 ();
 sg13g2_decap_8 FILLER_35_2907 ();
 sg13g2_decap_4 FILLER_35_2914 ();
 sg13g2_decap_8 FILLER_35_2940 ();
 sg13g2_fill_2 FILLER_35_2947 ();
 sg13g2_decap_8 FILLER_35_2956 ();
 sg13g2_decap_8 FILLER_35_2963 ();
 sg13g2_decap_8 FILLER_35_3002 ();
 sg13g2_decap_4 FILLER_35_3009 ();
 sg13g2_fill_1 FILLER_35_3013 ();
 sg13g2_decap_4 FILLER_35_3034 ();
 sg13g2_fill_1 FILLER_35_3043 ();
 sg13g2_decap_8 FILLER_35_3053 ();
 sg13g2_fill_2 FILLER_35_3060 ();
 sg13g2_fill_2 FILLER_35_3090 ();
 sg13g2_fill_1 FILLER_35_3092 ();
 sg13g2_fill_1 FILLER_35_3101 ();
 sg13g2_fill_2 FILLER_35_3121 ();
 sg13g2_decap_8 FILLER_35_3134 ();
 sg13g2_decap_8 FILLER_35_3141 ();
 sg13g2_decap_4 FILLER_35_3180 ();
 sg13g2_fill_2 FILLER_35_3184 ();
 sg13g2_fill_2 FILLER_35_3192 ();
 sg13g2_decap_8 FILLER_35_3207 ();
 sg13g2_decap_8 FILLER_35_3214 ();
 sg13g2_decap_4 FILLER_35_3221 ();
 sg13g2_fill_1 FILLER_35_3225 ();
 sg13g2_decap_8 FILLER_35_3254 ();
 sg13g2_decap_4 FILLER_35_3293 ();
 sg13g2_decap_8 FILLER_35_3302 ();
 sg13g2_decap_4 FILLER_35_3309 ();
 sg13g2_fill_2 FILLER_35_3313 ();
 sg13g2_fill_1 FILLER_35_3320 ();
 sg13g2_decap_8 FILLER_35_3337 ();
 sg13g2_decap_8 FILLER_35_3344 ();
 sg13g2_fill_2 FILLER_35_3351 ();
 sg13g2_decap_4 FILLER_35_3356 ();
 sg13g2_fill_2 FILLER_35_3360 ();
 sg13g2_fill_2 FILLER_35_3383 ();
 sg13g2_decap_8 FILLER_35_3390 ();
 sg13g2_fill_1 FILLER_35_3397 ();
 sg13g2_decap_4 FILLER_35_3406 ();
 sg13g2_fill_2 FILLER_35_3410 ();
 sg13g2_decap_8 FILLER_35_3440 ();
 sg13g2_fill_2 FILLER_35_3447 ();
 sg13g2_fill_1 FILLER_35_3449 ();
 sg13g2_fill_2 FILLER_35_3486 ();
 sg13g2_decap_8 FILLER_35_3492 ();
 sg13g2_decap_8 FILLER_35_3499 ();
 sg13g2_decap_8 FILLER_35_3506 ();
 sg13g2_decap_8 FILLER_35_3513 ();
 sg13g2_decap_8 FILLER_35_3520 ();
 sg13g2_decap_8 FILLER_35_3527 ();
 sg13g2_decap_8 FILLER_35_3534 ();
 sg13g2_decap_8 FILLER_35_3541 ();
 sg13g2_decap_8 FILLER_35_3548 ();
 sg13g2_decap_8 FILLER_35_3555 ();
 sg13g2_decap_8 FILLER_35_3562 ();
 sg13g2_decap_8 FILLER_35_3569 ();
 sg13g2_decap_4 FILLER_35_3576 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_95 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_decap_4 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_176 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_decap_4 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_decap_4 FILLER_36_248 ();
 sg13g2_fill_1 FILLER_36_252 ();
 sg13g2_decap_4 FILLER_36_257 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_4 FILLER_36_381 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_decap_4 FILLER_36_395 ();
 sg13g2_decap_4 FILLER_36_407 ();
 sg13g2_fill_1 FILLER_36_411 ();
 sg13g2_fill_2 FILLER_36_420 ();
 sg13g2_fill_1 FILLER_36_422 ();
 sg13g2_decap_4 FILLER_36_468 ();
 sg13g2_fill_2 FILLER_36_480 ();
 sg13g2_fill_2 FILLER_36_490 ();
 sg13g2_fill_1 FILLER_36_492 ();
 sg13g2_decap_4 FILLER_36_518 ();
 sg13g2_fill_2 FILLER_36_530 ();
 sg13g2_fill_1 FILLER_36_537 ();
 sg13g2_fill_1 FILLER_36_547 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_decap_8 FILLER_36_598 ();
 sg13g2_decap_8 FILLER_36_605 ();
 sg13g2_fill_2 FILLER_36_612 ();
 sg13g2_fill_1 FILLER_36_614 ();
 sg13g2_fill_1 FILLER_36_628 ();
 sg13g2_fill_2 FILLER_36_695 ();
 sg13g2_fill_1 FILLER_36_697 ();
 sg13g2_decap_8 FILLER_36_707 ();
 sg13g2_decap_4 FILLER_36_714 ();
 sg13g2_fill_1 FILLER_36_736 ();
 sg13g2_decap_8 FILLER_36_741 ();
 sg13g2_decap_4 FILLER_36_748 ();
 sg13g2_fill_1 FILLER_36_774 ();
 sg13g2_decap_8 FILLER_36_801 ();
 sg13g2_fill_2 FILLER_36_808 ();
 sg13g2_fill_1 FILLER_36_838 ();
 sg13g2_decap_4 FILLER_36_844 ();
 sg13g2_fill_2 FILLER_36_848 ();
 sg13g2_fill_2 FILLER_36_855 ();
 sg13g2_fill_1 FILLER_36_857 ();
 sg13g2_decap_4 FILLER_36_895 ();
 sg13g2_fill_1 FILLER_36_960 ();
 sg13g2_fill_2 FILLER_36_973 ();
 sg13g2_fill_2 FILLER_36_984 ();
 sg13g2_fill_2 FILLER_36_1075 ();
 sg13g2_fill_1 FILLER_36_1090 ();
 sg13g2_fill_1 FILLER_36_1113 ();
 sg13g2_fill_2 FILLER_36_1119 ();
 sg13g2_fill_1 FILLER_36_1125 ();
 sg13g2_fill_1 FILLER_36_1143 ();
 sg13g2_fill_2 FILLER_36_1177 ();
 sg13g2_fill_1 FILLER_36_1179 ();
 sg13g2_decap_4 FILLER_36_1212 ();
 sg13g2_fill_1 FILLER_36_1216 ();
 sg13g2_decap_4 FILLER_36_1269 ();
 sg13g2_fill_1 FILLER_36_1273 ();
 sg13g2_decap_4 FILLER_36_1311 ();
 sg13g2_fill_1 FILLER_36_1315 ();
 sg13g2_decap_8 FILLER_36_1368 ();
 sg13g2_decap_4 FILLER_36_1427 ();
 sg13g2_fill_1 FILLER_36_1459 ();
 sg13g2_fill_2 FILLER_36_1490 ();
 sg13g2_fill_1 FILLER_36_1492 ();
 sg13g2_decap_8 FILLER_36_1536 ();
 sg13g2_fill_1 FILLER_36_1543 ();
 sg13g2_fill_2 FILLER_36_1557 ();
 sg13g2_fill_1 FILLER_36_1559 ();
 sg13g2_decap_8 FILLER_36_1626 ();
 sg13g2_fill_1 FILLER_36_1633 ();
 sg13g2_decap_4 FILLER_36_1638 ();
 sg13g2_decap_4 FILLER_36_1654 ();
 sg13g2_fill_2 FILLER_36_1658 ();
 sg13g2_fill_2 FILLER_36_1675 ();
 sg13g2_fill_1 FILLER_36_1686 ();
 sg13g2_decap_4 FILLER_36_1709 ();
 sg13g2_fill_2 FILLER_36_1713 ();
 sg13g2_fill_2 FILLER_36_1719 ();
 sg13g2_fill_1 FILLER_36_1721 ();
 sg13g2_fill_2 FILLER_36_1740 ();
 sg13g2_fill_1 FILLER_36_1742 ();
 sg13g2_fill_2 FILLER_36_1759 ();
 sg13g2_fill_1 FILLER_36_1770 ();
 sg13g2_fill_1 FILLER_36_1776 ();
 sg13g2_decap_8 FILLER_36_1799 ();
 sg13g2_fill_2 FILLER_36_1806 ();
 sg13g2_fill_2 FILLER_36_1852 ();
 sg13g2_fill_1 FILLER_36_1854 ();
 sg13g2_decap_8 FILLER_36_1859 ();
 sg13g2_fill_2 FILLER_36_1866 ();
 sg13g2_fill_1 FILLER_36_1868 ();
 sg13g2_decap_8 FILLER_36_1877 ();
 sg13g2_fill_1 FILLER_36_1884 ();
 sg13g2_decap_4 FILLER_36_1889 ();
 sg13g2_decap_8 FILLER_36_1921 ();
 sg13g2_fill_2 FILLER_36_1928 ();
 sg13g2_fill_2 FILLER_36_1941 ();
 sg13g2_fill_1 FILLER_36_1984 ();
 sg13g2_decap_8 FILLER_36_1993 ();
 sg13g2_decap_4 FILLER_36_2000 ();
 sg13g2_fill_1 FILLER_36_2004 ();
 sg13g2_fill_1 FILLER_36_2022 ();
 sg13g2_decap_8 FILLER_36_2027 ();
 sg13g2_decap_8 FILLER_36_2034 ();
 sg13g2_fill_1 FILLER_36_2041 ();
 sg13g2_fill_2 FILLER_36_2063 ();
 sg13g2_fill_1 FILLER_36_2065 ();
 sg13g2_decap_8 FILLER_36_2094 ();
 sg13g2_decap_8 FILLER_36_2101 ();
 sg13g2_decap_8 FILLER_36_2108 ();
 sg13g2_fill_2 FILLER_36_2115 ();
 sg13g2_fill_1 FILLER_36_2117 ();
 sg13g2_decap_4 FILLER_36_2128 ();
 sg13g2_decap_4 FILLER_36_2159 ();
 sg13g2_fill_1 FILLER_36_2163 ();
 sg13g2_fill_2 FILLER_36_2192 ();
 sg13g2_fill_1 FILLER_36_2194 ();
 sg13g2_fill_2 FILLER_36_2204 ();
 sg13g2_decap_8 FILLER_36_2232 ();
 sg13g2_decap_4 FILLER_36_2239 ();
 sg13g2_decap_8 FILLER_36_2274 ();
 sg13g2_fill_1 FILLER_36_2294 ();
 sg13g2_decap_8 FILLER_36_2323 ();
 sg13g2_fill_2 FILLER_36_2330 ();
 sg13g2_fill_1 FILLER_36_2332 ();
 sg13g2_decap_8 FILLER_36_2376 ();
 sg13g2_decap_4 FILLER_36_2409 ();
 sg13g2_fill_1 FILLER_36_2413 ();
 sg13g2_fill_1 FILLER_36_2418 ();
 sg13g2_fill_2 FILLER_36_2456 ();
 sg13g2_fill_1 FILLER_36_2505 ();
 sg13g2_fill_2 FILLER_36_2515 ();
 sg13g2_fill_2 FILLER_36_2535 ();
 sg13g2_fill_2 FILLER_36_2550 ();
 sg13g2_fill_2 FILLER_36_2565 ();
 sg13g2_fill_1 FILLER_36_2567 ();
 sg13g2_decap_8 FILLER_36_2596 ();
 sg13g2_decap_4 FILLER_36_2603 ();
 sg13g2_decap_4 FILLER_36_2625 ();
 sg13g2_decap_8 FILLER_36_2670 ();
 sg13g2_fill_1 FILLER_36_2677 ();
 sg13g2_decap_8 FILLER_36_2687 ();
 sg13g2_decap_4 FILLER_36_2694 ();
 sg13g2_fill_1 FILLER_36_2730 ();
 sg13g2_decap_8 FILLER_36_2735 ();
 sg13g2_decap_8 FILLER_36_2742 ();
 sg13g2_decap_4 FILLER_36_2749 ();
 sg13g2_decap_4 FILLER_36_2761 ();
 sg13g2_fill_1 FILLER_36_2765 ();
 sg13g2_decap_4 FILLER_36_2782 ();
 sg13g2_decap_8 FILLER_36_2799 ();
 sg13g2_fill_2 FILLER_36_2806 ();
 sg13g2_fill_1 FILLER_36_2808 ();
 sg13g2_decap_4 FILLER_36_2841 ();
 sg13g2_fill_2 FILLER_36_2863 ();
 sg13g2_decap_8 FILLER_36_2892 ();
 sg13g2_decap_8 FILLER_36_2899 ();
 sg13g2_decap_4 FILLER_36_2906 ();
 sg13g2_fill_1 FILLER_36_2910 ();
 sg13g2_fill_2 FILLER_36_2939 ();
 sg13g2_fill_1 FILLER_36_2973 ();
 sg13g2_decap_8 FILLER_36_2990 ();
 sg13g2_decap_8 FILLER_36_2997 ();
 sg13g2_decap_8 FILLER_36_3004 ();
 sg13g2_decap_8 FILLER_36_3011 ();
 sg13g2_fill_1 FILLER_36_3018 ();
 sg13g2_fill_2 FILLER_36_3024 ();
 sg13g2_fill_2 FILLER_36_3033 ();
 sg13g2_decap_8 FILLER_36_3050 ();
 sg13g2_decap_8 FILLER_36_3057 ();
 sg13g2_decap_8 FILLER_36_3064 ();
 sg13g2_fill_1 FILLER_36_3071 ();
 sg13g2_decap_8 FILLER_36_3130 ();
 sg13g2_fill_2 FILLER_36_3150 ();
 sg13g2_fill_1 FILLER_36_3156 ();
 sg13g2_fill_1 FILLER_36_3169 ();
 sg13g2_decap_8 FILLER_36_3174 ();
 sg13g2_decap_4 FILLER_36_3227 ();
 sg13g2_fill_1 FILLER_36_3235 ();
 sg13g2_fill_1 FILLER_36_3244 ();
 sg13g2_fill_2 FILLER_36_3255 ();
 sg13g2_fill_1 FILLER_36_3257 ();
 sg13g2_decap_4 FILLER_36_3275 ();
 sg13g2_fill_2 FILLER_36_3279 ();
 sg13g2_fill_2 FILLER_36_3321 ();
 sg13g2_fill_2 FILLER_36_3366 ();
 sg13g2_fill_1 FILLER_36_3368 ();
 sg13g2_fill_2 FILLER_36_3397 ();
 sg13g2_decap_8 FILLER_36_3403 ();
 sg13g2_decap_4 FILLER_36_3410 ();
 sg13g2_fill_2 FILLER_36_3414 ();
 sg13g2_fill_1 FILLER_36_3428 ();
 sg13g2_fill_2 FILLER_36_3451 ();
 sg13g2_fill_1 FILLER_36_3453 ();
 sg13g2_decap_8 FILLER_36_3502 ();
 sg13g2_decap_8 FILLER_36_3509 ();
 sg13g2_decap_8 FILLER_36_3516 ();
 sg13g2_decap_8 FILLER_36_3523 ();
 sg13g2_decap_8 FILLER_36_3530 ();
 sg13g2_decap_8 FILLER_36_3537 ();
 sg13g2_decap_8 FILLER_36_3544 ();
 sg13g2_decap_8 FILLER_36_3551 ();
 sg13g2_decap_8 FILLER_36_3558 ();
 sg13g2_decap_8 FILLER_36_3565 ();
 sg13g2_decap_8 FILLER_36_3572 ();
 sg13g2_fill_1 FILLER_36_3579 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_117 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_fill_2 FILLER_37_131 ();
 sg13g2_fill_2 FILLER_37_169 ();
 sg13g2_decap_4 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_decap_4 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_226 ();
 sg13g2_decap_4 FILLER_37_246 ();
 sg13g2_decap_4 FILLER_37_275 ();
 sg13g2_fill_2 FILLER_37_279 ();
 sg13g2_decap_8 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_314 ();
 sg13g2_decap_8 FILLER_37_324 ();
 sg13g2_decap_4 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_356 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_410 ();
 sg13g2_decap_4 FILLER_37_417 ();
 sg13g2_fill_1 FILLER_37_421 ();
 sg13g2_decap_8 FILLER_37_435 ();
 sg13g2_decap_4 FILLER_37_442 ();
 sg13g2_decap_4 FILLER_37_472 ();
 sg13g2_fill_2 FILLER_37_486 ();
 sg13g2_decap_8 FILLER_37_493 ();
 sg13g2_decap_4 FILLER_37_500 ();
 sg13g2_fill_2 FILLER_37_504 ();
 sg13g2_decap_4 FILLER_37_511 ();
 sg13g2_fill_2 FILLER_37_523 ();
 sg13g2_fill_1 FILLER_37_525 ();
 sg13g2_fill_2 FILLER_37_553 ();
 sg13g2_fill_1 FILLER_37_555 ();
 sg13g2_decap_8 FILLER_37_593 ();
 sg13g2_decap_8 FILLER_37_600 ();
 sg13g2_decap_4 FILLER_37_607 ();
 sg13g2_fill_2 FILLER_37_628 ();
 sg13g2_fill_1 FILLER_37_630 ();
 sg13g2_decap_4 FILLER_37_644 ();
 sg13g2_fill_1 FILLER_37_648 ();
 sg13g2_fill_1 FILLER_37_654 ();
 sg13g2_fill_2 FILLER_37_659 ();
 sg13g2_fill_2 FILLER_37_683 ();
 sg13g2_fill_1 FILLER_37_685 ();
 sg13g2_decap_8 FILLER_37_717 ();
 sg13g2_fill_1 FILLER_37_724 ();
 sg13g2_fill_2 FILLER_37_733 ();
 sg13g2_fill_1 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_740 ();
 sg13g2_fill_1 FILLER_37_747 ();
 sg13g2_fill_2 FILLER_37_756 ();
 sg13g2_fill_2 FILLER_37_763 ();
 sg13g2_fill_2 FILLER_37_820 ();
 sg13g2_fill_1 FILLER_37_822 ();
 sg13g2_fill_2 FILLER_37_837 ();
 sg13g2_decap_4 FILLER_37_868 ();
 sg13g2_decap_4 FILLER_37_898 ();
 sg13g2_fill_1 FILLER_37_902 ();
 sg13g2_decap_8 FILLER_37_931 ();
 sg13g2_decap_8 FILLER_37_938 ();
 sg13g2_fill_2 FILLER_37_945 ();
 sg13g2_fill_1 FILLER_37_947 ();
 sg13g2_decap_4 FILLER_37_952 ();
 sg13g2_fill_1 FILLER_37_956 ();
 sg13g2_decap_4 FILLER_37_984 ();
 sg13g2_fill_2 FILLER_37_988 ();
 sg13g2_decap_8 FILLER_37_1009 ();
 sg13g2_decap_8 FILLER_37_1016 ();
 sg13g2_decap_8 FILLER_37_1023 ();
 sg13g2_decap_8 FILLER_37_1030 ();
 sg13g2_decap_4 FILLER_37_1037 ();
 sg13g2_decap_4 FILLER_37_1044 ();
 sg13g2_fill_1 FILLER_37_1048 ();
 sg13g2_fill_1 FILLER_37_1059 ();
 sg13g2_fill_2 FILLER_37_1073 ();
 sg13g2_fill_2 FILLER_37_1102 ();
 sg13g2_fill_1 FILLER_37_1104 ();
 sg13g2_decap_8 FILLER_37_1132 ();
 sg13g2_fill_2 FILLER_37_1139 ();
 sg13g2_fill_2 FILLER_37_1144 ();
 sg13g2_decap_8 FILLER_37_1165 ();
 sg13g2_decap_4 FILLER_37_1172 ();
 sg13g2_decap_8 FILLER_37_1252 ();
 sg13g2_fill_2 FILLER_37_1259 ();
 sg13g2_decap_4 FILLER_37_1265 ();
 sg13g2_decap_8 FILLER_37_1297 ();
 sg13g2_decap_4 FILLER_37_1317 ();
 sg13g2_fill_1 FILLER_37_1339 ();
 sg13g2_decap_4 FILLER_37_1345 ();
 sg13g2_decap_8 FILLER_37_1352 ();
 sg13g2_fill_2 FILLER_37_1359 ();
 sg13g2_fill_1 FILLER_37_1366 ();
 sg13g2_fill_2 FILLER_37_1388 ();
 sg13g2_decap_8 FILLER_37_1394 ();
 sg13g2_decap_4 FILLER_37_1401 ();
 sg13g2_fill_2 FILLER_37_1405 ();
 sg13g2_fill_2 FILLER_37_1433 ();
 sg13g2_fill_1 FILLER_37_1435 ();
 sg13g2_decap_4 FILLER_37_1440 ();
 sg13g2_decap_4 FILLER_37_1465 ();
 sg13g2_decap_4 FILLER_37_1483 ();
 sg13g2_fill_1 FILLER_37_1487 ();
 sg13g2_fill_1 FILLER_37_1500 ();
 sg13g2_decap_8 FILLER_37_1535 ();
 sg13g2_fill_1 FILLER_37_1565 ();
 sg13g2_decap_8 FILLER_37_1571 ();
 sg13g2_decap_8 FILLER_37_1578 ();
 sg13g2_fill_1 FILLER_37_1585 ();
 sg13g2_decap_8 FILLER_37_1599 ();
 sg13g2_decap_4 FILLER_37_1606 ();
 sg13g2_fill_2 FILLER_37_1610 ();
 sg13g2_decap_8 FILLER_37_1632 ();
 sg13g2_fill_2 FILLER_37_1746 ();
 sg13g2_fill_2 FILLER_37_1754 ();
 sg13g2_fill_1 FILLER_37_1756 ();
 sg13g2_fill_2 FILLER_37_1766 ();
 sg13g2_fill_1 FILLER_37_1768 ();
 sg13g2_decap_4 FILLER_37_1773 ();
 sg13g2_fill_1 FILLER_37_1777 ();
 sg13g2_fill_2 FILLER_37_1783 ();
 sg13g2_decap_4 FILLER_37_1821 ();
 sg13g2_fill_2 FILLER_37_1825 ();
 sg13g2_fill_2 FILLER_37_1845 ();
 sg13g2_fill_2 FILLER_37_1856 ();
 sg13g2_fill_2 FILLER_37_1866 ();
 sg13g2_decap_4 FILLER_37_1876 ();
 sg13g2_decap_8 FILLER_37_1908 ();
 sg13g2_decap_4 FILLER_37_1915 ();
 sg13g2_fill_1 FILLER_37_1919 ();
 sg13g2_decap_8 FILLER_37_1943 ();
 sg13g2_decap_8 FILLER_37_1950 ();
 sg13g2_fill_2 FILLER_37_1957 ();
 sg13g2_fill_1 FILLER_37_1959 ();
 sg13g2_decap_8 FILLER_37_1986 ();
 sg13g2_decap_8 FILLER_37_1993 ();
 sg13g2_decap_4 FILLER_37_2000 ();
 sg13g2_fill_2 FILLER_37_2022 ();
 sg13g2_decap_4 FILLER_37_2030 ();
 sg13g2_fill_1 FILLER_37_2034 ();
 sg13g2_fill_1 FILLER_37_2038 ();
 sg13g2_decap_8 FILLER_37_2048 ();
 sg13g2_fill_2 FILLER_37_2055 ();
 sg13g2_fill_1 FILLER_37_2062 ();
 sg13g2_fill_2 FILLER_37_2083 ();
 sg13g2_fill_1 FILLER_37_2085 ();
 sg13g2_fill_1 FILLER_37_2094 ();
 sg13g2_fill_1 FILLER_37_2111 ();
 sg13g2_decap_4 FILLER_37_2131 ();
 sg13g2_fill_1 FILLER_37_2135 ();
 sg13g2_decap_4 FILLER_37_2156 ();
 sg13g2_fill_2 FILLER_37_2160 ();
 sg13g2_fill_2 FILLER_37_2187 ();
 sg13g2_decap_4 FILLER_37_2230 ();
 sg13g2_fill_2 FILLER_37_2234 ();
 sg13g2_fill_2 FILLER_37_2249 ();
 sg13g2_fill_1 FILLER_37_2292 ();
 sg13g2_decap_4 FILLER_37_2325 ();
 sg13g2_fill_1 FILLER_37_2329 ();
 sg13g2_decap_4 FILLER_37_2340 ();
 sg13g2_decap_4 FILLER_37_2350 ();
 sg13g2_decap_8 FILLER_37_2358 ();
 sg13g2_fill_2 FILLER_37_2365 ();
 sg13g2_fill_1 FILLER_37_2371 ();
 sg13g2_decap_4 FILLER_37_2381 ();
 sg13g2_fill_1 FILLER_37_2385 ();
 sg13g2_decap_8 FILLER_37_2425 ();
 sg13g2_fill_1 FILLER_37_2432 ();
 sg13g2_decap_8 FILLER_37_2442 ();
 sg13g2_fill_1 FILLER_37_2449 ();
 sg13g2_decap_8 FILLER_37_2474 ();
 sg13g2_decap_4 FILLER_37_2481 ();
 sg13g2_fill_2 FILLER_37_2531 ();
 sg13g2_fill_1 FILLER_37_2541 ();
 sg13g2_decap_8 FILLER_37_2570 ();
 sg13g2_decap_4 FILLER_37_2577 ();
 sg13g2_fill_1 FILLER_37_2581 ();
 sg13g2_decap_8 FILLER_37_2594 ();
 sg13g2_fill_1 FILLER_37_2601 ();
 sg13g2_fill_2 FILLER_37_2615 ();
 sg13g2_decap_8 FILLER_37_2625 ();
 sg13g2_decap_4 FILLER_37_2640 ();
 sg13g2_fill_1 FILLER_37_2644 ();
 sg13g2_decap_8 FILLER_37_2696 ();
 sg13g2_fill_1 FILLER_37_2707 ();
 sg13g2_fill_2 FILLER_37_2721 ();
 sg13g2_fill_2 FILLER_37_2736 ();
 sg13g2_fill_1 FILLER_37_2738 ();
 sg13g2_fill_2 FILLER_37_2743 ();
 sg13g2_fill_1 FILLER_37_2745 ();
 sg13g2_fill_2 FILLER_37_2768 ();
 sg13g2_decap_8 FILLER_37_2807 ();
 sg13g2_fill_2 FILLER_37_2818 ();
 sg13g2_fill_2 FILLER_37_2832 ();
 sg13g2_fill_1 FILLER_37_2834 ();
 sg13g2_decap_8 FILLER_37_2840 ();
 sg13g2_decap_4 FILLER_37_2883 ();
 sg13g2_decap_4 FILLER_37_2900 ();
 sg13g2_fill_1 FILLER_37_2904 ();
 sg13g2_fill_2 FILLER_37_2922 ();
 sg13g2_fill_1 FILLER_37_2933 ();
 sg13g2_fill_1 FILLER_37_2939 ();
 sg13g2_fill_1 FILLER_37_2944 ();
 sg13g2_fill_1 FILLER_37_2963 ();
 sg13g2_fill_1 FILLER_37_3009 ();
 sg13g2_fill_1 FILLER_37_3033 ();
 sg13g2_fill_2 FILLER_37_3043 ();
 sg13g2_fill_1 FILLER_37_3045 ();
 sg13g2_fill_2 FILLER_37_3059 ();
 sg13g2_fill_1 FILLER_37_3090 ();
 sg13g2_decap_4 FILLER_37_3104 ();
 sg13g2_decap_8 FILLER_37_3136 ();
 sg13g2_fill_1 FILLER_37_3143 ();
 sg13g2_fill_2 FILLER_37_3163 ();
 sg13g2_decap_4 FILLER_37_3193 ();
 sg13g2_fill_1 FILLER_37_3197 ();
 sg13g2_decap_8 FILLER_37_3211 ();
 sg13g2_decap_8 FILLER_37_3218 ();
 sg13g2_fill_2 FILLER_37_3225 ();
 sg13g2_fill_1 FILLER_37_3227 ();
 sg13g2_fill_2 FILLER_37_3257 ();
 sg13g2_fill_1 FILLER_37_3259 ();
 sg13g2_fill_2 FILLER_37_3266 ();
 sg13g2_fill_1 FILLER_37_3268 ();
 sg13g2_decap_4 FILLER_37_3282 ();
 sg13g2_fill_2 FILLER_37_3299 ();
 sg13g2_fill_1 FILLER_37_3304 ();
 sg13g2_fill_1 FILLER_37_3314 ();
 sg13g2_decap_8 FILLER_37_3383 ();
 sg13g2_decap_4 FILLER_37_3390 ();
 sg13g2_fill_2 FILLER_37_3421 ();
 sg13g2_fill_1 FILLER_37_3423 ();
 sg13g2_fill_2 FILLER_37_3449 ();
 sg13g2_fill_1 FILLER_37_3451 ();
 sg13g2_fill_1 FILLER_37_3465 ();
 sg13g2_decap_8 FILLER_37_3525 ();
 sg13g2_decap_8 FILLER_37_3532 ();
 sg13g2_decap_8 FILLER_37_3539 ();
 sg13g2_decap_8 FILLER_37_3546 ();
 sg13g2_decap_8 FILLER_37_3553 ();
 sg13g2_decap_8 FILLER_37_3560 ();
 sg13g2_decap_8 FILLER_37_3567 ();
 sg13g2_decap_4 FILLER_37_3574 ();
 sg13g2_fill_2 FILLER_37_3578 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_fill_2 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_decap_8 FILLER_38_191 ();
 sg13g2_decap_4 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_217 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_259 ();
 sg13g2_decap_4 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_decap_4 FILLER_38_378 ();
 sg13g2_fill_2 FILLER_38_395 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_fill_1 FILLER_38_411 ();
 sg13g2_fill_2 FILLER_38_421 ();
 sg13g2_fill_1 FILLER_38_423 ();
 sg13g2_fill_1 FILLER_38_480 ();
 sg13g2_decap_4 FILLER_38_490 ();
 sg13g2_fill_2 FILLER_38_494 ();
 sg13g2_fill_2 FILLER_38_502 ();
 sg13g2_fill_1 FILLER_38_504 ();
 sg13g2_fill_2 FILLER_38_516 ();
 sg13g2_fill_1 FILLER_38_518 ();
 sg13g2_decap_8 FILLER_38_529 ();
 sg13g2_fill_1 FILLER_38_536 ();
 sg13g2_fill_2 FILLER_38_551 ();
 sg13g2_fill_2 FILLER_38_557 ();
 sg13g2_fill_1 FILLER_38_559 ();
 sg13g2_fill_2 FILLER_38_578 ();
 sg13g2_decap_4 FILLER_38_585 ();
 sg13g2_fill_1 FILLER_38_589 ();
 sg13g2_fill_1 FILLER_38_640 ();
 sg13g2_decap_4 FILLER_38_653 ();
 sg13g2_decap_4 FILLER_38_662 ();
 sg13g2_fill_1 FILLER_38_694 ();
 sg13g2_fill_1 FILLER_38_722 ();
 sg13g2_fill_1 FILLER_38_728 ();
 sg13g2_fill_1 FILLER_38_736 ();
 sg13g2_decap_8 FILLER_38_740 ();
 sg13g2_fill_1 FILLER_38_747 ();
 sg13g2_fill_1 FILLER_38_776 ();
 sg13g2_fill_2 FILLER_38_794 ();
 sg13g2_fill_1 FILLER_38_796 ();
 sg13g2_decap_4 FILLER_38_801 ();
 sg13g2_fill_2 FILLER_38_805 ();
 sg13g2_decap_4 FILLER_38_852 ();
 sg13g2_fill_2 FILLER_38_856 ();
 sg13g2_decap_8 FILLER_38_869 ();
 sg13g2_fill_2 FILLER_38_876 ();
 sg13g2_fill_1 FILLER_38_878 ();
 sg13g2_decap_8 FILLER_38_894 ();
 sg13g2_fill_1 FILLER_38_901 ();
 sg13g2_decap_8 FILLER_38_922 ();
 sg13g2_decap_4 FILLER_38_929 ();
 sg13g2_fill_1 FILLER_38_933 ();
 sg13g2_fill_1 FILLER_38_942 ();
 sg13g2_decap_8 FILLER_38_971 ();
 sg13g2_decap_4 FILLER_38_978 ();
 sg13g2_fill_2 FILLER_38_1001 ();
 sg13g2_fill_2 FILLER_38_1011 ();
 sg13g2_fill_2 FILLER_38_1017 ();
 sg13g2_fill_1 FILLER_38_1019 ();
 sg13g2_fill_2 FILLER_38_1037 ();
 sg13g2_fill_1 FILLER_38_1039 ();
 sg13g2_decap_4 FILLER_38_1058 ();
 sg13g2_fill_1 FILLER_38_1062 ();
 sg13g2_fill_2 FILLER_38_1076 ();
 sg13g2_fill_1 FILLER_38_1078 ();
 sg13g2_fill_2 FILLER_38_1088 ();
 sg13g2_fill_2 FILLER_38_1165 ();
 sg13g2_fill_1 FILLER_38_1193 ();
 sg13g2_decap_8 FILLER_38_1198 ();
 sg13g2_fill_1 FILLER_38_1205 ();
 sg13g2_fill_2 FILLER_38_1219 ();
 sg13g2_fill_1 FILLER_38_1221 ();
 sg13g2_fill_2 FILLER_38_1239 ();
 sg13g2_fill_1 FILLER_38_1241 ();
 sg13g2_fill_2 FILLER_38_1254 ();
 sg13g2_fill_1 FILLER_38_1256 ();
 sg13g2_fill_1 FILLER_38_1270 ();
 sg13g2_fill_1 FILLER_38_1302 ();
 sg13g2_decap_8 FILLER_38_1327 ();
 sg13g2_fill_1 FILLER_38_1334 ();
 sg13g2_decap_4 FILLER_38_1346 ();
 sg13g2_decap_8 FILLER_38_1382 ();
 sg13g2_fill_1 FILLER_38_1389 ();
 sg13g2_decap_8 FILLER_38_1396 ();
 sg13g2_decap_8 FILLER_38_1403 ();
 sg13g2_decap_4 FILLER_38_1410 ();
 sg13g2_fill_1 FILLER_38_1414 ();
 sg13g2_decap_4 FILLER_38_1436 ();
 sg13g2_decap_4 FILLER_38_1447 ();
 sg13g2_fill_1 FILLER_38_1451 ();
 sg13g2_decap_8 FILLER_38_1474 ();
 sg13g2_decap_4 FILLER_38_1481 ();
 sg13g2_fill_1 FILLER_38_1485 ();
 sg13g2_fill_2 FILLER_38_1496 ();
 sg13g2_fill_1 FILLER_38_1498 ();
 sg13g2_fill_1 FILLER_38_1507 ();
 sg13g2_fill_2 FILLER_38_1511 ();
 sg13g2_fill_1 FILLER_38_1513 ();
 sg13g2_fill_2 FILLER_38_1538 ();
 sg13g2_fill_1 FILLER_38_1540 ();
 sg13g2_decap_8 FILLER_38_1576 ();
 sg13g2_fill_1 FILLER_38_1583 ();
 sg13g2_decap_4 FILLER_38_1605 ();
 sg13g2_fill_1 FILLER_38_1609 ();
 sg13g2_decap_8 FILLER_38_1635 ();
 sg13g2_fill_2 FILLER_38_1642 ();
 sg13g2_decap_8 FILLER_38_1648 ();
 sg13g2_decap_8 FILLER_38_1655 ();
 sg13g2_fill_2 FILLER_38_1678 ();
 sg13g2_fill_1 FILLER_38_1706 ();
 sg13g2_decap_4 FILLER_38_1724 ();
 sg13g2_decap_8 FILLER_38_1736 ();
 sg13g2_fill_1 FILLER_38_1743 ();
 sg13g2_fill_2 FILLER_38_1748 ();
 sg13g2_decap_4 FILLER_38_1786 ();
 sg13g2_fill_2 FILLER_38_1790 ();
 sg13g2_decap_4 FILLER_38_1807 ();
 sg13g2_fill_2 FILLER_38_1811 ();
 sg13g2_decap_4 FILLER_38_1817 ();
 sg13g2_fill_1 FILLER_38_1821 ();
 sg13g2_decap_4 FILLER_38_1838 ();
 sg13g2_fill_2 FILLER_38_1842 ();
 sg13g2_fill_2 FILLER_38_1860 ();
 sg13g2_decap_8 FILLER_38_1875 ();
 sg13g2_fill_2 FILLER_38_1882 ();
 sg13g2_fill_1 FILLER_38_1884 ();
 sg13g2_decap_8 FILLER_38_1907 ();
 sg13g2_decap_4 FILLER_38_1914 ();
 sg13g2_fill_1 FILLER_38_1918 ();
 sg13g2_fill_2 FILLER_38_1932 ();
 sg13g2_fill_1 FILLER_38_1934 ();
 sg13g2_decap_8 FILLER_38_1957 ();
 sg13g2_fill_2 FILLER_38_1964 ();
 sg13g2_fill_1 FILLER_38_1966 ();
 sg13g2_fill_1 FILLER_38_2013 ();
 sg13g2_decap_4 FILLER_38_2034 ();
 sg13g2_fill_1 FILLER_38_2038 ();
 sg13g2_fill_1 FILLER_38_2047 ();
 sg13g2_decap_4 FILLER_38_2102 ();
 sg13g2_decap_8 FILLER_38_2124 ();
 sg13g2_decap_4 FILLER_38_2131 ();
 sg13g2_fill_2 FILLER_38_2135 ();
 sg13g2_fill_2 FILLER_38_2165 ();
 sg13g2_decap_8 FILLER_38_2203 ();
 sg13g2_fill_1 FILLER_38_2232 ();
 sg13g2_decap_8 FILLER_38_2249 ();
 sg13g2_decap_8 FILLER_38_2260 ();
 sg13g2_decap_8 FILLER_38_2267 ();
 sg13g2_fill_2 FILLER_38_2274 ();
 sg13g2_fill_1 FILLER_38_2276 ();
 sg13g2_fill_2 FILLER_38_2290 ();
 sg13g2_fill_2 FILLER_38_2318 ();
 sg13g2_fill_1 FILLER_38_2320 ();
 sg13g2_decap_4 FILLER_38_2350 ();
 sg13g2_fill_1 FILLER_38_2354 ();
 sg13g2_decap_8 FILLER_38_2363 ();
 sg13g2_fill_1 FILLER_38_2374 ();
 sg13g2_decap_8 FILLER_38_2379 ();
 sg13g2_fill_2 FILLER_38_2403 ();
 sg13g2_fill_1 FILLER_38_2405 ();
 sg13g2_decap_4 FILLER_38_2410 ();
 sg13g2_fill_2 FILLER_38_2414 ();
 sg13g2_decap_4 FILLER_38_2429 ();
 sg13g2_fill_2 FILLER_38_2441 ();
 sg13g2_fill_2 FILLER_38_2451 ();
 sg13g2_fill_2 FILLER_38_2474 ();
 sg13g2_fill_2 FILLER_38_2481 ();
 sg13g2_fill_1 FILLER_38_2483 ();
 sg13g2_decap_8 FILLER_38_2492 ();
 sg13g2_decap_4 FILLER_38_2499 ();
 sg13g2_decap_8 FILLER_38_2507 ();
 sg13g2_fill_1 FILLER_38_2514 ();
 sg13g2_fill_2 FILLER_38_2521 ();
 sg13g2_fill_1 FILLER_38_2523 ();
 sg13g2_decap_4 FILLER_38_2529 ();
 sg13g2_fill_1 FILLER_38_2533 ();
 sg13g2_decap_4 FILLER_38_2542 ();
 sg13g2_fill_2 FILLER_38_2546 ();
 sg13g2_decap_4 FILLER_38_2552 ();
 sg13g2_fill_1 FILLER_38_2556 ();
 sg13g2_fill_1 FILLER_38_2561 ();
 sg13g2_decap_8 FILLER_38_2579 ();
 sg13g2_fill_2 FILLER_38_2586 ();
 sg13g2_fill_1 FILLER_38_2598 ();
 sg13g2_decap_4 FILLER_38_2626 ();
 sg13g2_fill_1 FILLER_38_2630 ();
 sg13g2_fill_1 FILLER_38_2637 ();
 sg13g2_fill_1 FILLER_38_2651 ();
 sg13g2_decap_4 FILLER_38_2657 ();
 sg13g2_decap_8 FILLER_38_2669 ();
 sg13g2_decap_8 FILLER_38_2676 ();
 sg13g2_decap_8 FILLER_38_2697 ();
 sg13g2_decap_4 FILLER_38_2704 ();
 sg13g2_fill_2 FILLER_38_2721 ();
 sg13g2_fill_1 FILLER_38_2723 ();
 sg13g2_fill_2 FILLER_38_2733 ();
 sg13g2_fill_1 FILLER_38_2752 ();
 sg13g2_fill_2 FILLER_38_2761 ();
 sg13g2_fill_1 FILLER_38_2763 ();
 sg13g2_decap_8 FILLER_38_2772 ();
 sg13g2_fill_2 FILLER_38_2779 ();
 sg13g2_fill_1 FILLER_38_2794 ();
 sg13g2_fill_1 FILLER_38_2845 ();
 sg13g2_fill_1 FILLER_38_2853 ();
 sg13g2_decap_8 FILLER_38_2863 ();
 sg13g2_fill_1 FILLER_38_2870 ();
 sg13g2_decap_4 FILLER_38_2878 ();
 sg13g2_fill_2 FILLER_38_2882 ();
 sg13g2_decap_8 FILLER_38_2894 ();
 sg13g2_decap_8 FILLER_38_2901 ();
 sg13g2_fill_2 FILLER_38_2908 ();
 sg13g2_fill_1 FILLER_38_2910 ();
 sg13g2_fill_1 FILLER_38_2998 ();
 sg13g2_fill_2 FILLER_38_3011 ();
 sg13g2_fill_1 FILLER_38_3080 ();
 sg13g2_decap_4 FILLER_38_3095 ();
 sg13g2_fill_1 FILLER_38_3121 ();
 sg13g2_decap_8 FILLER_38_3130 ();
 sg13g2_decap_4 FILLER_38_3137 ();
 sg13g2_decap_4 FILLER_38_3158 ();
 sg13g2_fill_2 FILLER_38_3162 ();
 sg13g2_fill_2 FILLER_38_3173 ();
 sg13g2_decap_4 FILLER_38_3192 ();
 sg13g2_fill_1 FILLER_38_3196 ();
 sg13g2_fill_1 FILLER_38_3271 ();
 sg13g2_decap_8 FILLER_38_3300 ();
 sg13g2_decap_4 FILLER_38_3307 ();
 sg13g2_fill_2 FILLER_38_3332 ();
 sg13g2_fill_2 FILLER_38_3339 ();
 sg13g2_decap_8 FILLER_38_3346 ();
 sg13g2_decap_8 FILLER_38_3353 ();
 sg13g2_decap_4 FILLER_38_3360 ();
 sg13g2_decap_4 FILLER_38_3368 ();
 sg13g2_fill_2 FILLER_38_3372 ();
 sg13g2_decap_8 FILLER_38_3378 ();
 sg13g2_fill_1 FILLER_38_3385 ();
 sg13g2_decap_4 FILLER_38_3399 ();
 sg13g2_fill_1 FILLER_38_3403 ();
 sg13g2_fill_2 FILLER_38_3421 ();
 sg13g2_fill_2 FILLER_38_3446 ();
 sg13g2_fill_1 FILLER_38_3448 ();
 sg13g2_fill_2 FILLER_38_3458 ();
 sg13g2_fill_1 FILLER_38_3506 ();
 sg13g2_decap_8 FILLER_38_3516 ();
 sg13g2_decap_8 FILLER_38_3523 ();
 sg13g2_decap_8 FILLER_38_3530 ();
 sg13g2_decap_8 FILLER_38_3537 ();
 sg13g2_decap_8 FILLER_38_3544 ();
 sg13g2_decap_8 FILLER_38_3551 ();
 sg13g2_decap_8 FILLER_38_3558 ();
 sg13g2_decap_8 FILLER_38_3565 ();
 sg13g2_decap_8 FILLER_38_3572 ();
 sg13g2_fill_1 FILLER_38_3579 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_4 FILLER_39_105 ();
 sg13g2_fill_2 FILLER_39_109 ();
 sg13g2_fill_2 FILLER_39_138 ();
 sg13g2_fill_2 FILLER_39_162 ();
 sg13g2_decap_4 FILLER_39_168 ();
 sg13g2_fill_2 FILLER_39_172 ();
 sg13g2_fill_2 FILLER_39_179 ();
 sg13g2_fill_1 FILLER_39_181 ();
 sg13g2_decap_8 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_193 ();
 sg13g2_fill_1 FILLER_39_195 ();
 sg13g2_fill_2 FILLER_39_205 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_decap_4 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_247 ();
 sg13g2_fill_1 FILLER_39_283 ();
 sg13g2_decap_4 FILLER_39_302 ();
 sg13g2_fill_1 FILLER_39_306 ();
 sg13g2_decap_8 FILLER_39_327 ();
 sg13g2_decap_4 FILLER_39_334 ();
 sg13g2_fill_2 FILLER_39_343 ();
 sg13g2_fill_2 FILLER_39_367 ();
 sg13g2_fill_1 FILLER_39_369 ();
 sg13g2_fill_2 FILLER_39_431 ();
 sg13g2_fill_1 FILLER_39_433 ();
 sg13g2_fill_2 FILLER_39_439 ();
 sg13g2_decap_8 FILLER_39_466 ();
 sg13g2_decap_8 FILLER_39_473 ();
 sg13g2_decap_4 FILLER_39_480 ();
 sg13g2_fill_2 FILLER_39_520 ();
 sg13g2_decap_8 FILLER_39_527 ();
 sg13g2_decap_4 FILLER_39_534 ();
 sg13g2_fill_1 FILLER_39_544 ();
 sg13g2_fill_2 FILLER_39_558 ();
 sg13g2_fill_1 FILLER_39_573 ();
 sg13g2_fill_1 FILLER_39_635 ();
 sg13g2_fill_1 FILLER_39_641 ();
 sg13g2_fill_2 FILLER_39_662 ();
 sg13g2_fill_2 FILLER_39_669 ();
 sg13g2_fill_2 FILLER_39_693 ();
 sg13g2_fill_1 FILLER_39_695 ();
 sg13g2_fill_1 FILLER_39_710 ();
 sg13g2_decap_4 FILLER_39_747 ();
 sg13g2_fill_2 FILLER_39_751 ();
 sg13g2_decap_8 FILLER_39_757 ();
 sg13g2_decap_8 FILLER_39_764 ();
 sg13g2_fill_2 FILLER_39_771 ();
 sg13g2_fill_1 FILLER_39_773 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_fill_2 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_fill_2 FILLER_39_807 ();
 sg13g2_fill_2 FILLER_39_824 ();
 sg13g2_decap_8 FILLER_39_830 ();
 sg13g2_fill_2 FILLER_39_837 ();
 sg13g2_fill_1 FILLER_39_839 ();
 sg13g2_fill_1 FILLER_39_845 ();
 sg13g2_fill_2 FILLER_39_851 ();
 sg13g2_decap_4 FILLER_39_859 ();
 sg13g2_fill_1 FILLER_39_863 ();
 sg13g2_fill_1 FILLER_39_883 ();
 sg13g2_fill_2 FILLER_39_893 ();
 sg13g2_fill_1 FILLER_39_895 ();
 sg13g2_fill_1 FILLER_39_900 ();
 sg13g2_decap_8 FILLER_39_928 ();
 sg13g2_decap_4 FILLER_39_935 ();
 sg13g2_fill_2 FILLER_39_939 ();
 sg13g2_decap_8 FILLER_39_955 ();
 sg13g2_decap_8 FILLER_39_970 ();
 sg13g2_decap_4 FILLER_39_977 ();
 sg13g2_fill_2 FILLER_39_1006 ();
 sg13g2_decap_4 FILLER_39_1057 ();
 sg13g2_fill_2 FILLER_39_1061 ();
 sg13g2_fill_2 FILLER_39_1076 ();
 sg13g2_decap_8 FILLER_39_1092 ();
 sg13g2_fill_1 FILLER_39_1099 ();
 sg13g2_fill_2 FILLER_39_1113 ();
 sg13g2_fill_1 FILLER_39_1115 ();
 sg13g2_fill_2 FILLER_39_1125 ();
 sg13g2_decap_8 FILLER_39_1157 ();
 sg13g2_decap_4 FILLER_39_1164 ();
 sg13g2_decap_4 FILLER_39_1185 ();
 sg13g2_decap_8 FILLER_39_1239 ();
 sg13g2_decap_4 FILLER_39_1246 ();
 sg13g2_fill_1 FILLER_39_1250 ();
 sg13g2_decap_8 FILLER_39_1256 ();
 sg13g2_decap_8 FILLER_39_1263 ();
 sg13g2_fill_2 FILLER_39_1270 ();
 sg13g2_fill_1 FILLER_39_1272 ();
 sg13g2_fill_1 FILLER_39_1279 ();
 sg13g2_decap_8 FILLER_39_1288 ();
 sg13g2_decap_8 FILLER_39_1303 ();
 sg13g2_decap_4 FILLER_39_1310 ();
 sg13g2_fill_2 FILLER_39_1317 ();
 sg13g2_decap_8 FILLER_39_1324 ();
 sg13g2_decap_8 FILLER_39_1355 ();
 sg13g2_fill_2 FILLER_39_1362 ();
 sg13g2_fill_1 FILLER_39_1364 ();
 sg13g2_decap_8 FILLER_39_1406 ();
 sg13g2_fill_1 FILLER_39_1426 ();
 sg13g2_decap_8 FILLER_39_1452 ();
 sg13g2_fill_1 FILLER_39_1459 ();
 sg13g2_decap_8 FILLER_39_1468 ();
 sg13g2_fill_2 FILLER_39_1483 ();
 sg13g2_fill_1 FILLER_39_1485 ();
 sg13g2_decap_8 FILLER_39_1502 ();
 sg13g2_fill_1 FILLER_39_1509 ();
 sg13g2_decap_4 FILLER_39_1520 ();
 sg13g2_fill_2 FILLER_39_1524 ();
 sg13g2_fill_2 FILLER_39_1531 ();
 sg13g2_fill_2 FILLER_39_1542 ();
 sg13g2_fill_1 FILLER_39_1544 ();
 sg13g2_decap_4 FILLER_39_1564 ();
 sg13g2_fill_2 FILLER_39_1568 ();
 sg13g2_decap_4 FILLER_39_1610 ();
 sg13g2_fill_1 FILLER_39_1618 ();
 sg13g2_fill_2 FILLER_39_1632 ();
 sg13g2_fill_1 FILLER_39_1634 ();
 sg13g2_decap_4 FILLER_39_1640 ();
 sg13g2_decap_8 FILLER_39_1662 ();
 sg13g2_fill_2 FILLER_39_1669 ();
 sg13g2_fill_1 FILLER_39_1671 ();
 sg13g2_decap_4 FILLER_39_1694 ();
 sg13g2_fill_1 FILLER_39_1698 ();
 sg13g2_decap_4 FILLER_39_1704 ();
 sg13g2_decap_4 FILLER_39_1729 ();
 sg13g2_fill_2 FILLER_39_1733 ();
 sg13g2_decap_8 FILLER_39_1743 ();
 sg13g2_decap_4 FILLER_39_1750 ();
 sg13g2_fill_1 FILLER_39_1754 ();
 sg13g2_decap_8 FILLER_39_1759 ();
 sg13g2_decap_4 FILLER_39_1766 ();
 sg13g2_fill_1 FILLER_39_1770 ();
 sg13g2_decap_4 FILLER_39_1781 ();
 sg13g2_fill_2 FILLER_39_1785 ();
 sg13g2_fill_2 FILLER_39_1802 ();
 sg13g2_decap_8 FILLER_39_1816 ();
 sg13g2_decap_4 FILLER_39_1823 ();
 sg13g2_fill_1 FILLER_39_1827 ();
 sg13g2_decap_8 FILLER_39_1845 ();
 sg13g2_decap_4 FILLER_39_1852 ();
 sg13g2_fill_1 FILLER_39_1856 ();
 sg13g2_fill_2 FILLER_39_1863 ();
 sg13g2_decap_8 FILLER_39_1869 ();
 sg13g2_decap_8 FILLER_39_1876 ();
 sg13g2_fill_2 FILLER_39_1883 ();
 sg13g2_fill_1 FILLER_39_1910 ();
 sg13g2_decap_4 FILLER_39_1937 ();
 sg13g2_decap_4 FILLER_39_1972 ();
 sg13g2_fill_2 FILLER_39_1976 ();
 sg13g2_decap_8 FILLER_39_1989 ();
 sg13g2_fill_1 FILLER_39_1996 ();
 sg13g2_fill_1 FILLER_39_2001 ();
 sg13g2_decap_4 FILLER_39_2008 ();
 sg13g2_decap_8 FILLER_39_2045 ();
 sg13g2_decap_8 FILLER_39_2061 ();
 sg13g2_decap_8 FILLER_39_2068 ();
 sg13g2_decap_4 FILLER_39_2075 ();
 sg13g2_decap_8 FILLER_39_2083 ();
 sg13g2_fill_2 FILLER_39_2090 ();
 sg13g2_fill_1 FILLER_39_2092 ();
 sg13g2_fill_1 FILLER_39_2129 ();
 sg13g2_decap_8 FILLER_39_2133 ();
 sg13g2_decap_4 FILLER_39_2140 ();
 sg13g2_fill_2 FILLER_39_2149 ();
 sg13g2_fill_1 FILLER_39_2151 ();
 sg13g2_decap_8 FILLER_39_2156 ();
 sg13g2_decap_4 FILLER_39_2168 ();
 sg13g2_fill_1 FILLER_39_2172 ();
 sg13g2_decap_8 FILLER_39_2177 ();
 sg13g2_decap_8 FILLER_39_2184 ();
 sg13g2_decap_8 FILLER_39_2191 ();
 sg13g2_decap_8 FILLER_39_2211 ();
 sg13g2_decap_4 FILLER_39_2218 ();
 sg13g2_decap_8 FILLER_39_2236 ();
 sg13g2_decap_4 FILLER_39_2248 ();
 sg13g2_decap_4 FILLER_39_2291 ();
 sg13g2_fill_2 FILLER_39_2295 ();
 sg13g2_decap_8 FILLER_39_2327 ();
 sg13g2_fill_2 FILLER_39_2334 ();
 sg13g2_fill_1 FILLER_39_2336 ();
 sg13g2_decap_8 FILLER_39_2350 ();
 sg13g2_fill_2 FILLER_39_2357 ();
 sg13g2_fill_1 FILLER_39_2359 ();
 sg13g2_fill_2 FILLER_39_2368 ();
 sg13g2_fill_2 FILLER_39_2407 ();
 sg13g2_fill_1 FILLER_39_2409 ();
 sg13g2_fill_2 FILLER_39_2423 ();
 sg13g2_fill_1 FILLER_39_2425 ();
 sg13g2_fill_1 FILLER_39_2432 ();
 sg13g2_decap_8 FILLER_39_2448 ();
 sg13g2_fill_2 FILLER_39_2455 ();
 sg13g2_decap_4 FILLER_39_2483 ();
 sg13g2_fill_2 FILLER_39_2487 ();
 sg13g2_fill_2 FILLER_39_2506 ();
 sg13g2_fill_2 FILLER_39_2519 ();
 sg13g2_fill_1 FILLER_39_2521 ();
 sg13g2_decap_4 FILLER_39_2546 ();
 sg13g2_decap_4 FILLER_39_2577 ();
 sg13g2_fill_1 FILLER_39_2581 ();
 sg13g2_fill_1 FILLER_39_2590 ();
 sg13g2_fill_1 FILLER_39_2596 ();
 sg13g2_fill_2 FILLER_39_2608 ();
 sg13g2_fill_1 FILLER_39_2610 ();
 sg13g2_fill_2 FILLER_39_2619 ();
 sg13g2_fill_1 FILLER_39_2621 ();
 sg13g2_decap_8 FILLER_39_2630 ();
 sg13g2_decap_8 FILLER_39_2637 ();
 sg13g2_decap_4 FILLER_39_2644 ();
 sg13g2_fill_2 FILLER_39_2677 ();
 sg13g2_fill_1 FILLER_39_2679 ();
 sg13g2_decap_8 FILLER_39_2698 ();
 sg13g2_decap_4 FILLER_39_2705 ();
 sg13g2_fill_2 FILLER_39_2709 ();
 sg13g2_fill_1 FILLER_39_2728 ();
 sg13g2_fill_2 FILLER_39_2753 ();
 sg13g2_fill_1 FILLER_39_2755 ();
 sg13g2_fill_2 FILLER_39_2761 ();
 sg13g2_fill_1 FILLER_39_2763 ();
 sg13g2_fill_2 FILLER_39_2784 ();
 sg13g2_decap_8 FILLER_39_2812 ();
 sg13g2_fill_2 FILLER_39_2819 ();
 sg13g2_fill_2 FILLER_39_2829 ();
 sg13g2_fill_1 FILLER_39_2831 ();
 sg13g2_fill_1 FILLER_39_2848 ();
 sg13g2_decap_8 FILLER_39_2903 ();
 sg13g2_decap_4 FILLER_39_2918 ();
 sg13g2_fill_2 FILLER_39_2922 ();
 sg13g2_fill_2 FILLER_39_2937 ();
 sg13g2_fill_1 FILLER_39_2944 ();
 sg13g2_decap_8 FILLER_39_2953 ();
 sg13g2_decap_8 FILLER_39_2960 ();
 sg13g2_decap_8 FILLER_39_2967 ();
 sg13g2_decap_4 FILLER_39_2974 ();
 sg13g2_fill_2 FILLER_39_3018 ();
 sg13g2_fill_2 FILLER_39_3028 ();
 sg13g2_fill_2 FILLER_39_3047 ();
 sg13g2_decap_8 FILLER_39_3057 ();
 sg13g2_decap_8 FILLER_39_3064 ();
 sg13g2_fill_2 FILLER_39_3071 ();
 sg13g2_fill_1 FILLER_39_3080 ();
 sg13g2_fill_1 FILLER_39_3094 ();
 sg13g2_decap_8 FILLER_39_3143 ();
 sg13g2_fill_1 FILLER_39_3150 ();
 sg13g2_decap_8 FILLER_39_3170 ();
 sg13g2_decap_4 FILLER_39_3177 ();
 sg13g2_decap_4 FILLER_39_3189 ();
 sg13g2_fill_2 FILLER_39_3193 ();
 sg13g2_fill_2 FILLER_39_3200 ();
 sg13g2_decap_4 FILLER_39_3216 ();
 sg13g2_decap_4 FILLER_39_3230 ();
 sg13g2_fill_2 FILLER_39_3249 ();
 sg13g2_fill_1 FILLER_39_3251 ();
 sg13g2_fill_2 FILLER_39_3285 ();
 sg13g2_fill_2 FILLER_39_3295 ();
 sg13g2_fill_2 FILLER_39_3303 ();
 sg13g2_fill_1 FILLER_39_3305 ();
 sg13g2_fill_2 FILLER_39_3316 ();
 sg13g2_fill_2 FILLER_39_3323 ();
 sg13g2_fill_1 FILLER_39_3325 ();
 sg13g2_fill_1 FILLER_39_3373 ();
 sg13g2_fill_2 FILLER_39_3424 ();
 sg13g2_decap_8 FILLER_39_3443 ();
 sg13g2_fill_1 FILLER_39_3450 ();
 sg13g2_fill_2 FILLER_39_3461 ();
 sg13g2_fill_1 FILLER_39_3487 ();
 sg13g2_fill_2 FILLER_39_3497 ();
 sg13g2_decap_8 FILLER_39_3516 ();
 sg13g2_decap_8 FILLER_39_3523 ();
 sg13g2_decap_8 FILLER_39_3530 ();
 sg13g2_decap_8 FILLER_39_3537 ();
 sg13g2_decap_8 FILLER_39_3544 ();
 sg13g2_decap_8 FILLER_39_3551 ();
 sg13g2_decap_8 FILLER_39_3558 ();
 sg13g2_decap_8 FILLER_39_3565 ();
 sg13g2_decap_8 FILLER_39_3572 ();
 sg13g2_fill_1 FILLER_39_3579 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_fill_1 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_226 ();
 sg13g2_fill_2 FILLER_40_233 ();
 sg13g2_fill_1 FILLER_40_235 ();
 sg13g2_decap_8 FILLER_40_241 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_fill_2 FILLER_40_270 ();
 sg13g2_fill_1 FILLER_40_272 ();
 sg13g2_fill_1 FILLER_40_280 ();
 sg13g2_fill_2 FILLER_40_296 ();
 sg13g2_fill_2 FILLER_40_320 ();
 sg13g2_decap_8 FILLER_40_331 ();
 sg13g2_fill_2 FILLER_40_338 ();
 sg13g2_fill_1 FILLER_40_340 ();
 sg13g2_fill_2 FILLER_40_381 ();
 sg13g2_fill_2 FILLER_40_419 ();
 sg13g2_fill_1 FILLER_40_421 ();
 sg13g2_decap_4 FILLER_40_506 ();
 sg13g2_decap_8 FILLER_40_580 ();
 sg13g2_decap_4 FILLER_40_587 ();
 sg13g2_fill_2 FILLER_40_596 ();
 sg13g2_fill_1 FILLER_40_598 ();
 sg13g2_fill_2 FILLER_40_611 ();
 sg13g2_decap_8 FILLER_40_631 ();
 sg13g2_decap_8 FILLER_40_638 ();
 sg13g2_decap_4 FILLER_40_645 ();
 sg13g2_fill_2 FILLER_40_653 ();
 sg13g2_decap_8 FILLER_40_664 ();
 sg13g2_fill_1 FILLER_40_671 ();
 sg13g2_fill_2 FILLER_40_699 ();
 sg13g2_fill_1 FILLER_40_701 ();
 sg13g2_decap_8 FILLER_40_746 ();
 sg13g2_fill_2 FILLER_40_796 ();
 sg13g2_fill_2 FILLER_40_832 ();
 sg13g2_fill_1 FILLER_40_863 ();
 sg13g2_decap_4 FILLER_40_882 ();
 sg13g2_decap_8 FILLER_40_905 ();
 sg13g2_fill_1 FILLER_40_912 ();
 sg13g2_decap_8 FILLER_40_922 ();
 sg13g2_decap_4 FILLER_40_929 ();
 sg13g2_fill_1 FILLER_40_950 ();
 sg13g2_decap_8 FILLER_40_977 ();
 sg13g2_fill_2 FILLER_40_1023 ();
 sg13g2_fill_2 FILLER_40_1043 ();
 sg13g2_fill_1 FILLER_40_1045 ();
 sg13g2_decap_8 FILLER_40_1059 ();
 sg13g2_decap_8 FILLER_40_1066 ();
 sg13g2_decap_8 FILLER_40_1073 ();
 sg13g2_fill_1 FILLER_40_1107 ();
 sg13g2_fill_2 FILLER_40_1126 ();
 sg13g2_fill_1 FILLER_40_1128 ();
 sg13g2_fill_2 FILLER_40_1169 ();
 sg13g2_fill_1 FILLER_40_1171 ();
 sg13g2_fill_2 FILLER_40_1200 ();
 sg13g2_fill_1 FILLER_40_1202 ();
 sg13g2_decap_4 FILLER_40_1216 ();
 sg13g2_fill_1 FILLER_40_1220 ();
 sg13g2_fill_2 FILLER_40_1244 ();
 sg13g2_fill_1 FILLER_40_1246 ();
 sg13g2_decap_8 FILLER_40_1264 ();
 sg13g2_fill_1 FILLER_40_1271 ();
 sg13g2_decap_8 FILLER_40_1297 ();
 sg13g2_fill_1 FILLER_40_1304 ();
 sg13g2_decap_4 FILLER_40_1327 ();
 sg13g2_fill_1 FILLER_40_1331 ();
 sg13g2_fill_2 FILLER_40_1337 ();
 sg13g2_decap_8 FILLER_40_1348 ();
 sg13g2_decap_4 FILLER_40_1355 ();
 sg13g2_fill_1 FILLER_40_1359 ();
 sg13g2_fill_2 FILLER_40_1377 ();
 sg13g2_fill_1 FILLER_40_1379 ();
 sg13g2_decap_8 FILLER_40_1385 ();
 sg13g2_fill_2 FILLER_40_1397 ();
 sg13g2_fill_1 FILLER_40_1399 ();
 sg13g2_decap_8 FILLER_40_1409 ();
 sg13g2_decap_8 FILLER_40_1416 ();
 sg13g2_decap_4 FILLER_40_1423 ();
 sg13g2_fill_1 FILLER_40_1427 ();
 sg13g2_fill_1 FILLER_40_1441 ();
 sg13g2_fill_1 FILLER_40_1472 ();
 sg13g2_fill_2 FILLER_40_1489 ();
 sg13g2_decap_8 FILLER_40_1507 ();
 sg13g2_fill_2 FILLER_40_1514 ();
 sg13g2_decap_4 FILLER_40_1520 ();
 sg13g2_decap_8 FILLER_40_1559 ();
 sg13g2_fill_1 FILLER_40_1566 ();
 sg13g2_decap_4 FILLER_40_1590 ();
 sg13g2_decap_8 FILLER_40_1606 ();
 sg13g2_decap_4 FILLER_40_1613 ();
 sg13g2_fill_2 FILLER_40_1617 ();
 sg13g2_fill_2 FILLER_40_1627 ();
 sg13g2_fill_2 FILLER_40_1683 ();
 sg13g2_decap_4 FILLER_40_1712 ();
 sg13g2_decap_4 FILLER_40_1725 ();
 sg13g2_decap_8 FILLER_40_1741 ();
 sg13g2_fill_1 FILLER_40_1748 ();
 sg13g2_decap_4 FILLER_40_1771 ();
 sg13g2_fill_2 FILLER_40_1791 ();
 sg13g2_decap_8 FILLER_40_1821 ();
 sg13g2_fill_2 FILLER_40_1828 ();
 sg13g2_fill_1 FILLER_40_1830 ();
 sg13g2_decap_8 FILLER_40_1852 ();
 sg13g2_fill_2 FILLER_40_1859 ();
 sg13g2_decap_8 FILLER_40_1887 ();
 sg13g2_decap_4 FILLER_40_1894 ();
 sg13g2_fill_1 FILLER_40_1898 ();
 sg13g2_decap_8 FILLER_40_1912 ();
 sg13g2_decap_4 FILLER_40_1919 ();
 sg13g2_fill_1 FILLER_40_1923 ();
 sg13g2_decap_8 FILLER_40_1937 ();
 sg13g2_fill_2 FILLER_40_1944 ();
 sg13g2_decap_8 FILLER_40_1962 ();
 sg13g2_fill_2 FILLER_40_1969 ();
 sg13g2_fill_1 FILLER_40_1971 ();
 sg13g2_fill_1 FILLER_40_1997 ();
 sg13g2_decap_4 FILLER_40_2017 ();
 sg13g2_fill_2 FILLER_40_2021 ();
 sg13g2_fill_1 FILLER_40_2055 ();
 sg13g2_decap_4 FILLER_40_2077 ();
 sg13g2_fill_2 FILLER_40_2081 ();
 sg13g2_fill_2 FILLER_40_2131 ();
 sg13g2_decap_8 FILLER_40_2181 ();
 sg13g2_decap_4 FILLER_40_2188 ();
 sg13g2_fill_2 FILLER_40_2192 ();
 sg13g2_fill_2 FILLER_40_2221 ();
 sg13g2_fill_1 FILLER_40_2223 ();
 sg13g2_decap_8 FILLER_40_2290 ();
 sg13g2_fill_2 FILLER_40_2297 ();
 sg13g2_decap_8 FILLER_40_2331 ();
 sg13g2_fill_1 FILLER_40_2338 ();
 sg13g2_fill_2 FILLER_40_2347 ();
 sg13g2_decap_8 FILLER_40_2371 ();
 sg13g2_fill_2 FILLER_40_2378 ();
 sg13g2_fill_1 FILLER_40_2380 ();
 sg13g2_fill_2 FILLER_40_2395 ();
 sg13g2_fill_1 FILLER_40_2397 ();
 sg13g2_decap_4 FILLER_40_2423 ();
 sg13g2_decap_8 FILLER_40_2453 ();
 sg13g2_fill_2 FILLER_40_2460 ();
 sg13g2_decap_4 FILLER_40_2486 ();
 sg13g2_decap_4 FILLER_40_2498 ();
 sg13g2_fill_1 FILLER_40_2502 ();
 sg13g2_fill_2 FILLER_40_2529 ();
 sg13g2_decap_4 FILLER_40_2585 ();
 sg13g2_fill_2 FILLER_40_2589 ();
 sg13g2_fill_2 FILLER_40_2614 ();
 sg13g2_decap_4 FILLER_40_2624 ();
 sg13g2_decap_4 FILLER_40_2641 ();
 sg13g2_fill_2 FILLER_40_2645 ();
 sg13g2_fill_2 FILLER_40_2655 ();
 sg13g2_decap_8 FILLER_40_2666 ();
 sg13g2_decap_4 FILLER_40_2673 ();
 sg13g2_decap_8 FILLER_40_2698 ();
 sg13g2_fill_1 FILLER_40_2705 ();
 sg13g2_decap_4 FILLER_40_2732 ();
 sg13g2_fill_2 FILLER_40_2762 ();
 sg13g2_fill_1 FILLER_40_2764 ();
 sg13g2_fill_2 FILLER_40_2780 ();
 sg13g2_decap_8 FILLER_40_2811 ();
 sg13g2_fill_2 FILLER_40_2818 ();
 sg13g2_fill_2 FILLER_40_2824 ();
 sg13g2_fill_1 FILLER_40_2826 ();
 sg13g2_fill_1 FILLER_40_2840 ();
 sg13g2_fill_2 FILLER_40_2863 ();
 sg13g2_fill_1 FILLER_40_2873 ();
 sg13g2_decap_4 FILLER_40_2896 ();
 sg13g2_fill_1 FILLER_40_2900 ();
 sg13g2_fill_2 FILLER_40_2910 ();
 sg13g2_fill_1 FILLER_40_2935 ();
 sg13g2_fill_2 FILLER_40_2953 ();
 sg13g2_fill_1 FILLER_40_2955 ();
 sg13g2_fill_2 FILLER_40_2960 ();
 sg13g2_fill_2 FILLER_40_2971 ();
 sg13g2_decap_4 FILLER_40_3001 ();
 sg13g2_decap_4 FILLER_40_3024 ();
 sg13g2_fill_2 FILLER_40_3098 ();
 sg13g2_fill_1 FILLER_40_3100 ();
 sg13g2_decap_8 FILLER_40_3113 ();
 sg13g2_fill_1 FILLER_40_3120 ();
 sg13g2_fill_1 FILLER_40_3125 ();
 sg13g2_decap_4 FILLER_40_3132 ();
 sg13g2_decap_8 FILLER_40_3142 ();
 sg13g2_decap_8 FILLER_40_3149 ();
 sg13g2_fill_2 FILLER_40_3156 ();
 sg13g2_decap_4 FILLER_40_3172 ();
 sg13g2_fill_1 FILLER_40_3176 ();
 sg13g2_fill_2 FILLER_40_3200 ();
 sg13g2_fill_2 FILLER_40_3209 ();
 sg13g2_decap_4 FILLER_40_3226 ();
 sg13g2_fill_2 FILLER_40_3241 ();
 sg13g2_fill_1 FILLER_40_3243 ();
 sg13g2_decap_4 FILLER_40_3249 ();
 sg13g2_fill_2 FILLER_40_3253 ();
 sg13g2_decap_8 FILLER_40_3265 ();
 sg13g2_decap_4 FILLER_40_3272 ();
 sg13g2_decap_4 FILLER_40_3298 ();
 sg13g2_fill_1 FILLER_40_3302 ();
 sg13g2_decap_8 FILLER_40_3308 ();
 sg13g2_decap_8 FILLER_40_3315 ();
 sg13g2_fill_1 FILLER_40_3322 ();
 sg13g2_decap_8 FILLER_40_3346 ();
 sg13g2_decap_8 FILLER_40_3366 ();
 sg13g2_decap_8 FILLER_40_3373 ();
 sg13g2_decap_8 FILLER_40_3380 ();
 sg13g2_decap_4 FILLER_40_3387 ();
 sg13g2_fill_1 FILLER_40_3391 ();
 sg13g2_decap_4 FILLER_40_3396 ();
 sg13g2_fill_2 FILLER_40_3400 ();
 sg13g2_fill_1 FILLER_40_3411 ();
 sg13g2_decap_8 FILLER_40_3443 ();
 sg13g2_decap_8 FILLER_40_3450 ();
 sg13g2_decap_4 FILLER_40_3457 ();
 sg13g2_fill_1 FILLER_40_3461 ();
 sg13g2_decap_4 FILLER_40_3490 ();
 sg13g2_decap_8 FILLER_40_3522 ();
 sg13g2_decap_8 FILLER_40_3529 ();
 sg13g2_decap_8 FILLER_40_3536 ();
 sg13g2_decap_8 FILLER_40_3543 ();
 sg13g2_decap_8 FILLER_40_3550 ();
 sg13g2_decap_8 FILLER_40_3557 ();
 sg13g2_decap_8 FILLER_40_3564 ();
 sg13g2_decap_8 FILLER_40_3571 ();
 sg13g2_fill_2 FILLER_40_3578 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_4 FILLER_41_119 ();
 sg13g2_fill_1 FILLER_41_123 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_fill_2 FILLER_41_152 ();
 sg13g2_fill_1 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_173 ();
 sg13g2_decap_4 FILLER_41_229 ();
 sg13g2_fill_1 FILLER_41_233 ();
 sg13g2_fill_2 FILLER_41_264 ();
 sg13g2_fill_1 FILLER_41_279 ();
 sg13g2_fill_2 FILLER_41_320 ();
 sg13g2_fill_1 FILLER_41_358 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_430 ();
 sg13g2_fill_2 FILLER_41_437 ();
 sg13g2_decap_8 FILLER_41_452 ();
 sg13g2_fill_2 FILLER_41_459 ();
 sg13g2_fill_1 FILLER_41_461 ();
 sg13g2_fill_2 FILLER_41_475 ();
 sg13g2_fill_1 FILLER_41_509 ();
 sg13g2_fill_2 FILLER_41_562 ();
 sg13g2_fill_1 FILLER_41_564 ();
 sg13g2_fill_2 FILLER_41_574 ();
 sg13g2_fill_1 FILLER_41_576 ();
 sg13g2_fill_2 FILLER_41_608 ();
 sg13g2_decap_4 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_740 ();
 sg13g2_fill_1 FILLER_41_747 ();
 sg13g2_decap_8 FILLER_41_762 ();
 sg13g2_decap_4 FILLER_41_769 ();
 sg13g2_fill_1 FILLER_41_773 ();
 sg13g2_fill_2 FILLER_41_778 ();
 sg13g2_fill_1 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_4 FILLER_41_805 ();
 sg13g2_fill_2 FILLER_41_809 ();
 sg13g2_fill_2 FILLER_41_816 ();
 sg13g2_fill_1 FILLER_41_823 ();
 sg13g2_decap_8 FILLER_41_837 ();
 sg13g2_fill_2 FILLER_41_844 ();
 sg13g2_fill_1 FILLER_41_846 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_4 FILLER_41_868 ();
 sg13g2_fill_2 FILLER_41_872 ();
 sg13g2_fill_2 FILLER_41_887 ();
 sg13g2_decap_8 FILLER_41_902 ();
 sg13g2_fill_2 FILLER_41_925 ();
 sg13g2_fill_1 FILLER_41_927 ();
 sg13g2_fill_1 FILLER_41_946 ();
 sg13g2_decap_4 FILLER_41_952 ();
 sg13g2_fill_2 FILLER_41_956 ();
 sg13g2_fill_2 FILLER_41_1004 ();
 sg13g2_fill_1 FILLER_41_1006 ();
 sg13g2_fill_2 FILLER_41_1034 ();
 sg13g2_decap_4 FILLER_41_1067 ();
 sg13g2_fill_2 FILLER_41_1098 ();
 sg13g2_fill_1 FILLER_41_1104 ();
 sg13g2_fill_2 FILLER_41_1110 ();
 sg13g2_decap_8 FILLER_41_1134 ();
 sg13g2_fill_1 FILLER_41_1150 ();
 sg13g2_fill_2 FILLER_41_1203 ();
 sg13g2_fill_1 FILLER_41_1231 ();
 sg13g2_fill_2 FILLER_41_1248 ();
 sg13g2_decap_4 FILLER_41_1255 ();
 sg13g2_decap_8 FILLER_41_1267 ();
 sg13g2_fill_2 FILLER_41_1282 ();
 sg13g2_decap_4 FILLER_41_1306 ();
 sg13g2_fill_2 FILLER_41_1334 ();
 sg13g2_fill_2 FILLER_41_1349 ();
 sg13g2_fill_2 FILLER_41_1356 ();
 sg13g2_fill_2 FILLER_41_1389 ();
 sg13g2_fill_2 FILLER_41_1411 ();
 sg13g2_decap_8 FILLER_41_1433 ();
 sg13g2_decap_8 FILLER_41_1440 ();
 sg13g2_fill_2 FILLER_41_1447 ();
 sg13g2_fill_1 FILLER_41_1449 ();
 sg13g2_fill_1 FILLER_41_1463 ();
 sg13g2_fill_2 FILLER_41_1477 ();
 sg13g2_decap_4 FILLER_41_1492 ();
 sg13g2_fill_2 FILLER_41_1496 ();
 sg13g2_fill_2 FILLER_41_1503 ();
 sg13g2_fill_1 FILLER_41_1505 ();
 sg13g2_decap_8 FILLER_41_1511 ();
 sg13g2_fill_2 FILLER_41_1522 ();
 sg13g2_fill_1 FILLER_41_1524 ();
 sg13g2_fill_2 FILLER_41_1539 ();
 sg13g2_fill_1 FILLER_41_1541 ();
 sg13g2_decap_4 FILLER_41_1565 ();
 sg13g2_decap_4 FILLER_41_1573 ();
 sg13g2_fill_1 FILLER_41_1577 ();
 sg13g2_fill_1 FILLER_41_1587 ();
 sg13g2_fill_1 FILLER_41_1598 ();
 sg13g2_fill_1 FILLER_41_1611 ();
 sg13g2_fill_1 FILLER_41_1621 ();
 sg13g2_decap_8 FILLER_41_1653 ();
 sg13g2_decap_8 FILLER_41_1660 ();
 sg13g2_decap_8 FILLER_41_1667 ();
 sg13g2_fill_1 FILLER_41_1674 ();
 sg13g2_fill_1 FILLER_41_1679 ();
 sg13g2_fill_2 FILLER_41_1689 ();
 sg13g2_decap_8 FILLER_41_1732 ();
 sg13g2_decap_4 FILLER_41_1739 ();
 sg13g2_decap_4 FILLER_41_1769 ();
 sg13g2_fill_2 FILLER_41_1773 ();
 sg13g2_fill_2 FILLER_41_1796 ();
 sg13g2_fill_1 FILLER_41_1798 ();
 sg13g2_fill_2 FILLER_41_1804 ();
 sg13g2_fill_1 FILLER_41_1806 ();
 sg13g2_decap_8 FILLER_41_1815 ();
 sg13g2_decap_4 FILLER_41_1847 ();
 sg13g2_fill_2 FILLER_41_1851 ();
 sg13g2_fill_1 FILLER_41_1869 ();
 sg13g2_fill_2 FILLER_41_1874 ();
 sg13g2_fill_2 FILLER_41_1894 ();
 sg13g2_fill_1 FILLER_41_1896 ();
 sg13g2_decap_8 FILLER_41_1938 ();
 sg13g2_decap_8 FILLER_41_1950 ();
 sg13g2_fill_2 FILLER_41_1957 ();
 sg13g2_fill_1 FILLER_41_1959 ();
 sg13g2_decap_4 FILLER_41_1964 ();
 sg13g2_fill_1 FILLER_41_1968 ();
 sg13g2_fill_1 FILLER_41_1983 ();
 sg13g2_fill_2 FILLER_41_1988 ();
 sg13g2_fill_1 FILLER_41_1990 ();
 sg13g2_fill_1 FILLER_41_2005 ();
 sg13g2_decap_4 FILLER_41_2044 ();
 sg13g2_decap_8 FILLER_41_2071 ();
 sg13g2_fill_1 FILLER_41_2078 ();
 sg13g2_fill_2 FILLER_41_2101 ();
 sg13g2_fill_1 FILLER_41_2103 ();
 sg13g2_decap_8 FILLER_41_2130 ();
 sg13g2_decap_4 FILLER_41_2137 ();
 sg13g2_fill_1 FILLER_41_2141 ();
 sg13g2_fill_2 FILLER_41_2152 ();
 sg13g2_fill_1 FILLER_41_2154 ();
 sg13g2_fill_1 FILLER_41_2159 ();
 sg13g2_decap_8 FILLER_41_2177 ();
 sg13g2_fill_2 FILLER_41_2184 ();
 sg13g2_fill_1 FILLER_41_2186 ();
 sg13g2_fill_2 FILLER_41_2236 ();
 sg13g2_decap_8 FILLER_41_2251 ();
 sg13g2_fill_2 FILLER_41_2294 ();
 sg13g2_fill_2 FILLER_41_2300 ();
 sg13g2_fill_1 FILLER_41_2302 ();
 sg13g2_fill_2 FILLER_41_2316 ();
 sg13g2_fill_1 FILLER_41_2332 ();
 sg13g2_fill_2 FILLER_41_2402 ();
 sg13g2_fill_1 FILLER_41_2404 ();
 sg13g2_fill_2 FILLER_41_2424 ();
 sg13g2_decap_4 FILLER_41_2443 ();
 sg13g2_decap_8 FILLER_41_2451 ();
 sg13g2_fill_1 FILLER_41_2471 ();
 sg13g2_decap_8 FILLER_41_2480 ();
 sg13g2_decap_8 FILLER_41_2487 ();
 sg13g2_decap_8 FILLER_41_2494 ();
 sg13g2_fill_1 FILLER_41_2501 ();
 sg13g2_fill_1 FILLER_41_2520 ();
 sg13g2_decap_8 FILLER_41_2535 ();
 sg13g2_decap_4 FILLER_41_2542 ();
 sg13g2_fill_1 FILLER_41_2546 ();
 sg13g2_decap_8 FILLER_41_2556 ();
 sg13g2_fill_1 FILLER_41_2563 ();
 sg13g2_decap_4 FILLER_41_2568 ();
 sg13g2_fill_1 FILLER_41_2572 ();
 sg13g2_decap_8 FILLER_41_2578 ();
 sg13g2_decap_4 FILLER_41_2585 ();
 sg13g2_fill_1 FILLER_41_2589 ();
 sg13g2_decap_4 FILLER_41_2630 ();
 sg13g2_fill_1 FILLER_41_2634 ();
 sg13g2_decap_8 FILLER_41_2644 ();
 sg13g2_fill_2 FILLER_41_2651 ();
 sg13g2_fill_1 FILLER_41_2653 ();
 sg13g2_fill_2 FILLER_41_2670 ();
 sg13g2_fill_1 FILLER_41_2672 ();
 sg13g2_fill_1 FILLER_41_2678 ();
 sg13g2_fill_2 FILLER_41_2701 ();
 sg13g2_fill_1 FILLER_41_2703 ();
 sg13g2_decap_8 FILLER_41_2746 ();
 sg13g2_decap_4 FILLER_41_2753 ();
 sg13g2_fill_1 FILLER_41_2757 ();
 sg13g2_decap_8 FILLER_41_2776 ();
 sg13g2_fill_2 FILLER_41_2783 ();
 sg13g2_fill_1 FILLER_41_2785 ();
 sg13g2_decap_8 FILLER_41_2804 ();
 sg13g2_decap_4 FILLER_41_2811 ();
 sg13g2_fill_2 FILLER_41_2868 ();
 sg13g2_decap_8 FILLER_41_2918 ();
 sg13g2_decap_4 FILLER_41_2925 ();
 sg13g2_fill_2 FILLER_41_2929 ();
 sg13g2_decap_8 FILLER_41_2937 ();
 sg13g2_decap_4 FILLER_41_2944 ();
 sg13g2_fill_2 FILLER_41_2948 ();
 sg13g2_fill_2 FILLER_41_2978 ();
 sg13g2_decap_4 FILLER_41_2993 ();
 sg13g2_fill_1 FILLER_41_2997 ();
 sg13g2_fill_1 FILLER_41_3004 ();
 sg13g2_decap_8 FILLER_41_3019 ();
 sg13g2_decap_8 FILLER_41_3026 ();
 sg13g2_decap_4 FILLER_41_3033 ();
 sg13g2_fill_1 FILLER_41_3044 ();
 sg13g2_decap_8 FILLER_41_3050 ();
 sg13g2_decap_4 FILLER_41_3057 ();
 sg13g2_decap_4 FILLER_41_3065 ();
 sg13g2_fill_2 FILLER_41_3077 ();
 sg13g2_decap_8 FILLER_41_3106 ();
 sg13g2_fill_2 FILLER_41_3113 ();
 sg13g2_fill_1 FILLER_41_3115 ();
 sg13g2_fill_2 FILLER_41_3129 ();
 sg13g2_fill_1 FILLER_41_3131 ();
 sg13g2_fill_1 FILLER_41_3135 ();
 sg13g2_fill_1 FILLER_41_3144 ();
 sg13g2_fill_2 FILLER_41_3174 ();
 sg13g2_decap_4 FILLER_41_3190 ();
 sg13g2_fill_1 FILLER_41_3194 ();
 sg13g2_fill_2 FILLER_41_3224 ();
 sg13g2_fill_2 FILLER_41_3233 ();
 sg13g2_fill_1 FILLER_41_3261 ();
 sg13g2_fill_2 FILLER_41_3270 ();
 sg13g2_fill_1 FILLER_41_3272 ();
 sg13g2_fill_2 FILLER_41_3294 ();
 sg13g2_decap_8 FILLER_41_3315 ();
 sg13g2_fill_1 FILLER_41_3335 ();
 sg13g2_fill_1 FILLER_41_3357 ();
 sg13g2_decap_8 FILLER_41_3363 ();
 sg13g2_decap_4 FILLER_41_3370 ();
 sg13g2_fill_1 FILLER_41_3374 ();
 sg13g2_fill_1 FILLER_41_3384 ();
 sg13g2_fill_2 FILLER_41_3427 ();
 sg13g2_fill_1 FILLER_41_3429 ();
 sg13g2_fill_2 FILLER_41_3440 ();
 sg13g2_decap_4 FILLER_41_3447 ();
 sg13g2_fill_2 FILLER_41_3451 ();
 sg13g2_decap_4 FILLER_41_3459 ();
 sg13g2_fill_1 FILLER_41_3474 ();
 sg13g2_decap_8 FILLER_41_3479 ();
 sg13g2_decap_8 FILLER_41_3486 ();
 sg13g2_fill_1 FILLER_41_3493 ();
 sg13g2_decap_8 FILLER_41_3503 ();
 sg13g2_decap_8 FILLER_41_3510 ();
 sg13g2_decap_8 FILLER_41_3517 ();
 sg13g2_decap_8 FILLER_41_3524 ();
 sg13g2_decap_8 FILLER_41_3531 ();
 sg13g2_decap_8 FILLER_41_3538 ();
 sg13g2_decap_8 FILLER_41_3545 ();
 sg13g2_decap_8 FILLER_41_3552 ();
 sg13g2_decap_8 FILLER_41_3559 ();
 sg13g2_decap_8 FILLER_41_3566 ();
 sg13g2_decap_8 FILLER_41_3573 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_4 FILLER_42_105 ();
 sg13g2_fill_2 FILLER_42_136 ();
 sg13g2_fill_2 FILLER_42_196 ();
 sg13g2_decap_4 FILLER_42_214 ();
 sg13g2_fill_2 FILLER_42_218 ();
 sg13g2_decap_8 FILLER_42_225 ();
 sg13g2_fill_2 FILLER_42_232 ();
 sg13g2_fill_1 FILLER_42_234 ();
 sg13g2_decap_8 FILLER_42_302 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_fill_1 FILLER_42_317 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_fill_2 FILLER_42_342 ();
 sg13g2_fill_1 FILLER_42_418 ();
 sg13g2_fill_2 FILLER_42_428 ();
 sg13g2_fill_1 FILLER_42_430 ();
 sg13g2_fill_2 FILLER_42_469 ();
 sg13g2_fill_2 FILLER_42_485 ();
 sg13g2_fill_2 FILLER_42_500 ();
 sg13g2_fill_1 FILLER_42_502 ();
 sg13g2_fill_2 FILLER_42_539 ();
 sg13g2_fill_1 FILLER_42_541 ();
 sg13g2_fill_2 FILLER_42_574 ();
 sg13g2_fill_2 FILLER_42_608 ();
 sg13g2_fill_1 FILLER_42_624 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_fill_2 FILLER_42_651 ();
 sg13g2_fill_1 FILLER_42_653 ();
 sg13g2_decap_4 FILLER_42_668 ();
 sg13g2_fill_1 FILLER_42_672 ();
 sg13g2_fill_2 FILLER_42_719 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_fill_2 FILLER_42_812 ();
 sg13g2_decap_4 FILLER_42_840 ();
 sg13g2_fill_2 FILLER_42_849 ();
 sg13g2_decap_8 FILLER_42_856 ();
 sg13g2_fill_2 FILLER_42_863 ();
 sg13g2_fill_1 FILLER_42_865 ();
 sg13g2_decap_8 FILLER_42_871 ();
 sg13g2_decap_4 FILLER_42_878 ();
 sg13g2_fill_1 FILLER_42_882 ();
 sg13g2_decap_8 FILLER_42_896 ();
 sg13g2_decap_8 FILLER_42_903 ();
 sg13g2_decap_8 FILLER_42_926 ();
 sg13g2_fill_2 FILLER_42_933 ();
 sg13g2_decap_8 FILLER_42_941 ();
 sg13g2_decap_8 FILLER_42_948 ();
 sg13g2_decap_8 FILLER_42_955 ();
 sg13g2_decap_4 FILLER_42_962 ();
 sg13g2_fill_2 FILLER_42_966 ();
 sg13g2_decap_4 FILLER_42_1018 ();
 sg13g2_fill_2 FILLER_42_1027 ();
 sg13g2_fill_1 FILLER_42_1029 ();
 sg13g2_fill_2 FILLER_42_1035 ();
 sg13g2_fill_1 FILLER_42_1037 ();
 sg13g2_fill_2 FILLER_42_1043 ();
 sg13g2_fill_2 FILLER_42_1113 ();
 sg13g2_decap_8 FILLER_42_1142 ();
 sg13g2_decap_4 FILLER_42_1149 ();
 sg13g2_fill_2 FILLER_42_1153 ();
 sg13g2_fill_2 FILLER_42_1177 ();
 sg13g2_fill_2 FILLER_42_1199 ();
 sg13g2_decap_4 FILLER_42_1206 ();
 sg13g2_fill_2 FILLER_42_1210 ();
 sg13g2_fill_2 FILLER_42_1225 ();
 sg13g2_fill_2 FILLER_42_1272 ();
 sg13g2_fill_1 FILLER_42_1274 ();
 sg13g2_decap_4 FILLER_42_1280 ();
 sg13g2_decap_4 FILLER_42_1288 ();
 sg13g2_fill_2 FILLER_42_1297 ();
 sg13g2_fill_1 FILLER_42_1299 ();
 sg13g2_decap_4 FILLER_42_1321 ();
 sg13g2_fill_2 FILLER_42_1338 ();
 sg13g2_decap_4 FILLER_42_1371 ();
 sg13g2_fill_1 FILLER_42_1375 ();
 sg13g2_fill_1 FILLER_42_1397 ();
 sg13g2_decap_8 FILLER_42_1423 ();
 sg13g2_fill_1 FILLER_42_1556 ();
 sg13g2_fill_2 FILLER_42_1615 ();
 sg13g2_fill_1 FILLER_42_1617 ();
 sg13g2_decap_8 FILLER_42_1658 ();
 sg13g2_decap_4 FILLER_42_1665 ();
 sg13g2_fill_1 FILLER_42_1686 ();
 sg13g2_fill_1 FILLER_42_1691 ();
 sg13g2_decap_4 FILLER_42_1696 ();
 sg13g2_fill_2 FILLER_42_1719 ();
 sg13g2_fill_1 FILLER_42_1721 ();
 sg13g2_decap_4 FILLER_42_1775 ();
 sg13g2_fill_2 FILLER_42_1792 ();
 sg13g2_fill_2 FILLER_42_1802 ();
 sg13g2_decap_8 FILLER_42_1816 ();
 sg13g2_fill_2 FILLER_42_1823 ();
 sg13g2_decap_8 FILLER_42_1838 ();
 sg13g2_fill_2 FILLER_42_1845 ();
 sg13g2_decap_8 FILLER_42_1874 ();
 sg13g2_decap_8 FILLER_42_1881 ();
 sg13g2_decap_4 FILLER_42_1888 ();
 sg13g2_fill_2 FILLER_42_1892 ();
 sg13g2_decap_4 FILLER_42_1907 ();
 sg13g2_fill_1 FILLER_42_1911 ();
 sg13g2_decap_8 FILLER_42_2015 ();
 sg13g2_decap_4 FILLER_42_2022 ();
 sg13g2_decap_8 FILLER_42_2039 ();
 sg13g2_decap_8 FILLER_42_2046 ();
 sg13g2_decap_4 FILLER_42_2053 ();
 sg13g2_fill_2 FILLER_42_2057 ();
 sg13g2_decap_4 FILLER_42_2077 ();
 sg13g2_decap_8 FILLER_42_2099 ();
 sg13g2_fill_2 FILLER_42_2106 ();
 sg13g2_fill_1 FILLER_42_2108 ();
 sg13g2_decap_8 FILLER_42_2125 ();
 sg13g2_fill_2 FILLER_42_2132 ();
 sg13g2_decap_8 FILLER_42_2160 ();
 sg13g2_decap_8 FILLER_42_2167 ();
 sg13g2_decap_8 FILLER_42_2174 ();
 sg13g2_decap_8 FILLER_42_2181 ();
 sg13g2_fill_1 FILLER_42_2188 ();
 sg13g2_fill_2 FILLER_42_2230 ();
 sg13g2_decap_8 FILLER_42_2263 ();
 sg13g2_decap_4 FILLER_42_2270 ();
 sg13g2_fill_1 FILLER_42_2274 ();
 sg13g2_fill_2 FILLER_42_2351 ();
 sg13g2_fill_2 FILLER_42_2420 ();
 sg13g2_fill_2 FILLER_42_2435 ();
 sg13g2_decap_4 FILLER_42_2469 ();
 sg13g2_decap_4 FILLER_42_2513 ();
 sg13g2_fill_1 FILLER_42_2561 ();
 sg13g2_fill_2 FILLER_42_2579 ();
 sg13g2_decap_4 FILLER_42_2648 ();
 sg13g2_fill_1 FILLER_42_2652 ();
 sg13g2_fill_2 FILLER_42_2721 ();
 sg13g2_fill_2 FILLER_42_2732 ();
 sg13g2_fill_1 FILLER_42_2734 ();
 sg13g2_fill_1 FILLER_42_2748 ();
 sg13g2_fill_1 FILLER_42_2758 ();
 sg13g2_decap_4 FILLER_42_2773 ();
 sg13g2_fill_2 FILLER_42_2777 ();
 sg13g2_decap_4 FILLER_42_2783 ();
 sg13g2_fill_2 FILLER_42_2792 ();
 sg13g2_decap_4 FILLER_42_2807 ();
 sg13g2_fill_2 FILLER_42_2811 ();
 sg13g2_decap_8 FILLER_42_2826 ();
 sg13g2_decap_8 FILLER_42_2833 ();
 sg13g2_fill_1 FILLER_42_2840 ();
 sg13g2_decap_8 FILLER_42_2873 ();
 sg13g2_decap_4 FILLER_42_2880 ();
 sg13g2_fill_1 FILLER_42_2884 ();
 sg13g2_fill_2 FILLER_42_2922 ();
 sg13g2_fill_1 FILLER_42_2924 ();
 sg13g2_decap_4 FILLER_42_2946 ();
 sg13g2_decap_8 FILLER_42_2965 ();
 sg13g2_decap_8 FILLER_42_2989 ();
 sg13g2_fill_2 FILLER_42_2996 ();
 sg13g2_fill_2 FILLER_42_3024 ();
 sg13g2_fill_1 FILLER_42_3026 ();
 sg13g2_fill_2 FILLER_42_3032 ();
 sg13g2_fill_1 FILLER_42_3034 ();
 sg13g2_fill_1 FILLER_42_3060 ();
 sg13g2_decap_8 FILLER_42_3074 ();
 sg13g2_fill_1 FILLER_42_3081 ();
 sg13g2_fill_2 FILLER_42_3110 ();
 sg13g2_fill_2 FILLER_42_3145 ();
 sg13g2_decap_8 FILLER_42_3164 ();
 sg13g2_fill_2 FILLER_42_3171 ();
 sg13g2_fill_1 FILLER_42_3173 ();
 sg13g2_fill_2 FILLER_42_3195 ();
 sg13g2_fill_1 FILLER_42_3197 ();
 sg13g2_fill_2 FILLER_42_3211 ();
 sg13g2_decap_4 FILLER_42_3243 ();
 sg13g2_fill_1 FILLER_42_3262 ();
 sg13g2_decap_4 FILLER_42_3277 ();
 sg13g2_fill_2 FILLER_42_3281 ();
 sg13g2_decap_8 FILLER_42_3297 ();
 sg13g2_decap_4 FILLER_42_3304 ();
 sg13g2_fill_2 FILLER_42_3308 ();
 sg13g2_decap_8 FILLER_42_3328 ();
 sg13g2_fill_2 FILLER_42_3335 ();
 sg13g2_fill_2 FILLER_42_3345 ();
 sg13g2_fill_1 FILLER_42_3347 ();
 sg13g2_fill_1 FILLER_42_3362 ();
 sg13g2_fill_2 FILLER_42_3391 ();
 sg13g2_decap_8 FILLER_42_3397 ();
 sg13g2_decap_8 FILLER_42_3404 ();
 sg13g2_fill_2 FILLER_42_3440 ();
 sg13g2_fill_1 FILLER_42_3442 ();
 sg13g2_fill_2 FILLER_42_3457 ();
 sg13g2_fill_1 FILLER_42_3459 ();
 sg13g2_decap_8 FILLER_42_3511 ();
 sg13g2_decap_8 FILLER_42_3518 ();
 sg13g2_decap_8 FILLER_42_3525 ();
 sg13g2_decap_8 FILLER_42_3532 ();
 sg13g2_decap_8 FILLER_42_3539 ();
 sg13g2_decap_8 FILLER_42_3546 ();
 sg13g2_decap_8 FILLER_42_3553 ();
 sg13g2_decap_8 FILLER_42_3560 ();
 sg13g2_decap_8 FILLER_42_3567 ();
 sg13g2_decap_4 FILLER_42_3574 ();
 sg13g2_fill_2 FILLER_42_3578 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_4 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_116 ();
 sg13g2_fill_2 FILLER_43_188 ();
 sg13g2_fill_2 FILLER_43_195 ();
 sg13g2_fill_1 FILLER_43_228 ();
 sg13g2_fill_2 FILLER_43_260 ();
 sg13g2_fill_2 FILLER_43_271 ();
 sg13g2_fill_1 FILLER_43_273 ();
 sg13g2_fill_2 FILLER_43_287 ();
 sg13g2_fill_1 FILLER_43_289 ();
 sg13g2_fill_1 FILLER_43_295 ();
 sg13g2_fill_2 FILLER_43_300 ();
 sg13g2_fill_2 FILLER_43_418 ();
 sg13g2_fill_1 FILLER_43_420 ();
 sg13g2_fill_2 FILLER_43_440 ();
 sg13g2_fill_1 FILLER_43_442 ();
 sg13g2_fill_2 FILLER_43_479 ();
 sg13g2_fill_1 FILLER_43_481 ();
 sg13g2_decap_4 FILLER_43_508 ();
 sg13g2_fill_2 FILLER_43_512 ();
 sg13g2_decap_4 FILLER_43_541 ();
 sg13g2_fill_2 FILLER_43_555 ();
 sg13g2_fill_1 FILLER_43_557 ();
 sg13g2_decap_4 FILLER_43_580 ();
 sg13g2_fill_2 FILLER_43_593 ();
 sg13g2_fill_1 FILLER_43_595 ();
 sg13g2_decap_4 FILLER_43_648 ();
 sg13g2_fill_2 FILLER_43_670 ();
 sg13g2_fill_2 FILLER_43_677 ();
 sg13g2_decap_4 FILLER_43_697 ();
 sg13g2_fill_2 FILLER_43_710 ();
 sg13g2_decap_4 FILLER_43_742 ();
 sg13g2_fill_1 FILLER_43_746 ();
 sg13g2_decap_8 FILLER_43_793 ();
 sg13g2_fill_2 FILLER_43_800 ();
 sg13g2_decap_4 FILLER_43_829 ();
 sg13g2_fill_2 FILLER_43_866 ();
 sg13g2_decap_8 FILLER_43_923 ();
 sg13g2_fill_1 FILLER_43_960 ();
 sg13g2_fill_2 FILLER_43_988 ();
 sg13g2_fill_1 FILLER_43_1062 ();
 sg13g2_fill_2 FILLER_43_1072 ();
 sg13g2_fill_1 FILLER_43_1096 ();
 sg13g2_fill_1 FILLER_43_1110 ();
 sg13g2_fill_2 FILLER_43_1199 ();
 sg13g2_fill_1 FILLER_43_1201 ();
 sg13g2_fill_2 FILLER_43_1230 ();
 sg13g2_decap_4 FILLER_43_1237 ();
 sg13g2_fill_1 FILLER_43_1241 ();
 sg13g2_fill_2 FILLER_43_1245 ();
 sg13g2_decap_8 FILLER_43_1314 ();
 sg13g2_decap_4 FILLER_43_1321 ();
 sg13g2_fill_2 FILLER_43_1351 ();
 sg13g2_fill_1 FILLER_43_1353 ();
 sg13g2_fill_2 FILLER_43_1363 ();
 sg13g2_fill_2 FILLER_43_1374 ();
 sg13g2_decap_8 FILLER_43_1380 ();
 sg13g2_decap_8 FILLER_43_1387 ();
 sg13g2_fill_2 FILLER_43_1394 ();
 sg13g2_fill_1 FILLER_43_1423 ();
 sg13g2_decap_4 FILLER_43_1437 ();
 sg13g2_fill_2 FILLER_43_1441 ();
 sg13g2_fill_2 FILLER_43_1479 ();
 sg13g2_fill_1 FILLER_43_1481 ();
 sg13g2_decap_8 FILLER_43_1513 ();
 sg13g2_fill_1 FILLER_43_1520 ();
 sg13g2_decap_8 FILLER_43_1526 ();
 sg13g2_decap_8 FILLER_43_1533 ();
 sg13g2_fill_1 FILLER_43_1540 ();
 sg13g2_decap_4 FILLER_43_1545 ();
 sg13g2_decap_8 FILLER_43_1558 ();
 sg13g2_decap_8 FILLER_43_1565 ();
 sg13g2_fill_2 FILLER_43_1572 ();
 sg13g2_fill_2 FILLER_43_1588 ();
 sg13g2_fill_2 FILLER_43_1604 ();
 sg13g2_fill_1 FILLER_43_1606 ();
 sg13g2_fill_1 FILLER_43_1652 ();
 sg13g2_fill_1 FILLER_43_1681 ();
 sg13g2_fill_1 FILLER_43_1797 ();
 sg13g2_fill_1 FILLER_43_1816 ();
 sg13g2_decap_4 FILLER_43_1830 ();
 sg13g2_fill_1 FILLER_43_1834 ();
 sg13g2_decap_8 FILLER_43_1838 ();
 sg13g2_decap_8 FILLER_43_1845 ();
 sg13g2_fill_2 FILLER_43_1852 ();
 sg13g2_fill_1 FILLER_43_1854 ();
 sg13g2_fill_2 FILLER_43_1919 ();
 sg13g2_fill_1 FILLER_43_1921 ();
 sg13g2_fill_2 FILLER_43_1941 ();
 sg13g2_fill_1 FILLER_43_1943 ();
 sg13g2_decap_4 FILLER_43_1968 ();
 sg13g2_fill_2 FILLER_43_1972 ();
 sg13g2_decap_8 FILLER_43_1979 ();
 sg13g2_fill_2 FILLER_43_1986 ();
 sg13g2_fill_1 FILLER_43_1988 ();
 sg13g2_fill_1 FILLER_43_2054 ();
 sg13g2_decap_4 FILLER_43_2060 ();
 sg13g2_fill_1 FILLER_43_2064 ();
 sg13g2_decap_8 FILLER_43_2078 ();
 sg13g2_fill_2 FILLER_43_2085 ();
 sg13g2_fill_1 FILLER_43_2087 ();
 sg13g2_decap_4 FILLER_43_2107 ();
 sg13g2_fill_2 FILLER_43_2111 ();
 sg13g2_fill_2 FILLER_43_2139 ();
 sg13g2_decap_8 FILLER_43_2157 ();
 sg13g2_fill_2 FILLER_43_2210 ();
 sg13g2_fill_1 FILLER_43_2212 ();
 sg13g2_decap_8 FILLER_43_2245 ();
 sg13g2_fill_2 FILLER_43_2279 ();
 sg13g2_fill_1 FILLER_43_2281 ();
 sg13g2_fill_1 FILLER_43_2302 ();
 sg13g2_fill_2 FILLER_43_2338 ();
 sg13g2_fill_2 FILLER_43_2350 ();
 sg13g2_fill_1 FILLER_43_2385 ();
 sg13g2_decap_4 FILLER_43_2427 ();
 sg13g2_fill_1 FILLER_43_2431 ();
 sg13g2_decap_4 FILLER_43_2445 ();
 sg13g2_fill_1 FILLER_43_2449 ();
 sg13g2_decap_4 FILLER_43_2455 ();
 sg13g2_fill_2 FILLER_43_2468 ();
 sg13g2_fill_1 FILLER_43_2470 ();
 sg13g2_decap_8 FILLER_43_2485 ();
 sg13g2_fill_2 FILLER_43_2505 ();
 sg13g2_decap_4 FILLER_43_2524 ();
 sg13g2_decap_4 FILLER_43_2542 ();
 sg13g2_decap_8 FILLER_43_2582 ();
 sg13g2_decap_4 FILLER_43_2589 ();
 sg13g2_decap_8 FILLER_43_2654 ();
 sg13g2_fill_2 FILLER_43_2661 ();
 sg13g2_fill_1 FILLER_43_2663 ();
 sg13g2_fill_1 FILLER_43_2673 ();
 sg13g2_decap_8 FILLER_43_2678 ();
 sg13g2_decap_8 FILLER_43_2685 ();
 sg13g2_decap_8 FILLER_43_2692 ();
 sg13g2_fill_1 FILLER_43_2699 ();
 sg13g2_fill_1 FILLER_43_2705 ();
 sg13g2_decap_8 FILLER_43_2733 ();
 sg13g2_fill_1 FILLER_43_2740 ();
 sg13g2_decap_8 FILLER_43_2822 ();
 sg13g2_fill_2 FILLER_43_2829 ();
 sg13g2_fill_2 FILLER_43_2901 ();
 sg13g2_fill_1 FILLER_43_2924 ();
 sg13g2_fill_2 FILLER_43_2930 ();
 sg13g2_fill_1 FILLER_43_2932 ();
 sg13g2_decap_8 FILLER_43_2937 ();
 sg13g2_fill_2 FILLER_43_2944 ();
 sg13g2_fill_1 FILLER_43_2946 ();
 sg13g2_decap_8 FILLER_43_2991 ();
 sg13g2_decap_4 FILLER_43_2998 ();
 sg13g2_fill_1 FILLER_43_3002 ();
 sg13g2_fill_2 FILLER_43_3020 ();
 sg13g2_fill_1 FILLER_43_3022 ();
 sg13g2_decap_8 FILLER_43_3031 ();
 sg13g2_fill_1 FILLER_43_3038 ();
 sg13g2_decap_8 FILLER_43_3073 ();
 sg13g2_decap_8 FILLER_43_3080 ();
 sg13g2_decap_8 FILLER_43_3091 ();
 sg13g2_decap_8 FILLER_43_3098 ();
 sg13g2_decap_4 FILLER_43_3105 ();
 sg13g2_fill_1 FILLER_43_3109 ();
 sg13g2_decap_8 FILLER_43_3115 ();
 sg13g2_fill_2 FILLER_43_3175 ();
 sg13g2_fill_2 FILLER_43_3199 ();
 sg13g2_fill_1 FILLER_43_3201 ();
 sg13g2_fill_1 FILLER_43_3220 ();
 sg13g2_fill_2 FILLER_43_3234 ();
 sg13g2_fill_2 FILLER_43_3245 ();
 sg13g2_fill_1 FILLER_43_3247 ();
 sg13g2_decap_4 FILLER_43_3261 ();
 sg13g2_fill_2 FILLER_43_3265 ();
 sg13g2_decap_8 FILLER_43_3299 ();
 sg13g2_fill_1 FILLER_43_3313 ();
 sg13g2_decap_8 FILLER_43_3332 ();
 sg13g2_decap_4 FILLER_43_3339 ();
 sg13g2_fill_2 FILLER_43_3343 ();
 sg13g2_decap_4 FILLER_43_3361 ();
 sg13g2_fill_1 FILLER_43_3365 ();
 sg13g2_decap_8 FILLER_43_3393 ();
 sg13g2_decap_4 FILLER_43_3400 ();
 sg13g2_decap_4 FILLER_43_3430 ();
 sg13g2_fill_2 FILLER_43_3434 ();
 sg13g2_fill_1 FILLER_43_3440 ();
 sg13g2_fill_2 FILLER_43_3458 ();
 sg13g2_fill_1 FILLER_43_3460 ();
 sg13g2_decap_8 FILLER_43_3478 ();
 sg13g2_fill_2 FILLER_43_3485 ();
 sg13g2_fill_1 FILLER_43_3487 ();
 sg13g2_decap_8 FILLER_43_3492 ();
 sg13g2_decap_8 FILLER_43_3499 ();
 sg13g2_decap_8 FILLER_43_3506 ();
 sg13g2_decap_8 FILLER_43_3513 ();
 sg13g2_decap_8 FILLER_43_3520 ();
 sg13g2_decap_8 FILLER_43_3527 ();
 sg13g2_decap_8 FILLER_43_3534 ();
 sg13g2_decap_8 FILLER_43_3541 ();
 sg13g2_decap_8 FILLER_43_3548 ();
 sg13g2_decap_8 FILLER_43_3555 ();
 sg13g2_decap_8 FILLER_43_3562 ();
 sg13g2_decap_8 FILLER_43_3569 ();
 sg13g2_decap_4 FILLER_43_3576 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_4 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_101 ();
 sg13g2_decap_8 FILLER_44_108 ();
 sg13g2_decap_8 FILLER_44_115 ();
 sg13g2_fill_2 FILLER_44_144 ();
 sg13g2_decap_4 FILLER_44_155 ();
 sg13g2_fill_2 FILLER_44_159 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_208 ();
 sg13g2_fill_1 FILLER_44_210 ();
 sg13g2_fill_2 FILLER_44_220 ();
 sg13g2_fill_2 FILLER_44_404 ();
 sg13g2_fill_1 FILLER_44_419 ();
 sg13g2_fill_1 FILLER_44_465 ();
 sg13g2_decap_4 FILLER_44_526 ();
 sg13g2_fill_1 FILLER_44_530 ();
 sg13g2_fill_2 FILLER_44_541 ();
 sg13g2_fill_1 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_625 ();
 sg13g2_decap_4 FILLER_44_632 ();
 sg13g2_decap_8 FILLER_44_653 ();
 sg13g2_fill_2 FILLER_44_673 ();
 sg13g2_fill_1 FILLER_44_675 ();
 sg13g2_fill_2 FILLER_44_717 ();
 sg13g2_fill_1 FILLER_44_733 ();
 sg13g2_decap_4 FILLER_44_744 ();
 sg13g2_fill_1 FILLER_44_748 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_fill_2 FILLER_44_863 ();
 sg13g2_fill_1 FILLER_44_907 ();
 sg13g2_decap_4 FILLER_44_918 ();
 sg13g2_fill_1 FILLER_44_922 ();
 sg13g2_decap_8 FILLER_44_955 ();
 sg13g2_fill_1 FILLER_44_962 ();
 sg13g2_fill_2 FILLER_44_990 ();
 sg13g2_fill_1 FILLER_44_1014 ();
 sg13g2_fill_2 FILLER_44_1024 ();
 sg13g2_fill_2 FILLER_44_1084 ();
 sg13g2_fill_1 FILLER_44_1086 ();
 sg13g2_fill_1 FILLER_44_1118 ();
 sg13g2_decap_8 FILLER_44_1137 ();
 sg13g2_fill_1 FILLER_44_1144 ();
 sg13g2_fill_2 FILLER_44_1154 ();
 sg13g2_fill_2 FILLER_44_1189 ();
 sg13g2_fill_2 FILLER_44_1204 ();
 sg13g2_fill_1 FILLER_44_1215 ();
 sg13g2_fill_2 FILLER_44_1225 ();
 sg13g2_fill_1 FILLER_44_1236 ();
 sg13g2_decap_8 FILLER_44_1264 ();
 sg13g2_decap_8 FILLER_44_1271 ();
 sg13g2_decap_8 FILLER_44_1291 ();
 sg13g2_decap_4 FILLER_44_1298 ();
 sg13g2_fill_2 FILLER_44_1307 ();
 sg13g2_fill_1 FILLER_44_1309 ();
 sg13g2_fill_2 FILLER_44_1319 ();
 sg13g2_decap_4 FILLER_44_1334 ();
 sg13g2_fill_1 FILLER_44_1342 ();
 sg13g2_fill_1 FILLER_44_1370 ();
 sg13g2_fill_1 FILLER_44_1408 ();
 sg13g2_fill_2 FILLER_44_1504 ();
 sg13g2_fill_1 FILLER_44_1506 ();
 sg13g2_fill_1 FILLER_44_1549 ();
 sg13g2_decap_4 FILLER_44_1637 ();
 sg13g2_fill_1 FILLER_44_1641 ();
 sg13g2_fill_1 FILLER_44_1655 ();
 sg13g2_fill_2 FILLER_44_1666 ();
 sg13g2_fill_1 FILLER_44_1668 ();
 sg13g2_fill_2 FILLER_44_1724 ();
 sg13g2_decap_8 FILLER_44_1748 ();
 sg13g2_decap_4 FILLER_44_1765 ();
 sg13g2_fill_1 FILLER_44_1769 ();
 sg13g2_decap_4 FILLER_44_1815 ();
 sg13g2_fill_1 FILLER_44_1819 ();
 sg13g2_decap_8 FILLER_44_1848 ();
 sg13g2_decap_8 FILLER_44_1855 ();
 sg13g2_fill_2 FILLER_44_1862 ();
 sg13g2_decap_8 FILLER_44_1873 ();
 sg13g2_fill_2 FILLER_44_1880 ();
 sg13g2_decap_4 FILLER_44_1891 ();
 sg13g2_fill_1 FILLER_44_1895 ();
 sg13g2_fill_2 FILLER_44_1915 ();
 sg13g2_decap_4 FILLER_44_1935 ();
 sg13g2_fill_1 FILLER_44_1939 ();
 sg13g2_decap_4 FILLER_44_1986 ();
 sg13g2_fill_1 FILLER_44_2043 ();
 sg13g2_fill_2 FILLER_44_2072 ();
 sg13g2_fill_1 FILLER_44_2087 ();
 sg13g2_fill_1 FILLER_44_2101 ();
 sg13g2_fill_1 FILLER_44_2119 ();
 sg13g2_decap_4 FILLER_44_2148 ();
 sg13g2_fill_2 FILLER_44_2152 ();
 sg13g2_decap_4 FILLER_44_2228 ();
 sg13g2_fill_1 FILLER_44_2232 ();
 sg13g2_fill_1 FILLER_44_2264 ();
 sg13g2_fill_2 FILLER_44_2289 ();
 sg13g2_fill_2 FILLER_44_2345 ();
 sg13g2_fill_1 FILLER_44_2347 ();
 sg13g2_fill_2 FILLER_44_2401 ();
 sg13g2_fill_1 FILLER_44_2403 ();
 sg13g2_decap_4 FILLER_44_2436 ();
 sg13g2_fill_2 FILLER_44_2440 ();
 sg13g2_decap_4 FILLER_44_2447 ();
 sg13g2_fill_1 FILLER_44_2451 ();
 sg13g2_fill_2 FILLER_44_2488 ();
 sg13g2_fill_1 FILLER_44_2499 ();
 sg13g2_fill_2 FILLER_44_2514 ();
 sg13g2_decap_4 FILLER_44_2582 ();
 sg13g2_fill_2 FILLER_44_2600 ();
 sg13g2_fill_1 FILLER_44_2602 ();
 sg13g2_fill_2 FILLER_44_2612 ();
 sg13g2_fill_1 FILLER_44_2614 ();
 sg13g2_fill_2 FILLER_44_2624 ();
 sg13g2_decap_8 FILLER_44_2640 ();
 sg13g2_decap_8 FILLER_44_2647 ();
 sg13g2_fill_2 FILLER_44_2686 ();
 sg13g2_fill_1 FILLER_44_2688 ();
 sg13g2_fill_2 FILLER_44_2769 ();
 sg13g2_fill_1 FILLER_44_2771 ();
 sg13g2_fill_2 FILLER_44_2781 ();
 sg13g2_fill_1 FILLER_44_2783 ();
 sg13g2_fill_2 FILLER_44_2845 ();
 sg13g2_decap_4 FILLER_44_2984 ();
 sg13g2_fill_1 FILLER_44_2988 ();
 sg13g2_fill_1 FILLER_44_2998 ();
 sg13g2_decap_8 FILLER_44_3028 ();
 sg13g2_fill_2 FILLER_44_3035 ();
 sg13g2_fill_1 FILLER_44_3037 ();
 sg13g2_decap_4 FILLER_44_3051 ();
 sg13g2_fill_2 FILLER_44_3055 ();
 sg13g2_decap_8 FILLER_44_3066 ();
 sg13g2_fill_2 FILLER_44_3159 ();
 sg13g2_fill_1 FILLER_44_3161 ();
 sg13g2_fill_1 FILLER_44_3171 ();
 sg13g2_fill_2 FILLER_44_3213 ();
 sg13g2_decap_4 FILLER_44_3242 ();
 sg13g2_fill_2 FILLER_44_3246 ();
 sg13g2_fill_2 FILLER_44_3275 ();
 sg13g2_fill_1 FILLER_44_3277 ();
 sg13g2_fill_1 FILLER_44_3318 ();
 sg13g2_fill_2 FILLER_44_3346 ();
 sg13g2_fill_1 FILLER_44_3348 ();
 sg13g2_decap_8 FILLER_44_3389 ();
 sg13g2_decap_8 FILLER_44_3396 ();
 sg13g2_decap_4 FILLER_44_3403 ();
 sg13g2_fill_1 FILLER_44_3407 ();
 sg13g2_decap_8 FILLER_44_3482 ();
 sg13g2_decap_8 FILLER_44_3489 ();
 sg13g2_decap_8 FILLER_44_3496 ();
 sg13g2_decap_8 FILLER_44_3503 ();
 sg13g2_decap_8 FILLER_44_3510 ();
 sg13g2_decap_8 FILLER_44_3517 ();
 sg13g2_decap_8 FILLER_44_3524 ();
 sg13g2_decap_8 FILLER_44_3531 ();
 sg13g2_decap_8 FILLER_44_3538 ();
 sg13g2_decap_8 FILLER_44_3545 ();
 sg13g2_decap_8 FILLER_44_3552 ();
 sg13g2_decap_8 FILLER_44_3559 ();
 sg13g2_decap_8 FILLER_44_3566 ();
 sg13g2_decap_8 FILLER_44_3573 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_fill_2 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_149 ();
 sg13g2_decap_8 FILLER_45_155 ();
 sg13g2_decap_4 FILLER_45_162 ();
 sg13g2_fill_2 FILLER_45_166 ();
 sg13g2_fill_2 FILLER_45_173 ();
 sg13g2_fill_1 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_4 FILLER_45_238 ();
 sg13g2_fill_1 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_259 ();
 sg13g2_decap_4 FILLER_45_265 ();
 sg13g2_fill_2 FILLER_45_269 ();
 sg13g2_fill_2 FILLER_45_289 ();
 sg13g2_decap_4 FILLER_45_314 ();
 sg13g2_fill_1 FILLER_45_323 ();
 sg13g2_fill_2 FILLER_45_354 ();
 sg13g2_fill_1 FILLER_45_375 ();
 sg13g2_fill_1 FILLER_45_381 ();
 sg13g2_fill_1 FILLER_45_396 ();
 sg13g2_fill_2 FILLER_45_447 ();
 sg13g2_fill_1 FILLER_45_449 ();
 sg13g2_fill_2 FILLER_45_467 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_fill_2 FILLER_45_511 ();
 sg13g2_fill_2 FILLER_45_540 ();
 sg13g2_fill_2 FILLER_45_564 ();
 sg13g2_decap_4 FILLER_45_642 ();
 sg13g2_fill_2 FILLER_45_646 ();
 sg13g2_decap_4 FILLER_45_661 ();
 sg13g2_fill_2 FILLER_45_665 ();
 sg13g2_decap_4 FILLER_45_699 ();
 sg13g2_decap_4 FILLER_45_830 ();
 sg13g2_fill_2 FILLER_45_834 ();
 sg13g2_fill_1 FILLER_45_863 ();
 sg13g2_decap_8 FILLER_45_868 ();
 sg13g2_fill_2 FILLER_45_875 ();
 sg13g2_decap_4 FILLER_45_963 ();
 sg13g2_fill_2 FILLER_45_980 ();
 sg13g2_fill_2 FILLER_45_1056 ();
 sg13g2_decap_8 FILLER_45_1100 ();
 sg13g2_fill_1 FILLER_45_1107 ();
 sg13g2_decap_4 FILLER_45_1118 ();
 sg13g2_fill_2 FILLER_45_1207 ();
 sg13g2_fill_2 FILLER_45_1250 ();
 sg13g2_fill_1 FILLER_45_1252 ();
 sg13g2_fill_1 FILLER_45_1262 ();
 sg13g2_decap_4 FILLER_45_1295 ();
 sg13g2_fill_1 FILLER_45_1299 ();
 sg13g2_decap_4 FILLER_45_1327 ();
 sg13g2_fill_1 FILLER_45_1331 ();
 sg13g2_fill_1 FILLER_45_1351 ();
 sg13g2_decap_8 FILLER_45_1371 ();
 sg13g2_fill_1 FILLER_45_1378 ();
 sg13g2_decap_8 FILLER_45_1406 ();
 sg13g2_fill_2 FILLER_45_1413 ();
 sg13g2_fill_1 FILLER_45_1415 ();
 sg13g2_decap_4 FILLER_45_1435 ();
 sg13g2_fill_1 FILLER_45_1439 ();
 sg13g2_fill_2 FILLER_45_1477 ();
 sg13g2_fill_1 FILLER_45_1479 ();
 sg13g2_decap_4 FILLER_45_1494 ();
 sg13g2_fill_2 FILLER_45_1498 ();
 sg13g2_fill_1 FILLER_45_1510 ();
 sg13g2_fill_2 FILLER_45_1520 ();
 sg13g2_fill_1 FILLER_45_1522 ();
 sg13g2_fill_2 FILLER_45_1556 ();
 sg13g2_fill_1 FILLER_45_1582 ();
 sg13g2_fill_1 FILLER_45_1619 ();
 sg13g2_fill_2 FILLER_45_1629 ();
 sg13g2_fill_1 FILLER_45_1631 ();
 sg13g2_decap_4 FILLER_45_1672 ();
 sg13g2_fill_1 FILLER_45_1676 ();
 sg13g2_decap_4 FILLER_45_1695 ();
 sg13g2_decap_4 FILLER_45_1709 ();
 sg13g2_fill_2 FILLER_45_1755 ();
 sg13g2_fill_2 FILLER_45_1784 ();
 sg13g2_fill_1 FILLER_45_1791 ();
 sg13g2_fill_1 FILLER_45_1801 ();
 sg13g2_decap_8 FILLER_45_1811 ();
 sg13g2_decap_4 FILLER_45_1818 ();
 sg13g2_decap_4 FILLER_45_1825 ();
 sg13g2_fill_2 FILLER_45_1829 ();
 sg13g2_fill_2 FILLER_45_1858 ();
 sg13g2_fill_1 FILLER_45_1860 ();
 sg13g2_decap_8 FILLER_45_1888 ();
 sg13g2_fill_2 FILLER_45_1895 ();
 sg13g2_decap_4 FILLER_45_1929 ();
 sg13g2_fill_1 FILLER_45_1965 ();
 sg13g2_fill_2 FILLER_45_2020 ();
 sg13g2_fill_1 FILLER_45_2022 ();
 sg13g2_decap_8 FILLER_45_2087 ();
 sg13g2_fill_2 FILLER_45_2094 ();
 sg13g2_fill_2 FILLER_45_2123 ();
 sg13g2_fill_1 FILLER_45_2160 ();
 sg13g2_fill_2 FILLER_45_2179 ();
 sg13g2_decap_4 FILLER_45_2208 ();
 sg13g2_fill_2 FILLER_45_2312 ();
 sg13g2_fill_1 FILLER_45_2314 ();
 sg13g2_fill_2 FILLER_45_2328 ();
 sg13g2_fill_1 FILLER_45_2340 ();
 sg13g2_fill_1 FILLER_45_2354 ();
 sg13g2_fill_1 FILLER_45_2422 ();
 sg13g2_decap_8 FILLER_45_2456 ();
 sg13g2_decap_8 FILLER_45_2463 ();
 sg13g2_decap_8 FILLER_45_2470 ();
 sg13g2_fill_1 FILLER_45_2477 ();
 sg13g2_fill_1 FILLER_45_2550 ();
 sg13g2_fill_1 FILLER_45_2620 ();
 sg13g2_decap_4 FILLER_45_2653 ();
 sg13g2_fill_1 FILLER_45_2657 ();
 sg13g2_fill_2 FILLER_45_2663 ();
 sg13g2_fill_1 FILLER_45_2665 ();
 sg13g2_fill_2 FILLER_45_2670 ();
 sg13g2_decap_4 FILLER_45_2676 ();
 sg13g2_decap_4 FILLER_45_2689 ();
 sg13g2_fill_2 FILLER_45_2693 ();
 sg13g2_fill_1 FILLER_45_2735 ();
 sg13g2_fill_2 FILLER_45_2781 ();
 sg13g2_decap_8 FILLER_45_2810 ();
 sg13g2_fill_2 FILLER_45_2817 ();
 sg13g2_fill_2 FILLER_45_2845 ();
 sg13g2_fill_1 FILLER_45_2847 ();
 sg13g2_fill_1 FILLER_45_2922 ();
 sg13g2_decap_8 FILLER_45_2941 ();
 sg13g2_decap_4 FILLER_45_2948 ();
 sg13g2_decap_4 FILLER_45_2975 ();
 sg13g2_fill_1 FILLER_45_2979 ();
 sg13g2_fill_1 FILLER_45_3016 ();
 sg13g2_fill_2 FILLER_45_3044 ();
 sg13g2_fill_1 FILLER_45_3076 ();
 sg13g2_decap_4 FILLER_45_3104 ();
 sg13g2_fill_1 FILLER_45_3120 ();
 sg13g2_decap_8 FILLER_45_3157 ();
 sg13g2_decap_4 FILLER_45_3164 ();
 sg13g2_fill_1 FILLER_45_3168 ();
 sg13g2_decap_8 FILLER_45_3181 ();
 sg13g2_decap_8 FILLER_45_3188 ();
 sg13g2_decap_4 FILLER_45_3195 ();
 sg13g2_fill_1 FILLER_45_3239 ();
 sg13g2_fill_1 FILLER_45_3253 ();
 sg13g2_decap_8 FILLER_45_3259 ();
 sg13g2_decap_8 FILLER_45_3266 ();
 sg13g2_fill_1 FILLER_45_3273 ();
 sg13g2_decap_8 FILLER_45_3279 ();
 sg13g2_decap_4 FILLER_45_3286 ();
 sg13g2_fill_2 FILLER_45_3294 ();
 sg13g2_fill_2 FILLER_45_3315 ();
 sg13g2_decap_4 FILLER_45_3351 ();
 sg13g2_fill_2 FILLER_45_3355 ();
 sg13g2_decap_8 FILLER_45_3398 ();
 sg13g2_decap_8 FILLER_45_3405 ();
 sg13g2_decap_4 FILLER_45_3412 ();
 sg13g2_decap_8 FILLER_45_3425 ();
 sg13g2_decap_8 FILLER_45_3432 ();
 sg13g2_fill_1 FILLER_45_3439 ();
 sg13g2_decap_4 FILLER_45_3445 ();
 sg13g2_fill_1 FILLER_45_3449 ();
 sg13g2_decap_8 FILLER_45_3454 ();
 sg13g2_decap_8 FILLER_45_3461 ();
 sg13g2_decap_8 FILLER_45_3468 ();
 sg13g2_decap_8 FILLER_45_3475 ();
 sg13g2_decap_8 FILLER_45_3482 ();
 sg13g2_decap_8 FILLER_45_3489 ();
 sg13g2_decap_8 FILLER_45_3496 ();
 sg13g2_decap_8 FILLER_45_3503 ();
 sg13g2_decap_8 FILLER_45_3510 ();
 sg13g2_decap_8 FILLER_45_3517 ();
 sg13g2_decap_8 FILLER_45_3524 ();
 sg13g2_decap_8 FILLER_45_3531 ();
 sg13g2_decap_8 FILLER_45_3538 ();
 sg13g2_decap_8 FILLER_45_3545 ();
 sg13g2_decap_8 FILLER_45_3552 ();
 sg13g2_decap_8 FILLER_45_3559 ();
 sg13g2_decap_8 FILLER_45_3566 ();
 sg13g2_decap_8 FILLER_45_3573 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_fill_1 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_61 ();
 sg13g2_decap_8 FILLER_46_68 ();
 sg13g2_decap_8 FILLER_46_75 ();
 sg13g2_decap_8 FILLER_46_82 ();
 sg13g2_decap_4 FILLER_46_89 ();
 sg13g2_decap_8 FILLER_46_97 ();
 sg13g2_decap_8 FILLER_46_104 ();
 sg13g2_decap_8 FILLER_46_111 ();
 sg13g2_decap_8 FILLER_46_118 ();
 sg13g2_fill_2 FILLER_46_125 ();
 sg13g2_fill_2 FILLER_46_183 ();
 sg13g2_decap_4 FILLER_46_203 ();
 sg13g2_fill_2 FILLER_46_207 ();
 sg13g2_fill_1 FILLER_46_219 ();
 sg13g2_fill_1 FILLER_46_225 ();
 sg13g2_fill_1 FILLER_46_230 ();
 sg13g2_decap_8 FILLER_46_240 ();
 sg13g2_fill_1 FILLER_46_247 ();
 sg13g2_fill_2 FILLER_46_262 ();
 sg13g2_fill_1 FILLER_46_264 ();
 sg13g2_fill_2 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_339 ();
 sg13g2_fill_2 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_376 ();
 sg13g2_fill_2 FILLER_46_410 ();
 sg13g2_decap_8 FILLER_46_433 ();
 sg13g2_fill_1 FILLER_46_440 ();
 sg13g2_fill_2 FILLER_46_445 ();
 sg13g2_fill_1 FILLER_46_447 ();
 sg13g2_decap_4 FILLER_46_464 ();
 sg13g2_fill_2 FILLER_46_486 ();
 sg13g2_fill_1 FILLER_46_488 ();
 sg13g2_decap_4 FILLER_46_547 ();
 sg13g2_fill_2 FILLER_46_597 ();
 sg13g2_decap_4 FILLER_46_669 ();
 sg13g2_fill_2 FILLER_46_673 ();
 sg13g2_fill_1 FILLER_46_702 ();
 sg13g2_fill_2 FILLER_46_706 ();
 sg13g2_decap_4 FILLER_46_712 ();
 sg13g2_fill_1 FILLER_46_716 ();
 sg13g2_decap_8 FILLER_46_726 ();
 sg13g2_decap_4 FILLER_46_733 ();
 sg13g2_decap_8 FILLER_46_750 ();
 sg13g2_decap_4 FILLER_46_757 ();
 sg13g2_fill_1 FILLER_46_811 ();
 sg13g2_fill_1 FILLER_46_848 ();
 sg13g2_fill_1 FILLER_46_923 ();
 sg13g2_fill_1 FILLER_46_933 ();
 sg13g2_decap_4 FILLER_46_961 ();
 sg13g2_fill_1 FILLER_46_965 ();
 sg13g2_decap_8 FILLER_46_971 ();
 sg13g2_decap_4 FILLER_46_978 ();
 sg13g2_fill_2 FILLER_46_991 ();
 sg13g2_fill_1 FILLER_46_993 ();
 sg13g2_decap_8 FILLER_46_1034 ();
 sg13g2_fill_1 FILLER_46_1041 ();
 sg13g2_decap_8 FILLER_46_1074 ();
 sg13g2_fill_2 FILLER_46_1117 ();
 sg13g2_fill_2 FILLER_46_1146 ();
 sg13g2_fill_1 FILLER_46_1148 ();
 sg13g2_decap_8 FILLER_46_1208 ();
 sg13g2_decap_4 FILLER_46_1215 ();
 sg13g2_fill_1 FILLER_46_1219 ();
 sg13g2_fill_2 FILLER_46_1237 ();
 sg13g2_fill_1 FILLER_46_1239 ();
 sg13g2_decap_8 FILLER_46_1244 ();
 sg13g2_decap_8 FILLER_46_1251 ();
 sg13g2_fill_2 FILLER_46_1258 ();
 sg13g2_fill_1 FILLER_46_1260 ();
 sg13g2_fill_2 FILLER_46_1275 ();
 sg13g2_fill_1 FILLER_46_1277 ();
 sg13g2_decap_8 FILLER_46_1287 ();
 sg13g2_fill_2 FILLER_46_1294 ();
 sg13g2_fill_2 FILLER_46_1334 ();
 sg13g2_fill_1 FILLER_46_1336 ();
 sg13g2_fill_1 FILLER_46_1369 ();
 sg13g2_decap_4 FILLER_46_1439 ();
 sg13g2_fill_1 FILLER_46_1443 ();
 sg13g2_fill_2 FILLER_46_1508 ();
 sg13g2_fill_2 FILLER_46_1634 ();
 sg13g2_fill_1 FILLER_46_1636 ();
 sg13g2_fill_1 FILLER_46_1668 ();
 sg13g2_fill_1 FILLER_46_1678 ();
 sg13g2_decap_4 FILLER_46_1684 ();
 sg13g2_fill_2 FILLER_46_1688 ();
 sg13g2_fill_2 FILLER_46_1735 ();
 sg13g2_fill_1 FILLER_46_1737 ();
 sg13g2_fill_1 FILLER_46_1752 ();
 sg13g2_fill_1 FILLER_46_1766 ();
 sg13g2_fill_1 FILLER_46_1781 ();
 sg13g2_fill_1 FILLER_46_1819 ();
 sg13g2_decap_4 FILLER_46_1856 ();
 sg13g2_fill_2 FILLER_46_1860 ();
 sg13g2_decap_4 FILLER_46_1871 ();
 sg13g2_fill_1 FILLER_46_1888 ();
 sg13g2_decap_8 FILLER_46_1944 ();
 sg13g2_fill_1 FILLER_46_1951 ();
 sg13g2_decap_8 FILLER_46_1984 ();
 sg13g2_fill_1 FILLER_46_1991 ();
 sg13g2_fill_2 FILLER_46_2011 ();
 sg13g2_fill_1 FILLER_46_2031 ();
 sg13g2_fill_2 FILLER_46_2059 ();
 sg13g2_fill_1 FILLER_46_2061 ();
 sg13g2_decap_4 FILLER_46_2094 ();
 sg13g2_fill_2 FILLER_46_2134 ();
 sg13g2_fill_1 FILLER_46_2136 ();
 sg13g2_decap_8 FILLER_46_2206 ();
 sg13g2_decap_4 FILLER_46_2213 ();
 sg13g2_fill_2 FILLER_46_2217 ();
 sg13g2_fill_2 FILLER_46_2264 ();
 sg13g2_fill_2 FILLER_46_2289 ();
 sg13g2_fill_1 FILLER_46_2301 ();
 sg13g2_fill_2 FILLER_46_2307 ();
 sg13g2_fill_1 FILLER_46_2385 ();
 sg13g2_decap_4 FILLER_46_2432 ();
 sg13g2_fill_2 FILLER_46_2450 ();
 sg13g2_decap_8 FILLER_46_2492 ();
 sg13g2_decap_8 FILLER_46_2499 ();
 sg13g2_fill_2 FILLER_46_2506 ();
 sg13g2_decap_4 FILLER_46_2530 ();
 sg13g2_fill_2 FILLER_46_2534 ();
 sg13g2_decap_4 FILLER_46_2597 ();
 sg13g2_fill_1 FILLER_46_2619 ();
 sg13g2_fill_2 FILLER_46_2652 ();
 sg13g2_fill_1 FILLER_46_2654 ();
 sg13g2_fill_2 FILLER_46_2736 ();
 sg13g2_fill_2 FILLER_46_2769 ();
 sg13g2_fill_1 FILLER_46_2771 ();
 sg13g2_fill_1 FILLER_46_2795 ();
 sg13g2_fill_1 FILLER_46_2800 ();
 sg13g2_fill_2 FILLER_46_2834 ();
 sg13g2_fill_1 FILLER_46_2836 ();
 sg13g2_fill_2 FILLER_46_2869 ();
 sg13g2_fill_1 FILLER_46_2871 ();
 sg13g2_decap_8 FILLER_46_2939 ();
 sg13g2_fill_2 FILLER_46_2946 ();
 sg13g2_fill_1 FILLER_46_2948 ();
 sg13g2_fill_1 FILLER_46_2966 ();
 sg13g2_fill_2 FILLER_46_2994 ();
 sg13g2_fill_1 FILLER_46_2996 ();
 sg13g2_fill_1 FILLER_46_3039 ();
 sg13g2_decap_8 FILLER_46_3045 ();
 sg13g2_decap_8 FILLER_46_3052 ();
 sg13g2_decap_8 FILLER_46_3059 ();
 sg13g2_fill_2 FILLER_46_3088 ();
 sg13g2_fill_1 FILLER_46_3090 ();
 sg13g2_decap_4 FILLER_46_3118 ();
 sg13g2_fill_1 FILLER_46_3122 ();
 sg13g2_fill_2 FILLER_46_3167 ();
 sg13g2_fill_2 FILLER_46_3191 ();
 sg13g2_fill_1 FILLER_46_3193 ();
 sg13g2_fill_2 FILLER_46_3199 ();
 sg13g2_fill_2 FILLER_46_3217 ();
 sg13g2_fill_2 FILLER_46_3367 ();
 sg13g2_fill_1 FILLER_46_3391 ();
 sg13g2_decap_8 FILLER_46_3432 ();
 sg13g2_decap_8 FILLER_46_3439 ();
 sg13g2_decap_8 FILLER_46_3446 ();
 sg13g2_decap_8 FILLER_46_3453 ();
 sg13g2_decap_8 FILLER_46_3460 ();
 sg13g2_decap_8 FILLER_46_3467 ();
 sg13g2_decap_8 FILLER_46_3474 ();
 sg13g2_decap_8 FILLER_46_3481 ();
 sg13g2_decap_8 FILLER_46_3488 ();
 sg13g2_decap_8 FILLER_46_3495 ();
 sg13g2_decap_8 FILLER_46_3502 ();
 sg13g2_decap_8 FILLER_46_3509 ();
 sg13g2_decap_8 FILLER_46_3516 ();
 sg13g2_decap_8 FILLER_46_3523 ();
 sg13g2_decap_8 FILLER_46_3530 ();
 sg13g2_decap_8 FILLER_46_3537 ();
 sg13g2_decap_8 FILLER_46_3544 ();
 sg13g2_decap_8 FILLER_46_3551 ();
 sg13g2_decap_8 FILLER_46_3558 ();
 sg13g2_decap_8 FILLER_46_3565 ();
 sg13g2_decap_8 FILLER_46_3572 ();
 sg13g2_fill_1 FILLER_46_3579 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_49 ();
 sg13g2_fill_1 FILLER_47_51 ();
 sg13g2_fill_2 FILLER_47_79 ();
 sg13g2_fill_2 FILLER_47_85 ();
 sg13g2_fill_1 FILLER_47_87 ();
 sg13g2_fill_2 FILLER_47_115 ();
 sg13g2_fill_2 FILLER_47_145 ();
 sg13g2_fill_1 FILLER_47_147 ();
 sg13g2_decap_4 FILLER_47_157 ();
 sg13g2_decap_4 FILLER_47_180 ();
 sg13g2_decap_4 FILLER_47_188 ();
 sg13g2_fill_2 FILLER_47_192 ();
 sg13g2_decap_8 FILLER_47_199 ();
 sg13g2_fill_2 FILLER_47_206 ();
 sg13g2_fill_1 FILLER_47_208 ();
 sg13g2_fill_1 FILLER_47_268 ();
 sg13g2_fill_1 FILLER_47_274 ();
 sg13g2_fill_1 FILLER_47_291 ();
 sg13g2_fill_2 FILLER_47_334 ();
 sg13g2_fill_1 FILLER_47_345 ();
 sg13g2_fill_2 FILLER_47_351 ();
 sg13g2_fill_1 FILLER_47_353 ();
 sg13g2_fill_2 FILLER_47_358 ();
 sg13g2_fill_1 FILLER_47_360 ();
 sg13g2_fill_2 FILLER_47_370 ();
 sg13g2_fill_1 FILLER_47_372 ();
 sg13g2_fill_1 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_449 ();
 sg13g2_decap_8 FILLER_47_471 ();
 sg13g2_fill_2 FILLER_47_478 ();
 sg13g2_decap_8 FILLER_47_514 ();
 sg13g2_decap_8 FILLER_47_521 ();
 sg13g2_decap_4 FILLER_47_556 ();
 sg13g2_fill_2 FILLER_47_576 ();
 sg13g2_fill_2 FILLER_47_599 ();
 sg13g2_fill_2 FILLER_47_611 ();
 sg13g2_fill_1 FILLER_47_613 ();
 sg13g2_decap_4 FILLER_47_623 ();
 sg13g2_fill_2 FILLER_47_653 ();
 sg13g2_fill_1 FILLER_47_659 ();
 sg13g2_fill_2 FILLER_47_683 ();
 sg13g2_fill_1 FILLER_47_685 ();
 sg13g2_fill_2 FILLER_47_695 ();
 sg13g2_decap_4 FILLER_47_731 ();
 sg13g2_decap_4 FILLER_47_795 ();
 sg13g2_decap_4 FILLER_47_843 ();
 sg13g2_fill_1 FILLER_47_847 ();
 sg13g2_fill_1 FILLER_47_864 ();
 sg13g2_fill_2 FILLER_47_911 ();
 sg13g2_decap_4 FILLER_47_974 ();
 sg13g2_decap_8 FILLER_47_982 ();
 sg13g2_decap_4 FILLER_47_989 ();
 sg13g2_fill_2 FILLER_47_993 ();
 sg13g2_fill_1 FILLER_47_1000 ();
 sg13g2_fill_2 FILLER_47_1010 ();
 sg13g2_decap_4 FILLER_47_1044 ();
 sg13g2_decap_8 FILLER_47_1081 ();
 sg13g2_fill_1 FILLER_47_1088 ();
 sg13g2_decap_8 FILLER_47_1126 ();
 sg13g2_fill_2 FILLER_47_1133 ();
 sg13g2_decap_4 FILLER_47_1170 ();
 sg13g2_fill_2 FILLER_47_1205 ();
 sg13g2_fill_1 FILLER_47_1207 ();
 sg13g2_fill_2 FILLER_47_1264 ();
 sg13g2_fill_1 FILLER_47_1309 ();
 sg13g2_decap_8 FILLER_47_1354 ();
 sg13g2_decap_8 FILLER_47_1365 ();
 sg13g2_decap_8 FILLER_47_1372 ();
 sg13g2_decap_8 FILLER_47_1379 ();
 sg13g2_fill_1 FILLER_47_1386 ();
 sg13g2_fill_1 FILLER_47_1401 ();
 sg13g2_decap_8 FILLER_47_1406 ();
 sg13g2_decap_4 FILLER_47_1422 ();
 sg13g2_fill_1 FILLER_47_1426 ();
 sg13g2_fill_2 FILLER_47_1454 ();
 sg13g2_fill_1 FILLER_47_1473 ();
 sg13g2_decap_4 FILLER_47_1483 ();
 sg13g2_fill_1 FILLER_47_1487 ();
 sg13g2_fill_2 FILLER_47_1525 ();
 sg13g2_decap_8 FILLER_47_1545 ();
 sg13g2_fill_1 FILLER_47_1552 ();
 sg13g2_fill_2 FILLER_47_1562 ();
 sg13g2_decap_8 FILLER_47_1573 ();
 sg13g2_decap_8 FILLER_47_1580 ();
 sg13g2_decap_4 FILLER_47_1587 ();
 sg13g2_decap_4 FILLER_47_1622 ();
 sg13g2_fill_2 FILLER_47_1626 ();
 sg13g2_fill_2 FILLER_47_1656 ();
 sg13g2_decap_4 FILLER_47_1690 ();
 sg13g2_fill_2 FILLER_47_1694 ();
 sg13g2_decap_4 FILLER_47_1791 ();
 sg13g2_decap_8 FILLER_47_1800 ();
 sg13g2_fill_2 FILLER_47_1807 ();
 sg13g2_fill_1 FILLER_47_1809 ();
 sg13g2_decap_4 FILLER_47_1838 ();
 sg13g2_fill_2 FILLER_47_1842 ();
 sg13g2_decap_4 FILLER_47_1899 ();
 sg13g2_decap_4 FILLER_47_1918 ();
 sg13g2_fill_1 FILLER_47_1956 ();
 sg13g2_decap_8 FILLER_47_1961 ();
 sg13g2_fill_2 FILLER_47_1968 ();
 sg13g2_fill_1 FILLER_47_1970 ();
 sg13g2_fill_2 FILLER_47_2008 ();
 sg13g2_fill_1 FILLER_47_2010 ();
 sg13g2_decap_4 FILLER_47_2052 ();
 sg13g2_fill_2 FILLER_47_2091 ();
 sg13g2_decap_4 FILLER_47_2115 ();
 sg13g2_fill_1 FILLER_47_2119 ();
 sg13g2_decap_8 FILLER_47_2125 ();
 sg13g2_fill_2 FILLER_47_2132 ();
 sg13g2_fill_1 FILLER_47_2160 ();
 sg13g2_fill_2 FILLER_47_2174 ();
 sg13g2_fill_2 FILLER_47_2191 ();
 sg13g2_fill_1 FILLER_47_2202 ();
 sg13g2_decap_4 FILLER_47_2230 ();
 sg13g2_fill_1 FILLER_47_2234 ();
 sg13g2_fill_2 FILLER_47_2266 ();
 sg13g2_fill_1 FILLER_47_2268 ();
 sg13g2_fill_2 FILLER_47_2302 ();
 sg13g2_decap_8 FILLER_47_2313 ();
 sg13g2_decap_4 FILLER_47_2334 ();
 sg13g2_fill_2 FILLER_47_2360 ();
 sg13g2_fill_1 FILLER_47_2362 ();
 sg13g2_fill_2 FILLER_47_2382 ();
 sg13g2_fill_1 FILLER_47_2384 ();
 sg13g2_fill_1 FILLER_47_2395 ();
 sg13g2_decap_4 FILLER_47_2405 ();
 sg13g2_fill_1 FILLER_47_2409 ();
 sg13g2_fill_2 FILLER_47_2455 ();
 sg13g2_fill_2 FILLER_47_2470 ();
 sg13g2_decap_8 FILLER_47_2509 ();
 sg13g2_fill_2 FILLER_47_2544 ();
 sg13g2_decap_8 FILLER_47_2550 ();
 sg13g2_fill_2 FILLER_47_2557 ();
 sg13g2_fill_1 FILLER_47_2586 ();
 sg13g2_fill_2 FILLER_47_2628 ();
 sg13g2_fill_1 FILLER_47_2630 ();
 sg13g2_fill_2 FILLER_47_2658 ();
 sg13g2_fill_1 FILLER_47_2660 ();
 sg13g2_fill_2 FILLER_47_2692 ();
 sg13g2_fill_1 FILLER_47_2694 ();
 sg13g2_fill_2 FILLER_47_2745 ();
 sg13g2_decap_8 FILLER_47_2765 ();
 sg13g2_fill_2 FILLER_47_2872 ();
 sg13g2_decap_8 FILLER_47_2907 ();
 sg13g2_fill_2 FILLER_47_2923 ();
 sg13g2_fill_1 FILLER_47_2925 ();
 sg13g2_fill_2 FILLER_47_2966 ();
 sg13g2_fill_1 FILLER_47_2968 ();
 sg13g2_decap_4 FILLER_47_2983 ();
 sg13g2_fill_2 FILLER_47_2987 ();
 sg13g2_fill_2 FILLER_47_2999 ();
 sg13g2_decap_4 FILLER_47_3032 ();
 sg13g2_fill_2 FILLER_47_3051 ();
 sg13g2_fill_1 FILLER_47_3053 ();
 sg13g2_fill_1 FILLER_47_3091 ();
 sg13g2_fill_1 FILLER_47_3097 ();
 sg13g2_decap_8 FILLER_47_3108 ();
 sg13g2_decap_4 FILLER_47_3115 ();
 sg13g2_fill_2 FILLER_47_3119 ();
 sg13g2_fill_2 FILLER_47_3131 ();
 sg13g2_fill_1 FILLER_47_3133 ();
 sg13g2_fill_2 FILLER_47_3138 ();
 sg13g2_decap_4 FILLER_47_3213 ();
 sg13g2_decap_4 FILLER_47_3237 ();
 sg13g2_fill_2 FILLER_47_3241 ();
 sg13g2_fill_2 FILLER_47_3247 ();
 sg13g2_fill_1 FILLER_47_3249 ();
 sg13g2_decap_8 FILLER_47_3268 ();
 sg13g2_fill_2 FILLER_47_3275 ();
 sg13g2_fill_2 FILLER_47_3322 ();
 sg13g2_decap_8 FILLER_47_3375 ();
 sg13g2_fill_1 FILLER_47_3401 ();
 sg13g2_decap_4 FILLER_47_3411 ();
 sg13g2_decap_8 FILLER_47_3425 ();
 sg13g2_decap_8 FILLER_47_3432 ();
 sg13g2_decap_8 FILLER_47_3439 ();
 sg13g2_decap_8 FILLER_47_3446 ();
 sg13g2_decap_8 FILLER_47_3453 ();
 sg13g2_decap_8 FILLER_47_3460 ();
 sg13g2_decap_8 FILLER_47_3467 ();
 sg13g2_decap_8 FILLER_47_3474 ();
 sg13g2_decap_8 FILLER_47_3481 ();
 sg13g2_decap_8 FILLER_47_3488 ();
 sg13g2_decap_8 FILLER_47_3495 ();
 sg13g2_decap_8 FILLER_47_3502 ();
 sg13g2_decap_8 FILLER_47_3509 ();
 sg13g2_decap_8 FILLER_47_3516 ();
 sg13g2_decap_8 FILLER_47_3523 ();
 sg13g2_decap_8 FILLER_47_3530 ();
 sg13g2_decap_8 FILLER_47_3537 ();
 sg13g2_decap_8 FILLER_47_3544 ();
 sg13g2_decap_8 FILLER_47_3551 ();
 sg13g2_decap_8 FILLER_47_3558 ();
 sg13g2_decap_8 FILLER_47_3565 ();
 sg13g2_decap_8 FILLER_47_3572 ();
 sg13g2_fill_1 FILLER_47_3579 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_fill_2 FILLER_48_56 ();
 sg13g2_fill_1 FILLER_48_58 ();
 sg13g2_fill_2 FILLER_48_77 ();
 sg13g2_fill_1 FILLER_48_138 ();
 sg13g2_decap_4 FILLER_48_167 ();
 sg13g2_fill_1 FILLER_48_171 ();
 sg13g2_decap_8 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_207 ();
 sg13g2_fill_1 FILLER_48_212 ();
 sg13g2_fill_1 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_249 ();
 sg13g2_fill_2 FILLER_48_266 ();
 sg13g2_fill_1 FILLER_48_286 ();
 sg13g2_fill_2 FILLER_48_327 ();
 sg13g2_fill_2 FILLER_48_334 ();
 sg13g2_fill_1 FILLER_48_345 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_fill_1 FILLER_48_402 ();
 sg13g2_fill_1 FILLER_48_430 ();
 sg13g2_fill_2 FILLER_48_457 ();
 sg13g2_fill_2 FILLER_48_473 ();
 sg13g2_decap_4 FILLER_48_480 ();
 sg13g2_decap_8 FILLER_48_509 ();
 sg13g2_fill_1 FILLER_48_516 ();
 sg13g2_fill_2 FILLER_48_529 ();
 sg13g2_fill_1 FILLER_48_531 ();
 sg13g2_decap_4 FILLER_48_540 ();
 sg13g2_fill_2 FILLER_48_544 ();
 sg13g2_fill_1 FILLER_48_569 ();
 sg13g2_fill_2 FILLER_48_606 ();
 sg13g2_fill_1 FILLER_48_608 ();
 sg13g2_decap_4 FILLER_48_613 ();
 sg13g2_fill_2 FILLER_48_617 ();
 sg13g2_fill_1 FILLER_48_628 ();
 sg13g2_fill_2 FILLER_48_664 ();
 sg13g2_fill_1 FILLER_48_666 ();
 sg13g2_fill_1 FILLER_48_716 ();
 sg13g2_decap_4 FILLER_48_738 ();
 sg13g2_fill_1 FILLER_48_760 ();
 sg13g2_decap_4 FILLER_48_789 ();
 sg13g2_fill_1 FILLER_48_793 ();
 sg13g2_fill_1 FILLER_48_817 ();
 sg13g2_fill_2 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_848 ();
 sg13g2_decap_8 FILLER_48_855 ();
 sg13g2_fill_2 FILLER_48_901 ();
 sg13g2_decap_4 FILLER_48_913 ();
 sg13g2_fill_2 FILLER_48_917 ();
 sg13g2_decap_8 FILLER_48_925 ();
 sg13g2_fill_2 FILLER_48_932 ();
 sg13g2_fill_1 FILLER_48_955 ();
 sg13g2_decap_4 FILLER_48_964 ();
 sg13g2_fill_1 FILLER_48_968 ();
 sg13g2_fill_2 FILLER_48_1015 ();
 sg13g2_fill_1 FILLER_48_1017 ();
 sg13g2_fill_2 FILLER_48_1032 ();
 sg13g2_fill_1 FILLER_48_1056 ();
 sg13g2_fill_1 FILLER_48_1096 ();
 sg13g2_decap_8 FILLER_48_1131 ();
 sg13g2_decap_4 FILLER_48_1171 ();
 sg13g2_fill_1 FILLER_48_1254 ();
 sg13g2_fill_1 FILLER_48_1273 ();
 sg13g2_decap_8 FILLER_48_1388 ();
 sg13g2_fill_2 FILLER_48_1395 ();
 sg13g2_decap_4 FILLER_48_1431 ();
 sg13g2_fill_1 FILLER_48_1468 ();
 sg13g2_fill_1 FILLER_48_1474 ();
 sg13g2_decap_8 FILLER_48_1479 ();
 sg13g2_fill_2 FILLER_48_1486 ();
 sg13g2_decap_4 FILLER_48_1497 ();
 sg13g2_decap_4 FILLER_48_1532 ();
 sg13g2_decap_4 FILLER_48_1558 ();
 sg13g2_fill_2 FILLER_48_1576 ();
 sg13g2_decap_4 FILLER_48_1605 ();
 sg13g2_fill_1 FILLER_48_1609 ();
 sg13g2_fill_2 FILLER_48_1637 ();
 sg13g2_fill_1 FILLER_48_1639 ();
 sg13g2_fill_2 FILLER_48_1648 ();
 sg13g2_fill_1 FILLER_48_1650 ();
 sg13g2_fill_2 FILLER_48_1665 ();
 sg13g2_fill_2 FILLER_48_1680 ();
 sg13g2_fill_2 FILLER_48_1695 ();
 sg13g2_fill_1 FILLER_48_1716 ();
 sg13g2_fill_2 FILLER_48_1726 ();
 sg13g2_fill_2 FILLER_48_1756 ();
 sg13g2_fill_2 FILLER_48_1785 ();
 sg13g2_fill_2 FILLER_48_1796 ();
 sg13g2_fill_1 FILLER_48_1798 ();
 sg13g2_decap_4 FILLER_48_1808 ();
 sg13g2_fill_2 FILLER_48_1812 ();
 sg13g2_fill_1 FILLER_48_1827 ();
 sg13g2_fill_2 FILLER_48_1850 ();
 sg13g2_fill_1 FILLER_48_1852 ();
 sg13g2_decap_4 FILLER_48_1870 ();
 sg13g2_fill_2 FILLER_48_1874 ();
 sg13g2_fill_2 FILLER_48_1889 ();
 sg13g2_decap_4 FILLER_48_1903 ();
 sg13g2_fill_1 FILLER_48_1907 ();
 sg13g2_fill_1 FILLER_48_1942 ();
 sg13g2_fill_2 FILLER_48_1947 ();
 sg13g2_decap_4 FILLER_48_1961 ();
 sg13g2_fill_2 FILLER_48_1983 ();
 sg13g2_fill_1 FILLER_48_2043 ();
 sg13g2_decap_8 FILLER_48_2120 ();
 sg13g2_fill_2 FILLER_48_2127 ();
 sg13g2_fill_1 FILLER_48_2129 ();
 sg13g2_fill_1 FILLER_48_2170 ();
 sg13g2_fill_2 FILLER_48_2205 ();
 sg13g2_fill_1 FILLER_48_2207 ();
 sg13g2_fill_2 FILLER_48_2212 ();
 sg13g2_fill_1 FILLER_48_2214 ();
 sg13g2_fill_2 FILLER_48_2223 ();
 sg13g2_decap_4 FILLER_48_2259 ();
 sg13g2_fill_2 FILLER_48_2294 ();
 sg13g2_fill_1 FILLER_48_2296 ();
 sg13g2_fill_2 FILLER_48_2300 ();
 sg13g2_decap_4 FILLER_48_2329 ();
 sg13g2_decap_8 FILLER_48_2342 ();
 sg13g2_decap_4 FILLER_48_2349 ();
 sg13g2_fill_1 FILLER_48_2353 ();
 sg13g2_decap_8 FILLER_48_2422 ();
 sg13g2_fill_2 FILLER_48_2429 ();
 sg13g2_fill_1 FILLER_48_2431 ();
 sg13g2_fill_1 FILLER_48_2509 ();
 sg13g2_fill_1 FILLER_48_2513 ();
 sg13g2_fill_2 FILLER_48_2540 ();
 sg13g2_decap_4 FILLER_48_2555 ();
 sg13g2_fill_1 FILLER_48_2559 ();
 sg13g2_fill_1 FILLER_48_2579 ();
 sg13g2_fill_1 FILLER_48_2602 ();
 sg13g2_decap_8 FILLER_48_2639 ();
 sg13g2_fill_2 FILLER_48_2646 ();
 sg13g2_fill_1 FILLER_48_2717 ();
 sg13g2_decap_4 FILLER_48_2762 ();
 sg13g2_fill_2 FILLER_48_2766 ();
 sg13g2_fill_2 FILLER_48_2792 ();
 sg13g2_decap_8 FILLER_48_2813 ();
 sg13g2_fill_1 FILLER_48_2847 ();
 sg13g2_fill_1 FILLER_48_2890 ();
 sg13g2_decap_8 FILLER_48_2904 ();
 sg13g2_fill_2 FILLER_48_2911 ();
 sg13g2_decap_4 FILLER_48_2931 ();
 sg13g2_fill_1 FILLER_48_2935 ();
 sg13g2_decap_4 FILLER_48_2954 ();
 sg13g2_fill_1 FILLER_48_2958 ();
 sg13g2_fill_1 FILLER_48_2965 ();
 sg13g2_decap_8 FILLER_48_2989 ();
 sg13g2_fill_2 FILLER_48_3032 ();
 sg13g2_fill_1 FILLER_48_3034 ();
 sg13g2_fill_1 FILLER_48_3045 ();
 sg13g2_decap_4 FILLER_48_3059 ();
 sg13g2_fill_1 FILLER_48_3063 ();
 sg13g2_fill_2 FILLER_48_3068 ();
 sg13g2_decap_8 FILLER_48_3110 ();
 sg13g2_decap_4 FILLER_48_3117 ();
 sg13g2_fill_1 FILLER_48_3121 ();
 sg13g2_fill_2 FILLER_48_3150 ();
 sg13g2_fill_1 FILLER_48_3152 ();
 sg13g2_fill_1 FILLER_48_3167 ();
 sg13g2_fill_1 FILLER_48_3181 ();
 sg13g2_fill_2 FILLER_48_3195 ();
 sg13g2_fill_1 FILLER_48_3197 ();
 sg13g2_decap_4 FILLER_48_3221 ();
 sg13g2_fill_2 FILLER_48_3230 ();
 sg13g2_fill_1 FILLER_48_3232 ();
 sg13g2_fill_2 FILLER_48_3323 ();
 sg13g2_fill_1 FILLER_48_3325 ();
 sg13g2_fill_2 FILLER_48_3345 ();
 sg13g2_fill_1 FILLER_48_3347 ();
 sg13g2_fill_1 FILLER_48_3357 ();
 sg13g2_fill_1 FILLER_48_3418 ();
 sg13g2_decap_8 FILLER_48_3436 ();
 sg13g2_decap_8 FILLER_48_3443 ();
 sg13g2_decap_8 FILLER_48_3450 ();
 sg13g2_decap_8 FILLER_48_3457 ();
 sg13g2_decap_8 FILLER_48_3464 ();
 sg13g2_decap_8 FILLER_48_3471 ();
 sg13g2_decap_8 FILLER_48_3478 ();
 sg13g2_decap_8 FILLER_48_3485 ();
 sg13g2_decap_8 FILLER_48_3492 ();
 sg13g2_decap_8 FILLER_48_3499 ();
 sg13g2_decap_8 FILLER_48_3506 ();
 sg13g2_decap_8 FILLER_48_3513 ();
 sg13g2_decap_8 FILLER_48_3520 ();
 sg13g2_decap_8 FILLER_48_3527 ();
 sg13g2_decap_8 FILLER_48_3534 ();
 sg13g2_decap_8 FILLER_48_3541 ();
 sg13g2_decap_8 FILLER_48_3548 ();
 sg13g2_decap_8 FILLER_48_3555 ();
 sg13g2_decap_8 FILLER_48_3562 ();
 sg13g2_decap_8 FILLER_48_3569 ();
 sg13g2_decap_4 FILLER_48_3576 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_4 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_25 ();
 sg13g2_decap_4 FILLER_49_44 ();
 sg13g2_fill_1 FILLER_49_48 ();
 sg13g2_decap_4 FILLER_49_130 ();
 sg13g2_fill_1 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_143 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_fill_1 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_fill_2 FILLER_49_200 ();
 sg13g2_fill_1 FILLER_49_202 ();
 sg13g2_decap_4 FILLER_49_231 ();
 sg13g2_decap_4 FILLER_49_281 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_decap_4 FILLER_49_379 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_fill_2 FILLER_49_397 ();
 sg13g2_fill_1 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_fill_2 FILLER_49_424 ();
 sg13g2_fill_1 FILLER_49_426 ();
 sg13g2_fill_2 FILLER_49_464 ();
 sg13g2_decap_8 FILLER_49_478 ();
 sg13g2_decap_4 FILLER_49_485 ();
 sg13g2_fill_1 FILLER_49_489 ();
 sg13g2_fill_2 FILLER_49_502 ();
 sg13g2_fill_1 FILLER_49_504 ();
 sg13g2_fill_1 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_531 ();
 sg13g2_fill_1 FILLER_49_538 ();
 sg13g2_fill_1 FILLER_49_554 ();
 sg13g2_fill_2 FILLER_49_561 ();
 sg13g2_fill_1 FILLER_49_563 ();
 sg13g2_fill_1 FILLER_49_572 ();
 sg13g2_fill_2 FILLER_49_592 ();
 sg13g2_fill_1 FILLER_49_594 ();
 sg13g2_decap_4 FILLER_49_622 ();
 sg13g2_fill_2 FILLER_49_639 ();
 sg13g2_fill_1 FILLER_49_652 ();
 sg13g2_decap_4 FILLER_49_667 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_4 FILLER_49_686 ();
 sg13g2_fill_1 FILLER_49_690 ();
 sg13g2_fill_1 FILLER_49_720 ();
 sg13g2_fill_2 FILLER_49_729 ();
 sg13g2_fill_1 FILLER_49_744 ();
 sg13g2_fill_1 FILLER_49_750 ();
 sg13g2_fill_2 FILLER_49_759 ();
 sg13g2_fill_2 FILLER_49_790 ();
 sg13g2_fill_1 FILLER_49_792 ();
 sg13g2_fill_2 FILLER_49_806 ();
 sg13g2_fill_1 FILLER_49_808 ();
 sg13g2_decap_4 FILLER_49_845 ();
 sg13g2_fill_2 FILLER_49_849 ();
 sg13g2_fill_2 FILLER_49_882 ();
 sg13g2_fill_1 FILLER_49_884 ();
 sg13g2_fill_2 FILLER_49_960 ();
 sg13g2_fill_1 FILLER_49_962 ();
 sg13g2_fill_1 FILLER_49_991 ();
 sg13g2_decap_4 FILLER_49_1023 ();
 sg13g2_fill_1 FILLER_49_1027 ();
 sg13g2_decap_8 FILLER_49_1057 ();
 sg13g2_decap_4 FILLER_49_1083 ();
 sg13g2_fill_2 FILLER_49_1106 ();
 sg13g2_decap_4 FILLER_49_1120 ();
 sg13g2_fill_2 FILLER_49_1156 ();
 sg13g2_decap_8 FILLER_49_1167 ();
 sg13g2_fill_2 FILLER_49_1174 ();
 sg13g2_fill_1 FILLER_49_1176 ();
 sg13g2_decap_4 FILLER_49_1199 ();
 sg13g2_fill_2 FILLER_49_1203 ();
 sg13g2_fill_2 FILLER_49_1224 ();
 sg13g2_fill_2 FILLER_49_1235 ();
 sg13g2_fill_2 FILLER_49_1250 ();
 sg13g2_fill_2 FILLER_49_1290 ();
 sg13g2_fill_1 FILLER_49_1292 ();
 sg13g2_fill_2 FILLER_49_1313 ();
 sg13g2_decap_4 FILLER_49_1354 ();
 sg13g2_fill_1 FILLER_49_1362 ();
 sg13g2_decap_8 FILLER_49_1405 ();
 sg13g2_fill_2 FILLER_49_1412 ();
 sg13g2_decap_4 FILLER_49_1421 ();
 sg13g2_fill_2 FILLER_49_1425 ();
 sg13g2_fill_2 FILLER_49_1497 ();
 sg13g2_decap_8 FILLER_49_1502 ();
 sg13g2_decap_8 FILLER_49_1509 ();
 sg13g2_fill_1 FILLER_49_1516 ();
 sg13g2_decap_8 FILLER_49_1592 ();
 sg13g2_fill_1 FILLER_49_1599 ();
 sg13g2_decap_4 FILLER_49_1609 ();
 sg13g2_fill_2 FILLER_49_1613 ();
 sg13g2_decap_4 FILLER_49_1619 ();
 sg13g2_fill_1 FILLER_49_1623 ();
 sg13g2_fill_1 FILLER_49_1664 ();
 sg13g2_fill_2 FILLER_49_1673 ();
 sg13g2_fill_1 FILLER_49_1675 ();
 sg13g2_fill_2 FILLER_49_1687 ();
 sg13g2_fill_1 FILLER_49_1694 ();
 sg13g2_decap_8 FILLER_49_1698 ();
 sg13g2_fill_1 FILLER_49_1705 ();
 sg13g2_decap_4 FILLER_49_1727 ();
 sg13g2_fill_1 FILLER_49_1731 ();
 sg13g2_decap_4 FILLER_49_1753 ();
 sg13g2_fill_1 FILLER_49_1757 ();
 sg13g2_fill_2 FILLER_49_1773 ();
 sg13g2_fill_1 FILLER_49_1775 ();
 sg13g2_decap_4 FILLER_49_1819 ();
 sg13g2_fill_1 FILLER_49_1823 ();
 sg13g2_fill_1 FILLER_49_1888 ();
 sg13g2_decap_4 FILLER_49_1907 ();
 sg13g2_fill_2 FILLER_49_1911 ();
 sg13g2_decap_8 FILLER_49_1917 ();
 sg13g2_fill_1 FILLER_49_1937 ();
 sg13g2_fill_2 FILLER_49_1947 ();
 sg13g2_fill_2 FILLER_49_1957 ();
 sg13g2_decap_8 FILLER_49_1982 ();
 sg13g2_decap_8 FILLER_49_1989 ();
 sg13g2_decap_8 FILLER_49_1996 ();
 sg13g2_fill_1 FILLER_49_2003 ();
 sg13g2_fill_2 FILLER_49_2008 ();
 sg13g2_fill_2 FILLER_49_2042 ();
 sg13g2_fill_1 FILLER_49_2044 ();
 sg13g2_decap_4 FILLER_49_2075 ();
 sg13g2_fill_1 FILLER_49_2162 ();
 sg13g2_fill_1 FILLER_49_2167 ();
 sg13g2_fill_2 FILLER_49_2181 ();
 sg13g2_fill_1 FILLER_49_2207 ();
 sg13g2_decap_4 FILLER_49_2220 ();
 sg13g2_fill_1 FILLER_49_2224 ();
 sg13g2_decap_8 FILLER_49_2232 ();
 sg13g2_fill_1 FILLER_49_2239 ();
 sg13g2_decap_8 FILLER_49_2246 ();
 sg13g2_decap_4 FILLER_49_2253 ();
 sg13g2_fill_1 FILLER_49_2257 ();
 sg13g2_fill_2 FILLER_49_2284 ();
 sg13g2_fill_2 FILLER_49_2300 ();
 sg13g2_fill_1 FILLER_49_2302 ();
 sg13g2_decap_8 FILLER_49_2316 ();
 sg13g2_fill_1 FILLER_49_2323 ();
 sg13g2_fill_2 FILLER_49_2361 ();
 sg13g2_fill_2 FILLER_49_2399 ();
 sg13g2_fill_1 FILLER_49_2419 ();
 sg13g2_decap_8 FILLER_49_2426 ();
 sg13g2_decap_8 FILLER_49_2433 ();
 sg13g2_fill_1 FILLER_49_2440 ();
 sg13g2_fill_2 FILLER_49_2465 ();
 sg13g2_decap_4 FILLER_49_2520 ();
 sg13g2_fill_2 FILLER_49_2524 ();
 sg13g2_decap_8 FILLER_49_2567 ();
 sg13g2_fill_2 FILLER_49_2585 ();
 sg13g2_fill_1 FILLER_49_2587 ();
 sg13g2_decap_4 FILLER_49_2606 ();
 sg13g2_fill_1 FILLER_49_2610 ();
 sg13g2_fill_2 FILLER_49_2620 ();
 sg13g2_fill_1 FILLER_49_2632 ();
 sg13g2_decap_8 FILLER_49_2637 ();
 sg13g2_fill_2 FILLER_49_2644 ();
 sg13g2_fill_2 FILLER_49_2674 ();
 sg13g2_fill_2 FILLER_49_2681 ();
 sg13g2_fill_1 FILLER_49_2696 ();
 sg13g2_fill_2 FILLER_49_2730 ();
 sg13g2_fill_2 FILLER_49_2828 ();
 sg13g2_fill_1 FILLER_49_2830 ();
 sg13g2_decap_4 FILLER_49_2857 ();
 sg13g2_fill_1 FILLER_49_2861 ();
 sg13g2_fill_2 FILLER_49_2898 ();
 sg13g2_fill_2 FILLER_49_2936 ();
 sg13g2_decap_4 FILLER_49_2969 ();
 sg13g2_fill_1 FILLER_49_2973 ();
 sg13g2_fill_2 FILLER_49_2991 ();
 sg13g2_decap_4 FILLER_49_3002 ();
 sg13g2_fill_2 FILLER_49_3006 ();
 sg13g2_fill_2 FILLER_49_3044 ();
 sg13g2_fill_2 FILLER_49_3073 ();
 sg13g2_fill_2 FILLER_49_3103 ();
 sg13g2_fill_1 FILLER_49_3105 ();
 sg13g2_fill_2 FILLER_49_3139 ();
 sg13g2_fill_1 FILLER_49_3141 ();
 sg13g2_fill_2 FILLER_49_3175 ();
 sg13g2_fill_1 FILLER_49_3177 ();
 sg13g2_fill_2 FILLER_49_3228 ();
 sg13g2_fill_1 FILLER_49_3230 ();
 sg13g2_fill_2 FILLER_49_3245 ();
 sg13g2_fill_1 FILLER_49_3247 ();
 sg13g2_fill_2 FILLER_49_3296 ();
 sg13g2_fill_1 FILLER_49_3298 ();
 sg13g2_fill_2 FILLER_49_3340 ();
 sg13g2_fill_1 FILLER_49_3342 ();
 sg13g2_fill_2 FILLER_49_3370 ();
 sg13g2_decap_4 FILLER_49_3405 ();
 sg13g2_fill_2 FILLER_49_3409 ();
 sg13g2_fill_1 FILLER_49_3422 ();
 sg13g2_decap_8 FILLER_49_3451 ();
 sg13g2_decap_8 FILLER_49_3458 ();
 sg13g2_decap_8 FILLER_49_3465 ();
 sg13g2_decap_8 FILLER_49_3472 ();
 sg13g2_decap_8 FILLER_49_3479 ();
 sg13g2_decap_8 FILLER_49_3486 ();
 sg13g2_decap_8 FILLER_49_3493 ();
 sg13g2_decap_8 FILLER_49_3500 ();
 sg13g2_decap_8 FILLER_49_3507 ();
 sg13g2_decap_8 FILLER_49_3514 ();
 sg13g2_decap_8 FILLER_49_3521 ();
 sg13g2_decap_8 FILLER_49_3528 ();
 sg13g2_decap_8 FILLER_49_3535 ();
 sg13g2_decap_8 FILLER_49_3542 ();
 sg13g2_decap_8 FILLER_49_3549 ();
 sg13g2_decap_8 FILLER_49_3556 ();
 sg13g2_decap_8 FILLER_49_3563 ();
 sg13g2_decap_8 FILLER_49_3570 ();
 sg13g2_fill_2 FILLER_49_3577 ();
 sg13g2_fill_1 FILLER_49_3579 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_4 FILLER_50_14 ();
 sg13g2_fill_2 FILLER_50_18 ();
 sg13g2_decap_4 FILLER_50_62 ();
 sg13g2_fill_2 FILLER_50_83 ();
 sg13g2_decap_8 FILLER_50_130 ();
 sg13g2_decap_4 FILLER_50_137 ();
 sg13g2_decap_4 FILLER_50_197 ();
 sg13g2_decap_8 FILLER_50_228 ();
 sg13g2_decap_8 FILLER_50_235 ();
 sg13g2_decap_8 FILLER_50_242 ();
 sg13g2_fill_2 FILLER_50_267 ();
 sg13g2_fill_2 FILLER_50_278 ();
 sg13g2_decap_8 FILLER_50_314 ();
 sg13g2_decap_4 FILLER_50_321 ();
 sg13g2_decap_8 FILLER_50_334 ();
 sg13g2_decap_4 FILLER_50_341 ();
 sg13g2_fill_2 FILLER_50_345 ();
 sg13g2_decap_4 FILLER_50_387 ();
 sg13g2_fill_2 FILLER_50_391 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_1 FILLER_50_409 ();
 sg13g2_fill_1 FILLER_50_438 ();
 sg13g2_fill_1 FILLER_50_453 ();
 sg13g2_decap_8 FILLER_50_477 ();
 sg13g2_decap_4 FILLER_50_484 ();
 sg13g2_fill_1 FILLER_50_493 ();
 sg13g2_decap_8 FILLER_50_501 ();
 sg13g2_decap_8 FILLER_50_508 ();
 sg13g2_decap_4 FILLER_50_515 ();
 sg13g2_fill_2 FILLER_50_519 ();
 sg13g2_decap_8 FILLER_50_529 ();
 sg13g2_decap_8 FILLER_50_536 ();
 sg13g2_fill_1 FILLER_50_551 ();
 sg13g2_fill_1 FILLER_50_574 ();
 sg13g2_fill_1 FILLER_50_596 ();
 sg13g2_fill_1 FILLER_50_607 ();
 sg13g2_fill_2 FILLER_50_671 ();
 sg13g2_decap_4 FILLER_50_689 ();
 sg13g2_decap_4 FILLER_50_716 ();
 sg13g2_fill_1 FILLER_50_720 ();
 sg13g2_decap_4 FILLER_50_724 ();
 sg13g2_fill_2 FILLER_50_745 ();
 sg13g2_fill_1 FILLER_50_747 ();
 sg13g2_fill_2 FILLER_50_752 ();
 sg13g2_fill_1 FILLER_50_754 ();
 sg13g2_fill_1 FILLER_50_759 ();
 sg13g2_decap_4 FILLER_50_766 ();
 sg13g2_fill_2 FILLER_50_778 ();
 sg13g2_fill_1 FILLER_50_780 ();
 sg13g2_decap_8 FILLER_50_786 ();
 sg13g2_decap_8 FILLER_50_793 ();
 sg13g2_fill_1 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_811 ();
 sg13g2_fill_2 FILLER_50_818 ();
 sg13g2_fill_1 FILLER_50_820 ();
 sg13g2_fill_2 FILLER_50_824 ();
 sg13g2_decap_8 FILLER_50_846 ();
 sg13g2_decap_8 FILLER_50_853 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_fill_2 FILLER_50_896 ();
 sg13g2_decap_8 FILLER_50_907 ();
 sg13g2_decap_8 FILLER_50_917 ();
 sg13g2_fill_1 FILLER_50_928 ();
 sg13g2_decap_4 FILLER_50_939 ();
 sg13g2_fill_2 FILLER_50_943 ();
 sg13g2_fill_2 FILLER_50_959 ();
 sg13g2_decap_4 FILLER_50_976 ();
 sg13g2_fill_2 FILLER_50_980 ();
 sg13g2_fill_1 FILLER_50_991 ();
 sg13g2_fill_2 FILLER_50_1030 ();
 sg13g2_decap_4 FILLER_50_1057 ();
 sg13g2_decap_4 FILLER_50_1081 ();
 sg13g2_fill_1 FILLER_50_1085 ();
 sg13g2_decap_8 FILLER_50_1117 ();
 sg13g2_fill_2 FILLER_50_1173 ();
 sg13g2_decap_4 FILLER_50_1179 ();
 sg13g2_fill_2 FILLER_50_1183 ();
 sg13g2_fill_2 FILLER_50_1205 ();
 sg13g2_fill_1 FILLER_50_1207 ();
 sg13g2_fill_2 FILLER_50_1229 ();
 sg13g2_fill_1 FILLER_50_1251 ();
 sg13g2_fill_2 FILLER_50_1270 ();
 sg13g2_fill_1 FILLER_50_1272 ();
 sg13g2_fill_2 FILLER_50_1288 ();
 sg13g2_fill_1 FILLER_50_1290 ();
 sg13g2_decap_8 FILLER_50_1313 ();
 sg13g2_fill_2 FILLER_50_1320 ();
 sg13g2_fill_1 FILLER_50_1322 ();
 sg13g2_decap_4 FILLER_50_1334 ();
 sg13g2_fill_1 FILLER_50_1338 ();
 sg13g2_fill_1 FILLER_50_1344 ();
 sg13g2_fill_1 FILLER_50_1357 ();
 sg13g2_fill_2 FILLER_50_1364 ();
 sg13g2_fill_1 FILLER_50_1366 ();
 sg13g2_fill_1 FILLER_50_1391 ();
 sg13g2_fill_1 FILLER_50_1405 ();
 sg13g2_fill_1 FILLER_50_1411 ();
 sg13g2_fill_2 FILLER_50_1454 ();
 sg13g2_fill_2 FILLER_50_1474 ();
 sg13g2_fill_2 FILLER_50_1504 ();
 sg13g2_fill_2 FILLER_50_1518 ();
 sg13g2_fill_2 FILLER_50_1538 ();
 sg13g2_fill_1 FILLER_50_1540 ();
 sg13g2_decap_8 FILLER_50_1550 ();
 sg13g2_fill_2 FILLER_50_1557 ();
 sg13g2_fill_1 FILLER_50_1559 ();
 sg13g2_fill_1 FILLER_50_1566 ();
 sg13g2_decap_8 FILLER_50_1573 ();
 sg13g2_fill_1 FILLER_50_1596 ();
 sg13g2_decap_4 FILLER_50_1605 ();
 sg13g2_fill_2 FILLER_50_1609 ();
 sg13g2_fill_1 FILLER_50_1661 ();
 sg13g2_fill_2 FILLER_50_1682 ();
 sg13g2_fill_1 FILLER_50_1684 ();
 sg13g2_decap_8 FILLER_50_1698 ();
 sg13g2_fill_2 FILLER_50_1705 ();
 sg13g2_decap_8 FILLER_50_1728 ();
 sg13g2_fill_2 FILLER_50_1735 ();
 sg13g2_fill_1 FILLER_50_1746 ();
 sg13g2_fill_2 FILLER_50_1764 ();
 sg13g2_decap_4 FILLER_50_1775 ();
 sg13g2_fill_1 FILLER_50_1779 ();
 sg13g2_decap_8 FILLER_50_1818 ();
 sg13g2_decap_4 FILLER_50_1825 ();
 sg13g2_decap_8 FILLER_50_1833 ();
 sg13g2_decap_4 FILLER_50_1840 ();
 sg13g2_fill_1 FILLER_50_1850 ();
 sg13g2_fill_1 FILLER_50_1868 ();
 sg13g2_fill_2 FILLER_50_1878 ();
 sg13g2_decap_4 FILLER_50_1884 ();
 sg13g2_fill_1 FILLER_50_1900 ();
 sg13g2_fill_2 FILLER_50_1914 ();
 sg13g2_fill_2 FILLER_50_1930 ();
 sg13g2_fill_1 FILLER_50_1950 ();
 sg13g2_decap_4 FILLER_50_1987 ();
 sg13g2_fill_1 FILLER_50_1991 ();
 sg13g2_fill_2 FILLER_50_1998 ();
 sg13g2_fill_1 FILLER_50_2000 ();
 sg13g2_fill_2 FILLER_50_2015 ();
 sg13g2_fill_1 FILLER_50_2017 ();
 sg13g2_decap_8 FILLER_50_2042 ();
 sg13g2_decap_8 FILLER_50_2072 ();
 sg13g2_fill_2 FILLER_50_2079 ();
 sg13g2_fill_1 FILLER_50_2081 ();
 sg13g2_fill_1 FILLER_50_2110 ();
 sg13g2_fill_2 FILLER_50_2115 ();
 sg13g2_fill_2 FILLER_50_2142 ();
 sg13g2_fill_1 FILLER_50_2158 ();
 sg13g2_fill_1 FILLER_50_2192 ();
 sg13g2_fill_2 FILLER_50_2207 ();
 sg13g2_fill_1 FILLER_50_2209 ();
 sg13g2_fill_2 FILLER_50_2215 ();
 sg13g2_fill_1 FILLER_50_2234 ();
 sg13g2_fill_2 FILLER_50_2270 ();
 sg13g2_fill_1 FILLER_50_2285 ();
 sg13g2_decap_8 FILLER_50_2331 ();
 sg13g2_fill_1 FILLER_50_2338 ();
 sg13g2_decap_8 FILLER_50_2343 ();
 sg13g2_decap_8 FILLER_50_2350 ();
 sg13g2_decap_4 FILLER_50_2357 ();
 sg13g2_fill_1 FILLER_50_2361 ();
 sg13g2_fill_2 FILLER_50_2365 ();
 sg13g2_fill_2 FILLER_50_2412 ();
 sg13g2_fill_1 FILLER_50_2442 ();
 sg13g2_fill_1 FILLER_50_2480 ();
 sg13g2_fill_2 FILLER_50_2505 ();
 sg13g2_fill_2 FILLER_50_2582 ();
 sg13g2_decap_4 FILLER_50_2618 ();
 sg13g2_decap_8 FILLER_50_2693 ();
 sg13g2_decap_8 FILLER_50_2700 ();
 sg13g2_fill_1 FILLER_50_2707 ();
 sg13g2_decap_4 FILLER_50_2743 ();
 sg13g2_fill_1 FILLER_50_2778 ();
 sg13g2_fill_2 FILLER_50_2798 ();
 sg13g2_fill_2 FILLER_50_2896 ();
 sg13g2_fill_1 FILLER_50_2898 ();
 sg13g2_decap_8 FILLER_50_2904 ();
 sg13g2_decap_4 FILLER_50_2911 ();
 sg13g2_fill_1 FILLER_50_2915 ();
 sg13g2_decap_4 FILLER_50_2920 ();
 sg13g2_fill_1 FILLER_50_2924 ();
 sg13g2_decap_4 FILLER_50_2956 ();
 sg13g2_fill_2 FILLER_50_2960 ();
 sg13g2_decap_4 FILLER_50_3003 ();
 sg13g2_fill_1 FILLER_50_3007 ();
 sg13g2_fill_2 FILLER_50_3031 ();
 sg13g2_fill_1 FILLER_50_3042 ();
 sg13g2_decap_8 FILLER_50_3085 ();
 sg13g2_fill_1 FILLER_50_3101 ();
 sg13g2_fill_2 FILLER_50_3156 ();
 sg13g2_fill_1 FILLER_50_3158 ();
 sg13g2_decap_4 FILLER_50_3185 ();
 sg13g2_fill_2 FILLER_50_3189 ();
 sg13g2_fill_1 FILLER_50_3200 ();
 sg13g2_fill_1 FILLER_50_3215 ();
 sg13g2_fill_1 FILLER_50_3221 ();
 sg13g2_fill_1 FILLER_50_3226 ();
 sg13g2_fill_1 FILLER_50_3300 ();
 sg13g2_fill_1 FILLER_50_3329 ();
 sg13g2_fill_2 FILLER_50_3367 ();
 sg13g2_fill_2 FILLER_50_3391 ();
 sg13g2_fill_2 FILLER_50_3415 ();
 sg13g2_fill_1 FILLER_50_3417 ();
 sg13g2_decap_8 FILLER_50_3448 ();
 sg13g2_decap_8 FILLER_50_3483 ();
 sg13g2_decap_8 FILLER_50_3490 ();
 sg13g2_decap_8 FILLER_50_3497 ();
 sg13g2_decap_8 FILLER_50_3504 ();
 sg13g2_decap_8 FILLER_50_3511 ();
 sg13g2_decap_8 FILLER_50_3518 ();
 sg13g2_decap_8 FILLER_50_3525 ();
 sg13g2_decap_8 FILLER_50_3532 ();
 sg13g2_decap_8 FILLER_50_3539 ();
 sg13g2_decap_8 FILLER_50_3546 ();
 sg13g2_decap_8 FILLER_50_3553 ();
 sg13g2_decap_8 FILLER_50_3560 ();
 sg13g2_decap_8 FILLER_50_3567 ();
 sg13g2_decap_4 FILLER_50_3574 ();
 sg13g2_fill_2 FILLER_50_3578 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_4 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_29 ();
 sg13g2_fill_2 FILLER_51_36 ();
 sg13g2_fill_1 FILLER_51_38 ();
 sg13g2_decap_4 FILLER_51_43 ();
 sg13g2_fill_1 FILLER_51_47 ();
 sg13g2_decap_4 FILLER_51_64 ();
 sg13g2_fill_2 FILLER_51_86 ();
 sg13g2_fill_1 FILLER_51_93 ();
 sg13g2_decap_8 FILLER_51_104 ();
 sg13g2_decap_8 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_118 ();
 sg13g2_decap_4 FILLER_51_129 ();
 sg13g2_fill_2 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_151 ();
 sg13g2_fill_1 FILLER_51_162 ();
 sg13g2_fill_2 FILLER_51_183 ();
 sg13g2_fill_1 FILLER_51_217 ();
 sg13g2_fill_2 FILLER_51_233 ();
 sg13g2_fill_1 FILLER_51_235 ();
 sg13g2_decap_8 FILLER_51_287 ();
 sg13g2_decap_4 FILLER_51_294 ();
 sg13g2_fill_2 FILLER_51_305 ();
 sg13g2_fill_1 FILLER_51_363 ();
 sg13g2_fill_1 FILLER_51_373 ();
 sg13g2_fill_1 FILLER_51_414 ();
 sg13g2_fill_1 FILLER_51_419 ();
 sg13g2_fill_2 FILLER_51_424 ();
 sg13g2_fill_2 FILLER_51_449 ();
 sg13g2_decap_4 FILLER_51_459 ();
 sg13g2_fill_2 FILLER_51_463 ();
 sg13g2_decap_4 FILLER_51_473 ();
 sg13g2_fill_2 FILLER_51_477 ();
 sg13g2_decap_8 FILLER_51_484 ();
 sg13g2_fill_1 FILLER_51_491 ();
 sg13g2_decap_4 FILLER_51_525 ();
 sg13g2_decap_8 FILLER_51_545 ();
 sg13g2_decap_4 FILLER_51_589 ();
 sg13g2_fill_1 FILLER_51_593 ();
 sg13g2_decap_4 FILLER_51_622 ();
 sg13g2_fill_2 FILLER_51_626 ();
 sg13g2_fill_2 FILLER_51_638 ();
 sg13g2_fill_1 FILLER_51_640 ();
 sg13g2_fill_2 FILLER_51_650 ();
 sg13g2_fill_1 FILLER_51_657 ();
 sg13g2_fill_2 FILLER_51_673 ();
 sg13g2_decap_4 FILLER_51_693 ();
 sg13g2_fill_1 FILLER_51_697 ();
 sg13g2_fill_1 FILLER_51_722 ();
 sg13g2_fill_2 FILLER_51_757 ();
 sg13g2_fill_1 FILLER_51_759 ();
 sg13g2_fill_1 FILLER_51_778 ();
 sg13g2_fill_2 FILLER_51_791 ();
 sg13g2_decap_4 FILLER_51_819 ();
 sg13g2_fill_1 FILLER_51_823 ();
 sg13g2_decap_4 FILLER_51_831 ();
 sg13g2_fill_1 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_fill_1 FILLER_51_862 ();
 sg13g2_fill_1 FILLER_51_886 ();
 sg13g2_fill_1 FILLER_51_914 ();
 sg13g2_decap_8 FILLER_51_948 ();
 sg13g2_decap_8 FILLER_51_955 ();
 sg13g2_fill_2 FILLER_51_962 ();
 sg13g2_fill_1 FILLER_51_964 ();
 sg13g2_decap_8 FILLER_51_982 ();
 sg13g2_fill_2 FILLER_51_989 ();
 sg13g2_fill_1 FILLER_51_991 ();
 sg13g2_decap_4 FILLER_51_995 ();
 sg13g2_fill_1 FILLER_51_999 ();
 sg13g2_decap_8 FILLER_51_1027 ();
 sg13g2_fill_1 FILLER_51_1034 ();
 sg13g2_decap_4 FILLER_51_1051 ();
 sg13g2_fill_1 FILLER_51_1055 ();
 sg13g2_fill_2 FILLER_51_1061 ();
 sg13g2_fill_2 FILLER_51_1069 ();
 sg13g2_fill_1 FILLER_51_1071 ();
 sg13g2_decap_4 FILLER_51_1078 ();
 sg13g2_fill_1 FILLER_51_1082 ();
 sg13g2_fill_2 FILLER_51_1093 ();
 sg13g2_fill_1 FILLER_51_1095 ();
 sg13g2_fill_2 FILLER_51_1113 ();
 sg13g2_fill_1 FILLER_51_1134 ();
 sg13g2_fill_1 FILLER_51_1149 ();
 sg13g2_decap_4 FILLER_51_1163 ();
 sg13g2_fill_2 FILLER_51_1167 ();
 sg13g2_decap_8 FILLER_51_1197 ();
 sg13g2_decap_8 FILLER_51_1204 ();
 sg13g2_fill_1 FILLER_51_1224 ();
 sg13g2_fill_2 FILLER_51_1230 ();
 sg13g2_fill_1 FILLER_51_1232 ();
 sg13g2_decap_4 FILLER_51_1242 ();
 sg13g2_fill_1 FILLER_51_1246 ();
 sg13g2_decap_8 FILLER_51_1251 ();
 sg13g2_fill_2 FILLER_51_1258 ();
 sg13g2_fill_1 FILLER_51_1260 ();
 sg13g2_fill_2 FILLER_51_1269 ();
 sg13g2_fill_1 FILLER_51_1271 ();
 sg13g2_fill_1 FILLER_51_1282 ();
 sg13g2_decap_8 FILLER_51_1288 ();
 sg13g2_fill_2 FILLER_51_1295 ();
 sg13g2_fill_1 FILLER_51_1297 ();
 sg13g2_decap_8 FILLER_51_1303 ();
 sg13g2_decap_4 FILLER_51_1310 ();
 sg13g2_fill_1 FILLER_51_1318 ();
 sg13g2_fill_2 FILLER_51_1338 ();
 sg13g2_decap_8 FILLER_51_1354 ();
 sg13g2_fill_2 FILLER_51_1381 ();
 sg13g2_fill_2 FILLER_51_1396 ();
 sg13g2_decap_8 FILLER_51_1418 ();
 sg13g2_decap_8 FILLER_51_1425 ();
 sg13g2_fill_1 FILLER_51_1453 ();
 sg13g2_fill_2 FILLER_51_1476 ();
 sg13g2_fill_1 FILLER_51_1478 ();
 sg13g2_fill_2 FILLER_51_1490 ();
 sg13g2_decap_8 FILLER_51_1504 ();
 sg13g2_fill_1 FILLER_51_1511 ();
 sg13g2_fill_1 FILLER_51_1527 ();
 sg13g2_decap_4 FILLER_51_1548 ();
 sg13g2_fill_2 FILLER_51_1560 ();
 sg13g2_decap_4 FILLER_51_1603 ();
 sg13g2_fill_1 FILLER_51_1617 ();
 sg13g2_fill_1 FILLER_51_1623 ();
 sg13g2_fill_2 FILLER_51_1637 ();
 sg13g2_fill_2 FILLER_51_1653 ();
 sg13g2_decap_4 FILLER_51_1668 ();
 sg13g2_fill_1 FILLER_51_1672 ();
 sg13g2_fill_2 FILLER_51_1677 ();
 sg13g2_fill_1 FILLER_51_1679 ();
 sg13g2_fill_2 FILLER_51_1705 ();
 sg13g2_fill_1 FILLER_51_1707 ();
 sg13g2_decap_8 FILLER_51_1719 ();
 sg13g2_fill_2 FILLER_51_1726 ();
 sg13g2_fill_1 FILLER_51_1732 ();
 sg13g2_fill_1 FILLER_51_1745 ();
 sg13g2_fill_1 FILLER_51_1756 ();
 sg13g2_decap_8 FILLER_51_1780 ();
 sg13g2_decap_8 FILLER_51_1787 ();
 sg13g2_fill_1 FILLER_51_1815 ();
 sg13g2_decap_4 FILLER_51_1831 ();
 sg13g2_fill_1 FILLER_51_1835 ();
 sg13g2_decap_4 FILLER_51_1839 ();
 sg13g2_decap_8 FILLER_51_1849 ();
 sg13g2_fill_1 FILLER_51_1909 ();
 sg13g2_fill_1 FILLER_51_1959 ();
 sg13g2_fill_1 FILLER_51_1965 ();
 sg13g2_decap_4 FILLER_51_1970 ();
 sg13g2_fill_2 FILLER_51_1974 ();
 sg13g2_fill_1 FILLER_51_1981 ();
 sg13g2_decap_8 FILLER_51_1988 ();
 sg13g2_fill_1 FILLER_51_2014 ();
 sg13g2_fill_2 FILLER_51_2020 ();
 sg13g2_fill_1 FILLER_51_2022 ();
 sg13g2_fill_2 FILLER_51_2053 ();
 sg13g2_decap_8 FILLER_51_2059 ();
 sg13g2_fill_2 FILLER_51_2066 ();
 sg13g2_fill_2 FILLER_51_2095 ();
 sg13g2_decap_4 FILLER_51_2117 ();
 sg13g2_decap_4 FILLER_51_2140 ();
 sg13g2_decap_8 FILLER_51_2148 ();
 sg13g2_fill_2 FILLER_51_2155 ();
 sg13g2_fill_1 FILLER_51_2157 ();
 sg13g2_decap_4 FILLER_51_2170 ();
 sg13g2_decap_4 FILLER_51_2220 ();
 sg13g2_fill_2 FILLER_51_2224 ();
 sg13g2_decap_4 FILLER_51_2231 ();
 sg13g2_fill_2 FILLER_51_2235 ();
 sg13g2_decap_8 FILLER_51_2247 ();
 sg13g2_fill_2 FILLER_51_2254 ();
 sg13g2_fill_1 FILLER_51_2256 ();
 sg13g2_decap_8 FILLER_51_2280 ();
 sg13g2_decap_8 FILLER_51_2287 ();
 sg13g2_decap_8 FILLER_51_2294 ();
 sg13g2_fill_1 FILLER_51_2326 ();
 sg13g2_fill_1 FILLER_51_2389 ();
 sg13g2_fill_2 FILLER_51_2404 ();
 sg13g2_fill_2 FILLER_51_2440 ();
 sg13g2_fill_1 FILLER_51_2464 ();
 sg13g2_fill_2 FILLER_51_2473 ();
 sg13g2_fill_1 FILLER_51_2475 ();
 sg13g2_fill_2 FILLER_51_2501 ();
 sg13g2_fill_1 FILLER_51_2503 ();
 sg13g2_decap_8 FILLER_51_2518 ();
 sg13g2_fill_2 FILLER_51_2547 ();
 sg13g2_decap_4 FILLER_51_2573 ();
 sg13g2_fill_1 FILLER_51_2586 ();
 sg13g2_decap_8 FILLER_51_2606 ();
 sg13g2_decap_8 FILLER_51_2613 ();
 sg13g2_fill_2 FILLER_51_2620 ();
 sg13g2_fill_1 FILLER_51_2632 ();
 sg13g2_decap_8 FILLER_51_2636 ();
 sg13g2_fill_2 FILLER_51_2643 ();
 sg13g2_fill_2 FILLER_51_2672 ();
 sg13g2_fill_1 FILLER_51_2674 ();
 sg13g2_decap_4 FILLER_51_2721 ();
 sg13g2_fill_1 FILLER_51_2725 ();
 sg13g2_decap_8 FILLER_51_2793 ();
 sg13g2_fill_2 FILLER_51_2800 ();
 sg13g2_fill_1 FILLER_51_2802 ();
 sg13g2_decap_8 FILLER_51_2835 ();
 sg13g2_fill_1 FILLER_51_2842 ();
 sg13g2_fill_1 FILLER_51_2877 ();
 sg13g2_fill_1 FILLER_51_2892 ();
 sg13g2_fill_2 FILLER_51_2932 ();
 sg13g2_fill_1 FILLER_51_2940 ();
 sg13g2_fill_2 FILLER_51_2953 ();
 sg13g2_decap_4 FILLER_51_2975 ();
 sg13g2_fill_2 FILLER_51_2979 ();
 sg13g2_decap_4 FILLER_51_3012 ();
 sg13g2_fill_1 FILLER_51_3016 ();
 sg13g2_fill_2 FILLER_51_3044 ();
 sg13g2_fill_2 FILLER_51_3064 ();
 sg13g2_fill_2 FILLER_51_3143 ();
 sg13g2_decap_4 FILLER_51_3177 ();
 sg13g2_fill_1 FILLER_51_3181 ();
 sg13g2_fill_1 FILLER_51_3209 ();
 sg13g2_fill_2 FILLER_51_3219 ();
 sg13g2_decap_8 FILLER_51_3249 ();
 sg13g2_decap_4 FILLER_51_3256 ();
 sg13g2_fill_1 FILLER_51_3260 ();
 sg13g2_fill_1 FILLER_51_3311 ();
 sg13g2_fill_1 FILLER_51_3447 ();
 sg13g2_decap_4 FILLER_51_3454 ();
 sg13g2_fill_2 FILLER_51_3458 ();
 sg13g2_decap_8 FILLER_51_3464 ();
 sg13g2_decap_8 FILLER_51_3471 ();
 sg13g2_decap_4 FILLER_51_3478 ();
 sg13g2_fill_2 FILLER_51_3482 ();
 sg13g2_decap_4 FILLER_51_3500 ();
 sg13g2_decap_8 FILLER_51_3513 ();
 sg13g2_decap_8 FILLER_51_3520 ();
 sg13g2_decap_8 FILLER_51_3527 ();
 sg13g2_decap_8 FILLER_51_3534 ();
 sg13g2_decap_8 FILLER_51_3541 ();
 sg13g2_decap_8 FILLER_51_3548 ();
 sg13g2_decap_8 FILLER_51_3555 ();
 sg13g2_decap_8 FILLER_51_3562 ();
 sg13g2_decap_8 FILLER_51_3569 ();
 sg13g2_decap_4 FILLER_51_3576 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_9 ();
 sg13g2_fill_2 FILLER_52_38 ();
 sg13g2_decap_8 FILLER_52_50 ();
 sg13g2_fill_1 FILLER_52_76 ();
 sg13g2_decap_8 FILLER_52_103 ();
 sg13g2_fill_2 FILLER_52_110 ();
 sg13g2_decap_8 FILLER_52_129 ();
 sg13g2_decap_4 FILLER_52_136 ();
 sg13g2_fill_1 FILLER_52_140 ();
 sg13g2_fill_2 FILLER_52_165 ();
 sg13g2_decap_4 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_206 ();
 sg13g2_fill_2 FILLER_52_231 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_263 ();
 sg13g2_fill_2 FILLER_52_306 ();
 sg13g2_decap_8 FILLER_52_327 ();
 sg13g2_decap_4 FILLER_52_334 ();
 sg13g2_fill_2 FILLER_52_338 ();
 sg13g2_decap_8 FILLER_52_344 ();
 sg13g2_decap_8 FILLER_52_351 ();
 sg13g2_fill_2 FILLER_52_358 ();
 sg13g2_decap_8 FILLER_52_373 ();
 sg13g2_decap_4 FILLER_52_380 ();
 sg13g2_fill_1 FILLER_52_384 ();
 sg13g2_fill_2 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_397 ();
 sg13g2_fill_2 FILLER_52_404 ();
 sg13g2_decap_4 FILLER_52_454 ();
 sg13g2_fill_2 FILLER_52_458 ();
 sg13g2_fill_1 FILLER_52_468 ();
 sg13g2_fill_2 FILLER_52_482 ();
 sg13g2_fill_1 FILLER_52_484 ();
 sg13g2_fill_1 FILLER_52_507 ();
 sg13g2_fill_2 FILLER_52_517 ();
 sg13g2_decap_8 FILLER_52_541 ();
 sg13g2_fill_2 FILLER_52_548 ();
 sg13g2_fill_2 FILLER_52_614 ();
 sg13g2_fill_1 FILLER_52_616 ();
 sg13g2_decap_4 FILLER_52_625 ();
 sg13g2_fill_1 FILLER_52_629 ();
 sg13g2_decap_8 FILLER_52_634 ();
 sg13g2_fill_2 FILLER_52_641 ();
 sg13g2_fill_1 FILLER_52_652 ();
 sg13g2_fill_1 FILLER_52_659 ();
 sg13g2_decap_8 FILLER_52_668 ();
 sg13g2_fill_2 FILLER_52_675 ();
 sg13g2_decap_4 FILLER_52_692 ();
 sg13g2_fill_1 FILLER_52_696 ();
 sg13g2_fill_1 FILLER_52_716 ();
 sg13g2_fill_2 FILLER_52_726 ();
 sg13g2_decap_8 FILLER_52_755 ();
 sg13g2_fill_2 FILLER_52_762 ();
 sg13g2_fill_1 FILLER_52_764 ();
 sg13g2_fill_2 FILLER_52_808 ();
 sg13g2_decap_8 FILLER_52_818 ();
 sg13g2_fill_2 FILLER_52_825 ();
 sg13g2_fill_2 FILLER_52_835 ();
 sg13g2_decap_8 FILLER_52_845 ();
 sg13g2_fill_1 FILLER_52_855 ();
 sg13g2_decap_4 FILLER_52_861 ();
 sg13g2_fill_2 FILLER_52_865 ();
 sg13g2_fill_2 FILLER_52_880 ();
 sg13g2_fill_1 FILLER_52_915 ();
 sg13g2_fill_2 FILLER_52_934 ();
 sg13g2_fill_1 FILLER_52_936 ();
 sg13g2_fill_2 FILLER_52_942 ();
 sg13g2_fill_1 FILLER_52_944 ();
 sg13g2_fill_2 FILLER_52_953 ();
 sg13g2_fill_1 FILLER_52_955 ();
 sg13g2_decap_8 FILLER_52_974 ();
 sg13g2_fill_1 FILLER_52_981 ();
 sg13g2_decap_8 FILLER_52_1028 ();
 sg13g2_fill_1 FILLER_52_1035 ();
 sg13g2_decap_8 FILLER_52_1041 ();
 sg13g2_decap_4 FILLER_52_1048 ();
 sg13g2_fill_2 FILLER_52_1064 ();
 sg13g2_fill_2 FILLER_52_1093 ();
 sg13g2_fill_1 FILLER_52_1095 ();
 sg13g2_fill_1 FILLER_52_1123 ();
 sg13g2_fill_1 FILLER_52_1153 ();
 sg13g2_decap_4 FILLER_52_1162 ();
 sg13g2_fill_1 FILLER_52_1166 ();
 sg13g2_decap_4 FILLER_52_1180 ();
 sg13g2_fill_2 FILLER_52_1184 ();
 sg13g2_fill_2 FILLER_52_1190 ();
 sg13g2_fill_1 FILLER_52_1219 ();
 sg13g2_fill_2 FILLER_52_1241 ();
 sg13g2_fill_2 FILLER_52_1266 ();
 sg13g2_decap_8 FILLER_52_1280 ();
 sg13g2_fill_1 FILLER_52_1287 ();
 sg13g2_fill_2 FILLER_52_1314 ();
 sg13g2_fill_2 FILLER_52_1334 ();
 sg13g2_fill_2 FILLER_52_1341 ();
 sg13g2_fill_1 FILLER_52_1343 ();
 sg13g2_fill_1 FILLER_52_1356 ();
 sg13g2_fill_1 FILLER_52_1377 ();
 sg13g2_fill_2 FILLER_52_1386 ();
 sg13g2_decap_4 FILLER_52_1392 ();
 sg13g2_decap_4 FILLER_52_1401 ();
 sg13g2_fill_2 FILLER_52_1405 ();
 sg13g2_decap_4 FILLER_52_1462 ();
 sg13g2_fill_2 FILLER_52_1466 ();
 sg13g2_fill_1 FILLER_52_1485 ();
 sg13g2_fill_1 FILLER_52_1510 ();
 sg13g2_fill_2 FILLER_52_1531 ();
 sg13g2_fill_1 FILLER_52_1564 ();
 sg13g2_fill_1 FILLER_52_1577 ();
 sg13g2_decap_8 FILLER_52_1589 ();
 sg13g2_decap_8 FILLER_52_1596 ();
 sg13g2_decap_8 FILLER_52_1603 ();
 sg13g2_fill_2 FILLER_52_1610 ();
 sg13g2_fill_1 FILLER_52_1612 ();
 sg13g2_fill_1 FILLER_52_1623 ();
 sg13g2_decap_8 FILLER_52_1629 ();
 sg13g2_fill_2 FILLER_52_1644 ();
 sg13g2_fill_1 FILLER_52_1646 ();
 sg13g2_decap_8 FILLER_52_1651 ();
 sg13g2_decap_8 FILLER_52_1663 ();
 sg13g2_decap_4 FILLER_52_1670 ();
 sg13g2_fill_1 FILLER_52_1674 ();
 sg13g2_fill_2 FILLER_52_1690 ();
 sg13g2_decap_4 FILLER_52_1723 ();
 sg13g2_fill_2 FILLER_52_1727 ();
 sg13g2_fill_2 FILLER_52_1735 ();
 sg13g2_fill_1 FILLER_52_1737 ();
 sg13g2_fill_1 FILLER_52_1750 ();
 sg13g2_decap_8 FILLER_52_1757 ();
 sg13g2_fill_2 FILLER_52_1764 ();
 sg13g2_fill_2 FILLER_52_1770 ();
 sg13g2_decap_8 FILLER_52_1784 ();
 sg13g2_decap_4 FILLER_52_1791 ();
 sg13g2_fill_1 FILLER_52_1795 ();
 sg13g2_fill_2 FILLER_52_1809 ();
 sg13g2_decap_8 FILLER_52_1852 ();
 sg13g2_fill_2 FILLER_52_1859 ();
 sg13g2_decap_8 FILLER_52_1877 ();
 sg13g2_fill_2 FILLER_52_1884 ();
 sg13g2_decap_8 FILLER_52_1901 ();
 sg13g2_decap_8 FILLER_52_1908 ();
 sg13g2_decap_8 FILLER_52_1927 ();
 sg13g2_decap_4 FILLER_52_1934 ();
 sg13g2_fill_1 FILLER_52_1938 ();
 sg13g2_decap_4 FILLER_52_1962 ();
 sg13g2_decap_8 FILLER_52_1989 ();
 sg13g2_fill_2 FILLER_52_1996 ();
 sg13g2_fill_1 FILLER_52_1998 ();
 sg13g2_fill_2 FILLER_52_2004 ();
 sg13g2_fill_1 FILLER_52_2006 ();
 sg13g2_decap_8 FILLER_52_2020 ();
 sg13g2_decap_4 FILLER_52_2027 ();
 sg13g2_fill_1 FILLER_52_2031 ();
 sg13g2_fill_2 FILLER_52_2037 ();
 sg13g2_fill_1 FILLER_52_2039 ();
 sg13g2_fill_1 FILLER_52_2054 ();
 sg13g2_fill_2 FILLER_52_2064 ();
 sg13g2_fill_1 FILLER_52_2066 ();
 sg13g2_fill_2 FILLER_52_2072 ();
 sg13g2_fill_2 FILLER_52_2082 ();
 sg13g2_fill_2 FILLER_52_2099 ();
 sg13g2_fill_2 FILLER_52_2109 ();
 sg13g2_fill_1 FILLER_52_2111 ();
 sg13g2_decap_4 FILLER_52_2132 ();
 sg13g2_fill_1 FILLER_52_2136 ();
 sg13g2_decap_8 FILLER_52_2169 ();
 sg13g2_decap_4 FILLER_52_2198 ();
 sg13g2_fill_1 FILLER_52_2202 ();
 sg13g2_decap_8 FILLER_52_2211 ();
 sg13g2_fill_1 FILLER_52_2235 ();
 sg13g2_decap_8 FILLER_52_2255 ();
 sg13g2_decap_8 FILLER_52_2262 ();
 sg13g2_fill_2 FILLER_52_2269 ();
 sg13g2_decap_8 FILLER_52_2306 ();
 sg13g2_decap_8 FILLER_52_2313 ();
 sg13g2_fill_2 FILLER_52_2320 ();
 sg13g2_fill_1 FILLER_52_2322 ();
 sg13g2_fill_1 FILLER_52_2331 ();
 sg13g2_fill_2 FILLER_52_2349 ();
 sg13g2_fill_2 FILLER_52_2378 ();
 sg13g2_fill_1 FILLER_52_2380 ();
 sg13g2_decap_8 FILLER_52_2419 ();
 sg13g2_decap_4 FILLER_52_2426 ();
 sg13g2_fill_2 FILLER_52_2430 ();
 sg13g2_decap_4 FILLER_52_2447 ();
 sg13g2_decap_4 FILLER_52_2474 ();
 sg13g2_fill_2 FILLER_52_2497 ();
 sg13g2_fill_1 FILLER_52_2499 ();
 sg13g2_decap_4 FILLER_52_2512 ();
 sg13g2_decap_4 FILLER_52_2524 ();
 sg13g2_fill_1 FILLER_52_2536 ();
 sg13g2_decap_8 FILLER_52_2542 ();
 sg13g2_decap_8 FILLER_52_2549 ();
 sg13g2_decap_4 FILLER_52_2556 ();
 sg13g2_fill_2 FILLER_52_2579 ();
 sg13g2_fill_1 FILLER_52_2581 ();
 sg13g2_decap_4 FILLER_52_2605 ();
 sg13g2_fill_1 FILLER_52_2609 ();
 sg13g2_fill_2 FILLER_52_2635 ();
 sg13g2_fill_1 FILLER_52_2637 ();
 sg13g2_decap_8 FILLER_52_2681 ();
 sg13g2_fill_1 FILLER_52_2693 ();
 sg13g2_fill_1 FILLER_52_2703 ();
 sg13g2_decap_8 FILLER_52_2718 ();
 sg13g2_fill_2 FILLER_52_2725 ();
 sg13g2_decap_8 FILLER_52_2735 ();
 sg13g2_decap_8 FILLER_52_2742 ();
 sg13g2_fill_2 FILLER_52_2749 ();
 sg13g2_fill_1 FILLER_52_2751 ();
 sg13g2_fill_1 FILLER_52_2756 ();
 sg13g2_fill_2 FILLER_52_2772 ();
 sg13g2_decap_4 FILLER_52_2801 ();
 sg13g2_decap_8 FILLER_52_2817 ();
 sg13g2_decap_4 FILLER_52_2824 ();
 sg13g2_fill_1 FILLER_52_2828 ();
 sg13g2_decap_8 FILLER_52_2875 ();
 sg13g2_decap_4 FILLER_52_2882 ();
 sg13g2_fill_2 FILLER_52_2886 ();
 sg13g2_fill_2 FILLER_52_2900 ();
 sg13g2_decap_8 FILLER_52_2931 ();
 sg13g2_fill_1 FILLER_52_2938 ();
 sg13g2_decap_4 FILLER_52_2954 ();
 sg13g2_fill_2 FILLER_52_2958 ();
 sg13g2_fill_2 FILLER_52_2976 ();
 sg13g2_fill_2 FILLER_52_2987 ();
 sg13g2_fill_1 FILLER_52_2993 ();
 sg13g2_decap_4 FILLER_52_3021 ();
 sg13g2_fill_2 FILLER_52_3025 ();
 sg13g2_decap_4 FILLER_52_3031 ();
 sg13g2_fill_2 FILLER_52_3035 ();
 sg13g2_fill_1 FILLER_52_3046 ();
 sg13g2_fill_1 FILLER_52_3089 ();
 sg13g2_decap_4 FILLER_52_3103 ();
 sg13g2_fill_1 FILLER_52_3120 ();
 sg13g2_decap_8 FILLER_52_3175 ();
 sg13g2_decap_8 FILLER_52_3182 ();
 sg13g2_fill_1 FILLER_52_3189 ();
 sg13g2_fill_1 FILLER_52_3204 ();
 sg13g2_decap_8 FILLER_52_3218 ();
 sg13g2_fill_1 FILLER_52_3225 ();
 sg13g2_decap_4 FILLER_52_3239 ();
 sg13g2_fill_2 FILLER_52_3275 ();
 sg13g2_fill_1 FILLER_52_3277 ();
 sg13g2_fill_1 FILLER_52_3304 ();
 sg13g2_decap_4 FILLER_52_3336 ();
 sg13g2_decap_8 FILLER_52_3414 ();
 sg13g2_fill_2 FILLER_52_3438 ();
 sg13g2_fill_2 FILLER_52_3449 ();
 sg13g2_fill_1 FILLER_52_3451 ();
 sg13g2_fill_1 FILLER_52_3489 ();
 sg13g2_decap_8 FILLER_52_3518 ();
 sg13g2_decap_8 FILLER_52_3525 ();
 sg13g2_decap_8 FILLER_52_3532 ();
 sg13g2_decap_8 FILLER_52_3539 ();
 sg13g2_decap_8 FILLER_52_3546 ();
 sg13g2_decap_8 FILLER_52_3553 ();
 sg13g2_decap_8 FILLER_52_3560 ();
 sg13g2_decap_8 FILLER_52_3567 ();
 sg13g2_decap_4 FILLER_52_3574 ();
 sg13g2_fill_2 FILLER_52_3578 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_19 ();
 sg13g2_fill_1 FILLER_53_26 ();
 sg13g2_fill_1 FILLER_53_46 ();
 sg13g2_fill_2 FILLER_53_68 ();
 sg13g2_decap_4 FILLER_53_87 ();
 sg13g2_fill_1 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_138 ();
 sg13g2_decap_8 FILLER_53_163 ();
 sg13g2_fill_2 FILLER_53_170 ();
 sg13g2_decap_8 FILLER_53_181 ();
 sg13g2_fill_1 FILLER_53_188 ();
 sg13g2_decap_4 FILLER_53_207 ();
 sg13g2_fill_1 FILLER_53_211 ();
 sg13g2_fill_1 FILLER_53_225 ();
 sg13g2_fill_1 FILLER_53_238 ();
 sg13g2_decap_4 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_decap_8 FILLER_53_275 ();
 sg13g2_fill_2 FILLER_53_287 ();
 sg13g2_fill_1 FILLER_53_316 ();
 sg13g2_decap_8 FILLER_53_325 ();
 sg13g2_fill_2 FILLER_53_332 ();
 sg13g2_fill_1 FILLER_53_341 ();
 sg13g2_decap_4 FILLER_53_355 ();
 sg13g2_fill_1 FILLER_53_359 ();
 sg13g2_fill_2 FILLER_53_380 ();
 sg13g2_fill_1 FILLER_53_382 ();
 sg13g2_decap_8 FILLER_53_401 ();
 sg13g2_fill_2 FILLER_53_408 ();
 sg13g2_fill_1 FILLER_53_410 ();
 sg13g2_fill_2 FILLER_53_424 ();
 sg13g2_decap_4 FILLER_53_434 ();
 sg13g2_fill_1 FILLER_53_438 ();
 sg13g2_fill_1 FILLER_53_443 ();
 sg13g2_decap_4 FILLER_53_447 ();
 sg13g2_fill_1 FILLER_53_455 ();
 sg13g2_fill_2 FILLER_53_475 ();
 sg13g2_fill_1 FILLER_53_482 ();
 sg13g2_fill_1 FILLER_53_508 ();
 sg13g2_fill_1 FILLER_53_521 ();
 sg13g2_fill_1 FILLER_53_527 ();
 sg13g2_fill_2 FILLER_53_565 ();
 sg13g2_fill_1 FILLER_53_567 ();
 sg13g2_fill_2 FILLER_53_595 ();
 sg13g2_decap_8 FILLER_53_615 ();
 sg13g2_fill_2 FILLER_53_622 ();
 sg13g2_fill_1 FILLER_53_624 ();
 sg13g2_fill_2 FILLER_53_653 ();
 sg13g2_fill_1 FILLER_53_655 ();
 sg13g2_fill_1 FILLER_53_665 ();
 sg13g2_decap_4 FILLER_53_676 ();
 sg13g2_fill_2 FILLER_53_680 ();
 sg13g2_fill_2 FILLER_53_685 ();
 sg13g2_decap_8 FILLER_53_691 ();
 sg13g2_decap_8 FILLER_53_698 ();
 sg13g2_fill_1 FILLER_53_705 ();
 sg13g2_fill_2 FILLER_53_737 ();
 sg13g2_fill_1 FILLER_53_739 ();
 sg13g2_decap_4 FILLER_53_749 ();
 sg13g2_fill_1 FILLER_53_753 ();
 sg13g2_fill_2 FILLER_53_763 ();
 sg13g2_fill_1 FILLER_53_765 ();
 sg13g2_fill_1 FILLER_53_774 ();
 sg13g2_fill_2 FILLER_53_788 ();
 sg13g2_decap_8 FILLER_53_840 ();
 sg13g2_fill_2 FILLER_53_847 ();
 sg13g2_fill_1 FILLER_53_849 ();
 sg13g2_fill_1 FILLER_53_859 ();
 sg13g2_decap_8 FILLER_53_882 ();
 sg13g2_fill_2 FILLER_53_889 ();
 sg13g2_fill_1 FILLER_53_891 ();
 sg13g2_decap_8 FILLER_53_907 ();
 sg13g2_decap_8 FILLER_53_914 ();
 sg13g2_fill_1 FILLER_53_921 ();
 sg13g2_fill_1 FILLER_53_961 ();
 sg13g2_decap_4 FILLER_53_1009 ();
 sg13g2_decap_4 FILLER_53_1047 ();
 sg13g2_fill_2 FILLER_53_1051 ();
 sg13g2_fill_1 FILLER_53_1058 ();
 sg13g2_fill_2 FILLER_53_1090 ();
 sg13g2_fill_1 FILLER_53_1097 ();
 sg13g2_decap_8 FILLER_53_1106 ();
 sg13g2_decap_4 FILLER_53_1113 ();
 sg13g2_fill_1 FILLER_53_1117 ();
 sg13g2_fill_1 FILLER_53_1123 ();
 sg13g2_fill_1 FILLER_53_1180 ();
 sg13g2_decap_8 FILLER_53_1223 ();
 sg13g2_decap_4 FILLER_53_1230 ();
 sg13g2_decap_8 FILLER_53_1252 ();
 sg13g2_decap_8 FILLER_53_1259 ();
 sg13g2_fill_2 FILLER_53_1266 ();
 sg13g2_fill_1 FILLER_53_1268 ();
 sg13g2_decap_4 FILLER_53_1285 ();
 sg13g2_fill_2 FILLER_53_1289 ();
 sg13g2_fill_1 FILLER_53_1299 ();
 sg13g2_fill_1 FILLER_53_1310 ();
 sg13g2_fill_2 FILLER_53_1315 ();
 sg13g2_fill_1 FILLER_53_1317 ();
 sg13g2_decap_8 FILLER_53_1331 ();
 sg13g2_decap_4 FILLER_53_1338 ();
 sg13g2_fill_1 FILLER_53_1342 ();
 sg13g2_fill_2 FILLER_53_1347 ();
 sg13g2_decap_4 FILLER_53_1353 ();
 sg13g2_fill_2 FILLER_53_1402 ();
 sg13g2_fill_1 FILLER_53_1404 ();
 sg13g2_decap_4 FILLER_53_1418 ();
 sg13g2_fill_2 FILLER_53_1422 ();
 sg13g2_decap_8 FILLER_53_1429 ();
 sg13g2_fill_2 FILLER_53_1436 ();
 sg13g2_fill_1 FILLER_53_1438 ();
 sg13g2_decap_8 FILLER_53_1472 ();
 sg13g2_fill_1 FILLER_53_1479 ();
 sg13g2_fill_2 FILLER_53_1489 ();
 sg13g2_fill_1 FILLER_53_1496 ();
 sg13g2_decap_4 FILLER_53_1510 ();
 sg13g2_fill_1 FILLER_53_1514 ();
 sg13g2_fill_1 FILLER_53_1528 ();
 sg13g2_decap_4 FILLER_53_1534 ();
 sg13g2_decap_8 FILLER_53_1542 ();
 sg13g2_fill_2 FILLER_53_1549 ();
 sg13g2_fill_1 FILLER_53_1551 ();
 sg13g2_decap_4 FILLER_53_1565 ();
 sg13g2_fill_1 FILLER_53_1569 ();
 sg13g2_fill_1 FILLER_53_1587 ();
 sg13g2_decap_8 FILLER_53_1606 ();
 sg13g2_decap_8 FILLER_53_1613 ();
 sg13g2_decap_8 FILLER_53_1638 ();
 sg13g2_fill_1 FILLER_53_1645 ();
 sg13g2_decap_4 FILLER_53_1672 ();
 sg13g2_fill_2 FILLER_53_1694 ();
 sg13g2_fill_2 FILLER_53_1709 ();
 sg13g2_fill_1 FILLER_53_1716 ();
 sg13g2_decap_4 FILLER_53_1727 ();
 sg13g2_fill_2 FILLER_53_1740 ();
 sg13g2_fill_1 FILLER_53_1742 ();
 sg13g2_decap_8 FILLER_53_1756 ();
 sg13g2_decap_4 FILLER_53_1763 ();
 sg13g2_fill_1 FILLER_53_1767 ();
 sg13g2_decap_8 FILLER_53_1807 ();
 sg13g2_decap_8 FILLER_53_1877 ();
 sg13g2_decap_8 FILLER_53_1884 ();
 sg13g2_fill_2 FILLER_53_1891 ();
 sg13g2_decap_8 FILLER_53_1911 ();
 sg13g2_fill_2 FILLER_53_1923 ();
 sg13g2_fill_1 FILLER_53_1925 ();
 sg13g2_fill_2 FILLER_53_1930 ();
 sg13g2_fill_1 FILLER_53_1932 ();
 sg13g2_decap_8 FILLER_53_1942 ();
 sg13g2_decap_8 FILLER_53_1962 ();
 sg13g2_decap_8 FILLER_53_1969 ();
 sg13g2_decap_8 FILLER_53_1989 ();
 sg13g2_decap_8 FILLER_53_1996 ();
 sg13g2_fill_2 FILLER_53_2003 ();
 sg13g2_fill_1 FILLER_53_2041 ();
 sg13g2_fill_2 FILLER_53_2057 ();
 sg13g2_fill_1 FILLER_53_2059 ();
 sg13g2_decap_8 FILLER_53_2079 ();
 sg13g2_fill_1 FILLER_53_2086 ();
 sg13g2_decap_4 FILLER_53_2095 ();
 sg13g2_fill_2 FILLER_53_2121 ();
 sg13g2_decap_8 FILLER_53_2158 ();
 sg13g2_decap_4 FILLER_53_2165 ();
 sg13g2_decap_4 FILLER_53_2173 ();
 sg13g2_fill_2 FILLER_53_2177 ();
 sg13g2_fill_2 FILLER_53_2184 ();
 sg13g2_fill_1 FILLER_53_2186 ();
 sg13g2_fill_2 FILLER_53_2195 ();
 sg13g2_decap_8 FILLER_53_2215 ();
 sg13g2_decap_4 FILLER_53_2222 ();
 sg13g2_fill_2 FILLER_53_2226 ();
 sg13g2_fill_2 FILLER_53_2238 ();
 sg13g2_fill_1 FILLER_53_2240 ();
 sg13g2_decap_8 FILLER_53_2251 ();
 sg13g2_decap_8 FILLER_53_2266 ();
 sg13g2_decap_8 FILLER_53_2273 ();
 sg13g2_fill_1 FILLER_53_2316 ();
 sg13g2_decap_4 FILLER_53_2322 ();
 sg13g2_fill_2 FILLER_53_2350 ();
 sg13g2_fill_1 FILLER_53_2352 ();
 sg13g2_fill_2 FILLER_53_2398 ();
 sg13g2_fill_1 FILLER_53_2400 ();
 sg13g2_decap_8 FILLER_53_2422 ();
 sg13g2_decap_8 FILLER_53_2469 ();
 sg13g2_fill_2 FILLER_53_2476 ();
 sg13g2_decap_4 FILLER_53_2490 ();
 sg13g2_fill_1 FILLER_53_2494 ();
 sg13g2_decap_8 FILLER_53_2498 ();
 sg13g2_fill_2 FILLER_53_2505 ();
 sg13g2_fill_1 FILLER_53_2507 ();
 sg13g2_decap_4 FILLER_53_2514 ();
 sg13g2_fill_2 FILLER_53_2518 ();
 sg13g2_decap_8 FILLER_53_2534 ();
 sg13g2_decap_4 FILLER_53_2541 ();
 sg13g2_fill_1 FILLER_53_2545 ();
 sg13g2_fill_1 FILLER_53_2559 ();
 sg13g2_decap_8 FILLER_53_2580 ();
 sg13g2_decap_4 FILLER_53_2587 ();
 sg13g2_decap_4 FILLER_53_2609 ();
 sg13g2_fill_1 FILLER_53_2617 ();
 sg13g2_decap_8 FILLER_53_2628 ();
 sg13g2_fill_2 FILLER_53_2635 ();
 sg13g2_fill_1 FILLER_53_2637 ();
 sg13g2_fill_2 FILLER_53_2656 ();
 sg13g2_fill_1 FILLER_53_2675 ();
 sg13g2_fill_2 FILLER_53_2730 ();
 sg13g2_decap_8 FILLER_53_2743 ();
 sg13g2_fill_2 FILLER_53_2750 ();
 sg13g2_fill_2 FILLER_53_2772 ();
 sg13g2_fill_1 FILLER_53_2778 ();
 sg13g2_fill_2 FILLER_53_2785 ();
 sg13g2_decap_8 FILLER_53_2799 ();
 sg13g2_fill_2 FILLER_53_2806 ();
 sg13g2_fill_1 FILLER_53_2808 ();
 sg13g2_decap_4 FILLER_53_2815 ();
 sg13g2_fill_2 FILLER_53_2837 ();
 sg13g2_fill_1 FILLER_53_2839 ();
 sg13g2_fill_2 FILLER_53_2857 ();
 sg13g2_fill_1 FILLER_53_2859 ();
 sg13g2_decap_4 FILLER_53_2887 ();
 sg13g2_decap_8 FILLER_53_2920 ();
 sg13g2_decap_4 FILLER_53_2927 ();
 sg13g2_fill_1 FILLER_53_2931 ();
 sg13g2_fill_1 FILLER_53_2945 ();
 sg13g2_fill_2 FILLER_53_2950 ();
 sg13g2_decap_4 FILLER_53_2957 ();
 sg13g2_fill_1 FILLER_53_2976 ();
 sg13g2_fill_1 FILLER_53_2992 ();
 sg13g2_fill_2 FILLER_53_3002 ();
 sg13g2_decap_4 FILLER_53_3013 ();
 sg13g2_fill_2 FILLER_53_3054 ();
 sg13g2_fill_1 FILLER_53_3056 ();
 sg13g2_decap_8 FILLER_53_3061 ();
 sg13g2_fill_2 FILLER_53_3068 ();
 sg13g2_fill_2 FILLER_53_3079 ();
 sg13g2_decap_8 FILLER_53_3109 ();
 sg13g2_fill_2 FILLER_53_3116 ();
 sg13g2_fill_2 FILLER_53_3131 ();
 sg13g2_fill_1 FILLER_53_3133 ();
 sg13g2_fill_2 FILLER_53_3170 ();
 sg13g2_fill_2 FILLER_53_3207 ();
 sg13g2_fill_1 FILLER_53_3214 ();
 sg13g2_fill_2 FILLER_53_3232 ();
 sg13g2_fill_2 FILLER_53_3311 ();
 sg13g2_fill_1 FILLER_53_3313 ();
 sg13g2_fill_2 FILLER_53_3361 ();
 sg13g2_fill_1 FILLER_53_3363 ();
 sg13g2_fill_2 FILLER_53_3369 ();
 sg13g2_fill_1 FILLER_53_3395 ();
 sg13g2_decap_4 FILLER_53_3413 ();
 sg13g2_fill_2 FILLER_53_3417 ();
 sg13g2_fill_2 FILLER_53_3427 ();
 sg13g2_fill_1 FILLER_53_3433 ();
 sg13g2_fill_1 FILLER_53_3461 ();
 sg13g2_fill_2 FILLER_53_3489 ();
 sg13g2_decap_8 FILLER_53_3497 ();
 sg13g2_decap_8 FILLER_53_3504 ();
 sg13g2_decap_8 FILLER_53_3511 ();
 sg13g2_decap_8 FILLER_53_3518 ();
 sg13g2_decap_8 FILLER_53_3525 ();
 sg13g2_decap_8 FILLER_53_3532 ();
 sg13g2_decap_8 FILLER_53_3539 ();
 sg13g2_decap_8 FILLER_53_3546 ();
 sg13g2_decap_8 FILLER_53_3553 ();
 sg13g2_decap_8 FILLER_53_3560 ();
 sg13g2_decap_8 FILLER_53_3567 ();
 sg13g2_decap_4 FILLER_53_3574 ();
 sg13g2_fill_2 FILLER_53_3578 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_85 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_decap_8 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_109 ();
 sg13g2_fill_2 FILLER_54_140 ();
 sg13g2_decap_4 FILLER_54_155 ();
 sg13g2_decap_4 FILLER_54_172 ();
 sg13g2_decap_8 FILLER_54_186 ();
 sg13g2_fill_1 FILLER_54_193 ();
 sg13g2_fill_1 FILLER_54_228 ();
 sg13g2_decap_8 FILLER_54_238 ();
 sg13g2_fill_2 FILLER_54_245 ();
 sg13g2_fill_1 FILLER_54_247 ();
 sg13g2_fill_2 FILLER_54_252 ();
 sg13g2_fill_2 FILLER_54_262 ();
 sg13g2_fill_2 FILLER_54_272 ();
 sg13g2_decap_4 FILLER_54_286 ();
 sg13g2_fill_2 FILLER_54_295 ();
 sg13g2_fill_1 FILLER_54_297 ();
 sg13g2_decap_4 FILLER_54_319 ();
 sg13g2_fill_2 FILLER_54_367 ();
 sg13g2_fill_2 FILLER_54_378 ();
 sg13g2_fill_1 FILLER_54_380 ();
 sg13g2_fill_2 FILLER_54_385 ();
 sg13g2_fill_1 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_405 ();
 sg13g2_fill_1 FILLER_54_412 ();
 sg13g2_fill_1 FILLER_54_431 ();
 sg13g2_fill_1 FILLER_54_437 ();
 sg13g2_fill_2 FILLER_54_449 ();
 sg13g2_fill_2 FILLER_54_476 ();
 sg13g2_fill_2 FILLER_54_486 ();
 sg13g2_fill_2 FILLER_54_498 ();
 sg13g2_fill_1 FILLER_54_500 ();
 sg13g2_decap_4 FILLER_54_520 ();
 sg13g2_fill_1 FILLER_54_524 ();
 sg13g2_fill_2 FILLER_54_541 ();
 sg13g2_decap_8 FILLER_54_547 ();
 sg13g2_decap_8 FILLER_54_554 ();
 sg13g2_decap_8 FILLER_54_561 ();
 sg13g2_decap_4 FILLER_54_568 ();
 sg13g2_decap_4 FILLER_54_639 ();
 sg13g2_fill_2 FILLER_54_732 ();
 sg13g2_fill_2 FILLER_54_761 ();
 sg13g2_fill_1 FILLER_54_763 ();
 sg13g2_fill_2 FILLER_54_863 ();
 sg13g2_decap_4 FILLER_54_883 ();
 sg13g2_fill_2 FILLER_54_946 ();
 sg13g2_fill_1 FILLER_54_948 ();
 sg13g2_decap_8 FILLER_54_953 ();
 sg13g2_fill_1 FILLER_54_960 ();
 sg13g2_fill_2 FILLER_54_989 ();
 sg13g2_decap_8 FILLER_54_1009 ();
 sg13g2_fill_2 FILLER_54_1016 ();
 sg13g2_decap_8 FILLER_54_1027 ();
 sg13g2_decap_4 FILLER_54_1038 ();
 sg13g2_fill_2 FILLER_54_1042 ();
 sg13g2_decap_8 FILLER_54_1066 ();
 sg13g2_fill_2 FILLER_54_1073 ();
 sg13g2_fill_1 FILLER_54_1075 ();
 sg13g2_fill_2 FILLER_54_1084 ();
 sg13g2_fill_1 FILLER_54_1096 ();
 sg13g2_fill_1 FILLER_54_1102 ();
 sg13g2_fill_1 FILLER_54_1114 ();
 sg13g2_fill_2 FILLER_54_1122 ();
 sg13g2_fill_1 FILLER_54_1124 ();
 sg13g2_fill_1 FILLER_54_1130 ();
 sg13g2_fill_2 FILLER_54_1139 ();
 sg13g2_fill_1 FILLER_54_1141 ();
 sg13g2_fill_2 FILLER_54_1155 ();
 sg13g2_decap_8 FILLER_54_1161 ();
 sg13g2_fill_1 FILLER_54_1168 ();
 sg13g2_decap_4 FILLER_54_1178 ();
 sg13g2_fill_2 FILLER_54_1186 ();
 sg13g2_decap_4 FILLER_54_1201 ();
 sg13g2_fill_1 FILLER_54_1205 ();
 sg13g2_decap_8 FILLER_54_1222 ();
 sg13g2_decap_8 FILLER_54_1229 ();
 sg13g2_decap_4 FILLER_54_1236 ();
 sg13g2_fill_2 FILLER_54_1240 ();
 sg13g2_fill_2 FILLER_54_1247 ();
 sg13g2_decap_4 FILLER_54_1253 ();
 sg13g2_fill_1 FILLER_54_1257 ();
 sg13g2_fill_2 FILLER_54_1289 ();
 sg13g2_fill_2 FILLER_54_1304 ();
 sg13g2_fill_1 FILLER_54_1306 ();
 sg13g2_decap_4 FILLER_54_1329 ();
 sg13g2_fill_1 FILLER_54_1333 ();
 sg13g2_decap_4 FILLER_54_1380 ();
 sg13g2_fill_1 FILLER_54_1422 ();
 sg13g2_decap_4 FILLER_54_1454 ();
 sg13g2_fill_2 FILLER_54_1588 ();
 sg13g2_fill_2 FILLER_54_1617 ();
 sg13g2_fill_1 FILLER_54_1619 ();
 sg13g2_fill_2 FILLER_54_1669 ();
 sg13g2_fill_1 FILLER_54_1708 ();
 sg13g2_fill_2 FILLER_54_1717 ();
 sg13g2_fill_1 FILLER_54_1719 ();
 sg13g2_fill_1 FILLER_54_1737 ();
 sg13g2_fill_2 FILLER_54_1771 ();
 sg13g2_fill_2 FILLER_54_1782 ();
 sg13g2_fill_1 FILLER_54_1784 ();
 sg13g2_fill_1 FILLER_54_1811 ();
 sg13g2_decap_8 FILLER_54_1816 ();
 sg13g2_fill_2 FILLER_54_1823 ();
 sg13g2_fill_1 FILLER_54_1825 ();
 sg13g2_fill_1 FILLER_54_1840 ();
 sg13g2_decap_4 FILLER_54_1869 ();
 sg13g2_fill_2 FILLER_54_1873 ();
 sg13g2_fill_2 FILLER_54_1938 ();
 sg13g2_fill_1 FILLER_54_1940 ();
 sg13g2_decap_8 FILLER_54_2009 ();
 sg13g2_fill_2 FILLER_54_2016 ();
 sg13g2_decap_8 FILLER_54_2022 ();
 sg13g2_fill_1 FILLER_54_2029 ();
 sg13g2_fill_2 FILLER_54_2039 ();
 sg13g2_decap_8 FILLER_54_2072 ();
 sg13g2_decap_4 FILLER_54_2079 ();
 sg13g2_fill_2 FILLER_54_2083 ();
 sg13g2_fill_2 FILLER_54_2090 ();
 sg13g2_fill_1 FILLER_54_2141 ();
 sg13g2_fill_2 FILLER_54_2182 ();
 sg13g2_fill_1 FILLER_54_2184 ();
 sg13g2_decap_4 FILLER_54_2198 ();
 sg13g2_fill_2 FILLER_54_2202 ();
 sg13g2_decap_8 FILLER_54_2216 ();
 sg13g2_decap_4 FILLER_54_2223 ();
 sg13g2_fill_2 FILLER_54_2240 ();
 sg13g2_fill_1 FILLER_54_2242 ();
 sg13g2_fill_2 FILLER_54_2253 ();
 sg13g2_fill_1 FILLER_54_2255 ();
 sg13g2_decap_8 FILLER_54_2280 ();
 sg13g2_fill_1 FILLER_54_2287 ();
 sg13g2_decap_8 FILLER_54_2306 ();
 sg13g2_fill_2 FILLER_54_2382 ();
 sg13g2_decap_4 FILLER_54_2431 ();
 sg13g2_fill_1 FILLER_54_2435 ();
 sg13g2_decap_4 FILLER_54_2449 ();
 sg13g2_fill_1 FILLER_54_2453 ();
 sg13g2_fill_2 FILLER_54_2458 ();
 sg13g2_fill_1 FILLER_54_2460 ();
 sg13g2_decap_4 FILLER_54_2466 ();
 sg13g2_fill_2 FILLER_54_2470 ();
 sg13g2_fill_1 FILLER_54_2499 ();
 sg13g2_fill_1 FILLER_54_2516 ();
 sg13g2_decap_4 FILLER_54_2568 ();
 sg13g2_fill_2 FILLER_54_2595 ();
 sg13g2_fill_1 FILLER_54_2597 ();
 sg13g2_fill_2 FILLER_54_2614 ();
 sg13g2_decap_8 FILLER_54_2628 ();
 sg13g2_fill_2 FILLER_54_2635 ();
 sg13g2_fill_2 FILLER_54_2650 ();
 sg13g2_fill_1 FILLER_54_2652 ();
 sg13g2_decap_4 FILLER_54_2661 ();
 sg13g2_fill_1 FILLER_54_2665 ();
 sg13g2_decap_8 FILLER_54_2682 ();
 sg13g2_fill_1 FILLER_54_2689 ();
 sg13g2_fill_1 FILLER_54_2694 ();
 sg13g2_decap_8 FILLER_54_2704 ();
 sg13g2_fill_2 FILLER_54_2711 ();
 sg13g2_fill_1 FILLER_54_2713 ();
 sg13g2_fill_1 FILLER_54_2727 ();
 sg13g2_fill_1 FILLER_54_2751 ();
 sg13g2_fill_1 FILLER_54_2760 ();
 sg13g2_fill_1 FILLER_54_2771 ();
 sg13g2_decap_4 FILLER_54_2797 ();
 sg13g2_fill_2 FILLER_54_2801 ();
 sg13g2_fill_2 FILLER_54_2819 ();
 sg13g2_fill_1 FILLER_54_2821 ();
 sg13g2_fill_1 FILLER_54_2833 ();
 sg13g2_fill_2 FILLER_54_2842 ();
 sg13g2_fill_1 FILLER_54_2844 ();
 sg13g2_fill_1 FILLER_54_2853 ();
 sg13g2_decap_8 FILLER_54_2870 ();
 sg13g2_decap_4 FILLER_54_2877 ();
 sg13g2_decap_4 FILLER_54_2896 ();
 sg13g2_fill_1 FILLER_54_2906 ();
 sg13g2_decap_4 FILLER_54_2947 ();
 sg13g2_fill_2 FILLER_54_2970 ();
 sg13g2_fill_2 FILLER_54_2978 ();
 sg13g2_fill_2 FILLER_54_3009 ();
 sg13g2_fill_1 FILLER_54_3011 ();
 sg13g2_fill_1 FILLER_54_3019 ();
 sg13g2_fill_1 FILLER_54_3040 ();
 sg13g2_fill_1 FILLER_54_3045 ();
 sg13g2_decap_8 FILLER_54_3051 ();
 sg13g2_decap_4 FILLER_54_3058 ();
 sg13g2_fill_1 FILLER_54_3062 ();
 sg13g2_decap_4 FILLER_54_3068 ();
 sg13g2_fill_1 FILLER_54_3072 ();
 sg13g2_decap_8 FILLER_54_3086 ();
 sg13g2_fill_2 FILLER_54_3093 ();
 sg13g2_fill_1 FILLER_54_3095 ();
 sg13g2_fill_2 FILLER_54_3114 ();
 sg13g2_decap_8 FILLER_54_3133 ();
 sg13g2_fill_1 FILLER_54_3140 ();
 sg13g2_fill_2 FILLER_54_3158 ();
 sg13g2_decap_8 FILLER_54_3173 ();
 sg13g2_decap_4 FILLER_54_3180 ();
 sg13g2_fill_2 FILLER_54_3184 ();
 sg13g2_fill_2 FILLER_54_3195 ();
 sg13g2_fill_1 FILLER_54_3197 ();
 sg13g2_fill_1 FILLER_54_3239 ();
 sg13g2_fill_2 FILLER_54_3271 ();
 sg13g2_fill_1 FILLER_54_3273 ();
 sg13g2_fill_2 FILLER_54_3287 ();
 sg13g2_fill_1 FILLER_54_3289 ();
 sg13g2_fill_2 FILLER_54_3303 ();
 sg13g2_fill_2 FILLER_54_3390 ();
 sg13g2_decap_8 FILLER_54_3419 ();
 sg13g2_fill_1 FILLER_54_3426 ();
 sg13g2_fill_2 FILLER_54_3440 ();
 sg13g2_fill_1 FILLER_54_3442 ();
 sg13g2_fill_2 FILLER_54_3458 ();
 sg13g2_fill_1 FILLER_54_3460 ();
 sg13g2_decap_4 FILLER_54_3471 ();
 sg13g2_fill_1 FILLER_54_3483 ();
 sg13g2_decap_8 FILLER_54_3499 ();
 sg13g2_fill_2 FILLER_54_3506 ();
 sg13g2_fill_1 FILLER_54_3508 ();
 sg13g2_decap_8 FILLER_54_3513 ();
 sg13g2_decap_8 FILLER_54_3520 ();
 sg13g2_decap_8 FILLER_54_3527 ();
 sg13g2_decap_8 FILLER_54_3534 ();
 sg13g2_decap_8 FILLER_54_3541 ();
 sg13g2_decap_8 FILLER_54_3548 ();
 sg13g2_decap_8 FILLER_54_3555 ();
 sg13g2_decap_8 FILLER_54_3562 ();
 sg13g2_decap_8 FILLER_54_3569 ();
 sg13g2_decap_4 FILLER_54_3576 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_13 ();
 sg13g2_fill_2 FILLER_55_20 ();
 sg13g2_fill_1 FILLER_55_22 ();
 sg13g2_decap_4 FILLER_55_32 ();
 sg13g2_decap_4 FILLER_55_45 ();
 sg13g2_decap_4 FILLER_55_52 ();
 sg13g2_fill_2 FILLER_55_70 ();
 sg13g2_fill_1 FILLER_55_72 ();
 sg13g2_fill_2 FILLER_55_77 ();
 sg13g2_fill_2 FILLER_55_93 ();
 sg13g2_decap_4 FILLER_55_109 ();
 sg13g2_fill_2 FILLER_55_113 ();
 sg13g2_decap_8 FILLER_55_160 ();
 sg13g2_fill_2 FILLER_55_167 ();
 sg13g2_fill_2 FILLER_55_194 ();
 sg13g2_decap_8 FILLER_55_209 ();
 sg13g2_decap_8 FILLER_55_216 ();
 sg13g2_fill_1 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_264 ();
 sg13g2_fill_2 FILLER_55_288 ();
 sg13g2_fill_1 FILLER_55_290 ();
 sg13g2_fill_2 FILLER_55_295 ();
 sg13g2_fill_1 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_338 ();
 sg13g2_fill_1 FILLER_55_382 ();
 sg13g2_fill_2 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_423 ();
 sg13g2_decap_4 FILLER_55_445 ();
 sg13g2_fill_1 FILLER_55_449 ();
 sg13g2_fill_2 FILLER_55_454 ();
 sg13g2_fill_1 FILLER_55_456 ();
 sg13g2_fill_2 FILLER_55_465 ();
 sg13g2_fill_1 FILLER_55_467 ();
 sg13g2_fill_1 FILLER_55_478 ();
 sg13g2_decap_4 FILLER_55_489 ();
 sg13g2_fill_1 FILLER_55_493 ();
 sg13g2_fill_2 FILLER_55_499 ();
 sg13g2_decap_4 FILLER_55_509 ();
 sg13g2_fill_1 FILLER_55_513 ();
 sg13g2_decap_4 FILLER_55_558 ();
 sg13g2_fill_1 FILLER_55_562 ();
 sg13g2_decap_4 FILLER_55_595 ();
 sg13g2_fill_1 FILLER_55_622 ();
 sg13g2_decap_8 FILLER_55_641 ();
 sg13g2_fill_1 FILLER_55_648 ();
 sg13g2_decap_4 FILLER_55_663 ();
 sg13g2_fill_2 FILLER_55_667 ();
 sg13g2_decap_8 FILLER_55_679 ();
 sg13g2_decap_8 FILLER_55_686 ();
 sg13g2_decap_8 FILLER_55_693 ();
 sg13g2_fill_2 FILLER_55_700 ();
 sg13g2_fill_2 FILLER_55_716 ();
 sg13g2_decap_8 FILLER_55_736 ();
 sg13g2_decap_8 FILLER_55_743 ();
 sg13g2_fill_1 FILLER_55_750 ();
 sg13g2_decap_8 FILLER_55_787 ();
 sg13g2_fill_2 FILLER_55_794 ();
 sg13g2_fill_1 FILLER_55_796 ();
 sg13g2_fill_2 FILLER_55_815 ();
 sg13g2_fill_2 FILLER_55_844 ();
 sg13g2_fill_1 FILLER_55_846 ();
 sg13g2_fill_1 FILLER_55_856 ();
 sg13g2_decap_8 FILLER_55_883 ();
 sg13g2_fill_1 FILLER_55_930 ();
 sg13g2_decap_4 FILLER_55_958 ();
 sg13g2_fill_2 FILLER_55_962 ();
 sg13g2_decap_8 FILLER_55_977 ();
 sg13g2_decap_8 FILLER_55_984 ();
 sg13g2_decap_4 FILLER_55_991 ();
 sg13g2_decap_4 FILLER_55_1023 ();
 sg13g2_fill_2 FILLER_55_1027 ();
 sg13g2_decap_8 FILLER_55_1033 ();
 sg13g2_fill_2 FILLER_55_1040 ();
 sg13g2_fill_2 FILLER_55_1045 ();
 sg13g2_fill_1 FILLER_55_1092 ();
 sg13g2_fill_2 FILLER_55_1112 ();
 sg13g2_decap_8 FILLER_55_1123 ();
 sg13g2_decap_4 FILLER_55_1130 ();
 sg13g2_fill_1 FILLER_55_1134 ();
 sg13g2_fill_1 FILLER_55_1140 ();
 sg13g2_fill_2 FILLER_55_1195 ();
 sg13g2_fill_2 FILLER_55_1264 ();
 sg13g2_fill_1 FILLER_55_1266 ();
 sg13g2_fill_2 FILLER_55_1308 ();
 sg13g2_decap_8 FILLER_55_1350 ();
 sg13g2_decap_4 FILLER_55_1357 ();
 sg13g2_fill_2 FILLER_55_1361 ();
 sg13g2_fill_1 FILLER_55_1390 ();
 sg13g2_fill_2 FILLER_55_1418 ();
 sg13g2_fill_1 FILLER_55_1420 ();
 sg13g2_fill_2 FILLER_55_1498 ();
 sg13g2_fill_2 FILLER_55_1513 ();
 sg13g2_fill_2 FILLER_55_1524 ();
 sg13g2_fill_1 FILLER_55_1526 ();
 sg13g2_fill_1 FILLER_55_1531 ();
 sg13g2_fill_2 FILLER_55_1537 ();
 sg13g2_fill_2 FILLER_55_1589 ();
 sg13g2_fill_2 FILLER_55_1608 ();
 sg13g2_fill_2 FILLER_55_1623 ();
 sg13g2_fill_2 FILLER_55_1643 ();
 sg13g2_decap_4 FILLER_55_1672 ();
 sg13g2_decap_8 FILLER_55_1680 ();
 sg13g2_decap_4 FILLER_55_1687 ();
 sg13g2_fill_2 FILLER_55_1713 ();
 sg13g2_fill_2 FILLER_55_1724 ();
 sg13g2_decap_8 FILLER_55_1746 ();
 sg13g2_fill_1 FILLER_55_1757 ();
 sg13g2_fill_1 FILLER_55_1772 ();
 sg13g2_fill_1 FILLER_55_1805 ();
 sg13g2_fill_2 FILLER_55_1865 ();
 sg13g2_fill_1 FILLER_55_1867 ();
 sg13g2_decap_4 FILLER_55_1926 ();
 sg13g2_fill_1 FILLER_55_1930 ();
 sg13g2_decap_4 FILLER_55_1957 ();
 sg13g2_fill_1 FILLER_55_1961 ();
 sg13g2_decap_8 FILLER_55_1971 ();
 sg13g2_fill_1 FILLER_55_1978 ();
 sg13g2_decap_4 FILLER_55_1992 ();
 sg13g2_decap_4 FILLER_55_2030 ();
 sg13g2_fill_1 FILLER_55_2034 ();
 sg13g2_fill_1 FILLER_55_2057 ();
 sg13g2_decap_8 FILLER_55_2094 ();
 sg13g2_fill_2 FILLER_55_2101 ();
 sg13g2_fill_2 FILLER_55_2121 ();
 sg13g2_decap_8 FILLER_55_2176 ();
 sg13g2_decap_8 FILLER_55_2183 ();
 sg13g2_fill_1 FILLER_55_2190 ();
 sg13g2_fill_2 FILLER_55_2256 ();
 sg13g2_fill_1 FILLER_55_2258 ();
 sg13g2_fill_2 FILLER_55_2275 ();
 sg13g2_fill_1 FILLER_55_2277 ();
 sg13g2_fill_1 FILLER_55_2296 ();
 sg13g2_fill_1 FILLER_55_2305 ();
 sg13g2_fill_2 FILLER_55_2314 ();
 sg13g2_fill_1 FILLER_55_2325 ();
 sg13g2_fill_1 FILLER_55_2330 ();
 sg13g2_decap_4 FILLER_55_2344 ();
 sg13g2_fill_1 FILLER_55_2348 ();
 sg13g2_fill_2 FILLER_55_2396 ();
 sg13g2_fill_1 FILLER_55_2398 ();
 sg13g2_fill_2 FILLER_55_2413 ();
 sg13g2_fill_1 FILLER_55_2415 ();
 sg13g2_fill_1 FILLER_55_2438 ();
 sg13g2_fill_2 FILLER_55_2467 ();
 sg13g2_fill_1 FILLER_55_2469 ();
 sg13g2_fill_2 FILLER_55_2479 ();
 sg13g2_fill_1 FILLER_55_2481 ();
 sg13g2_fill_2 FILLER_55_2497 ();
 sg13g2_fill_2 FILLER_55_2512 ();
 sg13g2_fill_1 FILLER_55_2514 ();
 sg13g2_fill_2 FILLER_55_2524 ();
 sg13g2_fill_1 FILLER_55_2526 ();
 sg13g2_decap_8 FILLER_55_2531 ();
 sg13g2_decap_8 FILLER_55_2538 ();
 sg13g2_fill_2 FILLER_55_2545 ();
 sg13g2_fill_1 FILLER_55_2547 ();
 sg13g2_decap_4 FILLER_55_2561 ();
 sg13g2_fill_1 FILLER_55_2580 ();
 sg13g2_decap_4 FILLER_55_2656 ();
 sg13g2_decap_8 FILLER_55_2693 ();
 sg13g2_fill_1 FILLER_55_2700 ();
 sg13g2_fill_2 FILLER_55_2727 ();
 sg13g2_fill_1 FILLER_55_2729 ();
 sg13g2_decap_8 FILLER_55_2743 ();
 sg13g2_fill_1 FILLER_55_2754 ();
 sg13g2_fill_1 FILLER_55_2764 ();
 sg13g2_fill_2 FILLER_55_2770 ();
 sg13g2_fill_1 FILLER_55_2772 ();
 sg13g2_fill_2 FILLER_55_2796 ();
 sg13g2_decap_4 FILLER_55_2815 ();
 sg13g2_fill_1 FILLER_55_2849 ();
 sg13g2_fill_2 FILLER_55_2858 ();
 sg13g2_decap_8 FILLER_55_2877 ();
 sg13g2_fill_1 FILLER_55_2884 ();
 sg13g2_decap_8 FILLER_55_2898 ();
 sg13g2_fill_1 FILLER_55_2905 ();
 sg13g2_fill_2 FILLER_55_2911 ();
 sg13g2_fill_1 FILLER_55_2913 ();
 sg13g2_decap_8 FILLER_55_2918 ();
 sg13g2_decap_8 FILLER_55_2925 ();
 sg13g2_fill_1 FILLER_55_2932 ();
 sg13g2_decap_4 FILLER_55_2942 ();
 sg13g2_fill_2 FILLER_55_2964 ();
 sg13g2_fill_1 FILLER_55_2966 ();
 sg13g2_decap_8 FILLER_55_2976 ();
 sg13g2_fill_2 FILLER_55_2983 ();
 sg13g2_fill_1 FILLER_55_2996 ();
 sg13g2_decap_8 FILLER_55_3025 ();
 sg13g2_decap_4 FILLER_55_3032 ();
 sg13g2_decap_4 FILLER_55_3070 ();
 sg13g2_fill_1 FILLER_55_3074 ();
 sg13g2_fill_1 FILLER_55_3088 ();
 sg13g2_fill_2 FILLER_55_3102 ();
 sg13g2_fill_1 FILLER_55_3145 ();
 sg13g2_fill_1 FILLER_55_3151 ();
 sg13g2_fill_1 FILLER_55_3162 ();
 sg13g2_fill_1 FILLER_55_3208 ();
 sg13g2_fill_1 FILLER_55_3219 ();
 sg13g2_fill_1 FILLER_55_3233 ();
 sg13g2_fill_2 FILLER_55_3258 ();
 sg13g2_fill_1 FILLER_55_3260 ();
 sg13g2_decap_8 FILLER_55_3275 ();
 sg13g2_fill_2 FILLER_55_3295 ();
 sg13g2_fill_2 FILLER_55_3357 ();
 sg13g2_fill_1 FILLER_55_3359 ();
 sg13g2_fill_2 FILLER_55_3364 ();
 sg13g2_fill_1 FILLER_55_3366 ();
 sg13g2_fill_2 FILLER_55_3373 ();
 sg13g2_fill_2 FILLER_55_3384 ();
 sg13g2_decap_8 FILLER_55_3397 ();
 sg13g2_fill_2 FILLER_55_3404 ();
 sg13g2_decap_8 FILLER_55_3417 ();
 sg13g2_decap_8 FILLER_55_3424 ();
 sg13g2_decap_4 FILLER_55_3450 ();
 sg13g2_fill_2 FILLER_55_3454 ();
 sg13g2_fill_1 FILLER_55_3461 ();
 sg13g2_fill_1 FILLER_55_3503 ();
 sg13g2_decap_8 FILLER_55_3532 ();
 sg13g2_decap_8 FILLER_55_3539 ();
 sg13g2_decap_8 FILLER_55_3546 ();
 sg13g2_decap_8 FILLER_55_3553 ();
 sg13g2_decap_8 FILLER_55_3560 ();
 sg13g2_decap_8 FILLER_55_3567 ();
 sg13g2_decap_4 FILLER_55_3574 ();
 sg13g2_fill_2 FILLER_55_3578 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_34 ();
 sg13g2_fill_1 FILLER_56_38 ();
 sg13g2_fill_1 FILLER_56_43 ();
 sg13g2_fill_2 FILLER_56_49 ();
 sg13g2_fill_1 FILLER_56_56 ();
 sg13g2_fill_2 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_67 ();
 sg13g2_fill_1 FILLER_56_78 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_4 FILLER_56_91 ();
 sg13g2_fill_1 FILLER_56_95 ();
 sg13g2_decap_4 FILLER_56_101 ();
 sg13g2_fill_2 FILLER_56_105 ();
 sg13g2_fill_2 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_159 ();
 sg13g2_decap_8 FILLER_56_173 ();
 sg13g2_fill_1 FILLER_56_180 ();
 sg13g2_decap_8 FILLER_56_208 ();
 sg13g2_decap_8 FILLER_56_215 ();
 sg13g2_decap_4 FILLER_56_222 ();
 sg13g2_fill_1 FILLER_56_226 ();
 sg13g2_fill_2 FILLER_56_240 ();
 sg13g2_fill_1 FILLER_56_242 ();
 sg13g2_fill_2 FILLER_56_248 ();
 sg13g2_fill_1 FILLER_56_250 ();
 sg13g2_fill_2 FILLER_56_283 ();
 sg13g2_fill_1 FILLER_56_285 ();
 sg13g2_fill_1 FILLER_56_323 ();
 sg13g2_decap_8 FILLER_56_352 ();
 sg13g2_fill_2 FILLER_56_359 ();
 sg13g2_fill_2 FILLER_56_379 ();
 sg13g2_fill_1 FILLER_56_409 ();
 sg13g2_fill_1 FILLER_56_418 ();
 sg13g2_fill_1 FILLER_56_425 ();
 sg13g2_fill_2 FILLER_56_430 ();
 sg13g2_fill_2 FILLER_56_442 ();
 sg13g2_fill_1 FILLER_56_444 ();
 sg13g2_fill_1 FILLER_56_466 ();
 sg13g2_fill_2 FILLER_56_492 ();
 sg13g2_fill_1 FILLER_56_494 ();
 sg13g2_fill_1 FILLER_56_518 ();
 sg13g2_fill_1 FILLER_56_534 ();
 sg13g2_decap_4 FILLER_56_548 ();
 sg13g2_fill_1 FILLER_56_552 ();
 sg13g2_fill_2 FILLER_56_590 ();
 sg13g2_fill_1 FILLER_56_592 ();
 sg13g2_fill_2 FILLER_56_607 ();
 sg13g2_fill_2 FILLER_56_677 ();
 sg13g2_fill_1 FILLER_56_679 ();
 sg13g2_fill_2 FILLER_56_693 ();
 sg13g2_fill_2 FILLER_56_735 ();
 sg13g2_fill_1 FILLER_56_737 ();
 sg13g2_decap_4 FILLER_56_757 ();
 sg13g2_fill_1 FILLER_56_761 ();
 sg13g2_decap_4 FILLER_56_775 ();
 sg13g2_decap_4 FILLER_56_791 ();
 sg13g2_fill_2 FILLER_56_831 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_fill_2 FILLER_56_906 ();
 sg13g2_fill_2 FILLER_56_917 ();
 sg13g2_fill_2 FILLER_56_941 ();
 sg13g2_fill_1 FILLER_56_943 ();
 sg13g2_decap_8 FILLER_56_985 ();
 sg13g2_fill_1 FILLER_56_992 ();
 sg13g2_decap_8 FILLER_56_1012 ();
 sg13g2_fill_1 FILLER_56_1019 ();
 sg13g2_fill_2 FILLER_56_1033 ();
 sg13g2_fill_1 FILLER_56_1035 ();
 sg13g2_fill_1 FILLER_56_1059 ();
 sg13g2_decap_4 FILLER_56_1092 ();
 sg13g2_fill_1 FILLER_56_1096 ();
 sg13g2_fill_2 FILLER_56_1100 ();
 sg13g2_fill_1 FILLER_56_1102 ();
 sg13g2_decap_8 FILLER_56_1131 ();
 sg13g2_fill_2 FILLER_56_1138 ();
 sg13g2_decap_8 FILLER_56_1158 ();
 sg13g2_fill_1 FILLER_56_1165 ();
 sg13g2_decap_8 FILLER_56_1224 ();
 sg13g2_decap_4 FILLER_56_1231 ();
 sg13g2_fill_1 FILLER_56_1249 ();
 sg13g2_fill_1 FILLER_56_1327 ();
 sg13g2_fill_1 FILLER_56_1347 ();
 sg13g2_fill_2 FILLER_56_1358 ();
 sg13g2_fill_2 FILLER_56_1370 ();
 sg13g2_fill_1 FILLER_56_1372 ();
 sg13g2_decap_4 FILLER_56_1377 ();
 sg13g2_fill_1 FILLER_56_1403 ();
 sg13g2_fill_1 FILLER_56_1450 ();
 sg13g2_fill_1 FILLER_56_1478 ();
 sg13g2_decap_4 FILLER_56_1530 ();
 sg13g2_fill_2 FILLER_56_1616 ();
 sg13g2_fill_2 FILLER_56_1680 ();
 sg13g2_fill_1 FILLER_56_1696 ();
 sg13g2_fill_1 FILLER_56_1729 ();
 sg13g2_fill_2 FILLER_56_1785 ();
 sg13g2_decap_8 FILLER_56_1805 ();
 sg13g2_fill_1 FILLER_56_1812 ();
 sg13g2_decap_8 FILLER_56_1818 ();
 sg13g2_fill_2 FILLER_56_1825 ();
 sg13g2_fill_1 FILLER_56_1827 ();
 sg13g2_fill_1 FILLER_56_1858 ();
 sg13g2_decap_4 FILLER_56_1868 ();
 sg13g2_decap_4 FILLER_56_1894 ();
 sg13g2_fill_2 FILLER_56_1907 ();
 sg13g2_fill_2 FILLER_56_1914 ();
 sg13g2_decap_8 FILLER_56_1929 ();
 sg13g2_decap_8 FILLER_56_1963 ();
 sg13g2_decap_4 FILLER_56_2010 ();
 sg13g2_fill_2 FILLER_56_2014 ();
 sg13g2_fill_1 FILLER_56_2025 ();
 sg13g2_decap_4 FILLER_56_2044 ();
 sg13g2_fill_1 FILLER_56_2052 ();
 sg13g2_fill_2 FILLER_56_2094 ();
 sg13g2_fill_1 FILLER_56_2141 ();
 sg13g2_decap_8 FILLER_56_2196 ();
 sg13g2_decap_4 FILLER_56_2203 ();
 sg13g2_fill_2 FILLER_56_2207 ();
 sg13g2_fill_1 FILLER_56_2213 ();
 sg13g2_fill_2 FILLER_56_2257 ();
 sg13g2_fill_2 FILLER_56_2272 ();
 sg13g2_fill_1 FILLER_56_2274 ();
 sg13g2_fill_2 FILLER_56_2299 ();
 sg13g2_decap_4 FILLER_56_2329 ();
 sg13g2_fill_1 FILLER_56_2333 ();
 sg13g2_fill_1 FILLER_56_2347 ();
 sg13g2_decap_8 FILLER_56_2357 ();
 sg13g2_fill_2 FILLER_56_2364 ();
 sg13g2_fill_2 FILLER_56_2371 ();
 sg13g2_fill_1 FILLER_56_2373 ();
 sg13g2_fill_2 FILLER_56_2412 ();
 sg13g2_fill_1 FILLER_56_2414 ();
 sg13g2_fill_1 FILLER_56_2481 ();
 sg13g2_fill_2 FILLER_56_2510 ();
 sg13g2_fill_1 FILLER_56_2512 ();
 sg13g2_fill_2 FILLER_56_2526 ();
 sg13g2_fill_2 FILLER_56_2559 ();
 sg13g2_fill_2 FILLER_56_2566 ();
 sg13g2_decap_4 FILLER_56_2596 ();
 sg13g2_fill_2 FILLER_56_2600 ();
 sg13g2_decap_4 FILLER_56_2629 ();
 sg13g2_fill_1 FILLER_56_2637 ();
 sg13g2_decap_8 FILLER_56_2647 ();
 sg13g2_fill_1 FILLER_56_2654 ();
 sg13g2_decap_8 FILLER_56_2659 ();
 sg13g2_fill_2 FILLER_56_2698 ();
 sg13g2_fill_1 FILLER_56_2700 ();
 sg13g2_fill_2 FILLER_56_2729 ();
 sg13g2_fill_1 FILLER_56_2731 ();
 sg13g2_decap_4 FILLER_56_2736 ();
 sg13g2_fill_1 FILLER_56_2740 ();
 sg13g2_fill_1 FILLER_56_2769 ();
 sg13g2_fill_1 FILLER_56_2814 ();
 sg13g2_fill_2 FILLER_56_2820 ();
 sg13g2_fill_2 FILLER_56_2849 ();
 sg13g2_fill_1 FILLER_56_2851 ();
 sg13g2_fill_2 FILLER_56_2880 ();
 sg13g2_fill_1 FILLER_56_2882 ();
 sg13g2_fill_1 FILLER_56_2941 ();
 sg13g2_fill_1 FILLER_56_2951 ();
 sg13g2_fill_1 FILLER_56_2956 ();
 sg13g2_decap_4 FILLER_56_2995 ();
 sg13g2_fill_1 FILLER_56_2999 ();
 sg13g2_fill_1 FILLER_56_3028 ();
 sg13g2_decap_8 FILLER_56_3034 ();
 sg13g2_fill_2 FILLER_56_3041 ();
 sg13g2_fill_1 FILLER_56_3047 ();
 sg13g2_fill_2 FILLER_56_3062 ();
 sg13g2_fill_2 FILLER_56_3106 ();
 sg13g2_fill_1 FILLER_56_3108 ();
 sg13g2_decap_4 FILLER_56_3122 ();
 sg13g2_fill_1 FILLER_56_3126 ();
 sg13g2_fill_2 FILLER_56_3140 ();
 sg13g2_fill_2 FILLER_56_3160 ();
 sg13g2_fill_1 FILLER_56_3162 ();
 sg13g2_fill_1 FILLER_56_3168 ();
 sg13g2_fill_2 FILLER_56_3212 ();
 sg13g2_fill_1 FILLER_56_3214 ();
 sg13g2_fill_2 FILLER_56_3238 ();
 sg13g2_fill_2 FILLER_56_3294 ();
 sg13g2_decap_4 FILLER_56_3356 ();
 sg13g2_fill_2 FILLER_56_3360 ();
 sg13g2_fill_1 FILLER_56_3375 ();
 sg13g2_fill_2 FILLER_56_3399 ();
 sg13g2_fill_1 FILLER_56_3422 ();
 sg13g2_decap_8 FILLER_56_3445 ();
 sg13g2_decap_8 FILLER_56_3452 ();
 sg13g2_fill_2 FILLER_56_3459 ();
 sg13g2_fill_1 FILLER_56_3461 ();
 sg13g2_fill_1 FILLER_56_3467 ();
 sg13g2_decap_8 FILLER_56_3478 ();
 sg13g2_decap_8 FILLER_56_3485 ();
 sg13g2_fill_1 FILLER_56_3492 ();
 sg13g2_fill_2 FILLER_56_3497 ();
 sg13g2_fill_1 FILLER_56_3499 ();
 sg13g2_fill_2 FILLER_56_3513 ();
 sg13g2_fill_1 FILLER_56_3515 ();
 sg13g2_decap_8 FILLER_56_3525 ();
 sg13g2_decap_8 FILLER_56_3532 ();
 sg13g2_decap_8 FILLER_56_3539 ();
 sg13g2_decap_8 FILLER_56_3546 ();
 sg13g2_decap_8 FILLER_56_3553 ();
 sg13g2_decap_8 FILLER_56_3560 ();
 sg13g2_decap_8 FILLER_56_3567 ();
 sg13g2_decap_4 FILLER_56_3574 ();
 sg13g2_fill_2 FILLER_56_3578 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_36 ();
 sg13g2_fill_2 FILLER_57_54 ();
 sg13g2_fill_2 FILLER_57_83 ();
 sg13g2_fill_1 FILLER_57_85 ();
 sg13g2_fill_1 FILLER_57_96 ();
 sg13g2_decap_8 FILLER_57_149 ();
 sg13g2_decap_4 FILLER_57_224 ();
 sg13g2_fill_2 FILLER_57_246 ();
 sg13g2_fill_2 FILLER_57_261 ();
 sg13g2_fill_1 FILLER_57_313 ();
 sg13g2_decap_8 FILLER_57_318 ();
 sg13g2_fill_1 FILLER_57_325 ();
 sg13g2_fill_2 FILLER_57_343 ();
 sg13g2_fill_1 FILLER_57_345 ();
 sg13g2_fill_2 FILLER_57_373 ();
 sg13g2_fill_1 FILLER_57_416 ();
 sg13g2_decap_4 FILLER_57_448 ();
 sg13g2_fill_2 FILLER_57_479 ();
 sg13g2_fill_2 FILLER_57_494 ();
 sg13g2_fill_1 FILLER_57_496 ();
 sg13g2_fill_1 FILLER_57_501 ();
 sg13g2_decap_8 FILLER_57_508 ();
 sg13g2_fill_1 FILLER_57_515 ();
 sg13g2_decap_8 FILLER_57_550 ();
 sg13g2_decap_4 FILLER_57_557 ();
 sg13g2_fill_1 FILLER_57_600 ();
 sg13g2_decap_4 FILLER_57_610 ();
 sg13g2_fill_1 FILLER_57_622 ();
 sg13g2_fill_1 FILLER_57_627 ();
 sg13g2_decap_8 FILLER_57_633 ();
 sg13g2_decap_4 FILLER_57_640 ();
 sg13g2_decap_4 FILLER_57_666 ();
 sg13g2_decap_8 FILLER_57_701 ();
 sg13g2_fill_2 FILLER_57_708 ();
 sg13g2_fill_1 FILLER_57_710 ();
 sg13g2_fill_2 FILLER_57_756 ();
 sg13g2_fill_1 FILLER_57_758 ();
 sg13g2_fill_1 FILLER_57_777 ();
 sg13g2_fill_2 FILLER_57_805 ();
 sg13g2_fill_2 FILLER_57_816 ();
 sg13g2_fill_2 FILLER_57_869 ();
 sg13g2_fill_1 FILLER_57_871 ();
 sg13g2_fill_2 FILLER_57_885 ();
 sg13g2_fill_1 FILLER_57_887 ();
 sg13g2_fill_2 FILLER_57_920 ();
 sg13g2_fill_2 FILLER_57_927 ();
 sg13g2_fill_1 FILLER_57_929 ();
 sg13g2_fill_2 FILLER_57_966 ();
 sg13g2_fill_1 FILLER_57_968 ();
 sg13g2_decap_8 FILLER_57_1001 ();
 sg13g2_decap_4 FILLER_57_1008 ();
 sg13g2_fill_1 FILLER_57_1017 ();
 sg13g2_decap_4 FILLER_57_1065 ();
 sg13g2_fill_2 FILLER_57_1073 ();
 sg13g2_fill_1 FILLER_57_1075 ();
 sg13g2_decap_8 FILLER_57_1085 ();
 sg13g2_decap_4 FILLER_57_1092 ();
 sg13g2_fill_1 FILLER_57_1096 ();
 sg13g2_decap_4 FILLER_57_1168 ();
 sg13g2_fill_2 FILLER_57_1172 ();
 sg13g2_fill_2 FILLER_57_1188 ();
 sg13g2_fill_1 FILLER_57_1190 ();
 sg13g2_fill_2 FILLER_57_1196 ();
 sg13g2_fill_2 FILLER_57_1207 ();
 sg13g2_fill_1 FILLER_57_1209 ();
 sg13g2_fill_1 FILLER_57_1242 ();
 sg13g2_fill_1 FILLER_57_1261 ();
 sg13g2_decap_8 FILLER_57_1298 ();
 sg13g2_fill_2 FILLER_57_1305 ();
 sg13g2_fill_1 FILLER_57_1307 ();
 sg13g2_fill_1 FILLER_57_1357 ();
 sg13g2_fill_2 FILLER_57_1439 ();
 sg13g2_fill_2 FILLER_57_1468 ();
 sg13g2_decap_4 FILLER_57_1523 ();
 sg13g2_decap_4 FILLER_57_1531 ();
 sg13g2_fill_2 FILLER_57_1535 ();
 sg13g2_fill_2 FILLER_57_1542 ();
 sg13g2_fill_1 FILLER_57_1544 ();
 sg13g2_fill_1 FILLER_57_1634 ();
 sg13g2_fill_1 FILLER_57_1648 ();
 sg13g2_fill_1 FILLER_57_1677 ();
 sg13g2_fill_1 FILLER_57_1696 ();
 sg13g2_fill_1 FILLER_57_1710 ();
 sg13g2_fill_2 FILLER_57_1738 ();
 sg13g2_fill_1 FILLER_57_1740 ();
 sg13g2_fill_2 FILLER_57_1764 ();
 sg13g2_fill_2 FILLER_57_1859 ();
 sg13g2_decap_4 FILLER_57_1889 ();
 sg13g2_fill_1 FILLER_57_1893 ();
 sg13g2_fill_2 FILLER_57_1904 ();
 sg13g2_fill_1 FILLER_57_1906 ();
 sg13g2_fill_2 FILLER_57_1948 ();
 sg13g2_fill_1 FILLER_57_1950 ();
 sg13g2_fill_1 FILLER_57_1956 ();
 sg13g2_fill_2 FILLER_57_1993 ();
 sg13g2_fill_1 FILLER_57_1995 ();
 sg13g2_fill_1 FILLER_57_2071 ();
 sg13g2_decap_8 FILLER_57_2108 ();
 sg13g2_fill_2 FILLER_57_2115 ();
 sg13g2_fill_1 FILLER_57_2117 ();
 sg13g2_decap_4 FILLER_57_2158 ();
 sg13g2_fill_2 FILLER_57_2180 ();
 sg13g2_fill_1 FILLER_57_2182 ();
 sg13g2_fill_1 FILLER_57_2197 ();
 sg13g2_decap_8 FILLER_57_2224 ();
 sg13g2_decap_4 FILLER_57_2231 ();
 sg13g2_fill_2 FILLER_57_2235 ();
 sg13g2_fill_1 FILLER_57_2296 ();
 sg13g2_fill_2 FILLER_57_2306 ();
 sg13g2_fill_2 FILLER_57_2322 ();
 sg13g2_fill_1 FILLER_57_2324 ();
 sg13g2_decap_8 FILLER_57_2330 ();
 sg13g2_fill_1 FILLER_57_2337 ();
 sg13g2_fill_1 FILLER_57_2397 ();
 sg13g2_decap_8 FILLER_57_2420 ();
 sg13g2_decap_8 FILLER_57_2427 ();
 sg13g2_fill_1 FILLER_57_2461 ();
 sg13g2_fill_1 FILLER_57_2466 ();
 sg13g2_fill_2 FILLER_57_2476 ();
 sg13g2_fill_1 FILLER_57_2478 ();
 sg13g2_fill_1 FILLER_57_2497 ();
 sg13g2_fill_2 FILLER_57_2515 ();
 sg13g2_fill_2 FILLER_57_2571 ();
 sg13g2_decap_8 FILLER_57_2577 ();
 sg13g2_decap_4 FILLER_57_2584 ();
 sg13g2_fill_1 FILLER_57_2588 ();
 sg13g2_decap_4 FILLER_57_2611 ();
 sg13g2_fill_2 FILLER_57_2615 ();
 sg13g2_decap_8 FILLER_57_2635 ();
 sg13g2_fill_2 FILLER_57_2642 ();
 sg13g2_decap_4 FILLER_57_2666 ();
 sg13g2_fill_2 FILLER_57_2670 ();
 sg13g2_fill_2 FILLER_57_2676 ();
 sg13g2_fill_1 FILLER_57_2687 ();
 sg13g2_fill_2 FILLER_57_2710 ();
 sg13g2_fill_1 FILLER_57_2721 ();
 sg13g2_decap_8 FILLER_57_2739 ();
 sg13g2_fill_1 FILLER_57_2746 ();
 sg13g2_fill_2 FILLER_57_2751 ();
 sg13g2_decap_8 FILLER_57_2758 ();
 sg13g2_fill_1 FILLER_57_2811 ();
 sg13g2_fill_1 FILLER_57_2816 ();
 sg13g2_fill_1 FILLER_57_2834 ();
 sg13g2_fill_1 FILLER_57_2861 ();
 sg13g2_fill_1 FILLER_57_2875 ();
 sg13g2_decap_4 FILLER_57_2906 ();
 sg13g2_decap_8 FILLER_57_2955 ();
 sg13g2_decap_8 FILLER_57_2979 ();
 sg13g2_fill_2 FILLER_57_2986 ();
 sg13g2_fill_2 FILLER_57_3015 ();
 sg13g2_fill_2 FILLER_57_3058 ();
 sg13g2_fill_2 FILLER_57_3099 ();
 sg13g2_fill_2 FILLER_57_3111 ();
 sg13g2_fill_1 FILLER_57_3113 ();
 sg13g2_fill_1 FILLER_57_3167 ();
 sg13g2_fill_1 FILLER_57_3177 ();
 sg13g2_fill_1 FILLER_57_3248 ();
 sg13g2_fill_1 FILLER_57_3276 ();
 sg13g2_fill_2 FILLER_57_3286 ();
 sg13g2_fill_1 FILLER_57_3288 ();
 sg13g2_fill_1 FILLER_57_3316 ();
 sg13g2_fill_2 FILLER_57_3327 ();
 sg13g2_decap_8 FILLER_57_3344 ();
 sg13g2_fill_1 FILLER_57_3351 ();
 sg13g2_decap_4 FILLER_57_3357 ();
 sg13g2_decap_8 FILLER_57_3395 ();
 sg13g2_fill_2 FILLER_57_3402 ();
 sg13g2_decap_8 FILLER_57_3417 ();
 sg13g2_decap_8 FILLER_57_3424 ();
 sg13g2_decap_8 FILLER_57_3450 ();
 sg13g2_decap_4 FILLER_57_3457 ();
 sg13g2_fill_1 FILLER_57_3474 ();
 sg13g2_decap_8 FILLER_57_3485 ();
 sg13g2_fill_2 FILLER_57_3495 ();
 sg13g2_decap_8 FILLER_57_3528 ();
 sg13g2_decap_8 FILLER_57_3535 ();
 sg13g2_decap_8 FILLER_57_3542 ();
 sg13g2_decap_8 FILLER_57_3549 ();
 sg13g2_decap_8 FILLER_57_3556 ();
 sg13g2_decap_8 FILLER_57_3563 ();
 sg13g2_decap_8 FILLER_57_3570 ();
 sg13g2_fill_2 FILLER_57_3577 ();
 sg13g2_fill_1 FILLER_57_3579 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_11 ();
 sg13g2_decap_8 FILLER_58_17 ();
 sg13g2_decap_8 FILLER_58_24 ();
 sg13g2_fill_2 FILLER_58_31 ();
 sg13g2_fill_1 FILLER_58_33 ();
 sg13g2_decap_4 FILLER_58_41 ();
 sg13g2_decap_4 FILLER_58_69 ();
 sg13g2_fill_2 FILLER_58_73 ();
 sg13g2_decap_8 FILLER_58_81 ();
 sg13g2_fill_1 FILLER_58_88 ();
 sg13g2_fill_2 FILLER_58_102 ();
 sg13g2_fill_1 FILLER_58_104 ();
 sg13g2_fill_2 FILLER_58_140 ();
 sg13g2_fill_1 FILLER_58_142 ();
 sg13g2_decap_4 FILLER_58_156 ();
 sg13g2_fill_2 FILLER_58_160 ();
 sg13g2_fill_1 FILLER_58_172 ();
 sg13g2_decap_8 FILLER_58_209 ();
 sg13g2_fill_2 FILLER_58_216 ();
 sg13g2_decap_4 FILLER_58_240 ();
 sg13g2_fill_1 FILLER_58_244 ();
 sg13g2_fill_1 FILLER_58_250 ();
 sg13g2_fill_2 FILLER_58_264 ();
 sg13g2_fill_1 FILLER_58_266 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_decap_4 FILLER_58_322 ();
 sg13g2_fill_2 FILLER_58_336 ();
 sg13g2_fill_1 FILLER_58_338 ();
 sg13g2_fill_2 FILLER_58_349 ();
 sg13g2_fill_1 FILLER_58_351 ();
 sg13g2_fill_1 FILLER_58_360 ();
 sg13g2_fill_2 FILLER_58_410 ();
 sg13g2_fill_1 FILLER_58_412 ();
 sg13g2_fill_1 FILLER_58_497 ();
 sg13g2_decap_4 FILLER_58_507 ();
 sg13g2_fill_2 FILLER_58_511 ();
 sg13g2_decap_4 FILLER_58_522 ();
 sg13g2_decap_8 FILLER_58_542 ();
 sg13g2_decap_8 FILLER_58_549 ();
 sg13g2_fill_2 FILLER_58_556 ();
 sg13g2_fill_2 FILLER_58_585 ();
 sg13g2_fill_1 FILLER_58_587 ();
 sg13g2_fill_1 FILLER_58_640 ();
 sg13g2_fill_1 FILLER_58_659 ();
 sg13g2_fill_1 FILLER_58_700 ();
 sg13g2_fill_1 FILLER_58_750 ();
 sg13g2_fill_1 FILLER_58_855 ();
 sg13g2_fill_2 FILLER_58_888 ();
 sg13g2_fill_1 FILLER_58_890 ();
 sg13g2_fill_2 FILLER_58_904 ();
 sg13g2_fill_2 FILLER_58_911 ();
 sg13g2_fill_1 FILLER_58_913 ();
 sg13g2_fill_2 FILLER_58_950 ();
 sg13g2_fill_1 FILLER_58_952 ();
 sg13g2_fill_2 FILLER_58_987 ();
 sg13g2_fill_2 FILLER_58_1030 ();
 sg13g2_fill_1 FILLER_58_1032 ();
 sg13g2_fill_1 FILLER_58_1195 ();
 sg13g2_fill_1 FILLER_58_1244 ();
 sg13g2_fill_1 FILLER_58_1268 ();
 sg13g2_fill_1 FILLER_58_1283 ();
 sg13g2_fill_1 FILLER_58_1294 ();
 sg13g2_fill_2 FILLER_58_1323 ();
 sg13g2_fill_1 FILLER_58_1325 ();
 sg13g2_fill_2 FILLER_58_1353 ();
 sg13g2_fill_2 FILLER_58_1489 ();
 sg13g2_fill_1 FILLER_58_1491 ();
 sg13g2_fill_1 FILLER_58_1505 ();
 sg13g2_fill_2 FILLER_58_1511 ();
 sg13g2_fill_1 FILLER_58_1513 ();
 sg13g2_decap_4 FILLER_58_1523 ();
 sg13g2_fill_2 FILLER_58_1621 ();
 sg13g2_fill_1 FILLER_58_1623 ();
 sg13g2_fill_1 FILLER_58_1656 ();
 sg13g2_fill_2 FILLER_58_1737 ();
 sg13g2_fill_1 FILLER_58_1739 ();
 sg13g2_fill_1 FILLER_58_1762 ();
 sg13g2_fill_2 FILLER_58_1783 ();
 sg13g2_fill_1 FILLER_58_1785 ();
 sg13g2_decap_4 FILLER_58_1813 ();
 sg13g2_decap_8 FILLER_58_1822 ();
 sg13g2_decap_4 FILLER_58_1829 ();
 sg13g2_fill_2 FILLER_58_1833 ();
 sg13g2_fill_2 FILLER_58_1853 ();
 sg13g2_fill_1 FILLER_58_1855 ();
 sg13g2_fill_2 FILLER_58_1860 ();
 sg13g2_fill_1 FILLER_58_1862 ();
 sg13g2_fill_2 FILLER_58_1946 ();
 sg13g2_fill_2 FILLER_58_1953 ();
 sg13g2_fill_1 FILLER_58_1955 ();
 sg13g2_fill_2 FILLER_58_1969 ();
 sg13g2_fill_2 FILLER_58_2001 ();
 sg13g2_fill_1 FILLER_58_2003 ();
 sg13g2_fill_2 FILLER_58_2024 ();
 sg13g2_fill_1 FILLER_58_2026 ();
 sg13g2_fill_2 FILLER_58_2036 ();
 sg13g2_fill_1 FILLER_58_2038 ();
 sg13g2_decap_4 FILLER_58_2056 ();
 sg13g2_fill_1 FILLER_58_2060 ();
 sg13g2_fill_2 FILLER_58_2087 ();
 sg13g2_fill_1 FILLER_58_2115 ();
 sg13g2_decap_4 FILLER_58_2211 ();
 sg13g2_fill_2 FILLER_58_2254 ();
 sg13g2_fill_2 FILLER_58_2310 ();
 sg13g2_fill_2 FILLER_58_2336 ();
 sg13g2_fill_1 FILLER_58_2338 ();
 sg13g2_decap_8 FILLER_58_2358 ();
 sg13g2_decap_4 FILLER_58_2365 ();
 sg13g2_fill_2 FILLER_58_2369 ();
 sg13g2_fill_2 FILLER_58_2384 ();
 sg13g2_decap_4 FILLER_58_2395 ();
 sg13g2_fill_2 FILLER_58_2412 ();
 sg13g2_fill_1 FILLER_58_2414 ();
 sg13g2_fill_2 FILLER_58_2526 ();
 sg13g2_fill_2 FILLER_58_2541 ();
 sg13g2_fill_1 FILLER_58_2543 ();
 sg13g2_fill_2 FILLER_58_2577 ();
 sg13g2_fill_1 FILLER_58_2579 ();
 sg13g2_decap_4 FILLER_58_2585 ();
 sg13g2_decap_8 FILLER_58_2594 ();
 sg13g2_decap_8 FILLER_58_2601 ();
 sg13g2_fill_1 FILLER_58_2608 ();
 sg13g2_fill_2 FILLER_58_2619 ();
 sg13g2_fill_1 FILLER_58_2621 ();
 sg13g2_fill_2 FILLER_58_2654 ();
 sg13g2_fill_1 FILLER_58_2656 ();
 sg13g2_fill_1 FILLER_58_2716 ();
 sg13g2_fill_1 FILLER_58_2726 ();
 sg13g2_decap_4 FILLER_58_2760 ();
 sg13g2_fill_1 FILLER_58_2764 ();
 sg13g2_fill_2 FILLER_58_2779 ();
 sg13g2_fill_1 FILLER_58_2781 ();
 sg13g2_fill_1 FILLER_58_2799 ();
 sg13g2_fill_2 FILLER_58_2805 ();
 sg13g2_fill_1 FILLER_58_2807 ();
 sg13g2_fill_2 FILLER_58_2848 ();
 sg13g2_fill_2 FILLER_58_2864 ();
 sg13g2_fill_2 FILLER_58_2879 ();
 sg13g2_fill_2 FILLER_58_2891 ();
 sg13g2_decap_4 FILLER_58_2929 ();
 sg13g2_fill_1 FILLER_58_2933 ();
 sg13g2_decap_8 FILLER_58_2975 ();
 sg13g2_decap_4 FILLER_58_2982 ();
 sg13g2_fill_1 FILLER_58_2986 ();
 sg13g2_fill_1 FILLER_58_2996 ();
 sg13g2_fill_1 FILLER_58_3006 ();
 sg13g2_fill_1 FILLER_58_3028 ();
 sg13g2_decap_8 FILLER_58_3066 ();
 sg13g2_fill_1 FILLER_58_3106 ();
 sg13g2_fill_2 FILLER_58_3122 ();
 sg13g2_fill_1 FILLER_58_3146 ();
 sg13g2_fill_2 FILLER_58_3170 ();
 sg13g2_fill_1 FILLER_58_3181 ();
 sg13g2_fill_1 FILLER_58_3195 ();
 sg13g2_fill_2 FILLER_58_3251 ();
 sg13g2_fill_1 FILLER_58_3253 ();
 sg13g2_fill_2 FILLER_58_3285 ();
 sg13g2_fill_1 FILLER_58_3287 ();
 sg13g2_decap_4 FILLER_58_3375 ();
 sg13g2_fill_1 FILLER_58_3379 ();
 sg13g2_fill_1 FILLER_58_3406 ();
 sg13g2_decap_8 FILLER_58_3413 ();
 sg13g2_decap_4 FILLER_58_3420 ();
 sg13g2_fill_2 FILLER_58_3424 ();
 sg13g2_fill_1 FILLER_58_3440 ();
 sg13g2_decap_8 FILLER_58_3451 ();
 sg13g2_fill_1 FILLER_58_3458 ();
 sg13g2_fill_2 FILLER_58_3463 ();
 sg13g2_fill_2 FILLER_58_3473 ();
 sg13g2_fill_2 FILLER_58_3483 ();
 sg13g2_decap_8 FILLER_58_3544 ();
 sg13g2_decap_8 FILLER_58_3551 ();
 sg13g2_decap_8 FILLER_58_3558 ();
 sg13g2_decap_8 FILLER_58_3565 ();
 sg13g2_decap_8 FILLER_58_3572 ();
 sg13g2_fill_1 FILLER_58_3579 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_2 ();
 sg13g2_fill_1 FILLER_59_57 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_fill_1 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_76 ();
 sg13g2_fill_1 FILLER_59_110 ();
 sg13g2_fill_2 FILLER_59_174 ();
 sg13g2_fill_1 FILLER_59_176 ();
 sg13g2_fill_1 FILLER_59_246 ();
 sg13g2_fill_1 FILLER_59_275 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_decap_4 FILLER_59_308 ();
 sg13g2_fill_2 FILLER_59_325 ();
 sg13g2_fill_2 FILLER_59_337 ();
 sg13g2_fill_1 FILLER_59_339 ();
 sg13g2_fill_2 FILLER_59_376 ();
 sg13g2_decap_4 FILLER_59_400 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_fill_2 FILLER_59_462 ();
 sg13g2_fill_1 FILLER_59_464 ();
 sg13g2_fill_1 FILLER_59_492 ();
 sg13g2_fill_2 FILLER_59_602 ();
 sg13g2_fill_1 FILLER_59_604 ();
 sg13g2_decap_4 FILLER_59_633 ();
 sg13g2_fill_1 FILLER_59_667 ();
 sg13g2_fill_2 FILLER_59_697 ();
 sg13g2_fill_2 FILLER_59_744 ();
 sg13g2_fill_1 FILLER_59_746 ();
 sg13g2_fill_1 FILLER_59_788 ();
 sg13g2_fill_2 FILLER_59_816 ();
 sg13g2_fill_1 FILLER_59_818 ();
 sg13g2_fill_2 FILLER_59_833 ();
 sg13g2_fill_2 FILLER_59_863 ();
 sg13g2_decap_8 FILLER_59_879 ();
 sg13g2_fill_2 FILLER_59_891 ();
 sg13g2_fill_1 FILLER_59_893 ();
 sg13g2_fill_2 FILLER_59_935 ();
 sg13g2_fill_1 FILLER_59_937 ();
 sg13g2_fill_1 FILLER_59_947 ();
 sg13g2_fill_2 FILLER_59_958 ();
 sg13g2_fill_1 FILLER_59_965 ();
 sg13g2_fill_2 FILLER_59_971 ();
 sg13g2_fill_2 FILLER_59_978 ();
 sg13g2_fill_1 FILLER_59_980 ();
 sg13g2_decap_8 FILLER_59_985 ();
 sg13g2_decap_8 FILLER_59_992 ();
 sg13g2_fill_2 FILLER_59_999 ();
 sg13g2_fill_2 FILLER_59_1010 ();
 sg13g2_fill_1 FILLER_59_1012 ();
 sg13g2_fill_1 FILLER_59_1032 ();
 sg13g2_fill_1 FILLER_59_1051 ();
 sg13g2_fill_2 FILLER_59_1079 ();
 sg13g2_fill_2 FILLER_59_1117 ();
 sg13g2_decap_4 FILLER_59_1164 ();
 sg13g2_fill_2 FILLER_59_1196 ();
 sg13g2_fill_2 FILLER_59_1244 ();
 sg13g2_fill_1 FILLER_59_1280 ();
 sg13g2_fill_2 FILLER_59_1305 ();
 sg13g2_fill_2 FILLER_59_1325 ();
 sg13g2_fill_1 FILLER_59_1363 ();
 sg13g2_decap_8 FILLER_59_1404 ();
 sg13g2_decap_8 FILLER_59_1411 ();
 sg13g2_fill_1 FILLER_59_1418 ();
 sg13g2_decap_4 FILLER_59_1441 ();
 sg13g2_fill_1 FILLER_59_1458 ();
 sg13g2_fill_1 FILLER_59_1491 ();
 sg13g2_fill_2 FILLER_59_1497 ();
 sg13g2_fill_1 FILLER_59_1499 ();
 sg13g2_fill_2 FILLER_59_1556 ();
 sg13g2_fill_2 FILLER_59_1612 ();
 sg13g2_fill_1 FILLER_59_1614 ();
 sg13g2_fill_2 FILLER_59_1668 ();
 sg13g2_fill_2 FILLER_59_1683 ();
 sg13g2_fill_1 FILLER_59_1685 ();
 sg13g2_fill_2 FILLER_59_1728 ();
 sg13g2_fill_2 FILLER_59_1794 ();
 sg13g2_fill_1 FILLER_59_1796 ();
 sg13g2_fill_1 FILLER_59_1839 ();
 sg13g2_fill_2 FILLER_59_1867 ();
 sg13g2_fill_2 FILLER_59_1923 ();
 sg13g2_fill_2 FILLER_59_1943 ();
 sg13g2_fill_1 FILLER_59_1945 ();
 sg13g2_fill_2 FILLER_59_1987 ();
 sg13g2_fill_2 FILLER_59_2007 ();
 sg13g2_fill_2 FILLER_59_2023 ();
 sg13g2_fill_1 FILLER_59_2025 ();
 sg13g2_fill_2 FILLER_59_2058 ();
 sg13g2_fill_1 FILLER_59_2060 ();
 sg13g2_decap_8 FILLER_59_2094 ();
 sg13g2_fill_1 FILLER_59_2177 ();
 sg13g2_fill_2 FILLER_59_2202 ();
 sg13g2_fill_2 FILLER_59_2277 ();
 sg13g2_fill_2 FILLER_59_2288 ();
 sg13g2_fill_1 FILLER_59_2290 ();
 sg13g2_fill_1 FILLER_59_2313 ();
 sg13g2_fill_2 FILLER_59_2346 ();
 sg13g2_fill_2 FILLER_59_2394 ();
 sg13g2_fill_1 FILLER_59_2396 ();
 sg13g2_fill_2 FILLER_59_2424 ();
 sg13g2_fill_1 FILLER_59_2440 ();
 sg13g2_fill_2 FILLER_59_2459 ();
 sg13g2_fill_1 FILLER_59_2470 ();
 sg13g2_fill_1 FILLER_59_2495 ();
 sg13g2_fill_2 FILLER_59_2515 ();
 sg13g2_fill_1 FILLER_59_2649 ();
 sg13g2_fill_2 FILLER_59_2716 ();
 sg13g2_fill_1 FILLER_59_2718 ();
 sg13g2_fill_1 FILLER_59_2746 ();
 sg13g2_decap_8 FILLER_59_2784 ();
 sg13g2_fill_1 FILLER_59_2827 ();
 sg13g2_fill_2 FILLER_59_2837 ();
 sg13g2_fill_1 FILLER_59_2839 ();
 sg13g2_fill_2 FILLER_59_2868 ();
 sg13g2_fill_1 FILLER_59_2902 ();
 sg13g2_decap_8 FILLER_59_2908 ();
 sg13g2_fill_2 FILLER_59_2939 ();
 sg13g2_fill_1 FILLER_59_2941 ();
 sg13g2_fill_2 FILLER_59_2952 ();
 sg13g2_fill_1 FILLER_59_2954 ();
 sg13g2_fill_2 FILLER_59_3075 ();
 sg13g2_fill_1 FILLER_59_3077 ();
 sg13g2_fill_1 FILLER_59_3095 ();
 sg13g2_fill_1 FILLER_59_3101 ();
 sg13g2_fill_2 FILLER_59_3157 ();
 sg13g2_fill_1 FILLER_59_3196 ();
 sg13g2_fill_2 FILLER_59_3256 ();
 sg13g2_fill_1 FILLER_59_3258 ();
 sg13g2_decap_8 FILLER_59_3285 ();
 sg13g2_fill_1 FILLER_59_3292 ();
 sg13g2_fill_1 FILLER_59_3325 ();
 sg13g2_fill_1 FILLER_59_3335 ();
 sg13g2_decap_4 FILLER_59_3359 ();
 sg13g2_fill_2 FILLER_59_3363 ();
 sg13g2_decap_4 FILLER_59_3391 ();
 sg13g2_fill_1 FILLER_59_3395 ();
 sg13g2_decap_4 FILLER_59_3419 ();
 sg13g2_fill_1 FILLER_59_3430 ();
 sg13g2_decap_4 FILLER_59_3453 ();
 sg13g2_decap_4 FILLER_59_3463 ();
 sg13g2_fill_1 FILLER_59_3467 ();
 sg13g2_fill_2 FILLER_59_3487 ();
 sg13g2_fill_1 FILLER_59_3489 ();
 sg13g2_decap_4 FILLER_59_3517 ();
 sg13g2_fill_1 FILLER_59_3521 ();
 sg13g2_decap_8 FILLER_59_3526 ();
 sg13g2_decap_8 FILLER_59_3533 ();
 sg13g2_decap_8 FILLER_59_3540 ();
 sg13g2_decap_8 FILLER_59_3547 ();
 sg13g2_decap_8 FILLER_59_3554 ();
 sg13g2_decap_8 FILLER_59_3561 ();
 sg13g2_decap_8 FILLER_59_3568 ();
 sg13g2_decap_4 FILLER_59_3575 ();
 sg13g2_fill_1 FILLER_59_3579 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_fill_2 FILLER_60_51 ();
 sg13g2_fill_1 FILLER_60_53 ();
 sg13g2_decap_4 FILLER_60_83 ();
 sg13g2_decap_4 FILLER_60_96 ();
 sg13g2_fill_1 FILLER_60_100 ();
 sg13g2_fill_2 FILLER_60_136 ();
 sg13g2_fill_2 FILLER_60_148 ();
 sg13g2_fill_1 FILLER_60_169 ();
 sg13g2_fill_2 FILLER_60_206 ();
 sg13g2_fill_1 FILLER_60_208 ();
 sg13g2_fill_2 FILLER_60_226 ();
 sg13g2_fill_2 FILLER_60_251 ();
 sg13g2_fill_2 FILLER_60_280 ();
 sg13g2_fill_2 FILLER_60_310 ();
 sg13g2_decap_4 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_370 ();
 sg13g2_fill_1 FILLER_60_445 ();
 sg13g2_decap_8 FILLER_60_494 ();
 sg13g2_decap_8 FILLER_60_501 ();
 sg13g2_fill_1 FILLER_60_508 ();
 sg13g2_fill_1 FILLER_60_554 ();
 sg13g2_decap_8 FILLER_60_568 ();
 sg13g2_decap_8 FILLER_60_575 ();
 sg13g2_decap_4 FILLER_60_591 ();
 sg13g2_fill_1 FILLER_60_595 ();
 sg13g2_fill_1 FILLER_60_637 ();
 sg13g2_fill_2 FILLER_60_651 ();
 sg13g2_fill_1 FILLER_60_703 ();
 sg13g2_fill_2 FILLER_60_802 ();
 sg13g2_fill_1 FILLER_60_824 ();
 sg13g2_fill_2 FILLER_60_838 ();
 sg13g2_fill_2 FILLER_60_944 ();
 sg13g2_fill_2 FILLER_60_1047 ();
 sg13g2_fill_1 FILLER_60_1086 ();
 sg13g2_fill_2 FILLER_60_1100 ();
 sg13g2_fill_1 FILLER_60_1102 ();
 sg13g2_fill_2 FILLER_60_1133 ();
 sg13g2_fill_1 FILLER_60_1190 ();
 sg13g2_fill_2 FILLER_60_1196 ();
 sg13g2_decap_4 FILLER_60_1229 ();
 sg13g2_fill_1 FILLER_60_1265 ();
 sg13g2_fill_1 FILLER_60_1298 ();
 sg13g2_fill_2 FILLER_60_1335 ();
 sg13g2_fill_1 FILLER_60_1337 ();
 sg13g2_fill_2 FILLER_60_1383 ();
 sg13g2_fill_1 FILLER_60_1385 ();
 sg13g2_fill_1 FILLER_60_1391 ();
 sg13g2_fill_1 FILLER_60_1420 ();
 sg13g2_decap_4 FILLER_60_1434 ();
 sg13g2_fill_1 FILLER_60_1438 ();
 sg13g2_fill_1 FILLER_60_1444 ();
 sg13g2_fill_1 FILLER_60_1486 ();
 sg13g2_fill_2 FILLER_60_1501 ();
 sg13g2_fill_1 FILLER_60_1503 ();
 sg13g2_fill_2 FILLER_60_1518 ();
 sg13g2_fill_2 FILLER_60_1533 ();
 sg13g2_fill_1 FILLER_60_1535 ();
 sg13g2_fill_2 FILLER_60_1549 ();
 sg13g2_fill_1 FILLER_60_1551 ();
 sg13g2_fill_2 FILLER_60_1597 ();
 sg13g2_fill_1 FILLER_60_1599 ();
 sg13g2_fill_2 FILLER_60_1661 ();
 sg13g2_decap_4 FILLER_60_1705 ();
 sg13g2_fill_2 FILLER_60_1733 ();
 sg13g2_fill_2 FILLER_60_1763 ();
 sg13g2_fill_1 FILLER_60_1792 ();
 sg13g2_fill_1 FILLER_60_1802 ();
 sg13g2_decap_8 FILLER_60_1825 ();
 sg13g2_decap_4 FILLER_60_1832 ();
 sg13g2_decap_8 FILLER_60_1846 ();
 sg13g2_fill_1 FILLER_60_1853 ();
 sg13g2_fill_1 FILLER_60_1863 ();
 sg13g2_fill_1 FILLER_60_1886 ();
 sg13g2_fill_2 FILLER_60_1896 ();
 sg13g2_fill_1 FILLER_60_1898 ();
 sg13g2_fill_1 FILLER_60_1904 ();
 sg13g2_fill_1 FILLER_60_1933 ();
 sg13g2_fill_1 FILLER_60_1939 ();
 sg13g2_fill_2 FILLER_60_1949 ();
 sg13g2_fill_1 FILLER_60_1951 ();
 sg13g2_fill_1 FILLER_60_1961 ();
 sg13g2_fill_1 FILLER_60_2008 ();
 sg13g2_decap_8 FILLER_60_2036 ();
 sg13g2_fill_2 FILLER_60_2043 ();
 sg13g2_fill_1 FILLER_60_2045 ();
 sg13g2_fill_1 FILLER_60_2060 ();
 sg13g2_fill_2 FILLER_60_2099 ();
 sg13g2_fill_1 FILLER_60_2101 ();
 sg13g2_fill_2 FILLER_60_2130 ();
 sg13g2_fill_1 FILLER_60_2132 ();
 sg13g2_fill_2 FILLER_60_2160 ();
 sg13g2_fill_2 FILLER_60_2194 ();
 sg13g2_fill_1 FILLER_60_2223 ();
 sg13g2_decap_4 FILLER_60_2233 ();
 sg13g2_fill_2 FILLER_60_2282 ();
 sg13g2_fill_1 FILLER_60_2284 ();
 sg13g2_fill_1 FILLER_60_2298 ();
 sg13g2_fill_1 FILLER_60_2312 ();
 sg13g2_fill_2 FILLER_60_2322 ();
 sg13g2_fill_1 FILLER_60_2352 ();
 sg13g2_decap_4 FILLER_60_2366 ();
 sg13g2_fill_2 FILLER_60_2370 ();
 sg13g2_fill_2 FILLER_60_2454 ();
 sg13g2_fill_1 FILLER_60_2456 ();
 sg13g2_fill_2 FILLER_60_2485 ();
 sg13g2_decap_8 FILLER_60_2492 ();
 sg13g2_fill_1 FILLER_60_2499 ();
 sg13g2_decap_4 FILLER_60_2579 ();
 sg13g2_fill_1 FILLER_60_2598 ();
 sg13g2_fill_2 FILLER_60_2618 ();
 sg13g2_fill_2 FILLER_60_2652 ();
 sg13g2_fill_1 FILLER_60_2718 ();
 sg13g2_decap_4 FILLER_60_2756 ();
 sg13g2_fill_2 FILLER_60_2769 ();
 sg13g2_fill_1 FILLER_60_2771 ();
 sg13g2_decap_8 FILLER_60_2790 ();
 sg13g2_decap_4 FILLER_60_2797 ();
 sg13g2_fill_1 FILLER_60_2801 ();
 sg13g2_fill_1 FILLER_60_2811 ();
 sg13g2_fill_1 FILLER_60_2845 ();
 sg13g2_fill_1 FILLER_60_2859 ();
 sg13g2_decap_4 FILLER_60_2898 ();
 sg13g2_decap_8 FILLER_60_2930 ();
 sg13g2_fill_2 FILLER_60_2937 ();
 sg13g2_fill_2 FILLER_60_2944 ();
 sg13g2_fill_1 FILLER_60_2946 ();
 sg13g2_decap_4 FILLER_60_2969 ();
 sg13g2_fill_2 FILLER_60_3169 ();
 sg13g2_fill_1 FILLER_60_3171 ();
 sg13g2_fill_1 FILLER_60_3219 ();
 sg13g2_fill_1 FILLER_60_3229 ();
 sg13g2_fill_2 FILLER_60_3234 ();
 sg13g2_decap_4 FILLER_60_3272 ();
 sg13g2_fill_2 FILLER_60_3330 ();
 sg13g2_fill_1 FILLER_60_3332 ();
 sg13g2_decap_8 FILLER_60_3361 ();
 sg13g2_decap_4 FILLER_60_3368 ();
 sg13g2_fill_1 FILLER_60_3372 ();
 sg13g2_decap_4 FILLER_60_3401 ();
 sg13g2_fill_1 FILLER_60_3405 ();
 sg13g2_decap_4 FILLER_60_3414 ();
 sg13g2_fill_1 FILLER_60_3418 ();
 sg13g2_fill_2 FILLER_60_3433 ();
 sg13g2_decap_8 FILLER_60_3448 ();
 sg13g2_decap_8 FILLER_60_3455 ();
 sg13g2_fill_2 FILLER_60_3462 ();
 sg13g2_fill_1 FILLER_60_3464 ();
 sg13g2_fill_2 FILLER_60_3478 ();
 sg13g2_fill_2 FILLER_60_3505 ();
 sg13g2_decap_8 FILLER_60_3544 ();
 sg13g2_decap_8 FILLER_60_3551 ();
 sg13g2_decap_8 FILLER_60_3558 ();
 sg13g2_decap_8 FILLER_60_3565 ();
 sg13g2_decap_8 FILLER_60_3572 ();
 sg13g2_fill_1 FILLER_60_3579 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_15 ();
 sg13g2_fill_2 FILLER_61_22 ();
 sg13g2_fill_1 FILLER_61_46 ();
 sg13g2_fill_1 FILLER_61_51 ();
 sg13g2_decap_8 FILLER_61_59 ();
 sg13g2_decap_8 FILLER_61_66 ();
 sg13g2_fill_2 FILLER_61_73 ();
 sg13g2_fill_1 FILLER_61_75 ();
 sg13g2_fill_1 FILLER_61_80 ();
 sg13g2_fill_1 FILLER_61_109 ();
 sg13g2_fill_2 FILLER_61_191 ();
 sg13g2_decap_8 FILLER_61_303 ();
 sg13g2_decap_8 FILLER_61_310 ();
 sg13g2_decap_4 FILLER_61_317 ();
 sg13g2_fill_2 FILLER_61_345 ();
 sg13g2_fill_1 FILLER_61_347 ();
 sg13g2_fill_2 FILLER_61_361 ();
 sg13g2_fill_2 FILLER_61_372 ();
 sg13g2_fill_1 FILLER_61_374 ();
 sg13g2_fill_2 FILLER_61_389 ();
 sg13g2_fill_2 FILLER_61_414 ();
 sg13g2_fill_1 FILLER_61_416 ();
 sg13g2_fill_2 FILLER_61_421 ();
 sg13g2_fill_1 FILLER_61_423 ();
 sg13g2_decap_8 FILLER_61_437 ();
 sg13g2_decap_8 FILLER_61_444 ();
 sg13g2_fill_2 FILLER_61_451 ();
 sg13g2_fill_1 FILLER_61_453 ();
 sg13g2_fill_1 FILLER_61_465 ();
 sg13g2_decap_8 FILLER_61_476 ();
 sg13g2_decap_8 FILLER_61_483 ();
 sg13g2_fill_2 FILLER_61_517 ();
 sg13g2_decap_8 FILLER_61_533 ();
 sg13g2_decap_8 FILLER_61_540 ();
 sg13g2_fill_2 FILLER_61_551 ();
 sg13g2_fill_1 FILLER_61_553 ();
 sg13g2_decap_8 FILLER_61_591 ();
 sg13g2_decap_8 FILLER_61_598 ();
 sg13g2_fill_2 FILLER_61_605 ();
 sg13g2_fill_1 FILLER_61_617 ();
 sg13g2_fill_2 FILLER_61_641 ();
 sg13g2_fill_1 FILLER_61_643 ();
 sg13g2_fill_1 FILLER_61_727 ();
 sg13g2_fill_1 FILLER_61_741 ();
 sg13g2_fill_2 FILLER_61_779 ();
 sg13g2_fill_1 FILLER_61_794 ();
 sg13g2_fill_1 FILLER_61_827 ();
 sg13g2_fill_1 FILLER_61_836 ();
 sg13g2_fill_2 FILLER_61_841 ();
 sg13g2_fill_1 FILLER_61_871 ();
 sg13g2_decap_4 FILLER_61_882 ();
 sg13g2_fill_2 FILLER_61_944 ();
 sg13g2_fill_1 FILLER_61_946 ();
 sg13g2_decap_8 FILLER_61_979 ();
 sg13g2_fill_1 FILLER_61_986 ();
 sg13g2_fill_2 FILLER_61_1023 ();
 sg13g2_fill_1 FILLER_61_1025 ();
 sg13g2_fill_1 FILLER_61_1068 ();
 sg13g2_fill_1 FILLER_61_1105 ();
 sg13g2_fill_2 FILLER_61_1153 ();
 sg13g2_fill_2 FILLER_61_1174 ();
 sg13g2_fill_1 FILLER_61_1176 ();
 sg13g2_fill_1 FILLER_61_1190 ();
 sg13g2_decap_8 FILLER_61_1228 ();
 sg13g2_decap_4 FILLER_61_1235 ();
 sg13g2_fill_2 FILLER_61_1262 ();
 sg13g2_fill_1 FILLER_61_1264 ();
 sg13g2_decap_4 FILLER_61_1302 ();
 sg13g2_decap_4 FILLER_61_1316 ();
 sg13g2_decap_4 FILLER_61_1371 ();
 sg13g2_fill_2 FILLER_61_1375 ();
 sg13g2_decap_4 FILLER_61_1387 ();
 sg13g2_fill_1 FILLER_61_1391 ();
 sg13g2_decap_4 FILLER_61_1410 ();
 sg13g2_fill_2 FILLER_61_1414 ();
 sg13g2_fill_2 FILLER_61_1429 ();
 sg13g2_fill_1 FILLER_61_1431 ();
 sg13g2_decap_4 FILLER_61_1459 ();
 sg13g2_fill_1 FILLER_61_1489 ();
 sg13g2_fill_2 FILLER_61_1527 ();
 sg13g2_fill_1 FILLER_61_1529 ();
 sg13g2_fill_1 FILLER_61_1583 ();
 sg13g2_fill_2 FILLER_61_1612 ();
 sg13g2_decap_4 FILLER_61_1623 ();
 sg13g2_fill_1 FILLER_61_1655 ();
 sg13g2_fill_2 FILLER_61_1661 ();
 sg13g2_fill_2 FILLER_61_1676 ();
 sg13g2_fill_2 FILLER_61_1687 ();
 sg13g2_fill_2 FILLER_61_1730 ();
 sg13g2_fill_1 FILLER_61_1732 ();
 sg13g2_decap_8 FILLER_61_1773 ();
 sg13g2_fill_1 FILLER_61_1830 ();
 sg13g2_fill_2 FILLER_61_1841 ();
 sg13g2_fill_1 FILLER_61_1843 ();
 sg13g2_decap_8 FILLER_61_1871 ();
 sg13g2_fill_1 FILLER_61_2021 ();
 sg13g2_decap_4 FILLER_61_2086 ();
 sg13g2_decap_4 FILLER_61_2225 ();
 sg13g2_decap_8 FILLER_61_2238 ();
 sg13g2_fill_2 FILLER_61_2274 ();
 sg13g2_fill_2 FILLER_61_2304 ();
 sg13g2_fill_1 FILLER_61_2306 ();
 sg13g2_decap_4 FILLER_61_2363 ();
 sg13g2_decap_8 FILLER_61_2412 ();
 sg13g2_decap_8 FILLER_61_2478 ();
 sg13g2_fill_2 FILLER_61_2485 ();
 sg13g2_decap_4 FILLER_61_2545 ();
 sg13g2_fill_2 FILLER_61_2566 ();
 sg13g2_decap_4 FILLER_61_2595 ();
 sg13g2_fill_2 FILLER_61_2599 ();
 sg13g2_fill_2 FILLER_61_2628 ();
 sg13g2_fill_2 FILLER_61_2639 ();
 sg13g2_fill_1 FILLER_61_2655 ();
 sg13g2_decap_4 FILLER_61_2683 ();
 sg13g2_decap_8 FILLER_61_2691 ();
 sg13g2_fill_1 FILLER_61_2698 ();
 sg13g2_fill_2 FILLER_61_2713 ();
 sg13g2_fill_2 FILLER_61_2802 ();
 sg13g2_fill_1 FILLER_61_2804 ();
 sg13g2_fill_1 FILLER_61_2814 ();
 sg13g2_decap_4 FILLER_61_2868 ();
 sg13g2_decap_8 FILLER_61_2914 ();
 sg13g2_fill_1 FILLER_61_2921 ();
 sg13g2_fill_1 FILLER_61_2935 ();
 sg13g2_decap_4 FILLER_61_2985 ();
 sg13g2_fill_1 FILLER_61_3022 ();
 sg13g2_decap_4 FILLER_61_3050 ();
 sg13g2_decap_8 FILLER_61_3059 ();
 sg13g2_decap_4 FILLER_61_3066 ();
 sg13g2_fill_1 FILLER_61_3070 ();
 sg13g2_fill_2 FILLER_61_3084 ();
 sg13g2_fill_1 FILLER_61_3086 ();
 sg13g2_fill_2 FILLER_61_3096 ();
 sg13g2_decap_8 FILLER_61_3127 ();
 sg13g2_fill_1 FILLER_61_3134 ();
 sg13g2_fill_1 FILLER_61_3246 ();
 sg13g2_fill_1 FILLER_61_3329 ();
 sg13g2_fill_1 FILLER_61_3373 ();
 sg13g2_decap_8 FILLER_61_3412 ();
 sg13g2_decap_4 FILLER_61_3427 ();
 sg13g2_fill_2 FILLER_61_3431 ();
 sg13g2_decap_4 FILLER_61_3451 ();
 sg13g2_fill_1 FILLER_61_3455 ();
 sg13g2_decap_4 FILLER_61_3463 ();
 sg13g2_fill_1 FILLER_61_3467 ();
 sg13g2_fill_2 FILLER_61_3482 ();
 sg13g2_fill_2 FILLER_61_3491 ();
 sg13g2_fill_1 FILLER_61_3493 ();
 sg13g2_decap_8 FILLER_61_3525 ();
 sg13g2_decap_8 FILLER_61_3532 ();
 sg13g2_decap_8 FILLER_61_3539 ();
 sg13g2_decap_8 FILLER_61_3546 ();
 sg13g2_decap_8 FILLER_61_3553 ();
 sg13g2_decap_8 FILLER_61_3560 ();
 sg13g2_decap_8 FILLER_61_3567 ();
 sg13g2_decap_4 FILLER_61_3574 ();
 sg13g2_fill_2 FILLER_61_3578 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_1 FILLER_62_64 ();
 sg13g2_fill_2 FILLER_62_74 ();
 sg13g2_fill_1 FILLER_62_76 ();
 sg13g2_decap_4 FILLER_62_82 ();
 sg13g2_decap_4 FILLER_62_95 ();
 sg13g2_fill_2 FILLER_62_99 ();
 sg13g2_fill_1 FILLER_62_128 ();
 sg13g2_fill_1 FILLER_62_152 ();
 sg13g2_fill_1 FILLER_62_167 ();
 sg13g2_decap_4 FILLER_62_193 ();
 sg13g2_fill_2 FILLER_62_197 ();
 sg13g2_decap_8 FILLER_62_235 ();
 sg13g2_decap_8 FILLER_62_242 ();
 sg13g2_decap_4 FILLER_62_249 ();
 sg13g2_fill_2 FILLER_62_281 ();
 sg13g2_decap_8 FILLER_62_292 ();
 sg13g2_decap_4 FILLER_62_299 ();
 sg13g2_decap_4 FILLER_62_307 ();
 sg13g2_fill_1 FILLER_62_311 ();
 sg13g2_fill_2 FILLER_62_384 ();
 sg13g2_fill_1 FILLER_62_386 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_fill_2 FILLER_62_434 ();
 sg13g2_fill_2 FILLER_62_468 ();
 sg13g2_fill_1 FILLER_62_470 ();
 sg13g2_fill_2 FILLER_62_498 ();
 sg13g2_fill_1 FILLER_62_500 ();
 sg13g2_fill_1 FILLER_62_515 ();
 sg13g2_decap_8 FILLER_62_520 ();
 sg13g2_decap_8 FILLER_62_555 ();
 sg13g2_decap_4 FILLER_62_562 ();
 sg13g2_fill_1 FILLER_62_566 ();
 sg13g2_fill_2 FILLER_62_657 ();
 sg13g2_fill_1 FILLER_62_696 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_fill_1 FILLER_62_721 ();
 sg13g2_fill_2 FILLER_62_813 ();
 sg13g2_decap_4 FILLER_62_870 ();
 sg13g2_decap_4 FILLER_62_910 ();
 sg13g2_fill_1 FILLER_62_914 ();
 sg13g2_decap_4 FILLER_62_952 ();
 sg13g2_decap_8 FILLER_62_978 ();
 sg13g2_decap_8 FILLER_62_985 ();
 sg13g2_decap_8 FILLER_62_992 ();
 sg13g2_fill_2 FILLER_62_1014 ();
 sg13g2_fill_1 FILLER_62_1016 ();
 sg13g2_decap_8 FILLER_62_1044 ();
 sg13g2_decap_8 FILLER_62_1144 ();
 sg13g2_fill_1 FILLER_62_1151 ();
 sg13g2_fill_1 FILLER_62_1165 ();
 sg13g2_fill_2 FILLER_62_1212 ();
 sg13g2_decap_8 FILLER_62_1223 ();
 sg13g2_decap_4 FILLER_62_1230 ();
 sg13g2_fill_1 FILLER_62_1234 ();
 sg13g2_decap_8 FILLER_62_1262 ();
 sg13g2_fill_1 FILLER_62_1269 ();
 sg13g2_decap_4 FILLER_62_1306 ();
 sg13g2_fill_1 FILLER_62_1310 ();
 sg13g2_decap_4 FILLER_62_1382 ();
 sg13g2_fill_2 FILLER_62_1423 ();
 sg13g2_decap_4 FILLER_62_1453 ();
 sg13g2_fill_1 FILLER_62_1457 ();
 sg13g2_decap_4 FILLER_62_1523 ();
 sg13g2_fill_2 FILLER_62_1582 ();
 sg13g2_fill_1 FILLER_62_1584 ();
 sg13g2_fill_2 FILLER_62_1636 ();
 sg13g2_decap_4 FILLER_62_1734 ();
 sg13g2_decap_4 FILLER_62_1751 ();
 sg13g2_fill_1 FILLER_62_1755 ();
 sg13g2_fill_1 FILLER_62_1802 ();
 sg13g2_fill_2 FILLER_62_1808 ();
 sg13g2_fill_2 FILLER_62_1820 ();
 sg13g2_decap_8 FILLER_62_1831 ();
 sg13g2_fill_1 FILLER_62_1838 ();
 sg13g2_decap_4 FILLER_62_1875 ();
 sg13g2_decap_4 FILLER_62_1924 ();
 sg13g2_fill_1 FILLER_62_1982 ();
 sg13g2_decap_4 FILLER_62_2011 ();
 sg13g2_fill_1 FILLER_62_2015 ();
 sg13g2_fill_2 FILLER_62_2020 ();
 sg13g2_decap_4 FILLER_62_2035 ();
 sg13g2_fill_1 FILLER_62_2052 ();
 sg13g2_decap_4 FILLER_62_2071 ();
 sg13g2_fill_1 FILLER_62_2119 ();
 sg13g2_fill_1 FILLER_62_2130 ();
 sg13g2_decap_8 FILLER_62_2144 ();
 sg13g2_fill_1 FILLER_62_2151 ();
 sg13g2_fill_2 FILLER_62_2175 ();
 sg13g2_fill_1 FILLER_62_2177 ();
 sg13g2_fill_2 FILLER_62_2191 ();
 sg13g2_fill_1 FILLER_62_2193 ();
 sg13g2_fill_2 FILLER_62_2209 ();
 sg13g2_fill_1 FILLER_62_2211 ();
 sg13g2_fill_1 FILLER_62_2239 ();
 sg13g2_fill_2 FILLER_62_2272 ();
 sg13g2_fill_1 FILLER_62_2274 ();
 sg13g2_fill_1 FILLER_62_2331 ();
 sg13g2_decap_8 FILLER_62_2342 ();
 sg13g2_fill_1 FILLER_62_2349 ();
 sg13g2_decap_4 FILLER_62_2360 ();
 sg13g2_fill_2 FILLER_62_2364 ();
 sg13g2_fill_1 FILLER_62_2415 ();
 sg13g2_fill_2 FILLER_62_2472 ();
 sg13g2_fill_1 FILLER_62_2474 ();
 sg13g2_decap_8 FILLER_62_2494 ();
 sg13g2_decap_8 FILLER_62_2510 ();
 sg13g2_fill_2 FILLER_62_2517 ();
 sg13g2_fill_1 FILLER_62_2519 ();
 sg13g2_decap_4 FILLER_62_2607 ();
 sg13g2_fill_2 FILLER_62_2611 ();
 sg13g2_fill_2 FILLER_62_2659 ();
 sg13g2_fill_2 FILLER_62_2689 ();
 sg13g2_fill_2 FILLER_62_2718 ();
 sg13g2_fill_1 FILLER_62_2747 ();
 sg13g2_fill_2 FILLER_62_2785 ();
 sg13g2_fill_2 FILLER_62_2819 ();
 sg13g2_decap_4 FILLER_62_2834 ();
 sg13g2_fill_2 FILLER_62_2838 ();
 sg13g2_decap_4 FILLER_62_2885 ();
 sg13g2_fill_2 FILLER_62_2889 ();
 sg13g2_fill_1 FILLER_62_2924 ();
 sg13g2_decap_4 FILLER_62_2930 ();
 sg13g2_decap_8 FILLER_62_2957 ();
 sg13g2_fill_1 FILLER_62_2964 ();
 sg13g2_fill_2 FILLER_62_2975 ();
 sg13g2_fill_2 FILLER_62_3014 ();
 sg13g2_fill_1 FILLER_62_3016 ();
 sg13g2_decap_4 FILLER_62_3026 ();
 sg13g2_decap_8 FILLER_62_3040 ();
 sg13g2_fill_1 FILLER_62_3047 ();
 sg13g2_decap_4 FILLER_62_3107 ();
 sg13g2_fill_2 FILLER_62_3138 ();
 sg13g2_decap_8 FILLER_62_3178 ();
 sg13g2_fill_1 FILLER_62_3185 ();
 sg13g2_fill_1 FILLER_62_3311 ();
 sg13g2_fill_2 FILLER_62_3318 ();
 sg13g2_fill_1 FILLER_62_3320 ();
 sg13g2_fill_1 FILLER_62_3343 ();
 sg13g2_fill_1 FILLER_62_3425 ();
 sg13g2_fill_2 FILLER_62_3450 ();
 sg13g2_fill_1 FILLER_62_3452 ();
 sg13g2_decap_8 FILLER_62_3496 ();
 sg13g2_decap_8 FILLER_62_3507 ();
 sg13g2_decap_8 FILLER_62_3523 ();
 sg13g2_decap_8 FILLER_62_3530 ();
 sg13g2_decap_8 FILLER_62_3537 ();
 sg13g2_decap_8 FILLER_62_3544 ();
 sg13g2_decap_8 FILLER_62_3551 ();
 sg13g2_decap_8 FILLER_62_3558 ();
 sg13g2_decap_8 FILLER_62_3565 ();
 sg13g2_decap_8 FILLER_62_3572 ();
 sg13g2_fill_1 FILLER_62_3579 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_35 ();
 sg13g2_fill_1 FILLER_63_45 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_4 FILLER_63_77 ();
 sg13g2_fill_2 FILLER_63_125 ();
 sg13g2_fill_1 FILLER_63_172 ();
 sg13g2_fill_2 FILLER_63_228 ();
 sg13g2_fill_1 FILLER_63_230 ();
 sg13g2_fill_2 FILLER_63_355 ();
 sg13g2_fill_1 FILLER_63_389 ();
 sg13g2_fill_1 FILLER_63_422 ();
 sg13g2_fill_2 FILLER_63_442 ();
 sg13g2_fill_2 FILLER_63_471 ();
 sg13g2_fill_1 FILLER_63_473 ();
 sg13g2_fill_1 FILLER_63_483 ();
 sg13g2_fill_2 FILLER_63_493 ();
 sg13g2_fill_1 FILLER_63_495 ();
 sg13g2_fill_2 FILLER_63_565 ();
 sg13g2_fill_2 FILLER_63_608 ();
 sg13g2_fill_2 FILLER_63_623 ();
 sg13g2_fill_1 FILLER_63_625 ();
 sg13g2_fill_2 FILLER_63_653 ();
 sg13g2_fill_1 FILLER_63_655 ();
 sg13g2_decap_8 FILLER_63_761 ();
 sg13g2_fill_1 FILLER_63_768 ();
 sg13g2_fill_2 FILLER_63_791 ();
 sg13g2_fill_1 FILLER_63_793 ();
 sg13g2_fill_2 FILLER_63_853 ();
 sg13g2_decap_8 FILLER_63_865 ();
 sg13g2_decap_4 FILLER_63_872 ();
 sg13g2_decap_8 FILLER_63_885 ();
 sg13g2_fill_2 FILLER_63_892 ();
 sg13g2_fill_1 FILLER_63_894 ();
 sg13g2_fill_2 FILLER_63_932 ();
 sg13g2_fill_1 FILLER_63_934 ();
 sg13g2_fill_2 FILLER_63_1018 ();
 sg13g2_fill_2 FILLER_63_1047 ();
 sg13g2_fill_2 FILLER_63_1106 ();
 sg13g2_fill_2 FILLER_63_1136 ();
 sg13g2_fill_1 FILLER_63_1138 ();
 sg13g2_fill_2 FILLER_63_1152 ();
 sg13g2_fill_1 FILLER_63_1154 ();
 sg13g2_decap_4 FILLER_63_1187 ();
 sg13g2_fill_2 FILLER_63_1209 ();
 sg13g2_decap_8 FILLER_63_1270 ();
 sg13g2_fill_2 FILLER_63_1290 ();
 sg13g2_fill_2 FILLER_63_1316 ();
 sg13g2_fill_1 FILLER_63_1318 ();
 sg13g2_decap_8 FILLER_63_1341 ();
 sg13g2_fill_1 FILLER_63_1348 ();
 sg13g2_decap_8 FILLER_63_1362 ();
 sg13g2_decap_4 FILLER_63_1378 ();
 sg13g2_fill_1 FILLER_63_1382 ();
 sg13g2_decap_8 FILLER_63_1420 ();
 sg13g2_fill_2 FILLER_63_1427 ();
 sg13g2_decap_8 FILLER_63_1456 ();
 sg13g2_fill_1 FILLER_63_1463 ();
 sg13g2_fill_2 FILLER_63_1477 ();
 sg13g2_fill_1 FILLER_63_1506 ();
 sg13g2_decap_4 FILLER_63_1565 ();
 sg13g2_fill_1 FILLER_63_1596 ();
 sg13g2_decap_8 FILLER_63_1629 ();
 sg13g2_fill_1 FILLER_63_1668 ();
 sg13g2_fill_1 FILLER_63_1701 ();
 sg13g2_decap_8 FILLER_63_1729 ();
 sg13g2_fill_1 FILLER_63_1736 ();
 sg13g2_fill_2 FILLER_63_1787 ();
 sg13g2_fill_1 FILLER_63_1789 ();
 sg13g2_decap_4 FILLER_63_1803 ();
 sg13g2_fill_2 FILLER_63_1831 ();
 sg13g2_fill_1 FILLER_63_1849 ();
 sg13g2_fill_2 FILLER_63_1872 ();
 sg13g2_fill_1 FILLER_63_1874 ();
 sg13g2_fill_1 FILLER_63_1917 ();
 sg13g2_fill_1 FILLER_63_1947 ();
 sg13g2_decap_4 FILLER_63_1970 ();
 sg13g2_fill_1 FILLER_63_1974 ();
 sg13g2_decap_8 FILLER_63_1992 ();
 sg13g2_decap_8 FILLER_63_1999 ();
 sg13g2_fill_2 FILLER_63_2006 ();
 sg13g2_decap_4 FILLER_63_2045 ();
 sg13g2_decap_4 FILLER_63_2077 ();
 sg13g2_fill_1 FILLER_63_2081 ();
 sg13g2_fill_2 FILLER_63_2121 ();
 sg13g2_fill_1 FILLER_63_2123 ();
 sg13g2_fill_1 FILLER_63_2178 ();
 sg13g2_decap_4 FILLER_63_2243 ();
 sg13g2_fill_2 FILLER_63_2247 ();
 sg13g2_fill_1 FILLER_63_2317 ();
 sg13g2_fill_1 FILLER_63_2458 ();
 sg13g2_fill_2 FILLER_63_2513 ();
 sg13g2_fill_1 FILLER_63_2515 ();
 sg13g2_fill_2 FILLER_63_2579 ();
 sg13g2_fill_1 FILLER_63_2581 ();
 sg13g2_fill_2 FILLER_63_2597 ();
 sg13g2_fill_2 FILLER_63_2658 ();
 sg13g2_fill_1 FILLER_63_2660 ();
 sg13g2_decap_8 FILLER_63_2674 ();
 sg13g2_decap_8 FILLER_63_2681 ();
 sg13g2_fill_2 FILLER_63_2698 ();
 sg13g2_fill_1 FILLER_63_2709 ();
 sg13g2_decap_8 FILLER_63_2747 ();
 sg13g2_decap_4 FILLER_63_2754 ();
 sg13g2_fill_1 FILLER_63_2767 ();
 sg13g2_fill_2 FILLER_63_2786 ();
 sg13g2_decap_4 FILLER_63_2847 ();
 sg13g2_decap_4 FILLER_63_2891 ();
 sg13g2_fill_1 FILLER_63_2895 ();
 sg13g2_fill_1 FILLER_63_2932 ();
 sg13g2_decap_4 FILLER_63_2943 ();
 sg13g2_fill_1 FILLER_63_2947 ();
 sg13g2_fill_2 FILLER_63_2975 ();
 sg13g2_fill_1 FILLER_63_2981 ();
 sg13g2_fill_2 FILLER_63_3013 ();
 sg13g2_fill_1 FILLER_63_3052 ();
 sg13g2_fill_1 FILLER_63_3072 ();
 sg13g2_fill_2 FILLER_63_3114 ();
 sg13g2_fill_1 FILLER_63_3116 ();
 sg13g2_fill_2 FILLER_63_3145 ();
 sg13g2_fill_1 FILLER_63_3147 ();
 sg13g2_fill_2 FILLER_63_3202 ();
 sg13g2_fill_1 FILLER_63_3204 ();
 sg13g2_decap_8 FILLER_63_3236 ();
 sg13g2_decap_4 FILLER_63_3270 ();
 sg13g2_fill_2 FILLER_63_3300 ();
 sg13g2_fill_1 FILLER_63_3302 ();
 sg13g2_fill_1 FILLER_63_3308 ();
 sg13g2_fill_1 FILLER_63_3332 ();
 sg13g2_decap_8 FILLER_63_3339 ();
 sg13g2_decap_8 FILLER_63_3346 ();
 sg13g2_fill_1 FILLER_63_3353 ();
 sg13g2_fill_2 FILLER_63_3371 ();
 sg13g2_fill_1 FILLER_63_3382 ();
 sg13g2_fill_2 FILLER_63_3400 ();
 sg13g2_decap_4 FILLER_63_3419 ();
 sg13g2_fill_2 FILLER_63_3429 ();
 sg13g2_decap_8 FILLER_63_3481 ();
 sg13g2_decap_8 FILLER_63_3488 ();
 sg13g2_decap_8 FILLER_63_3495 ();
 sg13g2_decap_8 FILLER_63_3502 ();
 sg13g2_decap_8 FILLER_63_3509 ();
 sg13g2_decap_8 FILLER_63_3516 ();
 sg13g2_decap_8 FILLER_63_3523 ();
 sg13g2_decap_8 FILLER_63_3530 ();
 sg13g2_decap_8 FILLER_63_3537 ();
 sg13g2_decap_8 FILLER_63_3544 ();
 sg13g2_decap_8 FILLER_63_3551 ();
 sg13g2_decap_8 FILLER_63_3558 ();
 sg13g2_decap_8 FILLER_63_3565 ();
 sg13g2_decap_8 FILLER_63_3572 ();
 sg13g2_fill_1 FILLER_63_3579 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_11 ();
 sg13g2_decap_8 FILLER_64_17 ();
 sg13g2_fill_1 FILLER_64_33 ();
 sg13g2_fill_2 FILLER_64_59 ();
 sg13g2_decap_8 FILLER_64_66 ();
 sg13g2_fill_2 FILLER_64_73 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_fill_2 FILLER_64_107 ();
 sg13g2_fill_1 FILLER_64_109 ();
 sg13g2_fill_1 FILLER_64_150 ();
 sg13g2_fill_1 FILLER_64_164 ();
 sg13g2_decap_4 FILLER_64_269 ();
 sg13g2_fill_1 FILLER_64_273 ();
 sg13g2_fill_1 FILLER_64_284 ();
 sg13g2_fill_2 FILLER_64_303 ();
 sg13g2_fill_1 FILLER_64_305 ();
 sg13g2_fill_2 FILLER_64_333 ();
 sg13g2_fill_1 FILLER_64_335 ();
 sg13g2_fill_1 FILLER_64_406 ();
 sg13g2_decap_4 FILLER_64_444 ();
 sg13g2_decap_4 FILLER_64_461 ();
 sg13g2_fill_2 FILLER_64_493 ();
 sg13g2_fill_2 FILLER_64_510 ();
 sg13g2_fill_2 FILLER_64_525 ();
 sg13g2_fill_1 FILLER_64_527 ();
 sg13g2_fill_2 FILLER_64_580 ();
 sg13g2_fill_1 FILLER_64_582 ();
 sg13g2_fill_2 FILLER_64_597 ();
 sg13g2_fill_1 FILLER_64_604 ();
 sg13g2_fill_2 FILLER_64_610 ();
 sg13g2_fill_1 FILLER_64_612 ();
 sg13g2_decap_4 FILLER_64_652 ();
 sg13g2_fill_2 FILLER_64_721 ();
 sg13g2_fill_1 FILLER_64_723 ();
 sg13g2_decap_4 FILLER_64_734 ();
 sg13g2_fill_2 FILLER_64_738 ();
 sg13g2_decap_8 FILLER_64_808 ();
 sg13g2_decap_8 FILLER_64_915 ();
 sg13g2_decap_8 FILLER_64_922 ();
 sg13g2_decap_4 FILLER_64_929 ();
 sg13g2_decap_4 FILLER_64_979 ();
 sg13g2_fill_2 FILLER_64_1010 ();
 sg13g2_decap_8 FILLER_64_1025 ();
 sg13g2_decap_4 FILLER_64_1032 ();
 sg13g2_decap_4 FILLER_64_1049 ();
 sg13g2_fill_2 FILLER_64_1053 ();
 sg13g2_decap_4 FILLER_64_1093 ();
 sg13g2_fill_1 FILLER_64_1125 ();
 sg13g2_fill_2 FILLER_64_1148 ();
 sg13g2_decap_8 FILLER_64_1155 ();
 sg13g2_fill_1 FILLER_64_1162 ();
 sg13g2_decap_4 FILLER_64_1176 ();
 sg13g2_fill_1 FILLER_64_1180 ();
 sg13g2_decap_4 FILLER_64_1257 ();
 sg13g2_fill_1 FILLER_64_1261 ();
 sg13g2_fill_2 FILLER_64_1290 ();
 sg13g2_fill_2 FILLER_64_1301 ();
 sg13g2_decap_4 FILLER_64_1322 ();
 sg13g2_fill_1 FILLER_64_1326 ();
 sg13g2_fill_2 FILLER_64_1391 ();
 sg13g2_fill_1 FILLER_64_1393 ();
 sg13g2_decap_4 FILLER_64_1445 ();
 sg13g2_fill_2 FILLER_64_1449 ();
 sg13g2_fill_2 FILLER_64_1486 ();
 sg13g2_fill_1 FILLER_64_1488 ();
 sg13g2_fill_1 FILLER_64_1522 ();
 sg13g2_fill_1 FILLER_64_1532 ();
 sg13g2_fill_2 FILLER_64_1565 ();
 sg13g2_fill_1 FILLER_64_1567 ();
 sg13g2_decap_8 FILLER_64_1640 ();
 sg13g2_fill_1 FILLER_64_1647 ();
 sg13g2_fill_1 FILLER_64_1680 ();
 sg13g2_decap_8 FILLER_64_1708 ();
 sg13g2_fill_2 FILLER_64_1715 ();
 sg13g2_fill_1 FILLER_64_1717 ();
 sg13g2_fill_1 FILLER_64_1728 ();
 sg13g2_decap_4 FILLER_64_1760 ();
 sg13g2_decap_4 FILLER_64_1798 ();
 sg13g2_fill_1 FILLER_64_1802 ();
 sg13g2_decap_4 FILLER_64_1844 ();
 sg13g2_fill_1 FILLER_64_1912 ();
 sg13g2_fill_2 FILLER_64_1950 ();
 sg13g2_fill_1 FILLER_64_2019 ();
 sg13g2_decap_8 FILLER_64_2033 ();
 sg13g2_decap_8 FILLER_64_2114 ();
 sg13g2_fill_2 FILLER_64_2121 ();
 sg13g2_decap_4 FILLER_64_2132 ();
 sg13g2_fill_2 FILLER_64_2136 ();
 sg13g2_decap_8 FILLER_64_2147 ();
 sg13g2_decap_8 FILLER_64_2154 ();
 sg13g2_decap_4 FILLER_64_2161 ();
 sg13g2_fill_2 FILLER_64_2165 ();
 sg13g2_decap_4 FILLER_64_2198 ();
 sg13g2_fill_2 FILLER_64_2211 ();
 sg13g2_fill_1 FILLER_64_2213 ();
 sg13g2_decap_4 FILLER_64_2236 ();
 sg13g2_fill_2 FILLER_64_2295 ();
 sg13g2_fill_1 FILLER_64_2297 ();
 sg13g2_fill_2 FILLER_64_2344 ();
 sg13g2_fill_1 FILLER_64_2346 ();
 sg13g2_fill_2 FILLER_64_2370 ();
 sg13g2_fill_2 FILLER_64_2412 ();
 sg13g2_decap_8 FILLER_64_2436 ();
 sg13g2_fill_2 FILLER_64_2479 ();
 sg13g2_fill_1 FILLER_64_2481 ();
 sg13g2_decap_8 FILLER_64_2505 ();
 sg13g2_fill_1 FILLER_64_2512 ();
 sg13g2_fill_1 FILLER_64_2545 ();
 sg13g2_fill_2 FILLER_64_2559 ();
 sg13g2_fill_1 FILLER_64_2561 ();
 sg13g2_fill_1 FILLER_64_2595 ();
 sg13g2_fill_2 FILLER_64_2605 ();
 sg13g2_fill_1 FILLER_64_2607 ();
 sg13g2_decap_4 FILLER_64_2621 ();
 sg13g2_decap_4 FILLER_64_2794 ();
 sg13g2_fill_2 FILLER_64_2824 ();
 sg13g2_fill_1 FILLER_64_2826 ();
 sg13g2_decap_8 FILLER_64_2832 ();
 sg13g2_fill_1 FILLER_64_2839 ();
 sg13g2_decap_4 FILLER_64_2853 ();
 sg13g2_fill_2 FILLER_64_2857 ();
 sg13g2_decap_8 FILLER_64_2872 ();
 sg13g2_fill_2 FILLER_64_2906 ();
 sg13g2_fill_1 FILLER_64_2908 ();
 sg13g2_decap_4 FILLER_64_3013 ();
 sg13g2_fill_1 FILLER_64_3017 ();
 sg13g2_fill_2 FILLER_64_3031 ();
 sg13g2_fill_2 FILLER_64_3047 ();
 sg13g2_fill_1 FILLER_64_3049 ();
 sg13g2_decap_4 FILLER_64_3077 ();
 sg13g2_fill_1 FILLER_64_3081 ();
 sg13g2_decap_8 FILLER_64_3112 ();
 sg13g2_fill_2 FILLER_64_3119 ();
 sg13g2_fill_1 FILLER_64_3121 ();
 sg13g2_fill_1 FILLER_64_3158 ();
 sg13g2_fill_2 FILLER_64_3173 ();
 sg13g2_fill_1 FILLER_64_3175 ();
 sg13g2_fill_1 FILLER_64_3198 ();
 sg13g2_fill_2 FILLER_64_3221 ();
 sg13g2_fill_1 FILLER_64_3254 ();
 sg13g2_fill_2 FILLER_64_3269 ();
 sg13g2_fill_1 FILLER_64_3271 ();
 sg13g2_fill_1 FILLER_64_3321 ();
 sg13g2_decap_4 FILLER_64_3328 ();
 sg13g2_decap_8 FILLER_64_3337 ();
 sg13g2_fill_2 FILLER_64_3344 ();
 sg13g2_fill_1 FILLER_64_3346 ();
 sg13g2_fill_1 FILLER_64_3373 ();
 sg13g2_decap_4 FILLER_64_3393 ();
 sg13g2_fill_1 FILLER_64_3397 ();
 sg13g2_decap_4 FILLER_64_3432 ();
 sg13g2_fill_2 FILLER_64_3436 ();
 sg13g2_decap_8 FILLER_64_3466 ();
 sg13g2_decap_8 FILLER_64_3473 ();
 sg13g2_decap_8 FILLER_64_3480 ();
 sg13g2_decap_8 FILLER_64_3487 ();
 sg13g2_decap_8 FILLER_64_3494 ();
 sg13g2_decap_8 FILLER_64_3501 ();
 sg13g2_decap_8 FILLER_64_3508 ();
 sg13g2_decap_8 FILLER_64_3515 ();
 sg13g2_decap_8 FILLER_64_3522 ();
 sg13g2_decap_8 FILLER_64_3529 ();
 sg13g2_decap_8 FILLER_64_3536 ();
 sg13g2_decap_8 FILLER_64_3543 ();
 sg13g2_decap_8 FILLER_64_3550 ();
 sg13g2_decap_8 FILLER_64_3557 ();
 sg13g2_decap_8 FILLER_64_3564 ();
 sg13g2_decap_8 FILLER_64_3571 ();
 sg13g2_fill_2 FILLER_64_3578 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_48 ();
 sg13g2_fill_2 FILLER_65_61 ();
 sg13g2_fill_2 FILLER_65_71 ();
 sg13g2_fill_2 FILLER_65_104 ();
 sg13g2_fill_1 FILLER_65_106 ();
 sg13g2_fill_1 FILLER_65_147 ();
 sg13g2_fill_1 FILLER_65_224 ();
 sg13g2_fill_2 FILLER_65_251 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_fill_2 FILLER_65_298 ();
 sg13g2_fill_1 FILLER_65_300 ();
 sg13g2_fill_2 FILLER_65_319 ();
 sg13g2_fill_1 FILLER_65_321 ();
 sg13g2_fill_2 FILLER_65_348 ();
 sg13g2_fill_2 FILLER_65_363 ();
 sg13g2_fill_1 FILLER_65_365 ();
 sg13g2_fill_2 FILLER_65_392 ();
 sg13g2_fill_1 FILLER_65_394 ();
 sg13g2_decap_4 FILLER_65_438 ();
 sg13g2_decap_8 FILLER_65_459 ();
 sg13g2_decap_4 FILLER_65_466 ();
 sg13g2_fill_2 FILLER_65_498 ();
 sg13g2_fill_1 FILLER_65_514 ();
 sg13g2_decap_8 FILLER_65_530 ();
 sg13g2_decap_4 FILLER_65_537 ();
 sg13g2_fill_1 FILLER_65_541 ();
 sg13g2_fill_2 FILLER_65_549 ();
 sg13g2_fill_1 FILLER_65_551 ();
 sg13g2_decap_8 FILLER_65_561 ();
 sg13g2_decap_4 FILLER_65_568 ();
 sg13g2_fill_1 FILLER_65_572 ();
 sg13g2_fill_2 FILLER_65_590 ();
 sg13g2_fill_1 FILLER_65_592 ();
 sg13g2_decap_8 FILLER_65_628 ();
 sg13g2_decap_4 FILLER_65_635 ();
 sg13g2_fill_1 FILLER_65_639 ();
 sg13g2_fill_2 FILLER_65_653 ();
 sg13g2_fill_2 FILLER_65_674 ();
 sg13g2_decap_4 FILLER_65_685 ();
 sg13g2_fill_1 FILLER_65_729 ();
 sg13g2_fill_2 FILLER_65_766 ();
 sg13g2_fill_1 FILLER_65_780 ();
 sg13g2_fill_1 FILLER_65_790 ();
 sg13g2_fill_2 FILLER_65_800 ();
 sg13g2_fill_2 FILLER_65_847 ();
 sg13g2_fill_1 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_65_891 ();
 sg13g2_fill_1 FILLER_65_898 ();
 sg13g2_decap_4 FILLER_65_945 ();
 sg13g2_fill_1 FILLER_65_949 ();
 sg13g2_fill_2 FILLER_65_968 ();
 sg13g2_fill_1 FILLER_65_970 ();
 sg13g2_fill_2 FILLER_65_981 ();
 sg13g2_fill_1 FILLER_65_983 ();
 sg13g2_fill_2 FILLER_65_997 ();
 sg13g2_fill_1 FILLER_65_999 ();
 sg13g2_decap_4 FILLER_65_1041 ();
 sg13g2_fill_2 FILLER_65_1049 ();
 sg13g2_fill_2 FILLER_65_1075 ();
 sg13g2_fill_2 FILLER_65_1105 ();
 sg13g2_fill_1 FILLER_65_1134 ();
 sg13g2_fill_1 FILLER_65_1148 ();
 sg13g2_fill_2 FILLER_65_1162 ();
 sg13g2_fill_1 FILLER_65_1218 ();
 sg13g2_fill_2 FILLER_65_1223 ();
 sg13g2_fill_1 FILLER_65_1225 ();
 sg13g2_fill_1 FILLER_65_1230 ();
 sg13g2_fill_2 FILLER_65_1254 ();
 sg13g2_decap_4 FILLER_65_1271 ();
 sg13g2_fill_1 FILLER_65_1275 ();
 sg13g2_fill_2 FILLER_65_1298 ();
 sg13g2_fill_1 FILLER_65_1342 ();
 sg13g2_fill_2 FILLER_65_1367 ();
 sg13g2_fill_2 FILLER_65_1432 ();
 sg13g2_decap_8 FILLER_65_1485 ();
 sg13g2_decap_4 FILLER_65_1492 ();
 sg13g2_fill_2 FILLER_65_1496 ();
 sg13g2_fill_2 FILLER_65_1516 ();
 sg13g2_fill_1 FILLER_65_1518 ();
 sg13g2_fill_2 FILLER_65_1545 ();
 sg13g2_decap_4 FILLER_65_1597 ();
 sg13g2_fill_1 FILLER_65_1619 ();
 sg13g2_fill_1 FILLER_65_1629 ();
 sg13g2_decap_4 FILLER_65_1652 ();
 sg13g2_fill_1 FILLER_65_1656 ();
 sg13g2_fill_2 FILLER_65_1679 ();
 sg13g2_fill_1 FILLER_65_1681 ();
 sg13g2_fill_2 FILLER_65_1695 ();
 sg13g2_fill_1 FILLER_65_1697 ();
 sg13g2_fill_2 FILLER_65_1730 ();
 sg13g2_decap_4 FILLER_65_1736 ();
 sg13g2_decap_4 FILLER_65_1753 ();
 sg13g2_fill_2 FILLER_65_1757 ();
 sg13g2_fill_1 FILLER_65_1770 ();
 sg13g2_fill_2 FILLER_65_1779 ();
 sg13g2_fill_1 FILLER_65_1781 ();
 sg13g2_fill_2 FILLER_65_1788 ();
 sg13g2_decap_4 FILLER_65_1807 ();
 sg13g2_fill_1 FILLER_65_1811 ();
 sg13g2_decap_4 FILLER_65_1825 ();
 sg13g2_fill_1 FILLER_65_1829 ();
 sg13g2_fill_1 FILLER_65_1852 ();
 sg13g2_fill_2 FILLER_65_1857 ();
 sg13g2_fill_1 FILLER_65_1859 ();
 sg13g2_decap_8 FILLER_65_1873 ();
 sg13g2_decap_8 FILLER_65_1880 ();
 sg13g2_fill_2 FILLER_65_1887 ();
 sg13g2_fill_1 FILLER_65_1889 ();
 sg13g2_fill_2 FILLER_65_1917 ();
 sg13g2_fill_1 FILLER_65_1919 ();
 sg13g2_decap_4 FILLER_65_1947 ();
 sg13g2_fill_1 FILLER_65_1951 ();
 sg13g2_decap_8 FILLER_65_1965 ();
 sg13g2_fill_2 FILLER_65_1991 ();
 sg13g2_decap_4 FILLER_65_2002 ();
 sg13g2_fill_1 FILLER_65_2036 ();
 sg13g2_fill_1 FILLER_65_2075 ();
 sg13g2_decap_4 FILLER_65_2139 ();
 sg13g2_fill_1 FILLER_65_2143 ();
 sg13g2_decap_4 FILLER_65_2149 ();
 sg13g2_fill_2 FILLER_65_2153 ();
 sg13g2_fill_1 FILLER_65_2181 ();
 sg13g2_decap_4 FILLER_65_2195 ();
 sg13g2_fill_1 FILLER_65_2225 ();
 sg13g2_decap_8 FILLER_65_2245 ();
 sg13g2_fill_2 FILLER_65_2274 ();
 sg13g2_decap_4 FILLER_65_2322 ();
 sg13g2_fill_2 FILLER_65_2326 ();
 sg13g2_fill_2 FILLER_65_2331 ();
 sg13g2_decap_4 FILLER_65_2338 ();
 sg13g2_fill_2 FILLER_65_2347 ();
 sg13g2_fill_1 FILLER_65_2362 ();
 sg13g2_decap_8 FILLER_65_2402 ();
 sg13g2_fill_1 FILLER_65_2409 ();
 sg13g2_fill_2 FILLER_65_2443 ();
 sg13g2_fill_1 FILLER_65_2445 ();
 sg13g2_fill_2 FILLER_65_2459 ();
 sg13g2_fill_1 FILLER_65_2470 ();
 sg13g2_fill_1 FILLER_65_2481 ();
 sg13g2_decap_4 FILLER_65_2500 ();
 sg13g2_fill_2 FILLER_65_2504 ();
 sg13g2_fill_1 FILLER_65_2563 ();
 sg13g2_fill_1 FILLER_65_2609 ();
 sg13g2_fill_2 FILLER_65_2615 ();
 sg13g2_fill_1 FILLER_65_2627 ();
 sg13g2_fill_2 FILLER_65_2656 ();
 sg13g2_decap_4 FILLER_65_2695 ();
 sg13g2_fill_1 FILLER_65_2717 ();
 sg13g2_decap_4 FILLER_65_2731 ();
 sg13g2_decap_4 FILLER_65_2758 ();
 sg13g2_fill_1 FILLER_65_2771 ();
 sg13g2_fill_2 FILLER_65_2798 ();
 sg13g2_fill_1 FILLER_65_2800 ();
 sg13g2_fill_1 FILLER_65_2879 ();
 sg13g2_fill_2 FILLER_65_2898 ();
 sg13g2_decap_8 FILLER_65_2919 ();
 sg13g2_fill_2 FILLER_65_2949 ();
 sg13g2_fill_2 FILLER_65_2964 ();
 sg13g2_fill_1 FILLER_65_2966 ();
 sg13g2_fill_2 FILLER_65_2998 ();
 sg13g2_fill_1 FILLER_65_3000 ();
 sg13g2_fill_1 FILLER_65_3066 ();
 sg13g2_fill_1 FILLER_65_3094 ();
 sg13g2_fill_2 FILLER_65_3119 ();
 sg13g2_fill_2 FILLER_65_3134 ();
 sg13g2_fill_1 FILLER_65_3136 ();
 sg13g2_decap_8 FILLER_65_3168 ();
 sg13g2_decap_4 FILLER_65_3188 ();
 sg13g2_fill_1 FILLER_65_3192 ();
 sg13g2_fill_2 FILLER_65_3220 ();
 sg13g2_fill_1 FILLER_65_3222 ();
 sg13g2_decap_8 FILLER_65_3251 ();
 sg13g2_fill_1 FILLER_65_3258 ();
 sg13g2_fill_2 FILLER_65_3303 ();
 sg13g2_fill_1 FILLER_65_3311 ();
 sg13g2_fill_1 FILLER_65_3321 ();
 sg13g2_fill_1 FILLER_65_3334 ();
 sg13g2_decap_8 FILLER_65_3349 ();
 sg13g2_decap_4 FILLER_65_3356 ();
 sg13g2_fill_2 FILLER_65_3360 ();
 sg13g2_decap_8 FILLER_65_3380 ();
 sg13g2_fill_2 FILLER_65_3387 ();
 sg13g2_fill_2 FILLER_65_3404 ();
 sg13g2_decap_8 FILLER_65_3430 ();
 sg13g2_decap_4 FILLER_65_3437 ();
 sg13g2_fill_1 FILLER_65_3441 ();
 sg13g2_decap_8 FILLER_65_3468 ();
 sg13g2_decap_8 FILLER_65_3475 ();
 sg13g2_decap_8 FILLER_65_3482 ();
 sg13g2_decap_8 FILLER_65_3489 ();
 sg13g2_decap_8 FILLER_65_3496 ();
 sg13g2_decap_8 FILLER_65_3503 ();
 sg13g2_decap_8 FILLER_65_3510 ();
 sg13g2_decap_8 FILLER_65_3517 ();
 sg13g2_decap_8 FILLER_65_3524 ();
 sg13g2_decap_8 FILLER_65_3531 ();
 sg13g2_decap_8 FILLER_65_3538 ();
 sg13g2_decap_8 FILLER_65_3545 ();
 sg13g2_decap_8 FILLER_65_3552 ();
 sg13g2_decap_8 FILLER_65_3559 ();
 sg13g2_decap_8 FILLER_65_3566 ();
 sg13g2_decap_8 FILLER_65_3573 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_20 ();
 sg13g2_fill_2 FILLER_66_36 ();
 sg13g2_fill_2 FILLER_66_41 ();
 sg13g2_decap_4 FILLER_66_48 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_fill_2 FILLER_66_77 ();
 sg13g2_fill_1 FILLER_66_162 ();
 sg13g2_decap_4 FILLER_66_190 ();
 sg13g2_fill_2 FILLER_66_194 ();
 sg13g2_fill_2 FILLER_66_261 ();
 sg13g2_decap_4 FILLER_66_283 ();
 sg13g2_fill_1 FILLER_66_306 ();
 sg13g2_fill_2 FILLER_66_332 ();
 sg13g2_fill_1 FILLER_66_342 ();
 sg13g2_fill_1 FILLER_66_394 ();
 sg13g2_fill_2 FILLER_66_424 ();
 sg13g2_fill_2 FILLER_66_480 ();
 sg13g2_decap_4 FILLER_66_503 ();
 sg13g2_fill_1 FILLER_66_507 ();
 sg13g2_decap_8 FILLER_66_535 ();
 sg13g2_fill_2 FILLER_66_542 ();
 sg13g2_decap_8 FILLER_66_560 ();
 sg13g2_decap_4 FILLER_66_595 ();
 sg13g2_fill_2 FILLER_66_603 ();
 sg13g2_fill_1 FILLER_66_651 ();
 sg13g2_fill_1 FILLER_66_712 ();
 sg13g2_fill_2 FILLER_66_801 ();
 sg13g2_fill_2 FILLER_66_831 ();
 sg13g2_fill_2 FILLER_66_846 ();
 sg13g2_fill_1 FILLER_66_848 ();
 sg13g2_decap_4 FILLER_66_867 ();
 sg13g2_fill_2 FILLER_66_871 ();
 sg13g2_fill_2 FILLER_66_878 ();
 sg13g2_fill_1 FILLER_66_880 ();
 sg13g2_fill_2 FILLER_66_887 ();
 sg13g2_decap_8 FILLER_66_894 ();
 sg13g2_fill_1 FILLER_66_901 ();
 sg13g2_decap_8 FILLER_66_906 ();
 sg13g2_decap_8 FILLER_66_913 ();
 sg13g2_fill_2 FILLER_66_920 ();
 sg13g2_decap_4 FILLER_66_926 ();
 sg13g2_fill_1 FILLER_66_935 ();
 sg13g2_decap_8 FILLER_66_953 ();
 sg13g2_decap_8 FILLER_66_960 ();
 sg13g2_fill_2 FILLER_66_967 ();
 sg13g2_fill_1 FILLER_66_969 ();
 sg13g2_fill_2 FILLER_66_1009 ();
 sg13g2_fill_1 FILLER_66_1030 ();
 sg13g2_decap_4 FILLER_66_1088 ();
 sg13g2_fill_2 FILLER_66_1092 ();
 sg13g2_fill_2 FILLER_66_1148 ();
 sg13g2_fill_2 FILLER_66_1176 ();
 sg13g2_fill_1 FILLER_66_1178 ();
 sg13g2_decap_8 FILLER_66_1204 ();
 sg13g2_fill_2 FILLER_66_1211 ();
 sg13g2_decap_4 FILLER_66_1227 ();
 sg13g2_fill_1 FILLER_66_1231 ();
 sg13g2_fill_2 FILLER_66_1259 ();
 sg13g2_fill_1 FILLER_66_1293 ();
 sg13g2_fill_2 FILLER_66_1300 ();
 sg13g2_fill_1 FILLER_66_1336 ();
 sg13g2_fill_1 FILLER_66_1341 ();
 sg13g2_fill_1 FILLER_66_1377 ();
 sg13g2_fill_2 FILLER_66_1410 ();
 sg13g2_decap_4 FILLER_66_1421 ();
 sg13g2_decap_4 FILLER_66_1457 ();
 sg13g2_fill_1 FILLER_66_1461 ();
 sg13g2_fill_2 FILLER_66_1515 ();
 sg13g2_decap_4 FILLER_66_1556 ();
 sg13g2_fill_2 FILLER_66_1574 ();
 sg13g2_decap_4 FILLER_66_1652 ();
 sg13g2_fill_2 FILLER_66_1669 ();
 sg13g2_fill_1 FILLER_66_1671 ();
 sg13g2_decap_4 FILLER_66_1678 ();
 sg13g2_fill_2 FILLER_66_1682 ();
 sg13g2_decap_4 FILLER_66_1755 ();
 sg13g2_fill_2 FILLER_66_1765 ();
 sg13g2_fill_1 FILLER_66_1773 ();
 sg13g2_decap_4 FILLER_66_1815 ();
 sg13g2_fill_1 FILLER_66_1819 ();
 sg13g2_decap_4 FILLER_66_1825 ();
 sg13g2_fill_1 FILLER_66_1844 ();
 sg13g2_decap_8 FILLER_66_1882 ();
 sg13g2_decap_8 FILLER_66_1889 ();
 sg13g2_fill_1 FILLER_66_1896 ();
 sg13g2_fill_2 FILLER_66_1952 ();
 sg13g2_fill_1 FILLER_66_1954 ();
 sg13g2_decap_8 FILLER_66_1968 ();
 sg13g2_fill_1 FILLER_66_1975 ();
 sg13g2_fill_1 FILLER_66_1998 ();
 sg13g2_fill_2 FILLER_66_2002 ();
 sg13g2_fill_2 FILLER_66_2020 ();
 sg13g2_fill_1 FILLER_66_2060 ();
 sg13g2_fill_2 FILLER_66_2105 ();
 sg13g2_fill_2 FILLER_66_2132 ();
 sg13g2_decap_8 FILLER_66_2149 ();
 sg13g2_decap_8 FILLER_66_2156 ();
 sg13g2_decap_4 FILLER_66_2163 ();
 sg13g2_fill_1 FILLER_66_2167 ();
 sg13g2_fill_1 FILLER_66_2186 ();
 sg13g2_fill_2 FILLER_66_2223 ();
 sg13g2_fill_2 FILLER_66_2235 ();
 sg13g2_decap_4 FILLER_66_2247 ();
 sg13g2_fill_2 FILLER_66_2251 ();
 sg13g2_fill_1 FILLER_66_2270 ();
 sg13g2_fill_2 FILLER_66_2277 ();
 sg13g2_fill_2 FILLER_66_2288 ();
 sg13g2_fill_1 FILLER_66_2321 ();
 sg13g2_fill_2 FILLER_66_2356 ();
 sg13g2_fill_1 FILLER_66_2376 ();
 sg13g2_fill_2 FILLER_66_2411 ();
 sg13g2_fill_1 FILLER_66_2413 ();
 sg13g2_decap_8 FILLER_66_2433 ();
 sg13g2_decap_4 FILLER_66_2440 ();
 sg13g2_fill_2 FILLER_66_2444 ();
 sg13g2_decap_8 FILLER_66_2481 ();
 sg13g2_fill_2 FILLER_66_2488 ();
 sg13g2_fill_2 FILLER_66_2495 ();
 sg13g2_fill_1 FILLER_66_2497 ();
 sg13g2_fill_2 FILLER_66_2520 ();
 sg13g2_fill_1 FILLER_66_2522 ();
 sg13g2_fill_2 FILLER_66_2549 ();
 sg13g2_fill_1 FILLER_66_2551 ();
 sg13g2_fill_1 FILLER_66_2586 ();
 sg13g2_decap_8 FILLER_66_2615 ();
 sg13g2_decap_8 FILLER_66_2645 ();
 sg13g2_fill_2 FILLER_66_2652 ();
 sg13g2_fill_1 FILLER_66_2663 ();
 sg13g2_fill_2 FILLER_66_2668 ();
 sg13g2_fill_1 FILLER_66_2670 ();
 sg13g2_fill_2 FILLER_66_2675 ();
 sg13g2_fill_1 FILLER_66_2677 ();
 sg13g2_decap_8 FILLER_66_2687 ();
 sg13g2_decap_4 FILLER_66_2694 ();
 sg13g2_fill_1 FILLER_66_2698 ();
 sg13g2_decap_4 FILLER_66_2704 ();
 sg13g2_fill_1 FILLER_66_2708 ();
 sg13g2_fill_1 FILLER_66_2743 ();
 sg13g2_fill_2 FILLER_66_2772 ();
 sg13g2_decap_4 FILLER_66_2824 ();
 sg13g2_fill_1 FILLER_66_2828 ();
 sg13g2_fill_2 FILLER_66_2842 ();
 sg13g2_fill_1 FILLER_66_2844 ();
 sg13g2_fill_1 FILLER_66_2873 ();
 sg13g2_decap_8 FILLER_66_2877 ();
 sg13g2_decap_8 FILLER_66_2911 ();
 sg13g2_fill_2 FILLER_66_2918 ();
 sg13g2_fill_1 FILLER_66_2920 ();
 sg13g2_fill_1 FILLER_66_2949 ();
 sg13g2_fill_2 FILLER_66_2978 ();
 sg13g2_fill_1 FILLER_66_2993 ();
 sg13g2_fill_1 FILLER_66_3017 ();
 sg13g2_decap_8 FILLER_66_3046 ();
 sg13g2_decap_8 FILLER_66_3057 ();
 sg13g2_decap_8 FILLER_66_3064 ();
 sg13g2_decap_4 FILLER_66_3071 ();
 sg13g2_decap_4 FILLER_66_3146 ();
 sg13g2_fill_1 FILLER_66_3186 ();
 sg13g2_fill_1 FILLER_66_3200 ();
 sg13g2_fill_2 FILLER_66_3232 ();
 sg13g2_fill_1 FILLER_66_3240 ();
 sg13g2_decap_4 FILLER_66_3268 ();
 sg13g2_fill_2 FILLER_66_3276 ();
 sg13g2_fill_1 FILLER_66_3278 ();
 sg13g2_fill_2 FILLER_66_3320 ();
 sg13g2_fill_1 FILLER_66_3322 ();
 sg13g2_decap_8 FILLER_66_3352 ();
 sg13g2_decap_4 FILLER_66_3359 ();
 sg13g2_fill_2 FILLER_66_3384 ();
 sg13g2_fill_2 FILLER_66_3399 ();
 sg13g2_fill_1 FILLER_66_3401 ();
 sg13g2_fill_2 FILLER_66_3407 ();
 sg13g2_fill_1 FILLER_66_3409 ();
 sg13g2_fill_1 FILLER_66_3433 ();
 sg13g2_decap_8 FILLER_66_3461 ();
 sg13g2_decap_8 FILLER_66_3468 ();
 sg13g2_decap_8 FILLER_66_3475 ();
 sg13g2_decap_8 FILLER_66_3482 ();
 sg13g2_decap_8 FILLER_66_3489 ();
 sg13g2_decap_8 FILLER_66_3496 ();
 sg13g2_decap_8 FILLER_66_3503 ();
 sg13g2_decap_8 FILLER_66_3510 ();
 sg13g2_decap_8 FILLER_66_3517 ();
 sg13g2_decap_8 FILLER_66_3524 ();
 sg13g2_decap_8 FILLER_66_3531 ();
 sg13g2_decap_8 FILLER_66_3538 ();
 sg13g2_decap_8 FILLER_66_3545 ();
 sg13g2_decap_8 FILLER_66_3552 ();
 sg13g2_decap_8 FILLER_66_3559 ();
 sg13g2_decap_8 FILLER_66_3566 ();
 sg13g2_decap_8 FILLER_66_3573 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_4 FILLER_67_35 ();
 sg13g2_fill_2 FILLER_67_39 ();
 sg13g2_decap_8 FILLER_67_68 ();
 sg13g2_decap_8 FILLER_67_75 ();
 sg13g2_decap_8 FILLER_67_82 ();
 sg13g2_decap_8 FILLER_67_89 ();
 sg13g2_decap_4 FILLER_67_96 ();
 sg13g2_fill_1 FILLER_67_113 ();
 sg13g2_fill_2 FILLER_67_136 ();
 sg13g2_fill_2 FILLER_67_165 ();
 sg13g2_fill_1 FILLER_67_167 ();
 sg13g2_fill_2 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_242 ();
 sg13g2_fill_2 FILLER_67_264 ();
 sg13g2_fill_1 FILLER_67_280 ();
 sg13g2_fill_2 FILLER_67_298 ();
 sg13g2_fill_1 FILLER_67_300 ();
 sg13g2_fill_2 FILLER_67_358 ();
 sg13g2_fill_1 FILLER_67_360 ();
 sg13g2_fill_2 FILLER_67_374 ();
 sg13g2_fill_1 FILLER_67_376 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_67_435 ();
 sg13g2_fill_2 FILLER_67_455 ();
 sg13g2_fill_1 FILLER_67_457 ();
 sg13g2_fill_1 FILLER_67_464 ();
 sg13g2_fill_1 FILLER_67_494 ();
 sg13g2_decap_8 FILLER_67_500 ();
 sg13g2_decap_8 FILLER_67_507 ();
 sg13g2_fill_1 FILLER_67_514 ();
 sg13g2_fill_2 FILLER_67_520 ();
 sg13g2_fill_2 FILLER_67_526 ();
 sg13g2_fill_1 FILLER_67_528 ();
 sg13g2_fill_2 FILLER_67_533 ();
 sg13g2_fill_1 FILLER_67_535 ();
 sg13g2_decap_8 FILLER_67_556 ();
 sg13g2_fill_2 FILLER_67_563 ();
 sg13g2_decap_8 FILLER_67_587 ();
 sg13g2_fill_2 FILLER_67_594 ();
 sg13g2_fill_1 FILLER_67_596 ();
 sg13g2_decap_4 FILLER_67_614 ();
 sg13g2_fill_1 FILLER_67_618 ();
 sg13g2_decap_4 FILLER_67_632 ();
 sg13g2_fill_1 FILLER_67_645 ();
 sg13g2_decap_8 FILLER_67_674 ();
 sg13g2_decap_8 FILLER_67_681 ();
 sg13g2_decap_4 FILLER_67_688 ();
 sg13g2_fill_2 FILLER_67_692 ();
 sg13g2_fill_1 FILLER_67_726 ();
 sg13g2_fill_2 FILLER_67_795 ();
 sg13g2_fill_2 FILLER_67_812 ();
 sg13g2_fill_2 FILLER_67_832 ();
 sg13g2_fill_2 FILLER_67_925 ();
 sg13g2_decap_8 FILLER_67_992 ();
 sg13g2_fill_2 FILLER_67_999 ();
 sg13g2_fill_1 FILLER_67_1001 ();
 sg13g2_decap_8 FILLER_67_1052 ();
 sg13g2_fill_2 FILLER_67_1059 ();
 sg13g2_fill_1 FILLER_67_1061 ();
 sg13g2_fill_2 FILLER_67_1070 ();
 sg13g2_fill_1 FILLER_67_1072 ();
 sg13g2_fill_1 FILLER_67_1083 ();
 sg13g2_fill_2 FILLER_67_1111 ();
 sg13g2_fill_2 FILLER_67_1154 ();
 sg13g2_decap_4 FILLER_67_1184 ();
 sg13g2_fill_1 FILLER_67_1188 ();
 sg13g2_fill_1 FILLER_67_1216 ();
 sg13g2_fill_1 FILLER_67_1225 ();
 sg13g2_fill_2 FILLER_67_1276 ();
 sg13g2_fill_1 FILLER_67_1278 ();
 sg13g2_fill_2 FILLER_67_1296 ();
 sg13g2_fill_1 FILLER_67_1298 ();
 sg13g2_fill_2 FILLER_67_1307 ();
 sg13g2_fill_2 FILLER_67_1315 ();
 sg13g2_fill_2 FILLER_67_1344 ();
 sg13g2_fill_1 FILLER_67_1346 ();
 sg13g2_fill_1 FILLER_67_1362 ();
 sg13g2_decap_8 FILLER_67_1392 ();
 sg13g2_fill_1 FILLER_67_1399 ();
 sg13g2_fill_1 FILLER_67_1475 ();
 sg13g2_fill_2 FILLER_67_1491 ();
 sg13g2_fill_2 FILLER_67_1531 ();
 sg13g2_fill_2 FILLER_67_1598 ();
 sg13g2_decap_8 FILLER_67_1658 ();
 sg13g2_fill_2 FILLER_67_1665 ();
 sg13g2_fill_2 FILLER_67_1695 ();
 sg13g2_fill_1 FILLER_67_1716 ();
 sg13g2_decap_8 FILLER_67_1733 ();
 sg13g2_fill_2 FILLER_67_1740 ();
 sg13g2_fill_1 FILLER_67_1742 ();
 sg13g2_decap_4 FILLER_67_1780 ();
 sg13g2_decap_4 FILLER_67_1787 ();
 sg13g2_fill_1 FILLER_67_1791 ();
 sg13g2_decap_8 FILLER_67_1797 ();
 sg13g2_decap_4 FILLER_67_1804 ();
 sg13g2_fill_2 FILLER_67_1822 ();
 sg13g2_fill_1 FILLER_67_1824 ();
 sg13g2_fill_2 FILLER_67_1853 ();
 sg13g2_fill_1 FILLER_67_1855 ();
 sg13g2_decap_4 FILLER_67_1865 ();
 sg13g2_fill_2 FILLER_67_1913 ();
 sg13g2_fill_1 FILLER_67_1915 ();
 sg13g2_fill_1 FILLER_67_1921 ();
 sg13g2_decap_4 FILLER_67_1927 ();
 sg13g2_fill_1 FILLER_67_1957 ();
 sg13g2_fill_1 FILLER_67_2014 ();
 sg13g2_fill_1 FILLER_67_2052 ();
 sg13g2_fill_2 FILLER_67_2074 ();
 sg13g2_fill_1 FILLER_67_2076 ();
 sg13g2_fill_2 FILLER_67_2172 ();
 sg13g2_decap_4 FILLER_67_2202 ();
 sg13g2_fill_2 FILLER_67_2232 ();
 sg13g2_fill_1 FILLER_67_2234 ();
 sg13g2_fill_1 FILLER_67_2281 ();
 sg13g2_fill_2 FILLER_67_2304 ();
 sg13g2_fill_1 FILLER_67_2328 ();
 sg13g2_decap_8 FILLER_67_2351 ();
 sg13g2_decap_8 FILLER_67_2358 ();
 sg13g2_fill_2 FILLER_67_2371 ();
 sg13g2_fill_1 FILLER_67_2373 ();
 sg13g2_fill_2 FILLER_67_2401 ();
 sg13g2_fill_1 FILLER_67_2416 ();
 sg13g2_decap_4 FILLER_67_2448 ();
 sg13g2_fill_1 FILLER_67_2452 ();
 sg13g2_fill_2 FILLER_67_2459 ();
 sg13g2_fill_2 FILLER_67_2503 ();
 sg13g2_fill_1 FILLER_67_2505 ();
 sg13g2_fill_2 FILLER_67_2510 ();
 sg13g2_fill_1 FILLER_67_2512 ();
 sg13g2_fill_2 FILLER_67_2592 ();
 sg13g2_fill_2 FILLER_67_2609 ();
 sg13g2_fill_1 FILLER_67_2611 ();
 sg13g2_decap_4 FILLER_67_2625 ();
 sg13g2_fill_2 FILLER_67_2629 ();
 sg13g2_fill_2 FILLER_67_2734 ();
 sg13g2_fill_2 FILLER_67_2745 ();
 sg13g2_fill_2 FILLER_67_2756 ();
 sg13g2_fill_2 FILLER_67_2807 ();
 sg13g2_fill_1 FILLER_67_2809 ();
 sg13g2_fill_1 FILLER_67_2834 ();
 sg13g2_fill_2 FILLER_67_2839 ();
 sg13g2_fill_1 FILLER_67_2841 ();
 sg13g2_fill_1 FILLER_67_2864 ();
 sg13g2_fill_1 FILLER_67_2869 ();
 sg13g2_fill_2 FILLER_67_2893 ();
 sg13g2_fill_1 FILLER_67_2895 ();
 sg13g2_fill_2 FILLER_67_2924 ();
 sg13g2_fill_1 FILLER_67_2953 ();
 sg13g2_fill_2 FILLER_67_2976 ();
 sg13g2_fill_1 FILLER_67_2978 ();
 sg13g2_fill_1 FILLER_67_3007 ();
 sg13g2_fill_1 FILLER_67_3024 ();
 sg13g2_fill_1 FILLER_67_3076 ();
 sg13g2_fill_2 FILLER_67_3096 ();
 sg13g2_decap_4 FILLER_67_3141 ();
 sg13g2_fill_2 FILLER_67_3167 ();
 sg13g2_fill_1 FILLER_67_3169 ();
 sg13g2_decap_4 FILLER_67_3183 ();
 sg13g2_fill_2 FILLER_67_3187 ();
 sg13g2_fill_2 FILLER_67_3212 ();
 sg13g2_fill_1 FILLER_67_3254 ();
 sg13g2_decap_8 FILLER_67_3272 ();
 sg13g2_decap_4 FILLER_67_3279 ();
 sg13g2_fill_1 FILLER_67_3283 ();
 sg13g2_decap_4 FILLER_67_3288 ();
 sg13g2_fill_2 FILLER_67_3292 ();
 sg13g2_fill_1 FILLER_67_3306 ();
 sg13g2_decap_8 FILLER_67_3326 ();
 sg13g2_decap_8 FILLER_67_3347 ();
 sg13g2_decap_8 FILLER_67_3354 ();
 sg13g2_fill_2 FILLER_67_3361 ();
 sg13g2_decap_4 FILLER_67_3372 ();
 sg13g2_fill_2 FILLER_67_3376 ();
 sg13g2_decap_8 FILLER_67_3404 ();
 sg13g2_decap_8 FILLER_67_3416 ();
 sg13g2_fill_1 FILLER_67_3423 ();
 sg13g2_decap_8 FILLER_67_3428 ();
 sg13g2_decap_4 FILLER_67_3435 ();
 sg13g2_decap_8 FILLER_67_3443 ();
 sg13g2_decap_8 FILLER_67_3450 ();
 sg13g2_decap_8 FILLER_67_3457 ();
 sg13g2_decap_8 FILLER_67_3464 ();
 sg13g2_decap_8 FILLER_67_3471 ();
 sg13g2_decap_8 FILLER_67_3478 ();
 sg13g2_decap_8 FILLER_67_3485 ();
 sg13g2_decap_8 FILLER_67_3492 ();
 sg13g2_decap_8 FILLER_67_3499 ();
 sg13g2_decap_8 FILLER_67_3506 ();
 sg13g2_decap_8 FILLER_67_3513 ();
 sg13g2_decap_8 FILLER_67_3520 ();
 sg13g2_decap_8 FILLER_67_3527 ();
 sg13g2_decap_8 FILLER_67_3534 ();
 sg13g2_decap_8 FILLER_67_3541 ();
 sg13g2_decap_8 FILLER_67_3548 ();
 sg13g2_decap_8 FILLER_67_3555 ();
 sg13g2_decap_8 FILLER_67_3562 ();
 sg13g2_decap_8 FILLER_67_3569 ();
 sg13g2_decap_4 FILLER_67_3576 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_4 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_50 ();
 sg13g2_decap_8 FILLER_68_57 ();
 sg13g2_decap_8 FILLER_68_64 ();
 sg13g2_decap_8 FILLER_68_71 ();
 sg13g2_decap_8 FILLER_68_78 ();
 sg13g2_decap_8 FILLER_68_85 ();
 sg13g2_decap_8 FILLER_68_92 ();
 sg13g2_decap_4 FILLER_68_99 ();
 sg13g2_fill_2 FILLER_68_103 ();
 sg13g2_fill_2 FILLER_68_147 ();
 sg13g2_fill_2 FILLER_68_162 ();
 sg13g2_fill_2 FILLER_68_183 ();
 sg13g2_fill_1 FILLER_68_185 ();
 sg13g2_fill_2 FILLER_68_200 ();
 sg13g2_fill_2 FILLER_68_229 ();
 sg13g2_fill_1 FILLER_68_231 ();
 sg13g2_fill_2 FILLER_68_247 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_fill_1 FILLER_68_268 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_1 FILLER_68_316 ();
 sg13g2_fill_2 FILLER_68_365 ();
 sg13g2_fill_1 FILLER_68_367 ();
 sg13g2_fill_2 FILLER_68_408 ();
 sg13g2_fill_2 FILLER_68_419 ();
 sg13g2_fill_1 FILLER_68_430 ();
 sg13g2_fill_2 FILLER_68_437 ();
 sg13g2_fill_2 FILLER_68_445 ();
 sg13g2_decap_4 FILLER_68_494 ();
 sg13g2_fill_2 FILLER_68_498 ();
 sg13g2_fill_2 FILLER_68_512 ();
 sg13g2_fill_1 FILLER_68_514 ();
 sg13g2_fill_1 FILLER_68_521 ();
 sg13g2_fill_2 FILLER_68_543 ();
 sg13g2_fill_1 FILLER_68_545 ();
 sg13g2_fill_2 FILLER_68_551 ();
 sg13g2_decap_8 FILLER_68_563 ();
 sg13g2_fill_2 FILLER_68_570 ();
 sg13g2_fill_1 FILLER_68_572 ();
 sg13g2_fill_2 FILLER_68_578 ();
 sg13g2_fill_2 FILLER_68_634 ();
 sg13g2_fill_2 FILLER_68_646 ();
 sg13g2_fill_2 FILLER_68_658 ();
 sg13g2_fill_1 FILLER_68_669 ();
 sg13g2_fill_2 FILLER_68_698 ();
 sg13g2_fill_1 FILLER_68_700 ();
 sg13g2_fill_1 FILLER_68_706 ();
 sg13g2_fill_1 FILLER_68_786 ();
 sg13g2_fill_1 FILLER_68_810 ();
 sg13g2_decap_4 FILLER_68_839 ();
 sg13g2_fill_2 FILLER_68_856 ();
 sg13g2_fill_1 FILLER_68_858 ();
 sg13g2_fill_1 FILLER_68_865 ();
 sg13g2_decap_8 FILLER_68_870 ();
 sg13g2_decap_4 FILLER_68_877 ();
 sg13g2_fill_2 FILLER_68_881 ();
 sg13g2_fill_1 FILLER_68_905 ();
 sg13g2_fill_2 FILLER_68_915 ();
 sg13g2_fill_1 FILLER_68_917 ();
 sg13g2_fill_1 FILLER_68_931 ();
 sg13g2_fill_1 FILLER_68_941 ();
 sg13g2_decap_8 FILLER_68_958 ();
 sg13g2_fill_1 FILLER_68_971 ();
 sg13g2_decap_4 FILLER_68_1019 ();
 sg13g2_fill_2 FILLER_68_1039 ();
 sg13g2_fill_1 FILLER_68_1041 ();
 sg13g2_decap_8 FILLER_68_1050 ();
 sg13g2_fill_1 FILLER_68_1057 ();
 sg13g2_decap_4 FILLER_68_1078 ();
 sg13g2_fill_2 FILLER_68_1082 ();
 sg13g2_fill_2 FILLER_68_1105 ();
 sg13g2_fill_2 FILLER_68_1133 ();
 sg13g2_fill_1 FILLER_68_1135 ();
 sg13g2_fill_1 FILLER_68_1155 ();
 sg13g2_fill_2 FILLER_68_1184 ();
 sg13g2_fill_2 FILLER_68_1190 ();
 sg13g2_fill_1 FILLER_68_1192 ();
 sg13g2_decap_4 FILLER_68_1208 ();
 sg13g2_decap_8 FILLER_68_1220 ();
 sg13g2_decap_4 FILLER_68_1227 ();
 sg13g2_fill_1 FILLER_68_1231 ();
 sg13g2_fill_2 FILLER_68_1243 ();
 sg13g2_fill_1 FILLER_68_1245 ();
 sg13g2_decap_8 FILLER_68_1254 ();
 sg13g2_decap_4 FILLER_68_1261 ();
 sg13g2_fill_2 FILLER_68_1286 ();
 sg13g2_fill_1 FILLER_68_1288 ();
 sg13g2_decap_4 FILLER_68_1299 ();
 sg13g2_fill_1 FILLER_68_1303 ();
 sg13g2_fill_2 FILLER_68_1315 ();
 sg13g2_fill_1 FILLER_68_1317 ();
 sg13g2_fill_1 FILLER_68_1331 ();
 sg13g2_fill_2 FILLER_68_1349 ();
 sg13g2_fill_1 FILLER_68_1385 ();
 sg13g2_decap_4 FILLER_68_1398 ();
 sg13g2_fill_2 FILLER_68_1402 ();
 sg13g2_fill_2 FILLER_68_1416 ();
 sg13g2_fill_1 FILLER_68_1418 ();
 sg13g2_fill_1 FILLER_68_1446 ();
 sg13g2_fill_2 FILLER_68_1455 ();
 sg13g2_fill_1 FILLER_68_1457 ();
 sg13g2_fill_1 FILLER_68_1495 ();
 sg13g2_fill_2 FILLER_68_1506 ();
 sg13g2_fill_2 FILLER_68_1512 ();
 sg13g2_fill_2 FILLER_68_1536 ();
 sg13g2_fill_2 FILLER_68_1551 ();
 sg13g2_fill_1 FILLER_68_1572 ();
 sg13g2_decap_8 FILLER_68_1625 ();
 sg13g2_fill_2 FILLER_68_1636 ();
 sg13g2_fill_2 FILLER_68_1644 ();
 sg13g2_fill_2 FILLER_68_1681 ();
 sg13g2_fill_2 FILLER_68_1696 ();
 sg13g2_fill_1 FILLER_68_1715 ();
 sg13g2_fill_2 FILLER_68_1725 ();
 sg13g2_fill_1 FILLER_68_1727 ();
 sg13g2_fill_1 FILLER_68_1731 ();
 sg13g2_fill_2 FILLER_68_1736 ();
 sg13g2_fill_1 FILLER_68_1751 ();
 sg13g2_fill_1 FILLER_68_1770 ();
 sg13g2_fill_1 FILLER_68_1780 ();
 sg13g2_fill_2 FILLER_68_1819 ();
 sg13g2_decap_4 FILLER_68_1834 ();
 sg13g2_fill_1 FILLER_68_1858 ();
 sg13g2_decap_4 FILLER_68_1880 ();
 sg13g2_decap_4 FILLER_68_1925 ();
 sg13g2_fill_2 FILLER_68_1929 ();
 sg13g2_fill_1 FILLER_68_1945 ();
 sg13g2_decap_4 FILLER_68_1959 ();
 sg13g2_decap_4 FILLER_68_1967 ();
 sg13g2_fill_1 FILLER_68_1971 ();
 sg13g2_fill_1 FILLER_68_1991 ();
 sg13g2_fill_1 FILLER_68_2001 ();
 sg13g2_decap_4 FILLER_68_2092 ();
 sg13g2_fill_1 FILLER_68_2096 ();
 sg13g2_fill_1 FILLER_68_2119 ();
 sg13g2_decap_8 FILLER_68_2152 ();
 sg13g2_decap_4 FILLER_68_2159 ();
 sg13g2_fill_1 FILLER_68_2188 ();
 sg13g2_decap_4 FILLER_68_2192 ();
 sg13g2_fill_2 FILLER_68_2223 ();
 sg13g2_fill_1 FILLER_68_2225 ();
 sg13g2_decap_4 FILLER_68_2232 ();
 sg13g2_fill_2 FILLER_68_2248 ();
 sg13g2_fill_1 FILLER_68_2250 ();
 sg13g2_fill_2 FILLER_68_2389 ();
 sg13g2_fill_1 FILLER_68_2416 ();
 sg13g2_fill_2 FILLER_68_2428 ();
 sg13g2_fill_1 FILLER_68_2456 ();
 sg13g2_decap_4 FILLER_68_2486 ();
 sg13g2_fill_2 FILLER_68_2490 ();
 sg13g2_fill_2 FILLER_68_2526 ();
 sg13g2_fill_1 FILLER_68_2576 ();
 sg13g2_fill_2 FILLER_68_2609 ();
 sg13g2_fill_1 FILLER_68_2611 ();
 sg13g2_fill_2 FILLER_68_2633 ();
 sg13g2_fill_1 FILLER_68_2648 ();
 sg13g2_fill_1 FILLER_68_2671 ();
 sg13g2_decap_8 FILLER_68_2683 ();
 sg13g2_decap_8 FILLER_68_2690 ();
 sg13g2_decap_4 FILLER_68_2701 ();
 sg13g2_fill_1 FILLER_68_2705 ();
 sg13g2_fill_2 FILLER_68_2736 ();
 sg13g2_fill_1 FILLER_68_2746 ();
 sg13g2_fill_2 FILLER_68_2796 ();
 sg13g2_fill_2 FILLER_68_2826 ();
 sg13g2_fill_1 FILLER_68_2828 ();
 sg13g2_fill_1 FILLER_68_2857 ();
 sg13g2_fill_1 FILLER_68_2868 ();
 sg13g2_decap_8 FILLER_68_2915 ();
 sg13g2_fill_2 FILLER_68_2922 ();
 sg13g2_decap_8 FILLER_68_2961 ();
 sg13g2_fill_2 FILLER_68_2968 ();
 sg13g2_decap_8 FILLER_68_2983 ();
 sg13g2_decap_4 FILLER_68_2990 ();
 sg13g2_fill_2 FILLER_68_2994 ();
 sg13g2_decap_8 FILLER_68_3048 ();
 sg13g2_fill_2 FILLER_68_3055 ();
 sg13g2_decap_4 FILLER_68_3066 ();
 sg13g2_fill_2 FILLER_68_3070 ();
 sg13g2_fill_1 FILLER_68_3145 ();
 sg13g2_fill_2 FILLER_68_3188 ();
 sg13g2_fill_1 FILLER_68_3190 ();
 sg13g2_fill_2 FILLER_68_3252 ();
 sg13g2_fill_2 FILLER_68_3266 ();
 sg13g2_decap_8 FILLER_68_3281 ();
 sg13g2_fill_2 FILLER_68_3316 ();
 sg13g2_fill_2 FILLER_68_3340 ();
 sg13g2_decap_8 FILLER_68_3380 ();
 sg13g2_fill_1 FILLER_68_3387 ();
 sg13g2_fill_1 FILLER_68_3393 ();
 sg13g2_decap_8 FILLER_68_3412 ();
 sg13g2_fill_2 FILLER_68_3447 ();
 sg13g2_decap_8 FILLER_68_3453 ();
 sg13g2_decap_8 FILLER_68_3460 ();
 sg13g2_decap_8 FILLER_68_3467 ();
 sg13g2_decap_8 FILLER_68_3474 ();
 sg13g2_decap_8 FILLER_68_3481 ();
 sg13g2_decap_8 FILLER_68_3488 ();
 sg13g2_decap_8 FILLER_68_3495 ();
 sg13g2_decap_8 FILLER_68_3502 ();
 sg13g2_decap_8 FILLER_68_3509 ();
 sg13g2_decap_8 FILLER_68_3516 ();
 sg13g2_decap_8 FILLER_68_3523 ();
 sg13g2_decap_8 FILLER_68_3530 ();
 sg13g2_decap_8 FILLER_68_3537 ();
 sg13g2_decap_8 FILLER_68_3544 ();
 sg13g2_decap_8 FILLER_68_3551 ();
 sg13g2_decap_8 FILLER_68_3558 ();
 sg13g2_decap_8 FILLER_68_3565 ();
 sg13g2_decap_8 FILLER_68_3572 ();
 sg13g2_fill_1 FILLER_68_3579 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_4 FILLER_69_112 ();
 sg13g2_fill_2 FILLER_69_120 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_fill_1 FILLER_69_147 ();
 sg13g2_fill_2 FILLER_69_184 ();
 sg13g2_fill_1 FILLER_69_186 ();
 sg13g2_fill_2 FILLER_69_259 ();
 sg13g2_fill_1 FILLER_69_261 ();
 sg13g2_fill_2 FILLER_69_290 ();
 sg13g2_fill_2 FILLER_69_323 ();
 sg13g2_fill_1 FILLER_69_347 ();
 sg13g2_decap_8 FILLER_69_376 ();
 sg13g2_fill_1 FILLER_69_392 ();
 sg13g2_decap_4 FILLER_69_436 ();
 sg13g2_fill_1 FILLER_69_440 ();
 sg13g2_decap_4 FILLER_69_453 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_fill_2 FILLER_69_462 ();
 sg13g2_fill_1 FILLER_69_464 ();
 sg13g2_decap_8 FILLER_69_470 ();
 sg13g2_fill_1 FILLER_69_477 ();
 sg13g2_fill_1 FILLER_69_490 ();
 sg13g2_fill_1 FILLER_69_496 ();
 sg13g2_fill_2 FILLER_69_509 ();
 sg13g2_fill_1 FILLER_69_511 ();
 sg13g2_fill_1 FILLER_69_522 ();
 sg13g2_decap_8 FILLER_69_531 ();
 sg13g2_fill_1 FILLER_69_577 ();
 sg13g2_decap_4 FILLER_69_582 ();
 sg13g2_fill_2 FILLER_69_598 ();
 sg13g2_fill_1 FILLER_69_606 ();
 sg13g2_fill_2 FILLER_69_620 ();
 sg13g2_fill_1 FILLER_69_622 ();
 sg13g2_fill_2 FILLER_69_627 ();
 sg13g2_fill_1 FILLER_69_629 ();
 sg13g2_fill_2 FILLER_69_643 ();
 sg13g2_decap_4 FILLER_69_659 ();
 sg13g2_decap_4 FILLER_69_683 ();
 sg13g2_fill_2 FILLER_69_701 ();
 sg13g2_fill_2 FILLER_69_742 ();
 sg13g2_fill_1 FILLER_69_756 ();
 sg13g2_fill_2 FILLER_69_768 ();
 sg13g2_fill_1 FILLER_69_770 ();
 sg13g2_fill_2 FILLER_69_784 ();
 sg13g2_fill_2 FILLER_69_815 ();
 sg13g2_fill_2 FILLER_69_821 ();
 sg13g2_decap_4 FILLER_69_832 ();
 sg13g2_fill_1 FILLER_69_836 ();
 sg13g2_decap_4 FILLER_69_850 ();
 sg13g2_fill_2 FILLER_69_854 ();
 sg13g2_decap_4 FILLER_69_870 ();
 sg13g2_fill_1 FILLER_69_897 ();
 sg13g2_fill_2 FILLER_69_917 ();
 sg13g2_fill_1 FILLER_69_919 ();
 sg13g2_fill_2 FILLER_69_933 ();
 sg13g2_decap_8 FILLER_69_953 ();
 sg13g2_fill_1 FILLER_69_960 ();
 sg13g2_fill_1 FILLER_69_981 ();
 sg13g2_decap_8 FILLER_69_1004 ();
 sg13g2_fill_2 FILLER_69_1011 ();
 sg13g2_decap_8 FILLER_69_1023 ();
 sg13g2_decap_8 FILLER_69_1030 ();
 sg13g2_fill_1 FILLER_69_1037 ();
 sg13g2_fill_2 FILLER_69_1043 ();
 sg13g2_fill_1 FILLER_69_1053 ();
 sg13g2_decap_4 FILLER_69_1085 ();
 sg13g2_fill_2 FILLER_69_1089 ();
 sg13g2_decap_8 FILLER_69_1106 ();
 sg13g2_decap_4 FILLER_69_1113 ();
 sg13g2_fill_2 FILLER_69_1127 ();
 sg13g2_fill_1 FILLER_69_1129 ();
 sg13g2_fill_2 FILLER_69_1147 ();
 sg13g2_fill_2 FILLER_69_1180 ();
 sg13g2_fill_1 FILLER_69_1182 ();
 sg13g2_fill_2 FILLER_69_1200 ();
 sg13g2_fill_1 FILLER_69_1219 ();
 sg13g2_fill_2 FILLER_69_1248 ();
 sg13g2_fill_1 FILLER_69_1258 ();
 sg13g2_decap_8 FILLER_69_1307 ();
 sg13g2_fill_2 FILLER_69_1314 ();
 sg13g2_fill_2 FILLER_69_1334 ();
 sg13g2_fill_2 FILLER_69_1373 ();
 sg13g2_fill_1 FILLER_69_1375 ();
 sg13g2_fill_2 FILLER_69_1397 ();
 sg13g2_fill_1 FILLER_69_1409 ();
 sg13g2_decap_4 FILLER_69_1414 ();
 sg13g2_fill_1 FILLER_69_1446 ();
 sg13g2_fill_1 FILLER_69_1456 ();
 sg13g2_fill_1 FILLER_69_1486 ();
 sg13g2_fill_2 FILLER_69_1506 ();
 sg13g2_fill_1 FILLER_69_1564 ();
 sg13g2_fill_2 FILLER_69_1580 ();
 sg13g2_fill_2 FILLER_69_1594 ();
 sg13g2_fill_1 FILLER_69_1596 ();
 sg13g2_fill_2 FILLER_69_1610 ();
 sg13g2_fill_1 FILLER_69_1612 ();
 sg13g2_fill_1 FILLER_69_1619 ();
 sg13g2_decap_8 FILLER_69_1624 ();
 sg13g2_fill_1 FILLER_69_1631 ();
 sg13g2_decap_4 FILLER_69_1638 ();
 sg13g2_fill_2 FILLER_69_1642 ();
 sg13g2_fill_1 FILLER_69_1686 ();
 sg13g2_decap_4 FILLER_69_1715 ();
 sg13g2_fill_2 FILLER_69_1719 ();
 sg13g2_fill_2 FILLER_69_1759 ();
 sg13g2_fill_1 FILLER_69_1761 ();
 sg13g2_fill_1 FILLER_69_1776 ();
 sg13g2_decap_4 FILLER_69_1785 ();
 sg13g2_fill_2 FILLER_69_1789 ();
 sg13g2_decap_8 FILLER_69_1796 ();
 sg13g2_decap_8 FILLER_69_1808 ();
 sg13g2_decap_4 FILLER_69_1815 ();
 sg13g2_decap_4 FILLER_69_1824 ();
 sg13g2_fill_1 FILLER_69_1828 ();
 sg13g2_decap_8 FILLER_69_1837 ();
 sg13g2_fill_2 FILLER_69_1852 ();
 sg13g2_fill_2 FILLER_69_1865 ();
 sg13g2_fill_1 FILLER_69_1867 ();
 sg13g2_decap_4 FILLER_69_1896 ();
 sg13g2_fill_2 FILLER_69_1900 ();
 sg13g2_fill_1 FILLER_69_1909 ();
 sg13g2_fill_1 FILLER_69_2017 ();
 sg13g2_fill_2 FILLER_69_2130 ();
 sg13g2_fill_1 FILLER_69_2132 ();
 sg13g2_decap_8 FILLER_69_2169 ();
 sg13g2_fill_2 FILLER_69_2176 ();
 sg13g2_decap_8 FILLER_69_2211 ();
 sg13g2_fill_1 FILLER_69_2218 ();
 sg13g2_fill_1 FILLER_69_2274 ();
 sg13g2_fill_2 FILLER_69_2320 ();
 sg13g2_fill_1 FILLER_69_2322 ();
 sg13g2_fill_1 FILLER_69_2334 ();
 sg13g2_decap_8 FILLER_69_2339 ();
 sg13g2_decap_8 FILLER_69_2346 ();
 sg13g2_decap_4 FILLER_69_2353 ();
 sg13g2_fill_1 FILLER_69_2357 ();
 sg13g2_fill_2 FILLER_69_2377 ();
 sg13g2_fill_1 FILLER_69_2379 ();
 sg13g2_fill_2 FILLER_69_2393 ();
 sg13g2_fill_2 FILLER_69_2411 ();
 sg13g2_fill_2 FILLER_69_2435 ();
 sg13g2_fill_2 FILLER_69_2451 ();
 sg13g2_fill_1 FILLER_69_2474 ();
 sg13g2_fill_2 FILLER_69_2488 ();
 sg13g2_fill_2 FILLER_69_2506 ();
 sg13g2_fill_1 FILLER_69_2517 ();
 sg13g2_decap_4 FILLER_69_2544 ();
 sg13g2_fill_1 FILLER_69_2548 ();
 sg13g2_fill_1 FILLER_69_2576 ();
 sg13g2_fill_1 FILLER_69_2611 ();
 sg13g2_fill_1 FILLER_69_2632 ();
 sg13g2_fill_2 FILLER_69_2670 ();
 sg13g2_fill_2 FILLER_69_2679 ();
 sg13g2_decap_8 FILLER_69_2691 ();
 sg13g2_fill_2 FILLER_69_2733 ();
 sg13g2_fill_1 FILLER_69_2735 ();
 sg13g2_fill_1 FILLER_69_2759 ();
 sg13g2_fill_1 FILLER_69_2765 ();
 sg13g2_decap_4 FILLER_69_2799 ();
 sg13g2_decap_8 FILLER_69_2807 ();
 sg13g2_fill_2 FILLER_69_2818 ();
 sg13g2_fill_1 FILLER_69_2820 ();
 sg13g2_decap_8 FILLER_69_2838 ();
 sg13g2_fill_1 FILLER_69_2845 ();
 sg13g2_decap_8 FILLER_69_2877 ();
 sg13g2_fill_2 FILLER_69_2884 ();
 sg13g2_fill_1 FILLER_69_2886 ();
 sg13g2_decap_4 FILLER_69_2890 ();
 sg13g2_decap_8 FILLER_69_2900 ();
 sg13g2_fill_1 FILLER_69_2913 ();
 sg13g2_decap_4 FILLER_69_2920 ();
 sg13g2_fill_1 FILLER_69_2949 ();
 sg13g2_fill_2 FILLER_69_2969 ();
 sg13g2_fill_2 FILLER_69_3016 ();
 sg13g2_fill_1 FILLER_69_3018 ();
 sg13g2_decap_4 FILLER_69_3029 ();
 sg13g2_fill_1 FILLER_69_3033 ();
 sg13g2_decap_4 FILLER_69_3039 ();
 sg13g2_fill_1 FILLER_69_3043 ();
 sg13g2_fill_2 FILLER_69_3056 ();
 sg13g2_fill_1 FILLER_69_3058 ();
 sg13g2_decap_4 FILLER_69_3065 ();
 sg13g2_decap_8 FILLER_69_3080 ();
 sg13g2_fill_2 FILLER_69_3087 ();
 sg13g2_fill_2 FILLER_69_3099 ();
 sg13g2_fill_2 FILLER_69_3105 ();
 sg13g2_fill_2 FILLER_69_3114 ();
 sg13g2_fill_1 FILLER_69_3159 ();
 sg13g2_decap_4 FILLER_69_3166 ();
 sg13g2_fill_1 FILLER_69_3179 ();
 sg13g2_fill_2 FILLER_69_3199 ();
 sg13g2_decap_8 FILLER_69_3214 ();
 sg13g2_fill_1 FILLER_69_3227 ();
 sg13g2_fill_1 FILLER_69_3254 ();
 sg13g2_fill_1 FILLER_69_3268 ();
 sg13g2_fill_2 FILLER_69_3275 ();
 sg13g2_fill_1 FILLER_69_3277 ();
 sg13g2_fill_2 FILLER_69_3291 ();
 sg13g2_decap_8 FILLER_69_3297 ();
 sg13g2_decap_8 FILLER_69_3304 ();
 sg13g2_fill_2 FILLER_69_3311 ();
 sg13g2_fill_1 FILLER_69_3313 ();
 sg13g2_decap_4 FILLER_69_3323 ();
 sg13g2_fill_1 FILLER_69_3327 ();
 sg13g2_fill_2 FILLER_69_3350 ();
 sg13g2_fill_1 FILLER_69_3371 ();
 sg13g2_fill_2 FILLER_69_3403 ();
 sg13g2_fill_2 FILLER_69_3425 ();
 sg13g2_fill_1 FILLER_69_3427 ();
 sg13g2_decap_8 FILLER_69_3471 ();
 sg13g2_decap_8 FILLER_69_3478 ();
 sg13g2_decap_8 FILLER_69_3485 ();
 sg13g2_decap_8 FILLER_69_3492 ();
 sg13g2_decap_8 FILLER_69_3499 ();
 sg13g2_decap_8 FILLER_69_3506 ();
 sg13g2_decap_8 FILLER_69_3513 ();
 sg13g2_decap_8 FILLER_69_3520 ();
 sg13g2_decap_8 FILLER_69_3527 ();
 sg13g2_decap_8 FILLER_69_3534 ();
 sg13g2_decap_8 FILLER_69_3541 ();
 sg13g2_decap_8 FILLER_69_3548 ();
 sg13g2_decap_8 FILLER_69_3555 ();
 sg13g2_decap_8 FILLER_69_3562 ();
 sg13g2_decap_8 FILLER_69_3569 ();
 sg13g2_decap_4 FILLER_69_3576 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_fill_2 FILLER_70_140 ();
 sg13g2_fill_2 FILLER_70_169 ();
 sg13g2_fill_1 FILLER_70_171 ();
 sg13g2_fill_2 FILLER_70_201 ();
 sg13g2_fill_1 FILLER_70_203 ();
 sg13g2_fill_1 FILLER_70_231 ();
 sg13g2_fill_2 FILLER_70_241 ();
 sg13g2_fill_2 FILLER_70_320 ();
 sg13g2_fill_1 FILLER_70_322 ();
 sg13g2_fill_2 FILLER_70_336 ();
 sg13g2_fill_1 FILLER_70_351 ();
 sg13g2_fill_1 FILLER_70_356 ();
 sg13g2_decap_4 FILLER_70_371 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_fill_1 FILLER_70_420 ();
 sg13g2_fill_2 FILLER_70_425 ();
 sg13g2_fill_1 FILLER_70_440 ();
 sg13g2_decap_8 FILLER_70_453 ();
 sg13g2_fill_1 FILLER_70_514 ();
 sg13g2_decap_4 FILLER_70_530 ();
 sg13g2_fill_2 FILLER_70_534 ();
 sg13g2_fill_2 FILLER_70_549 ();
 sg13g2_decap_8 FILLER_70_564 ();
 sg13g2_fill_2 FILLER_70_571 ();
 sg13g2_decap_4 FILLER_70_621 ();
 sg13g2_fill_2 FILLER_70_625 ();
 sg13g2_decap_4 FILLER_70_653 ();
 sg13g2_decap_4 FILLER_70_662 ();
 sg13g2_fill_2 FILLER_70_671 ();
 sg13g2_fill_1 FILLER_70_673 ();
 sg13g2_fill_1 FILLER_70_678 ();
 sg13g2_decap_8 FILLER_70_682 ();
 sg13g2_fill_1 FILLER_70_689 ();
 sg13g2_decap_8 FILLER_70_712 ();
 sg13g2_decap_8 FILLER_70_719 ();
 sg13g2_fill_2 FILLER_70_769 ();
 sg13g2_decap_8 FILLER_70_774 ();
 sg13g2_fill_2 FILLER_70_787 ();
 sg13g2_fill_1 FILLER_70_803 ();
 sg13g2_fill_2 FILLER_70_819 ();
 sg13g2_fill_1 FILLER_70_829 ();
 sg13g2_fill_2 FILLER_70_869 ();
 sg13g2_fill_1 FILLER_70_871 ();
 sg13g2_fill_2 FILLER_70_886 ();
 sg13g2_fill_1 FILLER_70_908 ();
 sg13g2_fill_1 FILLER_70_921 ();
 sg13g2_fill_2 FILLER_70_927 ();
 sg13g2_fill_1 FILLER_70_929 ();
 sg13g2_fill_2 FILLER_70_935 ();
 sg13g2_fill_1 FILLER_70_948 ();
 sg13g2_fill_1 FILLER_70_967 ();
 sg13g2_fill_1 FILLER_70_997 ();
 sg13g2_decap_4 FILLER_70_1010 ();
 sg13g2_fill_1 FILLER_70_1014 ();
 sg13g2_decap_4 FILLER_70_1043 ();
 sg13g2_fill_1 FILLER_70_1059 ();
 sg13g2_fill_2 FILLER_70_1065 ();
 sg13g2_fill_1 FILLER_70_1067 ();
 sg13g2_decap_4 FILLER_70_1082 ();
 sg13g2_fill_1 FILLER_70_1086 ();
 sg13g2_fill_2 FILLER_70_1093 ();
 sg13g2_fill_1 FILLER_70_1095 ();
 sg13g2_decap_8 FILLER_70_1112 ();
 sg13g2_fill_2 FILLER_70_1119 ();
 sg13g2_fill_1 FILLER_70_1121 ();
 sg13g2_fill_2 FILLER_70_1134 ();
 sg13g2_fill_1 FILLER_70_1136 ();
 sg13g2_fill_2 FILLER_70_1156 ();
 sg13g2_fill_2 FILLER_70_1174 ();
 sg13g2_fill_1 FILLER_70_1198 ();
 sg13g2_fill_1 FILLER_70_1204 ();
 sg13g2_decap_8 FILLER_70_1219 ();
 sg13g2_fill_2 FILLER_70_1226 ();
 sg13g2_fill_1 FILLER_70_1228 ();
 sg13g2_fill_1 FILLER_70_1252 ();
 sg13g2_decap_4 FILLER_70_1258 ();
 sg13g2_fill_1 FILLER_70_1262 ();
 sg13g2_decap_8 FILLER_70_1279 ();
 sg13g2_decap_8 FILLER_70_1310 ();
 sg13g2_fill_2 FILLER_70_1317 ();
 sg13g2_fill_1 FILLER_70_1319 ();
 sg13g2_fill_1 FILLER_70_1341 ();
 sg13g2_fill_1 FILLER_70_1363 ();
 sg13g2_fill_1 FILLER_70_1382 ();
 sg13g2_decap_8 FILLER_70_1387 ();
 sg13g2_decap_4 FILLER_70_1394 ();
 sg13g2_fill_1 FILLER_70_1398 ();
 sg13g2_decap_4 FILLER_70_1404 ();
 sg13g2_fill_1 FILLER_70_1408 ();
 sg13g2_fill_2 FILLER_70_1430 ();
 sg13g2_fill_1 FILLER_70_1432 ();
 sg13g2_decap_8 FILLER_70_1443 ();
 sg13g2_decap_8 FILLER_70_1450 ();
 sg13g2_decap_4 FILLER_70_1457 ();
 sg13g2_decap_8 FILLER_70_1474 ();
 sg13g2_fill_2 FILLER_70_1481 ();
 sg13g2_fill_1 FILLER_70_1483 ();
 sg13g2_fill_1 FILLER_70_1501 ();
 sg13g2_decap_8 FILLER_70_1521 ();
 sg13g2_decap_8 FILLER_70_1528 ();
 sg13g2_fill_2 FILLER_70_1535 ();
 sg13g2_fill_2 FILLER_70_1570 ();
 sg13g2_fill_1 FILLER_70_1576 ();
 sg13g2_fill_2 FILLER_70_1592 ();
 sg13g2_decap_8 FILLER_70_1599 ();
 sg13g2_fill_2 FILLER_70_1606 ();
 sg13g2_fill_1 FILLER_70_1608 ();
 sg13g2_fill_2 FILLER_70_1643 ();
 sg13g2_decap_8 FILLER_70_1665 ();
 sg13g2_decap_4 FILLER_70_1680 ();
 sg13g2_fill_2 FILLER_70_1684 ();
 sg13g2_fill_2 FILLER_70_1710 ();
 sg13g2_decap_8 FILLER_70_1747 ();
 sg13g2_fill_1 FILLER_70_1754 ();
 sg13g2_fill_1 FILLER_70_1773 ();
 sg13g2_fill_2 FILLER_70_1784 ();
 sg13g2_decap_4 FILLER_70_1791 ();
 sg13g2_fill_1 FILLER_70_1795 ();
 sg13g2_fill_1 FILLER_70_1843 ();
 sg13g2_fill_2 FILLER_70_1850 ();
 sg13g2_fill_1 FILLER_70_1852 ();
 sg13g2_decap_8 FILLER_70_1856 ();
 sg13g2_fill_1 FILLER_70_1863 ();
 sg13g2_fill_2 FILLER_70_1868 ();
 sg13g2_decap_8 FILLER_70_1883 ();
 sg13g2_fill_1 FILLER_70_1890 ();
 sg13g2_fill_2 FILLER_70_1895 ();
 sg13g2_fill_2 FILLER_70_1912 ();
 sg13g2_fill_1 FILLER_70_1914 ();
 sg13g2_fill_2 FILLER_70_1928 ();
 sg13g2_fill_1 FILLER_70_1930 ();
 sg13g2_decap_8 FILLER_70_1940 ();
 sg13g2_fill_1 FILLER_70_1947 ();
 sg13g2_decap_8 FILLER_70_1958 ();
 sg13g2_decap_8 FILLER_70_1965 ();
 sg13g2_fill_2 FILLER_70_1972 ();
 sg13g2_fill_1 FILLER_70_1974 ();
 sg13g2_fill_2 FILLER_70_2027 ();
 sg13g2_fill_1 FILLER_70_2034 ();
 sg13g2_fill_2 FILLER_70_2040 ();
 sg13g2_fill_1 FILLER_70_2042 ();
 sg13g2_fill_1 FILLER_70_2065 ();
 sg13g2_decap_4 FILLER_70_2081 ();
 sg13g2_fill_1 FILLER_70_2085 ();
 sg13g2_fill_1 FILLER_70_2110 ();
 sg13g2_fill_2 FILLER_70_2142 ();
 sg13g2_fill_1 FILLER_70_2153 ();
 sg13g2_fill_2 FILLER_70_2162 ();
 sg13g2_fill_1 FILLER_70_2164 ();
 sg13g2_fill_2 FILLER_70_2173 ();
 sg13g2_fill_2 FILLER_70_2180 ();
 sg13g2_fill_1 FILLER_70_2182 ();
 sg13g2_decap_4 FILLER_70_2213 ();
 sg13g2_fill_1 FILLER_70_2217 ();
 sg13g2_fill_1 FILLER_70_2231 ();
 sg13g2_decap_8 FILLER_70_2238 ();
 sg13g2_decap_4 FILLER_70_2245 ();
 sg13g2_fill_2 FILLER_70_2249 ();
 sg13g2_fill_2 FILLER_70_2260 ();
 sg13g2_fill_2 FILLER_70_2275 ();
 sg13g2_fill_2 FILLER_70_2285 ();
 sg13g2_fill_2 FILLER_70_2313 ();
 sg13g2_fill_2 FILLER_70_2319 ();
 sg13g2_fill_1 FILLER_70_2321 ();
 sg13g2_fill_2 FILLER_70_2340 ();
 sg13g2_fill_2 FILLER_70_2383 ();
 sg13g2_fill_1 FILLER_70_2385 ();
 sg13g2_fill_1 FILLER_70_2391 ();
 sg13g2_fill_1 FILLER_70_2402 ();
 sg13g2_fill_1 FILLER_70_2407 ();
 sg13g2_fill_1 FILLER_70_2442 ();
 sg13g2_fill_2 FILLER_70_2465 ();
 sg13g2_decap_8 FILLER_70_2472 ();
 sg13g2_decap_4 FILLER_70_2479 ();
 sg13g2_fill_2 FILLER_70_2483 ();
 sg13g2_decap_4 FILLER_70_2492 ();
 sg13g2_fill_2 FILLER_70_2496 ();
 sg13g2_fill_1 FILLER_70_2507 ();
 sg13g2_decap_4 FILLER_70_2548 ();
 sg13g2_fill_2 FILLER_70_2552 ();
 sg13g2_fill_1 FILLER_70_2572 ();
 sg13g2_fill_2 FILLER_70_2593 ();
 sg13g2_decap_8 FILLER_70_2605 ();
 sg13g2_decap_8 FILLER_70_2612 ();
 sg13g2_fill_2 FILLER_70_2619 ();
 sg13g2_decap_8 FILLER_70_2626 ();
 sg13g2_fill_2 FILLER_70_2633 ();
 sg13g2_fill_1 FILLER_70_2635 ();
 sg13g2_decap_8 FILLER_70_2658 ();
 sg13g2_decap_4 FILLER_70_2665 ();
 sg13g2_fill_1 FILLER_70_2669 ();
 sg13g2_decap_8 FILLER_70_2688 ();
 sg13g2_fill_2 FILLER_70_2695 ();
 sg13g2_fill_1 FILLER_70_2706 ();
 sg13g2_decap_8 FILLER_70_2713 ();
 sg13g2_decap_8 FILLER_70_2724 ();
 sg13g2_fill_2 FILLER_70_2731 ();
 sg13g2_fill_1 FILLER_70_2733 ();
 sg13g2_decap_8 FILLER_70_2751 ();
 sg13g2_decap_4 FILLER_70_2773 ();
 sg13g2_fill_2 FILLER_70_2789 ();
 sg13g2_decap_8 FILLER_70_2802 ();
 sg13g2_fill_1 FILLER_70_2809 ();
 sg13g2_decap_4 FILLER_70_2838 ();
 sg13g2_fill_2 FILLER_70_2842 ();
 sg13g2_fill_2 FILLER_70_2849 ();
 sg13g2_fill_1 FILLER_70_2851 ();
 sg13g2_fill_2 FILLER_70_2870 ();
 sg13g2_fill_1 FILLER_70_2872 ();
 sg13g2_fill_1 FILLER_70_2882 ();
 sg13g2_fill_2 FILLER_70_2888 ();
 sg13g2_fill_1 FILLER_70_2890 ();
 sg13g2_decap_8 FILLER_70_2920 ();
 sg13g2_fill_2 FILLER_70_2927 ();
 sg13g2_fill_1 FILLER_70_2929 ();
 sg13g2_decap_4 FILLER_70_2963 ();
 sg13g2_decap_4 FILLER_70_2991 ();
 sg13g2_fill_1 FILLER_70_2995 ();
 sg13g2_fill_1 FILLER_70_3002 ();
 sg13g2_fill_2 FILLER_70_3008 ();
 sg13g2_fill_2 FILLER_70_3024 ();
 sg13g2_decap_8 FILLER_70_3056 ();
 sg13g2_decap_8 FILLER_70_3084 ();
 sg13g2_fill_1 FILLER_70_3091 ();
 sg13g2_fill_2 FILLER_70_3110 ();
 sg13g2_fill_1 FILLER_70_3112 ();
 sg13g2_decap_8 FILLER_70_3140 ();
 sg13g2_fill_1 FILLER_70_3147 ();
 sg13g2_fill_2 FILLER_70_3173 ();
 sg13g2_fill_1 FILLER_70_3175 ();
 sg13g2_fill_1 FILLER_70_3239 ();
 sg13g2_fill_2 FILLER_70_3244 ();
 sg13g2_fill_1 FILLER_70_3275 ();
 sg13g2_fill_2 FILLER_70_3284 ();
 sg13g2_fill_1 FILLER_70_3286 ();
 sg13g2_fill_1 FILLER_70_3315 ();
 sg13g2_decap_8 FILLER_70_3325 ();
 sg13g2_fill_1 FILLER_70_3332 ();
 sg13g2_decap_4 FILLER_70_3355 ();
 sg13g2_fill_2 FILLER_70_3359 ();
 sg13g2_decap_8 FILLER_70_3379 ();
 sg13g2_decap_4 FILLER_70_3386 ();
 sg13g2_fill_1 FILLER_70_3390 ();
 sg13g2_fill_1 FILLER_70_3405 ();
 sg13g2_fill_1 FILLER_70_3410 ();
 sg13g2_fill_2 FILLER_70_3416 ();
 sg13g2_fill_2 FILLER_70_3423 ();
 sg13g2_fill_1 FILLER_70_3425 ();
 sg13g2_decap_8 FILLER_70_3472 ();
 sg13g2_decap_8 FILLER_70_3479 ();
 sg13g2_decap_8 FILLER_70_3486 ();
 sg13g2_decap_8 FILLER_70_3493 ();
 sg13g2_decap_8 FILLER_70_3500 ();
 sg13g2_decap_8 FILLER_70_3507 ();
 sg13g2_decap_8 FILLER_70_3514 ();
 sg13g2_decap_8 FILLER_70_3521 ();
 sg13g2_decap_8 FILLER_70_3528 ();
 sg13g2_decap_8 FILLER_70_3535 ();
 sg13g2_decap_8 FILLER_70_3542 ();
 sg13g2_decap_8 FILLER_70_3549 ();
 sg13g2_decap_8 FILLER_70_3556 ();
 sg13g2_decap_8 FILLER_70_3563 ();
 sg13g2_decap_8 FILLER_70_3570 ();
 sg13g2_fill_2 FILLER_70_3577 ();
 sg13g2_fill_1 FILLER_70_3579 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_4 FILLER_71_147 ();
 sg13g2_fill_2 FILLER_71_151 ();
 sg13g2_fill_2 FILLER_71_207 ();
 sg13g2_fill_2 FILLER_71_254 ();
 sg13g2_fill_2 FILLER_71_303 ();
 sg13g2_fill_1 FILLER_71_342 ();
 sg13g2_fill_2 FILLER_71_397 ();
 sg13g2_fill_2 FILLER_71_414 ();
 sg13g2_decap_4 FILLER_71_429 ();
 sg13g2_fill_2 FILLER_71_433 ();
 sg13g2_decap_8 FILLER_71_448 ();
 sg13g2_decap_4 FILLER_71_455 ();
 sg13g2_fill_1 FILLER_71_459 ();
 sg13g2_decap_8 FILLER_71_469 ();
 sg13g2_decap_8 FILLER_71_476 ();
 sg13g2_fill_2 FILLER_71_483 ();
 sg13g2_decap_8 FILLER_71_503 ();
 sg13g2_decap_4 FILLER_71_510 ();
 sg13g2_decap_8 FILLER_71_529 ();
 sg13g2_fill_1 FILLER_71_536 ();
 sg13g2_decap_8 FILLER_71_556 ();
 sg13g2_fill_2 FILLER_71_563 ();
 sg13g2_fill_2 FILLER_71_573 ();
 sg13g2_fill_1 FILLER_71_575 ();
 sg13g2_decap_8 FILLER_71_587 ();
 sg13g2_decap_4 FILLER_71_594 ();
 sg13g2_fill_1 FILLER_71_598 ();
 sg13g2_fill_2 FILLER_71_629 ();
 sg13g2_fill_1 FILLER_71_642 ();
 sg13g2_fill_2 FILLER_71_670 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_decap_8 FILLER_71_697 ();
 sg13g2_fill_1 FILLER_71_704 ();
 sg13g2_decap_4 FILLER_71_711 ();
 sg13g2_fill_2 FILLER_71_715 ();
 sg13g2_fill_2 FILLER_71_737 ();
 sg13g2_fill_2 FILLER_71_748 ();
 sg13g2_decap_8 FILLER_71_768 ();
 sg13g2_decap_4 FILLER_71_775 ();
 sg13g2_fill_2 FILLER_71_779 ();
 sg13g2_decap_8 FILLER_71_789 ();
 sg13g2_fill_2 FILLER_71_796 ();
 sg13g2_fill_2 FILLER_71_817 ();
 sg13g2_fill_1 FILLER_71_819 ();
 sg13g2_fill_2 FILLER_71_825 ();
 sg13g2_fill_1 FILLER_71_827 ();
 sg13g2_fill_2 FILLER_71_833 ();
 sg13g2_fill_1 FILLER_71_835 ();
 sg13g2_decap_8 FILLER_71_865 ();
 sg13g2_decap_4 FILLER_71_872 ();
 sg13g2_fill_1 FILLER_71_876 ();
 sg13g2_decap_8 FILLER_71_901 ();
 sg13g2_fill_2 FILLER_71_912 ();
 sg13g2_decap_4 FILLER_71_961 ();
 sg13g2_fill_2 FILLER_71_975 ();
 sg13g2_fill_1 FILLER_71_977 ();
 sg13g2_decap_4 FILLER_71_991 ();
 sg13g2_decap_4 FILLER_71_1003 ();
 sg13g2_fill_1 FILLER_71_1007 ();
 sg13g2_decap_4 FILLER_71_1030 ();
 sg13g2_fill_2 FILLER_71_1051 ();
 sg13g2_fill_1 FILLER_71_1053 ();
 sg13g2_fill_2 FILLER_71_1080 ();
 sg13g2_decap_4 FILLER_71_1088 ();
 sg13g2_decap_4 FILLER_71_1116 ();
 sg13g2_fill_1 FILLER_71_1120 ();
 sg13g2_decap_8 FILLER_71_1127 ();
 sg13g2_fill_2 FILLER_71_1149 ();
 sg13g2_fill_1 FILLER_71_1151 ();
 sg13g2_fill_2 FILLER_71_1180 ();
 sg13g2_fill_1 FILLER_71_1182 ();
 sg13g2_fill_2 FILLER_71_1200 ();
 sg13g2_fill_1 FILLER_71_1202 ();
 sg13g2_decap_4 FILLER_71_1217 ();
 sg13g2_fill_1 FILLER_71_1221 ();
 sg13g2_fill_2 FILLER_71_1227 ();
 sg13g2_fill_1 FILLER_71_1229 ();
 sg13g2_decap_8 FILLER_71_1238 ();
 sg13g2_decap_4 FILLER_71_1245 ();
 sg13g2_fill_1 FILLER_71_1249 ();
 sg13g2_decap_8 FILLER_71_1267 ();
 sg13g2_decap_4 FILLER_71_1274 ();
 sg13g2_fill_1 FILLER_71_1278 ();
 sg13g2_fill_1 FILLER_71_1287 ();
 sg13g2_decap_4 FILLER_71_1295 ();
 sg13g2_fill_1 FILLER_71_1299 ();
 sg13g2_decap_8 FILLER_71_1314 ();
 sg13g2_decap_4 FILLER_71_1321 ();
 sg13g2_fill_1 FILLER_71_1353 ();
 sg13g2_fill_1 FILLER_71_1389 ();
 sg13g2_decap_8 FILLER_71_1408 ();
 sg13g2_fill_1 FILLER_71_1415 ();
 sg13g2_fill_2 FILLER_71_1424 ();
 sg13g2_fill_1 FILLER_71_1426 ();
 sg13g2_fill_2 FILLER_71_1440 ();
 sg13g2_fill_1 FILLER_71_1442 ();
 sg13g2_decap_8 FILLER_71_1451 ();
 sg13g2_decap_8 FILLER_71_1458 ();
 sg13g2_fill_1 FILLER_71_1465 ();
 sg13g2_fill_2 FILLER_71_1479 ();
 sg13g2_fill_1 FILLER_71_1481 ();
 sg13g2_fill_1 FILLER_71_1503 ();
 sg13g2_fill_1 FILLER_71_1510 ();
 sg13g2_decap_8 FILLER_71_1517 ();
 sg13g2_decap_4 FILLER_71_1524 ();
 sg13g2_fill_2 FILLER_71_1538 ();
 sg13g2_fill_1 FILLER_71_1540 ();
 sg13g2_fill_1 FILLER_71_1547 ();
 sg13g2_fill_2 FILLER_71_1562 ();
 sg13g2_fill_1 FILLER_71_1574 ();
 sg13g2_fill_2 FILLER_71_1579 ();
 sg13g2_fill_2 FILLER_71_1605 ();
 sg13g2_fill_1 FILLER_71_1607 ();
 sg13g2_decap_8 FILLER_71_1628 ();
 sg13g2_decap_8 FILLER_71_1635 ();
 sg13g2_decap_4 FILLER_71_1642 ();
 sg13g2_fill_1 FILLER_71_1646 ();
 sg13g2_decap_4 FILLER_71_1687 ();
 sg13g2_fill_1 FILLER_71_1691 ();
 sg13g2_fill_2 FILLER_71_1696 ();
 sg13g2_fill_1 FILLER_71_1707 ();
 sg13g2_fill_1 FILLER_71_1713 ();
 sg13g2_fill_1 FILLER_71_1729 ();
 sg13g2_fill_1 FILLER_71_1747 ();
 sg13g2_decap_4 FILLER_71_1756 ();
 sg13g2_fill_1 FILLER_71_1765 ();
 sg13g2_decap_4 FILLER_71_1774 ();
 sg13g2_fill_1 FILLER_71_1778 ();
 sg13g2_fill_2 FILLER_71_1785 ();
 sg13g2_fill_1 FILLER_71_1787 ();
 sg13g2_fill_1 FILLER_71_1808 ();
 sg13g2_fill_2 FILLER_71_1815 ();
 sg13g2_fill_1 FILLER_71_1817 ();
 sg13g2_fill_1 FILLER_71_1828 ();
 sg13g2_decap_8 FILLER_71_1834 ();
 sg13g2_fill_1 FILLER_71_1841 ();
 sg13g2_fill_2 FILLER_71_1856 ();
 sg13g2_fill_1 FILLER_71_1858 ();
 sg13g2_decap_4 FILLER_71_1915 ();
 sg13g2_fill_2 FILLER_71_1919 ();
 sg13g2_fill_2 FILLER_71_1927 ();
 sg13g2_fill_1 FILLER_71_1929 ();
 sg13g2_fill_1 FILLER_71_1936 ();
 sg13g2_decap_8 FILLER_71_1943 ();
 sg13g2_decap_8 FILLER_71_1962 ();
 sg13g2_decap_8 FILLER_71_1988 ();
 sg13g2_fill_1 FILLER_71_2030 ();
 sg13g2_fill_2 FILLER_71_2036 ();
 sg13g2_fill_2 FILLER_71_2058 ();
 sg13g2_decap_8 FILLER_71_2080 ();
 sg13g2_decap_4 FILLER_71_2087 ();
 sg13g2_fill_1 FILLER_71_2091 ();
 sg13g2_fill_1 FILLER_71_2112 ();
 sg13g2_fill_2 FILLER_71_2131 ();
 sg13g2_fill_1 FILLER_71_2133 ();
 sg13g2_decap_4 FILLER_71_2152 ();
 sg13g2_fill_2 FILLER_71_2156 ();
 sg13g2_decap_4 FILLER_71_2168 ();
 sg13g2_fill_2 FILLER_71_2185 ();
 sg13g2_fill_1 FILLER_71_2187 ();
 sg13g2_decap_8 FILLER_71_2204 ();
 sg13g2_decap_8 FILLER_71_2211 ();
 sg13g2_fill_2 FILLER_71_2231 ();
 sg13g2_fill_1 FILLER_71_2233 ();
 sg13g2_decap_8 FILLER_71_2285 ();
 sg13g2_fill_2 FILLER_71_2292 ();
 sg13g2_fill_2 FILLER_71_2311 ();
 sg13g2_fill_2 FILLER_71_2323 ();
 sg13g2_decap_8 FILLER_71_2333 ();
 sg13g2_decap_8 FILLER_71_2340 ();
 sg13g2_decap_8 FILLER_71_2351 ();
 sg13g2_fill_2 FILLER_71_2358 ();
 sg13g2_fill_1 FILLER_71_2360 ();
 sg13g2_fill_2 FILLER_71_2367 ();
 sg13g2_decap_4 FILLER_71_2413 ();
 sg13g2_fill_1 FILLER_71_2417 ();
 sg13g2_fill_2 FILLER_71_2431 ();
 sg13g2_decap_4 FILLER_71_2442 ();
 sg13g2_fill_1 FILLER_71_2446 ();
 sg13g2_fill_2 FILLER_71_2460 ();
 sg13g2_fill_1 FILLER_71_2462 ();
 sg13g2_fill_1 FILLER_71_2476 ();
 sg13g2_fill_1 FILLER_71_2511 ();
 sg13g2_fill_2 FILLER_71_2516 ();
 sg13g2_fill_1 FILLER_71_2518 ();
 sg13g2_fill_2 FILLER_71_2523 ();
 sg13g2_fill_2 FILLER_71_2539 ();
 sg13g2_decap_8 FILLER_71_2553 ();
 sg13g2_decap_4 FILLER_71_2628 ();
 sg13g2_fill_2 FILLER_71_2632 ();
 sg13g2_fill_2 FILLER_71_2642 ();
 sg13g2_fill_1 FILLER_71_2654 ();
 sg13g2_decap_4 FILLER_71_2663 ();
 sg13g2_decap_8 FILLER_71_2687 ();
 sg13g2_fill_2 FILLER_71_2694 ();
 sg13g2_fill_1 FILLER_71_2708 ();
 sg13g2_decap_8 FILLER_71_2721 ();
 sg13g2_fill_1 FILLER_71_2728 ();
 sg13g2_fill_2 FILLER_71_2746 ();
 sg13g2_decap_4 FILLER_71_2754 ();
 sg13g2_fill_1 FILLER_71_2758 ();
 sg13g2_decap_8 FILLER_71_2768 ();
 sg13g2_decap_4 FILLER_71_2775 ();
 sg13g2_fill_2 FILLER_71_2779 ();
 sg13g2_fill_2 FILLER_71_2800 ();
 sg13g2_decap_8 FILLER_71_2828 ();
 sg13g2_decap_8 FILLER_71_2835 ();
 sg13g2_decap_8 FILLER_71_2842 ();
 sg13g2_fill_1 FILLER_71_2849 ();
 sg13g2_fill_2 FILLER_71_2867 ();
 sg13g2_fill_1 FILLER_71_2869 ();
 sg13g2_decap_4 FILLER_71_2888 ();
 sg13g2_fill_2 FILLER_71_2892 ();
 sg13g2_decap_8 FILLER_71_2900 ();
 sg13g2_fill_1 FILLER_71_2907 ();
 sg13g2_decap_8 FILLER_71_2912 ();
 sg13g2_fill_2 FILLER_71_2919 ();
 sg13g2_decap_4 FILLER_71_2931 ();
 sg13g2_fill_2 FILLER_71_2950 ();
 sg13g2_fill_2 FILLER_71_2967 ();
 sg13g2_fill_1 FILLER_71_2982 ();
 sg13g2_fill_2 FILLER_71_3009 ();
 sg13g2_fill_1 FILLER_71_3011 ();
 sg13g2_fill_1 FILLER_71_3020 ();
 sg13g2_decap_4 FILLER_71_3030 ();
 sg13g2_fill_2 FILLER_71_3034 ();
 sg13g2_fill_2 FILLER_71_3041 ();
 sg13g2_fill_1 FILLER_71_3043 ();
 sg13g2_decap_8 FILLER_71_3053 ();
 sg13g2_decap_8 FILLER_71_3060 ();
 sg13g2_decap_8 FILLER_71_3082 ();
 sg13g2_decap_4 FILLER_71_3089 ();
 sg13g2_decap_4 FILLER_71_3101 ();
 sg13g2_fill_1 FILLER_71_3109 ();
 sg13g2_decap_8 FILLER_71_3115 ();
 sg13g2_decap_4 FILLER_71_3122 ();
 sg13g2_decap_8 FILLER_71_3136 ();
 sg13g2_decap_8 FILLER_71_3143 ();
 sg13g2_fill_2 FILLER_71_3159 ();
 sg13g2_decap_4 FILLER_71_3179 ();
 sg13g2_fill_1 FILLER_71_3183 ();
 sg13g2_fill_1 FILLER_71_3188 ();
 sg13g2_decap_4 FILLER_71_3194 ();
 sg13g2_fill_1 FILLER_71_3198 ();
 sg13g2_decap_8 FILLER_71_3205 ();
 sg13g2_fill_2 FILLER_71_3212 ();
 sg13g2_fill_1 FILLER_71_3214 ();
 sg13g2_fill_2 FILLER_71_3228 ();
 sg13g2_fill_1 FILLER_71_3230 ();
 sg13g2_fill_2 FILLER_71_3237 ();
 sg13g2_decap_8 FILLER_71_3242 ();
 sg13g2_fill_2 FILLER_71_3249 ();
 sg13g2_decap_4 FILLER_71_3269 ();
 sg13g2_decap_4 FILLER_71_3287 ();
 sg13g2_fill_1 FILLER_71_3291 ();
 sg13g2_fill_1 FILLER_71_3329 ();
 sg13g2_fill_2 FILLER_71_3344 ();
 sg13g2_fill_1 FILLER_71_3346 ();
 sg13g2_decap_4 FILLER_71_3360 ();
 sg13g2_fill_1 FILLER_71_3364 ();
 sg13g2_decap_4 FILLER_71_3384 ();
 sg13g2_fill_2 FILLER_71_3404 ();
 sg13g2_fill_2 FILLER_71_3419 ();
 sg13g2_fill_1 FILLER_71_3421 ();
 sg13g2_fill_2 FILLER_71_3434 ();
 sg13g2_decap_8 FILLER_71_3440 ();
 sg13g2_fill_2 FILLER_71_3447 ();
 sg13g2_fill_1 FILLER_71_3449 ();
 sg13g2_decap_8 FILLER_71_3463 ();
 sg13g2_decap_8 FILLER_71_3470 ();
 sg13g2_decap_8 FILLER_71_3477 ();
 sg13g2_decap_8 FILLER_71_3484 ();
 sg13g2_decap_8 FILLER_71_3491 ();
 sg13g2_decap_8 FILLER_71_3498 ();
 sg13g2_decap_8 FILLER_71_3505 ();
 sg13g2_decap_8 FILLER_71_3512 ();
 sg13g2_decap_8 FILLER_71_3519 ();
 sg13g2_decap_8 FILLER_71_3526 ();
 sg13g2_decap_8 FILLER_71_3533 ();
 sg13g2_decap_8 FILLER_71_3540 ();
 sg13g2_decap_8 FILLER_71_3547 ();
 sg13g2_decap_8 FILLER_71_3554 ();
 sg13g2_decap_8 FILLER_71_3561 ();
 sg13g2_decap_8 FILLER_71_3568 ();
 sg13g2_decap_4 FILLER_71_3575 ();
 sg13g2_fill_1 FILLER_71_3579 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_fill_1 FILLER_72_168 ();
 sg13g2_fill_2 FILLER_72_196 ();
 sg13g2_fill_2 FILLER_72_212 ();
 sg13g2_fill_1 FILLER_72_214 ();
 sg13g2_fill_2 FILLER_72_228 ();
 sg13g2_fill_2 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_292 ();
 sg13g2_fill_2 FILLER_72_375 ();
 sg13g2_fill_1 FILLER_72_377 ();
 sg13g2_fill_1 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_fill_2 FILLER_72_448 ();
 sg13g2_decap_8 FILLER_72_503 ();
 sg13g2_fill_2 FILLER_72_510 ();
 sg13g2_fill_1 FILLER_72_512 ();
 sg13g2_fill_1 FILLER_72_518 ();
 sg13g2_decap_4 FILLER_72_523 ();
 sg13g2_fill_1 FILLER_72_527 ();
 sg13g2_decap_4 FILLER_72_534 ();
 sg13g2_decap_8 FILLER_72_550 ();
 sg13g2_decap_4 FILLER_72_557 ();
 sg13g2_fill_2 FILLER_72_561 ();
 sg13g2_fill_2 FILLER_72_581 ();
 sg13g2_fill_2 FILLER_72_608 ();
 sg13g2_decap_4 FILLER_72_622 ();
 sg13g2_fill_1 FILLER_72_626 ();
 sg13g2_fill_2 FILLER_72_645 ();
 sg13g2_fill_1 FILLER_72_647 ();
 sg13g2_fill_1 FILLER_72_659 ();
 sg13g2_fill_1 FILLER_72_671 ();
 sg13g2_fill_2 FILLER_72_685 ();
 sg13g2_fill_1 FILLER_72_687 ();
 sg13g2_decap_8 FILLER_72_716 ();
 sg13g2_decap_4 FILLER_72_723 ();
 sg13g2_fill_1 FILLER_72_727 ();
 sg13g2_decap_8 FILLER_72_769 ();
 sg13g2_decap_4 FILLER_72_776 ();
 sg13g2_fill_1 FILLER_72_780 ();
 sg13g2_fill_1 FILLER_72_787 ();
 sg13g2_decap_4 FILLER_72_810 ();
 sg13g2_decap_8 FILLER_72_833 ();
 sg13g2_fill_2 FILLER_72_840 ();
 sg13g2_fill_1 FILLER_72_846 ();
 sg13g2_fill_1 FILLER_72_896 ();
 sg13g2_decap_8 FILLER_72_913 ();
 sg13g2_fill_2 FILLER_72_920 ();
 sg13g2_decap_8 FILLER_72_927 ();
 sg13g2_decap_4 FILLER_72_934 ();
 sg13g2_fill_2 FILLER_72_938 ();
 sg13g2_decap_8 FILLER_72_952 ();
 sg13g2_decap_8 FILLER_72_959 ();
 sg13g2_decap_4 FILLER_72_966 ();
 sg13g2_fill_1 FILLER_72_970 ();
 sg13g2_fill_2 FILLER_72_980 ();
 sg13g2_fill_1 FILLER_72_982 ();
 sg13g2_decap_8 FILLER_72_988 ();
 sg13g2_decap_4 FILLER_72_995 ();
 sg13g2_fill_2 FILLER_72_1013 ();
 sg13g2_decap_4 FILLER_72_1018 ();
 sg13g2_fill_2 FILLER_72_1022 ();
 sg13g2_decap_4 FILLER_72_1039 ();
 sg13g2_fill_2 FILLER_72_1043 ();
 sg13g2_fill_1 FILLER_72_1050 ();
 sg13g2_decap_4 FILLER_72_1079 ();
 sg13g2_fill_2 FILLER_72_1083 ();
 sg13g2_decap_8 FILLER_72_1089 ();
 sg13g2_decap_8 FILLER_72_1096 ();
 sg13g2_decap_4 FILLER_72_1103 ();
 sg13g2_fill_1 FILLER_72_1107 ();
 sg13g2_decap_8 FILLER_72_1114 ();
 sg13g2_fill_2 FILLER_72_1121 ();
 sg13g2_fill_1 FILLER_72_1123 ();
 sg13g2_decap_8 FILLER_72_1162 ();
 sg13g2_decap_4 FILLER_72_1169 ();
 sg13g2_fill_2 FILLER_72_1188 ();
 sg13g2_fill_1 FILLER_72_1190 ();
 sg13g2_decap_4 FILLER_72_1206 ();
 sg13g2_fill_2 FILLER_72_1218 ();
 sg13g2_fill_1 FILLER_72_1233 ();
 sg13g2_decap_8 FILLER_72_1252 ();
 sg13g2_decap_8 FILLER_72_1259 ();
 sg13g2_decap_8 FILLER_72_1266 ();
 sg13g2_decap_4 FILLER_72_1293 ();
 sg13g2_fill_2 FILLER_72_1297 ();
 sg13g2_decap_8 FILLER_72_1305 ();
 sg13g2_decap_8 FILLER_72_1312 ();
 sg13g2_fill_2 FILLER_72_1319 ();
 sg13g2_fill_1 FILLER_72_1321 ();
 sg13g2_fill_2 FILLER_72_1344 ();
 sg13g2_fill_1 FILLER_72_1346 ();
 sg13g2_fill_1 FILLER_72_1384 ();
 sg13g2_decap_4 FILLER_72_1389 ();
 sg13g2_fill_2 FILLER_72_1393 ();
 sg13g2_decap_8 FILLER_72_1400 ();
 sg13g2_decap_8 FILLER_72_1407 ();
 sg13g2_fill_1 FILLER_72_1423 ();
 sg13g2_fill_1 FILLER_72_1429 ();
 sg13g2_decap_8 FILLER_72_1458 ();
 sg13g2_fill_2 FILLER_72_1480 ();
 sg13g2_fill_1 FILLER_72_1482 ();
 sg13g2_fill_2 FILLER_72_1488 ();
 sg13g2_fill_1 FILLER_72_1490 ();
 sg13g2_fill_1 FILLER_72_1499 ();
 sg13g2_decap_8 FILLER_72_1512 ();
 sg13g2_decap_4 FILLER_72_1519 ();
 sg13g2_fill_1 FILLER_72_1535 ();
 sg13g2_decap_8 FILLER_72_1539 ();
 sg13g2_decap_4 FILLER_72_1546 ();
 sg13g2_fill_2 FILLER_72_1564 ();
 sg13g2_fill_2 FILLER_72_1571 ();
 sg13g2_fill_1 FILLER_72_1573 ();
 sg13g2_decap_4 FILLER_72_1597 ();
 sg13g2_fill_1 FILLER_72_1601 ();
 sg13g2_decap_8 FILLER_72_1616 ();
 sg13g2_fill_1 FILLER_72_1623 ();
 sg13g2_fill_2 FILLER_72_1637 ();
 sg13g2_decap_4 FILLER_72_1666 ();
 sg13g2_fill_1 FILLER_72_1670 ();
 sg13g2_fill_2 FILLER_72_1692 ();
 sg13g2_decap_4 FILLER_72_1725 ();
 sg13g2_decap_8 FILLER_72_1741 ();
 sg13g2_fill_2 FILLER_72_1748 ();
 sg13g2_decap_8 FILLER_72_1773 ();
 sg13g2_decap_4 FILLER_72_1780 ();
 sg13g2_fill_2 FILLER_72_1784 ();
 sg13g2_fill_2 FILLER_72_1792 ();
 sg13g2_decap_8 FILLER_72_1820 ();
 sg13g2_decap_4 FILLER_72_1827 ();
 sg13g2_decap_4 FILLER_72_1841 ();
 sg13g2_fill_1 FILLER_72_1845 ();
 sg13g2_fill_2 FILLER_72_1852 ();
 sg13g2_fill_1 FILLER_72_1854 ();
 sg13g2_decap_4 FILLER_72_1889 ();
 sg13g2_fill_1 FILLER_72_1893 ();
 sg13g2_fill_2 FILLER_72_1902 ();
 sg13g2_fill_2 FILLER_72_1928 ();
 sg13g2_decap_4 FILLER_72_1943 ();
 sg13g2_decap_8 FILLER_72_1966 ();
 sg13g2_decap_4 FILLER_72_1979 ();
 sg13g2_fill_1 FILLER_72_1983 ();
 sg13g2_fill_1 FILLER_72_1997 ();
 sg13g2_fill_2 FILLER_72_2009 ();
 sg13g2_decap_4 FILLER_72_2021 ();
 sg13g2_decap_4 FILLER_72_2060 ();
 sg13g2_decap_8 FILLER_72_2076 ();
 sg13g2_decap_8 FILLER_72_2083 ();
 sg13g2_decap_4 FILLER_72_2090 ();
 sg13g2_decap_4 FILLER_72_2126 ();
 sg13g2_decap_4 FILLER_72_2134 ();
 sg13g2_fill_1 FILLER_72_2148 ();
 sg13g2_decap_8 FILLER_72_2168 ();
 sg13g2_decap_8 FILLER_72_2208 ();
 sg13g2_fill_2 FILLER_72_2215 ();
 sg13g2_fill_1 FILLER_72_2217 ();
 sg13g2_fill_2 FILLER_72_2245 ();
 sg13g2_decap_4 FILLER_72_2255 ();
 sg13g2_decap_8 FILLER_72_2264 ();
 sg13g2_fill_1 FILLER_72_2271 ();
 sg13g2_decap_4 FILLER_72_2275 ();
 sg13g2_fill_1 FILLER_72_2313 ();
 sg13g2_decap_4 FILLER_72_2319 ();
 sg13g2_decap_4 FILLER_72_2328 ();
 sg13g2_fill_1 FILLER_72_2332 ();
 sg13g2_decap_8 FILLER_72_2339 ();
 sg13g2_decap_8 FILLER_72_2346 ();
 sg13g2_fill_2 FILLER_72_2353 ();
 sg13g2_fill_1 FILLER_72_2355 ();
 sg13g2_fill_1 FILLER_72_2375 ();
 sg13g2_fill_2 FILLER_72_2382 ();
 sg13g2_fill_1 FILLER_72_2384 ();
 sg13g2_fill_2 FILLER_72_2393 ();
 sg13g2_decap_8 FILLER_72_2409 ();
 sg13g2_fill_2 FILLER_72_2420 ();
 sg13g2_decap_4 FILLER_72_2426 ();
 sg13g2_fill_1 FILLER_72_2430 ();
 sg13g2_fill_1 FILLER_72_2441 ();
 sg13g2_fill_1 FILLER_72_2454 ();
 sg13g2_decap_8 FILLER_72_2473 ();
 sg13g2_fill_2 FILLER_72_2480 ();
 sg13g2_fill_2 FILLER_72_2502 ();
 sg13g2_decap_8 FILLER_72_2514 ();
 sg13g2_decap_4 FILLER_72_2521 ();
 sg13g2_fill_1 FILLER_72_2525 ();
 sg13g2_fill_1 FILLER_72_2530 ();
 sg13g2_fill_1 FILLER_72_2535 ();
 sg13g2_fill_2 FILLER_72_2541 ();
 sg13g2_fill_2 FILLER_72_2547 ();
 sg13g2_decap_4 FILLER_72_2561 ();
 sg13g2_fill_2 FILLER_72_2565 ();
 sg13g2_fill_2 FILLER_72_2573 ();
 sg13g2_decap_8 FILLER_72_2585 ();
 sg13g2_fill_1 FILLER_72_2592 ();
 sg13g2_decap_4 FILLER_72_2618 ();
 sg13g2_fill_2 FILLER_72_2622 ();
 sg13g2_decap_4 FILLER_72_2628 ();
 sg13g2_decap_8 FILLER_72_2637 ();
 sg13g2_fill_2 FILLER_72_2644 ();
 sg13g2_fill_1 FILLER_72_2664 ();
 sg13g2_decap_8 FILLER_72_2689 ();
 sg13g2_decap_4 FILLER_72_2696 ();
 sg13g2_fill_2 FILLER_72_2700 ();
 sg13g2_fill_1 FILLER_72_2720 ();
 sg13g2_decap_4 FILLER_72_2726 ();
 sg13g2_fill_1 FILLER_72_2730 ();
 sg13g2_decap_8 FILLER_72_2745 ();
 sg13g2_decap_4 FILLER_72_2752 ();
 sg13g2_fill_2 FILLER_72_2756 ();
 sg13g2_decap_8 FILLER_72_2768 ();
 sg13g2_decap_8 FILLER_72_2775 ();
 sg13g2_fill_1 FILLER_72_2790 ();
 sg13g2_fill_2 FILLER_72_2800 ();
 sg13g2_fill_1 FILLER_72_2802 ();
 sg13g2_fill_1 FILLER_72_2815 ();
 sg13g2_decap_8 FILLER_72_2835 ();
 sg13g2_decap_8 FILLER_72_2842 ();
 sg13g2_decap_8 FILLER_72_2849 ();
 sg13g2_decap_4 FILLER_72_2856 ();
 sg13g2_fill_1 FILLER_72_2860 ();
 sg13g2_fill_1 FILLER_72_2866 ();
 sg13g2_fill_1 FILLER_72_2878 ();
 sg13g2_decap_8 FILLER_72_2892 ();
 sg13g2_decap_4 FILLER_72_2899 ();
 sg13g2_fill_1 FILLER_72_2931 ();
 sg13g2_decap_8 FILLER_72_2947 ();
 sg13g2_decap_4 FILLER_72_2962 ();
 sg13g2_fill_1 FILLER_72_2966 ();
 sg13g2_fill_2 FILLER_72_2972 ();
 sg13g2_fill_1 FILLER_72_2978 ();
 sg13g2_decap_4 FILLER_72_2992 ();
 sg13g2_fill_2 FILLER_72_2996 ();
 sg13g2_decap_8 FILLER_72_3022 ();
 sg13g2_decap_8 FILLER_72_3057 ();
 sg13g2_fill_2 FILLER_72_3064 ();
 sg13g2_fill_1 FILLER_72_3066 ();
 sg13g2_decap_8 FILLER_72_3080 ();
 sg13g2_fill_1 FILLER_72_3087 ();
 sg13g2_fill_2 FILLER_72_3096 ();
 sg13g2_decap_4 FILLER_72_3141 ();
 sg13g2_fill_1 FILLER_72_3145 ();
 sg13g2_fill_2 FILLER_72_3175 ();
 sg13g2_fill_1 FILLER_72_3177 ();
 sg13g2_decap_8 FILLER_72_3211 ();
 sg13g2_decap_4 FILLER_72_3218 ();
 sg13g2_decap_8 FILLER_72_3226 ();
 sg13g2_decap_8 FILLER_72_3246 ();
 sg13g2_fill_1 FILLER_72_3253 ();
 sg13g2_decap_8 FILLER_72_3273 ();
 sg13g2_fill_2 FILLER_72_3280 ();
 sg13g2_decap_8 FILLER_72_3287 ();
 sg13g2_decap_8 FILLER_72_3294 ();
 sg13g2_decap_4 FILLER_72_3301 ();
 sg13g2_decap_4 FILLER_72_3309 ();
 sg13g2_fill_2 FILLER_72_3313 ();
 sg13g2_fill_2 FILLER_72_3321 ();
 sg13g2_decap_8 FILLER_72_3353 ();
 sg13g2_fill_2 FILLER_72_3377 ();
 sg13g2_fill_1 FILLER_72_3379 ();
 sg13g2_fill_2 FILLER_72_3390 ();
 sg13g2_fill_2 FILLER_72_3405 ();
 sg13g2_fill_1 FILLER_72_3415 ();
 sg13g2_fill_1 FILLER_72_3425 ();
 sg13g2_decap_8 FILLER_72_3463 ();
 sg13g2_decap_8 FILLER_72_3470 ();
 sg13g2_decap_8 FILLER_72_3477 ();
 sg13g2_decap_8 FILLER_72_3484 ();
 sg13g2_decap_8 FILLER_72_3491 ();
 sg13g2_decap_8 FILLER_72_3498 ();
 sg13g2_decap_8 FILLER_72_3505 ();
 sg13g2_decap_8 FILLER_72_3512 ();
 sg13g2_decap_8 FILLER_72_3519 ();
 sg13g2_decap_8 FILLER_72_3526 ();
 sg13g2_decap_8 FILLER_72_3533 ();
 sg13g2_decap_8 FILLER_72_3540 ();
 sg13g2_decap_8 FILLER_72_3547 ();
 sg13g2_decap_8 FILLER_72_3554 ();
 sg13g2_decap_8 FILLER_72_3561 ();
 sg13g2_decap_8 FILLER_72_3568 ();
 sg13g2_decap_4 FILLER_72_3575 ();
 sg13g2_fill_1 FILLER_72_3579 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_fill_2 FILLER_73_168 ();
 sg13g2_fill_1 FILLER_73_170 ();
 sg13g2_fill_2 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_248 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_decap_4 FILLER_73_259 ();
 sg13g2_fill_2 FILLER_73_263 ();
 sg13g2_decap_4 FILLER_73_314 ();
 sg13g2_fill_1 FILLER_73_318 ();
 sg13g2_fill_2 FILLER_73_346 ();
 sg13g2_decap_8 FILLER_73_368 ();
 sg13g2_fill_2 FILLER_73_375 ();
 sg13g2_fill_1 FILLER_73_377 ();
 sg13g2_fill_2 FILLER_73_391 ();
 sg13g2_fill_2 FILLER_73_434 ();
 sg13g2_decap_4 FILLER_73_441 ();
 sg13g2_fill_2 FILLER_73_445 ();
 sg13g2_fill_2 FILLER_73_452 ();
 sg13g2_decap_8 FILLER_73_478 ();
 sg13g2_decap_4 FILLER_73_485 ();
 sg13g2_fill_2 FILLER_73_502 ();
 sg13g2_fill_1 FILLER_73_504 ();
 sg13g2_decap_8 FILLER_73_530 ();
 sg13g2_decap_4 FILLER_73_537 ();
 sg13g2_fill_2 FILLER_73_541 ();
 sg13g2_fill_2 FILLER_73_567 ();
 sg13g2_fill_2 FILLER_73_578 ();
 sg13g2_fill_1 FILLER_73_580 ();
 sg13g2_fill_2 FILLER_73_594 ();
 sg13g2_fill_1 FILLER_73_596 ();
 sg13g2_fill_1 FILLER_73_621 ();
 sg13g2_fill_1 FILLER_73_626 ();
 sg13g2_fill_2 FILLER_73_632 ();
 sg13g2_fill_1 FILLER_73_634 ();
 sg13g2_decap_4 FILLER_73_648 ();
 sg13g2_fill_1 FILLER_73_670 ();
 sg13g2_decap_4 FILLER_73_674 ();
 sg13g2_fill_1 FILLER_73_678 ();
 sg13g2_decap_8 FILLER_73_691 ();
 sg13g2_fill_2 FILLER_73_698 ();
 sg13g2_decap_8 FILLER_73_704 ();
 sg13g2_decap_8 FILLER_73_711 ();
 sg13g2_fill_1 FILLER_73_722 ();
 sg13g2_fill_2 FILLER_73_747 ();
 sg13g2_fill_1 FILLER_73_749 ();
 sg13g2_fill_2 FILLER_73_758 ();
 sg13g2_fill_1 FILLER_73_764 ();
 sg13g2_fill_2 FILLER_73_783 ();
 sg13g2_fill_1 FILLER_73_785 ();
 sg13g2_decap_8 FILLER_73_792 ();
 sg13g2_fill_1 FILLER_73_799 ();
 sg13g2_fill_1 FILLER_73_809 ();
 sg13g2_decap_8 FILLER_73_820 ();
 sg13g2_decap_8 FILLER_73_827 ();
 sg13g2_decap_4 FILLER_73_834 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_8 FILLER_73_857 ();
 sg13g2_fill_2 FILLER_73_868 ();
 sg13g2_fill_1 FILLER_73_870 ();
 sg13g2_fill_1 FILLER_73_880 ();
 sg13g2_decap_4 FILLER_73_899 ();
 sg13g2_decap_4 FILLER_73_927 ();
 sg13g2_fill_2 FILLER_73_931 ();
 sg13g2_decap_4 FILLER_73_936 ();
 sg13g2_decap_8 FILLER_73_959 ();
 sg13g2_fill_2 FILLER_73_972 ();
 sg13g2_decap_8 FILLER_73_980 ();
 sg13g2_fill_2 FILLER_73_987 ();
 sg13g2_fill_1 FILLER_73_1005 ();
 sg13g2_fill_2 FILLER_73_1019 ();
 sg13g2_fill_1 FILLER_73_1021 ();
 sg13g2_fill_2 FILLER_73_1027 ();
 sg13g2_fill_1 FILLER_73_1029 ();
 sg13g2_fill_2 FILLER_73_1045 ();
 sg13g2_decap_4 FILLER_73_1051 ();
 sg13g2_fill_1 FILLER_73_1055 ();
 sg13g2_fill_2 FILLER_73_1064 ();
 sg13g2_fill_1 FILLER_73_1066 ();
 sg13g2_decap_8 FILLER_73_1072 ();
 sg13g2_decap_4 FILLER_73_1107 ();
 sg13g2_fill_2 FILLER_73_1111 ();
 sg13g2_decap_4 FILLER_73_1134 ();
 sg13g2_fill_1 FILLER_73_1138 ();
 sg13g2_decap_4 FILLER_73_1143 ();
 sg13g2_fill_2 FILLER_73_1147 ();
 sg13g2_decap_8 FILLER_73_1167 ();
 sg13g2_fill_2 FILLER_73_1174 ();
 sg13g2_fill_1 FILLER_73_1199 ();
 sg13g2_decap_8 FILLER_73_1205 ();
 sg13g2_fill_2 FILLER_73_1212 ();
 sg13g2_decap_4 FILLER_73_1226 ();
 sg13g2_fill_2 FILLER_73_1230 ();
 sg13g2_fill_1 FILLER_73_1245 ();
 sg13g2_decap_8 FILLER_73_1256 ();
 sg13g2_fill_2 FILLER_73_1263 ();
 sg13g2_fill_1 FILLER_73_1265 ();
 sg13g2_fill_2 FILLER_73_1276 ();
 sg13g2_fill_1 FILLER_73_1281 ();
 sg13g2_fill_2 FILLER_73_1287 ();
 sg13g2_fill_2 FILLER_73_1297 ();
 sg13g2_fill_1 FILLER_73_1299 ();
 sg13g2_fill_2 FILLER_73_1306 ();
 sg13g2_fill_1 FILLER_73_1308 ();
 sg13g2_decap_4 FILLER_73_1322 ();
 sg13g2_fill_1 FILLER_73_1326 ();
 sg13g2_fill_1 FILLER_73_1333 ();
 sg13g2_decap_4 FILLER_73_1368 ();
 sg13g2_fill_1 FILLER_73_1372 ();
 sg13g2_fill_2 FILLER_73_1378 ();
 sg13g2_fill_1 FILLER_73_1380 ();
 sg13g2_fill_2 FILLER_73_1401 ();
 sg13g2_decap_4 FILLER_73_1413 ();
 sg13g2_decap_4 FILLER_73_1422 ();
 sg13g2_fill_2 FILLER_73_1431 ();
 sg13g2_decap_8 FILLER_73_1438 ();
 sg13g2_decap_8 FILLER_73_1445 ();
 sg13g2_decap_8 FILLER_73_1452 ();
 sg13g2_decap_4 FILLER_73_1459 ();
 sg13g2_fill_1 FILLER_73_1463 ();
 sg13g2_fill_1 FILLER_73_1484 ();
 sg13g2_decap_8 FILLER_73_1490 ();
 sg13g2_decap_4 FILLER_73_1497 ();
 sg13g2_fill_2 FILLER_73_1501 ();
 sg13g2_decap_8 FILLER_73_1519 ();
 sg13g2_fill_2 FILLER_73_1526 ();
 sg13g2_fill_1 FILLER_73_1528 ();
 sg13g2_decap_8 FILLER_73_1542 ();
 sg13g2_decap_8 FILLER_73_1549 ();
 sg13g2_fill_2 FILLER_73_1566 ();
 sg13g2_fill_1 FILLER_73_1568 ();
 sg13g2_decap_4 FILLER_73_1585 ();
 sg13g2_fill_1 FILLER_73_1589 ();
 sg13g2_fill_1 FILLER_73_1596 ();
 sg13g2_fill_2 FILLER_73_1609 ();
 sg13g2_fill_1 FILLER_73_1615 ();
 sg13g2_decap_4 FILLER_73_1641 ();
 sg13g2_fill_1 FILLER_73_1645 ();
 sg13g2_decap_8 FILLER_73_1662 ();
 sg13g2_fill_2 FILLER_73_1669 ();
 sg13g2_fill_1 FILLER_73_1671 ();
 sg13g2_decap_8 FILLER_73_1689 ();
 sg13g2_decap_8 FILLER_73_1696 ();
 sg13g2_decap_8 FILLER_73_1703 ();
 sg13g2_decap_4 FILLER_73_1710 ();
 sg13g2_fill_1 FILLER_73_1725 ();
 sg13g2_decap_8 FILLER_73_1731 ();
 sg13g2_decap_8 FILLER_73_1738 ();
 sg13g2_fill_2 FILLER_73_1745 ();
 sg13g2_fill_1 FILLER_73_1747 ();
 sg13g2_decap_8 FILLER_73_1763 ();
 sg13g2_decap_4 FILLER_73_1770 ();
 sg13g2_fill_1 FILLER_73_1774 ();
 sg13g2_decap_4 FILLER_73_1789 ();
 sg13g2_decap_8 FILLER_73_1796 ();
 sg13g2_decap_4 FILLER_73_1803 ();
 sg13g2_decap_8 FILLER_73_1811 ();
 sg13g2_decap_8 FILLER_73_1818 ();
 sg13g2_decap_8 FILLER_73_1844 ();
 sg13g2_fill_1 FILLER_73_1851 ();
 sg13g2_fill_2 FILLER_73_1863 ();
 sg13g2_fill_1 FILLER_73_1872 ();
 sg13g2_fill_2 FILLER_73_1886 ();
 sg13g2_fill_1 FILLER_73_1888 ();
 sg13g2_fill_2 FILLER_73_1910 ();
 sg13g2_fill_1 FILLER_73_1912 ();
 sg13g2_fill_1 FILLER_73_1919 ();
 sg13g2_fill_1 FILLER_73_1933 ();
 sg13g2_decap_4 FILLER_73_1949 ();
 sg13g2_fill_1 FILLER_73_1953 ();
 sg13g2_decap_4 FILLER_73_1975 ();
 sg13g2_decap_8 FILLER_73_2003 ();
 sg13g2_decap_4 FILLER_73_2010 ();
 sg13g2_fill_1 FILLER_73_2022 ();
 sg13g2_decap_8 FILLER_73_2039 ();
 sg13g2_decap_8 FILLER_73_2046 ();
 sg13g2_fill_1 FILLER_73_2063 ();
 sg13g2_decap_8 FILLER_73_2068 ();
 sg13g2_decap_4 FILLER_73_2075 ();
 sg13g2_fill_1 FILLER_73_2079 ();
 sg13g2_fill_1 FILLER_73_2085 ();
 sg13g2_decap_8 FILLER_73_2094 ();
 sg13g2_decap_4 FILLER_73_2101 ();
 sg13g2_fill_1 FILLER_73_2105 ();
 sg13g2_fill_1 FILLER_73_2110 ();
 sg13g2_decap_8 FILLER_73_2116 ();
 sg13g2_decap_8 FILLER_73_2128 ();
 sg13g2_decap_8 FILLER_73_2135 ();
 sg13g2_decap_4 FILLER_73_2142 ();
 sg13g2_fill_1 FILLER_73_2173 ();
 sg13g2_fill_2 FILLER_73_2182 ();
 sg13g2_decap_4 FILLER_73_2211 ();
 sg13g2_fill_2 FILLER_73_2234 ();
 sg13g2_fill_1 FILLER_73_2236 ();
 sg13g2_fill_2 FILLER_73_2261 ();
 sg13g2_fill_1 FILLER_73_2263 ();
 sg13g2_fill_2 FILLER_73_2280 ();
 sg13g2_decap_8 FILLER_73_2290 ();
 sg13g2_decap_8 FILLER_73_2297 ();
 sg13g2_decap_4 FILLER_73_2304 ();
 sg13g2_fill_1 FILLER_73_2350 ();
 sg13g2_fill_2 FILLER_73_2384 ();
 sg13g2_fill_1 FILLER_73_2386 ();
 sg13g2_fill_2 FILLER_73_2407 ();
 sg13g2_fill_1 FILLER_73_2409 ();
 sg13g2_fill_1 FILLER_73_2414 ();
 sg13g2_decap_4 FILLER_73_2429 ();
 sg13g2_fill_2 FILLER_73_2439 ();
 sg13g2_decap_4 FILLER_73_2448 ();
 sg13g2_fill_1 FILLER_73_2452 ();
 sg13g2_decap_8 FILLER_73_2465 ();
 sg13g2_decap_8 FILLER_73_2472 ();
 sg13g2_decap_4 FILLER_73_2479 ();
 sg13g2_fill_1 FILLER_73_2488 ();
 sg13g2_fill_2 FILLER_73_2503 ();
 sg13g2_fill_1 FILLER_73_2505 ();
 sg13g2_fill_1 FILLER_73_2519 ();
 sg13g2_fill_2 FILLER_73_2528 ();
 sg13g2_decap_4 FILLER_73_2545 ();
 sg13g2_decap_8 FILLER_73_2561 ();
 sg13g2_decap_8 FILLER_73_2568 ();
 sg13g2_decap_8 FILLER_73_2575 ();
 sg13g2_decap_4 FILLER_73_2582 ();
 sg13g2_fill_1 FILLER_73_2586 ();
 sg13g2_decap_8 FILLER_73_2606 ();
 sg13g2_fill_1 FILLER_73_2613 ();
 sg13g2_decap_8 FILLER_73_2618 ();
 sg13g2_fill_2 FILLER_73_2625 ();
 sg13g2_fill_1 FILLER_73_2627 ();
 sg13g2_fill_2 FILLER_73_2633 ();
 sg13g2_fill_1 FILLER_73_2641 ();
 sg13g2_decap_4 FILLER_73_2647 ();
 sg13g2_fill_1 FILLER_73_2651 ();
 sg13g2_decap_8 FILLER_73_2661 ();
 sg13g2_decap_4 FILLER_73_2668 ();
 sg13g2_fill_2 FILLER_73_2672 ();
 sg13g2_decap_8 FILLER_73_2683 ();
 sg13g2_decap_8 FILLER_73_2690 ();
 sg13g2_decap_8 FILLER_73_2697 ();
 sg13g2_fill_1 FILLER_73_2704 ();
 sg13g2_decap_4 FILLER_73_2721 ();
 sg13g2_fill_2 FILLER_73_2730 ();
 sg13g2_fill_1 FILLER_73_2732 ();
 sg13g2_decap_8 FILLER_73_2740 ();
 sg13g2_fill_1 FILLER_73_2747 ();
 sg13g2_decap_4 FILLER_73_2773 ();
 sg13g2_fill_2 FILLER_73_2781 ();
 sg13g2_decap_8 FILLER_73_2802 ();
 sg13g2_decap_4 FILLER_73_2843 ();
 sg13g2_fill_1 FILLER_73_2847 ();
 sg13g2_decap_4 FILLER_73_2877 ();
 sg13g2_fill_2 FILLER_73_2881 ();
 sg13g2_decap_4 FILLER_73_2893 ();
 sg13g2_fill_2 FILLER_73_2914 ();
 sg13g2_fill_2 FILLER_73_2926 ();
 sg13g2_fill_1 FILLER_73_2928 ();
 sg13g2_decap_4 FILLER_73_2957 ();
 sg13g2_fill_2 FILLER_73_2966 ();
 sg13g2_fill_2 FILLER_73_2973 ();
 sg13g2_decap_8 FILLER_73_2993 ();
 sg13g2_fill_2 FILLER_73_3006 ();
 sg13g2_fill_1 FILLER_73_3008 ();
 sg13g2_decap_8 FILLER_73_3014 ();
 sg13g2_fill_2 FILLER_73_3032 ();
 sg13g2_fill_2 FILLER_73_3046 ();
 sg13g2_fill_1 FILLER_73_3053 ();
 sg13g2_fill_1 FILLER_73_3084 ();
 sg13g2_decap_8 FILLER_73_3093 ();
 sg13g2_fill_2 FILLER_73_3100 ();
 sg13g2_fill_1 FILLER_73_3102 ();
 sg13g2_decap_8 FILLER_73_3112 ();
 sg13g2_fill_2 FILLER_73_3119 ();
 sg13g2_decap_8 FILLER_73_3138 ();
 sg13g2_decap_8 FILLER_73_3145 ();
 sg13g2_fill_2 FILLER_73_3152 ();
 sg13g2_fill_1 FILLER_73_3154 ();
 sg13g2_decap_4 FILLER_73_3160 ();
 sg13g2_decap_8 FILLER_73_3173 ();
 sg13g2_fill_2 FILLER_73_3180 ();
 sg13g2_fill_2 FILLER_73_3191 ();
 sg13g2_fill_1 FILLER_73_3193 ();
 sg13g2_decap_4 FILLER_73_3202 ();
 sg13g2_decap_4 FILLER_73_3219 ();
 sg13g2_fill_2 FILLER_73_3223 ();
 sg13g2_fill_2 FILLER_73_3256 ();
 sg13g2_fill_1 FILLER_73_3273 ();
 sg13g2_fill_2 FILLER_73_3295 ();
 sg13g2_decap_8 FILLER_73_3382 ();
 sg13g2_fill_2 FILLER_73_3389 ();
 sg13g2_fill_1 FILLER_73_3423 ();
 sg13g2_fill_2 FILLER_73_3437 ();
 sg13g2_fill_1 FILLER_73_3439 ();
 sg13g2_fill_2 FILLER_73_3444 ();
 sg13g2_decap_8 FILLER_73_3455 ();
 sg13g2_decap_8 FILLER_73_3462 ();
 sg13g2_decap_8 FILLER_73_3469 ();
 sg13g2_decap_8 FILLER_73_3476 ();
 sg13g2_decap_8 FILLER_73_3483 ();
 sg13g2_decap_8 FILLER_73_3490 ();
 sg13g2_decap_8 FILLER_73_3497 ();
 sg13g2_decap_8 FILLER_73_3504 ();
 sg13g2_decap_8 FILLER_73_3511 ();
 sg13g2_decap_8 FILLER_73_3518 ();
 sg13g2_decap_8 FILLER_73_3525 ();
 sg13g2_decap_8 FILLER_73_3532 ();
 sg13g2_decap_8 FILLER_73_3539 ();
 sg13g2_decap_8 FILLER_73_3546 ();
 sg13g2_decap_8 FILLER_73_3553 ();
 sg13g2_decap_8 FILLER_73_3560 ();
 sg13g2_decap_8 FILLER_73_3567 ();
 sg13g2_decap_4 FILLER_73_3574 ();
 sg13g2_fill_2 FILLER_73_3578 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_4 FILLER_74_175 ();
 sg13g2_fill_2 FILLER_74_179 ();
 sg13g2_decap_8 FILLER_74_185 ();
 sg13g2_decap_8 FILLER_74_192 ();
 sg13g2_decap_8 FILLER_74_199 ();
 sg13g2_fill_1 FILLER_74_206 ();
 sg13g2_fill_2 FILLER_74_233 ();
 sg13g2_fill_1 FILLER_74_266 ();
 sg13g2_fill_1 FILLER_74_327 ();
 sg13g2_fill_1 FILLER_74_339 ();
 sg13g2_decap_4 FILLER_74_386 ();
 sg13g2_fill_1 FILLER_74_427 ();
 sg13g2_decap_4 FILLER_74_447 ();
 sg13g2_fill_1 FILLER_74_451 ();
 sg13g2_fill_2 FILLER_74_459 ();
 sg13g2_decap_8 FILLER_74_477 ();
 sg13g2_fill_2 FILLER_74_484 ();
 sg13g2_fill_1 FILLER_74_486 ();
 sg13g2_decap_4 FILLER_74_512 ();
 sg13g2_decap_8 FILLER_74_526 ();
 sg13g2_decap_4 FILLER_74_533 ();
 sg13g2_fill_2 FILLER_74_537 ();
 sg13g2_fill_2 FILLER_74_556 ();
 sg13g2_fill_1 FILLER_74_558 ();
 sg13g2_decap_4 FILLER_74_584 ();
 sg13g2_fill_1 FILLER_74_588 ();
 sg13g2_fill_1 FILLER_74_598 ();
 sg13g2_fill_1 FILLER_74_611 ();
 sg13g2_fill_2 FILLER_74_617 ();
 sg13g2_fill_1 FILLER_74_619 ();
 sg13g2_decap_8 FILLER_74_639 ();
 sg13g2_decap_8 FILLER_74_646 ();
 sg13g2_fill_2 FILLER_74_653 ();
 sg13g2_fill_2 FILLER_74_660 ();
 sg13g2_fill_1 FILLER_74_662 ();
 sg13g2_decap_4 FILLER_74_687 ();
 sg13g2_fill_2 FILLER_74_710 ();
 sg13g2_fill_1 FILLER_74_712 ();
 sg13g2_decap_8 FILLER_74_741 ();
 sg13g2_decap_4 FILLER_74_748 ();
 sg13g2_fill_2 FILLER_74_752 ();
 sg13g2_fill_1 FILLER_74_765 ();
 sg13g2_fill_1 FILLER_74_769 ();
 sg13g2_decap_4 FILLER_74_795 ();
 sg13g2_fill_2 FILLER_74_799 ();
 sg13g2_fill_1 FILLER_74_805 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_fill_2 FILLER_74_818 ();
 sg13g2_fill_1 FILLER_74_820 ();
 sg13g2_decap_4 FILLER_74_847 ();
 sg13g2_fill_2 FILLER_74_864 ();
 sg13g2_fill_2 FILLER_74_884 ();
 sg13g2_fill_1 FILLER_74_886 ();
 sg13g2_fill_2 FILLER_74_924 ();
 sg13g2_fill_1 FILLER_74_926 ();
 sg13g2_fill_1 FILLER_74_932 ();
 sg13g2_fill_2 FILLER_74_938 ();
 sg13g2_decap_4 FILLER_74_951 ();
 sg13g2_fill_2 FILLER_74_955 ();
 sg13g2_fill_2 FILLER_74_974 ();
 sg13g2_fill_1 FILLER_74_1000 ();
 sg13g2_decap_8 FILLER_74_1011 ();
 sg13g2_decap_8 FILLER_74_1043 ();
 sg13g2_decap_8 FILLER_74_1050 ();
 sg13g2_decap_8 FILLER_74_1066 ();
 sg13g2_decap_4 FILLER_74_1073 ();
 sg13g2_fill_1 FILLER_74_1077 ();
 sg13g2_fill_2 FILLER_74_1104 ();
 sg13g2_fill_1 FILLER_74_1106 ();
 sg13g2_decap_8 FILLER_74_1112 ();
 sg13g2_decap_4 FILLER_74_1127 ();
 sg13g2_fill_1 FILLER_74_1131 ();
 sg13g2_decap_4 FILLER_74_1137 ();
 sg13g2_decap_4 FILLER_74_1163 ();
 sg13g2_fill_2 FILLER_74_1185 ();
 sg13g2_fill_1 FILLER_74_1187 ();
 sg13g2_decap_4 FILLER_74_1200 ();
 sg13g2_fill_1 FILLER_74_1221 ();
 sg13g2_decap_8 FILLER_74_1233 ();
 sg13g2_fill_1 FILLER_74_1240 ();
 sg13g2_fill_2 FILLER_74_1249 ();
 sg13g2_fill_1 FILLER_74_1251 ();
 sg13g2_fill_1 FILLER_74_1265 ();
 sg13g2_decap_8 FILLER_74_1291 ();
 sg13g2_decap_4 FILLER_74_1298 ();
 sg13g2_fill_2 FILLER_74_1302 ();
 sg13g2_fill_1 FILLER_74_1323 ();
 sg13g2_decap_8 FILLER_74_1328 ();
 sg13g2_fill_2 FILLER_74_1335 ();
 sg13g2_fill_1 FILLER_74_1337 ();
 sg13g2_decap_8 FILLER_74_1344 ();
 sg13g2_decap_8 FILLER_74_1351 ();
 sg13g2_decap_8 FILLER_74_1358 ();
 sg13g2_decap_4 FILLER_74_1365 ();
 sg13g2_fill_1 FILLER_74_1381 ();
 sg13g2_decap_8 FILLER_74_1389 ();
 sg13g2_fill_2 FILLER_74_1396 ();
 sg13g2_decap_4 FILLER_74_1412 ();
 sg13g2_fill_2 FILLER_74_1419 ();
 sg13g2_decap_8 FILLER_74_1445 ();
 sg13g2_fill_2 FILLER_74_1452 ();
 sg13g2_fill_1 FILLER_74_1454 ();
 sg13g2_fill_2 FILLER_74_1468 ();
 sg13g2_fill_1 FILLER_74_1470 ();
 sg13g2_fill_1 FILLER_74_1481 ();
 sg13g2_fill_1 FILLER_74_1491 ();
 sg13g2_fill_2 FILLER_74_1497 ();
 sg13g2_fill_1 FILLER_74_1499 ();
 sg13g2_decap_4 FILLER_74_1517 ();
 sg13g2_fill_1 FILLER_74_1521 ();
 sg13g2_fill_1 FILLER_74_1542 ();
 sg13g2_decap_4 FILLER_74_1550 ();
 sg13g2_fill_1 FILLER_74_1554 ();
 sg13g2_fill_1 FILLER_74_1573 ();
 sg13g2_decap_4 FILLER_74_1594 ();
 sg13g2_decap_8 FILLER_74_1603 ();
 sg13g2_fill_1 FILLER_74_1610 ();
 sg13g2_decap_8 FILLER_74_1628 ();
 sg13g2_decap_4 FILLER_74_1639 ();
 sg13g2_fill_1 FILLER_74_1648 ();
 sg13g2_fill_2 FILLER_74_1662 ();
 sg13g2_fill_1 FILLER_74_1664 ();
 sg13g2_decap_8 FILLER_74_1695 ();
 sg13g2_decap_4 FILLER_74_1702 ();
 sg13g2_fill_2 FILLER_74_1715 ();
 sg13g2_fill_2 FILLER_74_1724 ();
 sg13g2_fill_1 FILLER_74_1726 ();
 sg13g2_fill_1 FILLER_74_1739 ();
 sg13g2_fill_2 FILLER_74_1755 ();
 sg13g2_fill_2 FILLER_74_1765 ();
 sg13g2_fill_2 FILLER_74_1805 ();
 sg13g2_decap_4 FILLER_74_1818 ();
 sg13g2_decap_4 FILLER_74_1846 ();
 sg13g2_decap_8 FILLER_74_1879 ();
 sg13g2_fill_2 FILLER_74_1886 ();
 sg13g2_fill_1 FILLER_74_1888 ();
 sg13g2_decap_8 FILLER_74_1902 ();
 sg13g2_decap_8 FILLER_74_1909 ();
 sg13g2_fill_2 FILLER_74_1941 ();
 sg13g2_fill_2 FILLER_74_1955 ();
 sg13g2_fill_1 FILLER_74_1957 ();
 sg13g2_decap_4 FILLER_74_1968 ();
 sg13g2_fill_2 FILLER_74_1972 ();
 sg13g2_fill_1 FILLER_74_1979 ();
 sg13g2_decap_4 FILLER_74_1988 ();
 sg13g2_fill_1 FILLER_74_1992 ();
 sg13g2_decap_8 FILLER_74_2005 ();
 sg13g2_fill_1 FILLER_74_2012 ();
 sg13g2_fill_2 FILLER_74_2052 ();
 sg13g2_fill_2 FILLER_74_2064 ();
 sg13g2_fill_1 FILLER_74_2066 ();
 sg13g2_fill_1 FILLER_74_2085 ();
 sg13g2_fill_1 FILLER_74_2102 ();
 sg13g2_fill_2 FILLER_74_2115 ();
 sg13g2_fill_1 FILLER_74_2117 ();
 sg13g2_fill_1 FILLER_74_2130 ();
 sg13g2_fill_2 FILLER_74_2144 ();
 sg13g2_decap_8 FILLER_74_2158 ();
 sg13g2_decap_8 FILLER_74_2165 ();
 sg13g2_decap_4 FILLER_74_2172 ();
 sg13g2_decap_8 FILLER_74_2183 ();
 sg13g2_decap_4 FILLER_74_2190 ();
 sg13g2_fill_1 FILLER_74_2194 ();
 sg13g2_fill_1 FILLER_74_2207 ();
 sg13g2_decap_4 FILLER_74_2213 ();
 sg13g2_fill_1 FILLER_74_2217 ();
 sg13g2_decap_8 FILLER_74_2231 ();
 sg13g2_fill_1 FILLER_74_2238 ();
 sg13g2_decap_4 FILLER_74_2251 ();
 sg13g2_decap_8 FILLER_74_2266 ();
 sg13g2_fill_2 FILLER_74_2273 ();
 sg13g2_fill_1 FILLER_74_2275 ();
 sg13g2_decap_8 FILLER_74_2282 ();
 sg13g2_decap_8 FILLER_74_2289 ();
 sg13g2_fill_2 FILLER_74_2296 ();
 sg13g2_fill_1 FILLER_74_2298 ();
 sg13g2_fill_1 FILLER_74_2304 ();
 sg13g2_fill_1 FILLER_74_2310 ();
 sg13g2_decap_4 FILLER_74_2316 ();
 sg13g2_fill_2 FILLER_74_2320 ();
 sg13g2_decap_8 FILLER_74_2338 ();
 sg13g2_decap_4 FILLER_74_2345 ();
 sg13g2_fill_2 FILLER_74_2349 ();
 sg13g2_decap_8 FILLER_74_2364 ();
 sg13g2_decap_8 FILLER_74_2371 ();
 sg13g2_decap_4 FILLER_74_2378 ();
 sg13g2_fill_2 FILLER_74_2392 ();
 sg13g2_decap_8 FILLER_74_2398 ();
 sg13g2_decap_8 FILLER_74_2405 ();
 sg13g2_fill_1 FILLER_74_2425 ();
 sg13g2_decap_4 FILLER_74_2450 ();
 sg13g2_fill_1 FILLER_74_2454 ();
 sg13g2_decap_8 FILLER_74_2472 ();
 sg13g2_fill_2 FILLER_74_2487 ();
 sg13g2_fill_1 FILLER_74_2494 ();
 sg13g2_decap_4 FILLER_74_2500 ();
 sg13g2_fill_1 FILLER_74_2504 ();
 sg13g2_fill_2 FILLER_74_2509 ();
 sg13g2_decap_8 FILLER_74_2516 ();
 sg13g2_decap_4 FILLER_74_2523 ();
 sg13g2_decap_8 FILLER_74_2542 ();
 sg13g2_fill_2 FILLER_74_2549 ();
 sg13g2_fill_1 FILLER_74_2551 ();
 sg13g2_fill_2 FILLER_74_2580 ();
 sg13g2_decap_8 FILLER_74_2601 ();
 sg13g2_fill_1 FILLER_74_2608 ();
 sg13g2_fill_2 FILLER_74_2645 ();
 sg13g2_decap_4 FILLER_74_2667 ();
 sg13g2_fill_2 FILLER_74_2671 ();
 sg13g2_fill_1 FILLER_74_2678 ();
 sg13g2_fill_1 FILLER_74_2683 ();
 sg13g2_decap_8 FILLER_74_2692 ();
 sg13g2_decap_4 FILLER_74_2699 ();
 sg13g2_fill_2 FILLER_74_2703 ();
 sg13g2_fill_2 FILLER_74_2728 ();
 sg13g2_fill_2 FILLER_74_2749 ();
 sg13g2_fill_1 FILLER_74_2751 ();
 sg13g2_decap_8 FILLER_74_2761 ();
 sg13g2_decap_4 FILLER_74_2768 ();
 sg13g2_fill_2 FILLER_74_2772 ();
 sg13g2_decap_8 FILLER_74_2797 ();
 sg13g2_decap_8 FILLER_74_2804 ();
 sg13g2_fill_2 FILLER_74_2811 ();
 sg13g2_fill_2 FILLER_74_2826 ();
 sg13g2_decap_8 FILLER_74_2842 ();
 sg13g2_decap_8 FILLER_74_2849 ();
 sg13g2_decap_8 FILLER_74_2856 ();
 sg13g2_decap_4 FILLER_74_2894 ();
 sg13g2_fill_1 FILLER_74_2898 ();
 sg13g2_fill_1 FILLER_74_2910 ();
 sg13g2_fill_2 FILLER_74_2945 ();
 sg13g2_fill_1 FILLER_74_2947 ();
 sg13g2_decap_4 FILLER_74_2953 ();
 sg13g2_decap_4 FILLER_74_2974 ();
 sg13g2_decap_8 FILLER_74_2990 ();
 sg13g2_fill_2 FILLER_74_2997 ();
 sg13g2_fill_1 FILLER_74_2999 ();
 sg13g2_fill_1 FILLER_74_3010 ();
 sg13g2_decap_8 FILLER_74_3054 ();
 sg13g2_fill_2 FILLER_74_3061 ();
 sg13g2_fill_1 FILLER_74_3063 ();
 sg13g2_fill_1 FILLER_74_3088 ();
 sg13g2_decap_4 FILLER_74_3097 ();
 sg13g2_decap_8 FILLER_74_3123 ();
 sg13g2_decap_8 FILLER_74_3134 ();
 sg13g2_fill_1 FILLER_74_3141 ();
 sg13g2_fill_2 FILLER_74_3148 ();
 sg13g2_decap_4 FILLER_74_3174 ();
 sg13g2_fill_2 FILLER_74_3178 ();
 sg13g2_fill_1 FILLER_74_3190 ();
 sg13g2_decap_8 FILLER_74_3200 ();
 sg13g2_fill_1 FILLER_74_3207 ();
 sg13g2_decap_8 FILLER_74_3225 ();
 sg13g2_fill_2 FILLER_74_3232 ();
 sg13g2_fill_1 FILLER_74_3234 ();
 sg13g2_decap_8 FILLER_74_3243 ();
 sg13g2_decap_4 FILLER_74_3250 ();
 sg13g2_fill_1 FILLER_74_3254 ();
 sg13g2_fill_2 FILLER_74_3265 ();
 sg13g2_fill_2 FILLER_74_3276 ();
 sg13g2_fill_1 FILLER_74_3278 ();
 sg13g2_fill_1 FILLER_74_3314 ();
 sg13g2_decap_4 FILLER_74_3324 ();
 sg13g2_fill_1 FILLER_74_3328 ();
 sg13g2_fill_2 FILLER_74_3369 ();
 sg13g2_decap_8 FILLER_74_3384 ();
 sg13g2_decap_4 FILLER_74_3391 ();
 sg13g2_fill_1 FILLER_74_3395 ();
 sg13g2_decap_8 FILLER_74_3400 ();
 sg13g2_decap_8 FILLER_74_3407 ();
 sg13g2_decap_8 FILLER_74_3414 ();
 sg13g2_decap_8 FILLER_74_3421 ();
 sg13g2_decap_8 FILLER_74_3428 ();
 sg13g2_decap_8 FILLER_74_3435 ();
 sg13g2_decap_8 FILLER_74_3442 ();
 sg13g2_decap_8 FILLER_74_3449 ();
 sg13g2_decap_8 FILLER_74_3456 ();
 sg13g2_decap_8 FILLER_74_3463 ();
 sg13g2_decap_8 FILLER_74_3470 ();
 sg13g2_decap_8 FILLER_74_3477 ();
 sg13g2_decap_8 FILLER_74_3484 ();
 sg13g2_decap_8 FILLER_74_3491 ();
 sg13g2_decap_8 FILLER_74_3498 ();
 sg13g2_decap_8 FILLER_74_3505 ();
 sg13g2_decap_8 FILLER_74_3512 ();
 sg13g2_decap_8 FILLER_74_3519 ();
 sg13g2_decap_8 FILLER_74_3526 ();
 sg13g2_decap_8 FILLER_74_3533 ();
 sg13g2_decap_8 FILLER_74_3540 ();
 sg13g2_decap_8 FILLER_74_3547 ();
 sg13g2_decap_8 FILLER_74_3554 ();
 sg13g2_decap_8 FILLER_74_3561 ();
 sg13g2_decap_8 FILLER_74_3568 ();
 sg13g2_decap_4 FILLER_74_3575 ();
 sg13g2_fill_1 FILLER_74_3579 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_4 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_230 ();
 sg13g2_decap_8 FILLER_75_237 ();
 sg13g2_decap_8 FILLER_75_244 ();
 sg13g2_decap_8 FILLER_75_251 ();
 sg13g2_decap_8 FILLER_75_258 ();
 sg13g2_fill_2 FILLER_75_265 ();
 sg13g2_fill_2 FILLER_75_276 ();
 sg13g2_fill_1 FILLER_75_278 ();
 sg13g2_fill_1 FILLER_75_297 ();
 sg13g2_fill_1 FILLER_75_320 ();
 sg13g2_fill_2 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_340 ();
 sg13g2_fill_2 FILLER_75_354 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_fill_1 FILLER_75_398 ();
 sg13g2_fill_1 FILLER_75_427 ();
 sg13g2_decap_8 FILLER_75_480 ();
 sg13g2_fill_2 FILLER_75_487 ();
 sg13g2_fill_1 FILLER_75_489 ();
 sg13g2_fill_2 FILLER_75_503 ();
 sg13g2_fill_1 FILLER_75_505 ();
 sg13g2_decap_4 FILLER_75_518 ();
 sg13g2_fill_2 FILLER_75_522 ();
 sg13g2_decap_4 FILLER_75_533 ();
 sg13g2_fill_1 FILLER_75_537 ();
 sg13g2_fill_2 FILLER_75_559 ();
 sg13g2_decap_8 FILLER_75_565 ();
 sg13g2_decap_8 FILLER_75_584 ();
 sg13g2_fill_2 FILLER_75_606 ();
 sg13g2_decap_8 FILLER_75_618 ();
 sg13g2_decap_8 FILLER_75_625 ();
 sg13g2_fill_1 FILLER_75_632 ();
 sg13g2_fill_2 FILLER_75_637 ();
 sg13g2_fill_1 FILLER_75_647 ();
 sg13g2_decap_4 FILLER_75_663 ();
 sg13g2_fill_1 FILLER_75_667 ();
 sg13g2_fill_2 FILLER_75_690 ();
 sg13g2_decap_8 FILLER_75_707 ();
 sg13g2_decap_8 FILLER_75_714 ();
 sg13g2_decap_4 FILLER_75_721 ();
 sg13g2_fill_1 FILLER_75_725 ();
 sg13g2_fill_2 FILLER_75_730 ();
 sg13g2_fill_1 FILLER_75_732 ();
 sg13g2_decap_8 FILLER_75_739 ();
 sg13g2_decap_4 FILLER_75_746 ();
 sg13g2_fill_2 FILLER_75_769 ();
 sg13g2_decap_4 FILLER_75_790 ();
 sg13g2_fill_2 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_814 ();
 sg13g2_decap_4 FILLER_75_821 ();
 sg13g2_fill_1 FILLER_75_825 ();
 sg13g2_fill_1 FILLER_75_831 ();
 sg13g2_decap_4 FILLER_75_840 ();
 sg13g2_fill_2 FILLER_75_844 ();
 sg13g2_fill_1 FILLER_75_854 ();
 sg13g2_fill_2 FILLER_75_867 ();
 sg13g2_fill_1 FILLER_75_869 ();
 sg13g2_decap_8 FILLER_75_878 ();
 sg13g2_decap_8 FILLER_75_885 ();
 sg13g2_decap_4 FILLER_75_896 ();
 sg13g2_fill_2 FILLER_75_900 ();
 sg13g2_fill_1 FILLER_75_905 ();
 sg13g2_fill_2 FILLER_75_912 ();
 sg13g2_fill_1 FILLER_75_914 ();
 sg13g2_fill_2 FILLER_75_930 ();
 sg13g2_fill_1 FILLER_75_932 ();
 sg13g2_decap_4 FILLER_75_955 ();
 sg13g2_fill_2 FILLER_75_964 ();
 sg13g2_decap_4 FILLER_75_971 ();
 sg13g2_decap_8 FILLER_75_980 ();
 sg13g2_fill_2 FILLER_75_1001 ();
 sg13g2_fill_2 FILLER_75_1015 ();
 sg13g2_fill_1 FILLER_75_1017 ();
 sg13g2_decap_4 FILLER_75_1039 ();
 sg13g2_fill_2 FILLER_75_1043 ();
 sg13g2_fill_2 FILLER_75_1073 ();
 sg13g2_fill_2 FILLER_75_1119 ();
 sg13g2_decap_8 FILLER_75_1134 ();
 sg13g2_decap_8 FILLER_75_1141 ();
 sg13g2_decap_8 FILLER_75_1148 ();
 sg13g2_fill_1 FILLER_75_1155 ();
 sg13g2_fill_2 FILLER_75_1176 ();
 sg13g2_fill_2 FILLER_75_1196 ();
 sg13g2_decap_4 FILLER_75_1216 ();
 sg13g2_decap_8 FILLER_75_1235 ();
 sg13g2_decap_8 FILLER_75_1242 ();
 sg13g2_fill_1 FILLER_75_1249 ();
 sg13g2_fill_1 FILLER_75_1263 ();
 sg13g2_decap_8 FILLER_75_1271 ();
 sg13g2_decap_4 FILLER_75_1278 ();
 sg13g2_decap_4 FILLER_75_1286 ();
 sg13g2_decap_4 FILLER_75_1302 ();
 sg13g2_fill_1 FILLER_75_1306 ();
 sg13g2_fill_2 FILLER_75_1310 ();
 sg13g2_fill_2 FILLER_75_1316 ();
 sg13g2_decap_4 FILLER_75_1331 ();
 sg13g2_fill_2 FILLER_75_1353 ();
 sg13g2_fill_2 FILLER_75_1360 ();
 sg13g2_fill_2 FILLER_75_1367 ();
 sg13g2_decap_8 FILLER_75_1380 ();
 sg13g2_decap_8 FILLER_75_1387 ();
 sg13g2_fill_2 FILLER_75_1394 ();
 sg13g2_fill_1 FILLER_75_1406 ();
 sg13g2_decap_8 FILLER_75_1411 ();
 sg13g2_decap_4 FILLER_75_1418 ();
 sg13g2_decap_8 FILLER_75_1441 ();
 sg13g2_fill_2 FILLER_75_1448 ();
 sg13g2_fill_2 FILLER_75_1478 ();
 sg13g2_fill_1 FILLER_75_1493 ();
 sg13g2_decap_8 FILLER_75_1509 ();
 sg13g2_decap_4 FILLER_75_1516 ();
 sg13g2_decap_4 FILLER_75_1534 ();
 sg13g2_decap_4 FILLER_75_1543 ();
 sg13g2_fill_1 FILLER_75_1547 ();
 sg13g2_fill_1 FILLER_75_1556 ();
 sg13g2_fill_2 FILLER_75_1590 ();
 sg13g2_decap_8 FILLER_75_1597 ();
 sg13g2_decap_8 FILLER_75_1604 ();
 sg13g2_fill_1 FILLER_75_1611 ();
 sg13g2_fill_2 FILLER_75_1625 ();
 sg13g2_fill_2 FILLER_75_1632 ();
 sg13g2_fill_1 FILLER_75_1642 ();
 sg13g2_decap_8 FILLER_75_1656 ();
 sg13g2_decap_8 FILLER_75_1663 ();
 sg13g2_fill_1 FILLER_75_1670 ();
 sg13g2_fill_2 FILLER_75_1686 ();
 sg13g2_fill_1 FILLER_75_1688 ();
 sg13g2_decap_8 FILLER_75_1729 ();
 sg13g2_decap_4 FILLER_75_1736 ();
 sg13g2_fill_1 FILLER_75_1740 ();
 sg13g2_fill_1 FILLER_75_1750 ();
 sg13g2_decap_8 FILLER_75_1758 ();
 sg13g2_decap_8 FILLER_75_1765 ();
 sg13g2_decap_4 FILLER_75_1772 ();
 sg13g2_fill_1 FILLER_75_1776 ();
 sg13g2_fill_1 FILLER_75_1782 ();
 sg13g2_decap_8 FILLER_75_1787 ();
 sg13g2_decap_4 FILLER_75_1794 ();
 sg13g2_fill_2 FILLER_75_1818 ();
 sg13g2_fill_1 FILLER_75_1820 ();
 sg13g2_decap_8 FILLER_75_1839 ();
 sg13g2_fill_2 FILLER_75_1846 ();
 sg13g2_fill_1 FILLER_75_1848 ();
 sg13g2_fill_1 FILLER_75_1858 ();
 sg13g2_decap_4 FILLER_75_1868 ();
 sg13g2_fill_2 FILLER_75_1872 ();
 sg13g2_decap_4 FILLER_75_1889 ();
 sg13g2_fill_2 FILLER_75_1893 ();
 sg13g2_fill_2 FILLER_75_1899 ();
 sg13g2_fill_1 FILLER_75_1901 ();
 sg13g2_fill_2 FILLER_75_1917 ();
 sg13g2_fill_1 FILLER_75_1923 ();
 sg13g2_decap_8 FILLER_75_1942 ();
 sg13g2_fill_2 FILLER_75_1974 ();
 sg13g2_fill_1 FILLER_75_1976 ();
 sg13g2_decap_8 FILLER_75_1998 ();
 sg13g2_decap_4 FILLER_75_2005 ();
 sg13g2_fill_2 FILLER_75_2009 ();
 sg13g2_fill_1 FILLER_75_2016 ();
 sg13g2_decap_4 FILLER_75_2050 ();
 sg13g2_decap_8 FILLER_75_2061 ();
 sg13g2_decap_8 FILLER_75_2068 ();
 sg13g2_fill_2 FILLER_75_2075 ();
 sg13g2_fill_1 FILLER_75_2077 ();
 sg13g2_fill_2 FILLER_75_2083 ();
 sg13g2_decap_8 FILLER_75_2092 ();
 sg13g2_decap_8 FILLER_75_2099 ();
 sg13g2_fill_2 FILLER_75_2106 ();
 sg13g2_decap_8 FILLER_75_2116 ();
 sg13g2_fill_2 FILLER_75_2123 ();
 sg13g2_fill_1 FILLER_75_2125 ();
 sg13g2_decap_8 FILLER_75_2141 ();
 sg13g2_decap_4 FILLER_75_2161 ();
 sg13g2_decap_8 FILLER_75_2183 ();
 sg13g2_fill_2 FILLER_75_2217 ();
 sg13g2_fill_1 FILLER_75_2219 ();
 sg13g2_fill_1 FILLER_75_2231 ();
 sg13g2_decap_8 FILLER_75_2243 ();
 sg13g2_decap_8 FILLER_75_2250 ();
 sg13g2_fill_2 FILLER_75_2257 ();
 sg13g2_fill_1 FILLER_75_2259 ();
 sg13g2_decap_8 FILLER_75_2264 ();
 sg13g2_fill_2 FILLER_75_2280 ();
 sg13g2_fill_1 FILLER_75_2285 ();
 sg13g2_fill_2 FILLER_75_2290 ();
 sg13g2_fill_1 FILLER_75_2292 ();
 sg13g2_decap_8 FILLER_75_2342 ();
 sg13g2_decap_8 FILLER_75_2362 ();
 sg13g2_decap_4 FILLER_75_2369 ();
 sg13g2_fill_2 FILLER_75_2373 ();
 sg13g2_fill_2 FILLER_75_2384 ();
 sg13g2_decap_4 FILLER_75_2398 ();
 sg13g2_decap_4 FILLER_75_2423 ();
 sg13g2_decap_8 FILLER_75_2449 ();
 sg13g2_fill_1 FILLER_75_2460 ();
 sg13g2_decap_8 FILLER_75_2471 ();
 sg13g2_fill_1 FILLER_75_2478 ();
 sg13g2_fill_2 FILLER_75_2502 ();
 sg13g2_fill_1 FILLER_75_2504 ();
 sg13g2_decap_4 FILLER_75_2540 ();
 sg13g2_fill_1 FILLER_75_2544 ();
 sg13g2_decap_4 FILLER_75_2553 ();
 sg13g2_decap_8 FILLER_75_2561 ();
 sg13g2_decap_8 FILLER_75_2568 ();
 sg13g2_fill_2 FILLER_75_2582 ();
 sg13g2_fill_1 FILLER_75_2584 ();
 sg13g2_fill_1 FILLER_75_2605 ();
 sg13g2_decap_4 FILLER_75_2610 ();
 sg13g2_decap_4 FILLER_75_2618 ();
 sg13g2_decap_8 FILLER_75_2645 ();
 sg13g2_decap_8 FILLER_75_2666 ();
 sg13g2_decap_8 FILLER_75_2673 ();
 sg13g2_fill_1 FILLER_75_2680 ();
 sg13g2_decap_4 FILLER_75_2696 ();
 sg13g2_fill_2 FILLER_75_2706 ();
 sg13g2_fill_2 FILLER_75_2724 ();
 sg13g2_fill_1 FILLER_75_2726 ();
 sg13g2_decap_8 FILLER_75_2744 ();
 sg13g2_decap_8 FILLER_75_2751 ();
 sg13g2_fill_1 FILLER_75_2758 ();
 sg13g2_fill_2 FILLER_75_2764 ();
 sg13g2_decap_8 FILLER_75_2775 ();
 sg13g2_fill_2 FILLER_75_2782 ();
 sg13g2_fill_2 FILLER_75_2799 ();
 sg13g2_fill_1 FILLER_75_2801 ();
 sg13g2_fill_2 FILLER_75_2842 ();
 sg13g2_fill_1 FILLER_75_2844 ();
 sg13g2_decap_8 FILLER_75_2849 ();
 sg13g2_decap_8 FILLER_75_2856 ();
 sg13g2_fill_2 FILLER_75_2900 ();
 sg13g2_fill_1 FILLER_75_2910 ();
 sg13g2_decap_8 FILLER_75_2948 ();
 sg13g2_decap_8 FILLER_75_2955 ();
 sg13g2_fill_2 FILLER_75_2962 ();
 sg13g2_fill_2 FILLER_75_2973 ();
 sg13g2_fill_1 FILLER_75_2975 ();
 sg13g2_fill_2 FILLER_75_3001 ();
 sg13g2_decap_8 FILLER_75_3034 ();
 sg13g2_fill_2 FILLER_75_3041 ();
 sg13g2_decap_8 FILLER_75_3059 ();
 sg13g2_fill_2 FILLER_75_3066 ();
 sg13g2_decap_8 FILLER_75_3080 ();
 sg13g2_decap_4 FILLER_75_3087 ();
 sg13g2_fill_2 FILLER_75_3091 ();
 sg13g2_decap_4 FILLER_75_3098 ();
 sg13g2_fill_2 FILLER_75_3102 ();
 sg13g2_fill_1 FILLER_75_3113 ();
 sg13g2_decap_8 FILLER_75_3126 ();
 sg13g2_decap_8 FILLER_75_3133 ();
 sg13g2_decap_4 FILLER_75_3140 ();
 sg13g2_fill_2 FILLER_75_3144 ();
 sg13g2_decap_8 FILLER_75_3168 ();
 sg13g2_decap_4 FILLER_75_3175 ();
 sg13g2_fill_1 FILLER_75_3179 ();
 sg13g2_fill_2 FILLER_75_3200 ();
 sg13g2_fill_1 FILLER_75_3202 ();
 sg13g2_decap_4 FILLER_75_3208 ();
 sg13g2_fill_1 FILLER_75_3212 ();
 sg13g2_fill_2 FILLER_75_3231 ();
 sg13g2_decap_8 FILLER_75_3274 ();
 sg13g2_decap_8 FILLER_75_3281 ();
 sg13g2_decap_8 FILLER_75_3288 ();
 sg13g2_decap_4 FILLER_75_3295 ();
 sg13g2_fill_1 FILLER_75_3299 ();
 sg13g2_fill_2 FILLER_75_3313 ();
 sg13g2_decap_8 FILLER_75_3387 ();
 sg13g2_decap_8 FILLER_75_3394 ();
 sg13g2_decap_8 FILLER_75_3401 ();
 sg13g2_decap_8 FILLER_75_3408 ();
 sg13g2_decap_8 FILLER_75_3415 ();
 sg13g2_decap_8 FILLER_75_3422 ();
 sg13g2_decap_8 FILLER_75_3429 ();
 sg13g2_decap_8 FILLER_75_3436 ();
 sg13g2_decap_8 FILLER_75_3443 ();
 sg13g2_decap_8 FILLER_75_3450 ();
 sg13g2_decap_8 FILLER_75_3457 ();
 sg13g2_decap_8 FILLER_75_3464 ();
 sg13g2_decap_8 FILLER_75_3471 ();
 sg13g2_decap_8 FILLER_75_3478 ();
 sg13g2_decap_8 FILLER_75_3485 ();
 sg13g2_decap_8 FILLER_75_3492 ();
 sg13g2_decap_8 FILLER_75_3499 ();
 sg13g2_decap_8 FILLER_75_3506 ();
 sg13g2_decap_8 FILLER_75_3513 ();
 sg13g2_decap_8 FILLER_75_3520 ();
 sg13g2_decap_8 FILLER_75_3527 ();
 sg13g2_decap_8 FILLER_75_3534 ();
 sg13g2_decap_8 FILLER_75_3541 ();
 sg13g2_decap_8 FILLER_75_3548 ();
 sg13g2_decap_8 FILLER_75_3555 ();
 sg13g2_decap_8 FILLER_75_3562 ();
 sg13g2_decap_8 FILLER_75_3569 ();
 sg13g2_decap_4 FILLER_75_3576 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_fill_1 FILLER_76_231 ();
 sg13g2_decap_4 FILLER_76_266 ();
 sg13g2_fill_1 FILLER_76_281 ();
 sg13g2_fill_1 FILLER_76_310 ();
 sg13g2_fill_1 FILLER_76_354 ();
 sg13g2_fill_2 FILLER_76_361 ();
 sg13g2_decap_4 FILLER_76_405 ();
 sg13g2_fill_2 FILLER_76_409 ();
 sg13g2_decap_8 FILLER_76_417 ();
 sg13g2_fill_2 FILLER_76_424 ();
 sg13g2_fill_1 FILLER_76_426 ();
 sg13g2_fill_1 FILLER_76_455 ();
 sg13g2_fill_2 FILLER_76_465 ();
 sg13g2_fill_2 FILLER_76_503 ();
 sg13g2_decap_8 FILLER_76_510 ();
 sg13g2_decap_4 FILLER_76_530 ();
 sg13g2_fill_2 FILLER_76_556 ();
 sg13g2_decap_4 FILLER_76_571 ();
 sg13g2_decap_4 FILLER_76_585 ();
 sg13g2_fill_2 FILLER_76_589 ();
 sg13g2_decap_8 FILLER_76_619 ();
 sg13g2_decap_4 FILLER_76_643 ();
 sg13g2_fill_1 FILLER_76_647 ();
 sg13g2_decap_8 FILLER_76_658 ();
 sg13g2_fill_2 FILLER_76_665 ();
 sg13g2_fill_1 FILLER_76_667 ();
 sg13g2_decap_4 FILLER_76_676 ();
 sg13g2_decap_4 FILLER_76_688 ();
 sg13g2_fill_1 FILLER_76_692 ();
 sg13g2_decap_8 FILLER_76_702 ();
 sg13g2_fill_2 FILLER_76_709 ();
 sg13g2_fill_1 FILLER_76_711 ();
 sg13g2_decap_4 FILLER_76_716 ();
 sg13g2_fill_1 FILLER_76_720 ();
 sg13g2_fill_2 FILLER_76_753 ();
 sg13g2_fill_1 FILLER_76_755 ();
 sg13g2_fill_2 FILLER_76_769 ();
 sg13g2_decap_4 FILLER_76_778 ();
 sg13g2_decap_4 FILLER_76_792 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_decap_4 FILLER_76_819 ();
 sg13g2_fill_2 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_846 ();
 sg13g2_fill_2 FILLER_76_853 ();
 sg13g2_fill_1 FILLER_76_855 ();
 sg13g2_decap_8 FILLER_76_861 ();
 sg13g2_decap_4 FILLER_76_868 ();
 sg13g2_fill_2 FILLER_76_872 ();
 sg13g2_fill_2 FILLER_76_902 ();
 sg13g2_fill_2 FILLER_76_918 ();
 sg13g2_fill_1 FILLER_76_920 ();
 sg13g2_decap_4 FILLER_76_947 ();
 sg13g2_decap_4 FILLER_76_973 ();
 sg13g2_decap_8 FILLER_76_1007 ();
 sg13g2_decap_4 FILLER_76_1014 ();
 sg13g2_fill_2 FILLER_76_1018 ();
 sg13g2_decap_4 FILLER_76_1058 ();
 sg13g2_fill_1 FILLER_76_1062 ();
 sg13g2_fill_2 FILLER_76_1079 ();
 sg13g2_decap_8 FILLER_76_1100 ();
 sg13g2_fill_2 FILLER_76_1107 ();
 sg13g2_fill_1 FILLER_76_1109 ();
 sg13g2_decap_4 FILLER_76_1117 ();
 sg13g2_fill_2 FILLER_76_1133 ();
 sg13g2_fill_2 FILLER_76_1158 ();
 sg13g2_decap_8 FILLER_76_1165 ();
 sg13g2_fill_1 FILLER_76_1172 ();
 sg13g2_decap_8 FILLER_76_1176 ();
 sg13g2_fill_2 FILLER_76_1183 ();
 sg13g2_fill_1 FILLER_76_1185 ();
 sg13g2_decap_8 FILLER_76_1194 ();
 sg13g2_decap_8 FILLER_76_1201 ();
 sg13g2_decap_8 FILLER_76_1225 ();
 sg13g2_decap_8 FILLER_76_1232 ();
 sg13g2_fill_1 FILLER_76_1264 ();
 sg13g2_fill_2 FILLER_76_1306 ();
 sg13g2_fill_2 FILLER_76_1326 ();
 sg13g2_fill_1 FILLER_76_1350 ();
 sg13g2_fill_2 FILLER_76_1360 ();
 sg13g2_decap_4 FILLER_76_1385 ();
 sg13g2_fill_1 FILLER_76_1389 ();
 sg13g2_decap_8 FILLER_76_1416 ();
 sg13g2_decap_8 FILLER_76_1444 ();
 sg13g2_decap_4 FILLER_76_1451 ();
 sg13g2_fill_1 FILLER_76_1459 ();
 sg13g2_fill_1 FILLER_76_1496 ();
 sg13g2_fill_1 FILLER_76_1506 ();
 sg13g2_decap_8 FILLER_76_1511 ();
 sg13g2_fill_2 FILLER_76_1518 ();
 sg13g2_fill_1 FILLER_76_1520 ();
 sg13g2_fill_1 FILLER_76_1526 ();
 sg13g2_fill_2 FILLER_76_1542 ();
 sg13g2_fill_2 FILLER_76_1578 ();
 sg13g2_decap_8 FILLER_76_1596 ();
 sg13g2_fill_1 FILLER_76_1603 ();
 sg13g2_decap_4 FILLER_76_1622 ();
 sg13g2_fill_2 FILLER_76_1642 ();
 sg13g2_fill_1 FILLER_76_1666 ();
 sg13g2_fill_1 FILLER_76_1693 ();
 sg13g2_decap_4 FILLER_76_1705 ();
 sg13g2_fill_1 FILLER_76_1750 ();
 sg13g2_fill_2 FILLER_76_1769 ();
 sg13g2_fill_1 FILLER_76_1771 ();
 sg13g2_decap_8 FILLER_76_1792 ();
 sg13g2_decap_8 FILLER_76_1799 ();
 sg13g2_decap_4 FILLER_76_1812 ();
 sg13g2_fill_2 FILLER_76_1816 ();
 sg13g2_decap_8 FILLER_76_1835 ();
 sg13g2_decap_8 FILLER_76_1947 ();
 sg13g2_fill_2 FILLER_76_1954 ();
 sg13g2_fill_1 FILLER_76_1956 ();
 sg13g2_fill_1 FILLER_76_1960 ();
 sg13g2_fill_1 FILLER_76_1970 ();
 sg13g2_decap_4 FILLER_76_1974 ();
 sg13g2_fill_1 FILLER_76_1978 ();
 sg13g2_decap_8 FILLER_76_1984 ();
 sg13g2_decap_8 FILLER_76_1991 ();
 sg13g2_fill_2 FILLER_76_2010 ();
 sg13g2_fill_1 FILLER_76_2012 ();
 sg13g2_decap_4 FILLER_76_2025 ();
 sg13g2_fill_1 FILLER_76_2029 ();
 sg13g2_fill_1 FILLER_76_2038 ();
 sg13g2_fill_1 FILLER_76_2087 ();
 sg13g2_decap_4 FILLER_76_2094 ();
 sg13g2_fill_2 FILLER_76_2127 ();
 sg13g2_fill_2 FILLER_76_2156 ();
 sg13g2_fill_1 FILLER_76_2158 ();
 sg13g2_fill_2 FILLER_76_2192 ();
 sg13g2_fill_2 FILLER_76_2197 ();
 sg13g2_fill_1 FILLER_76_2199 ();
 sg13g2_decap_4 FILLER_76_2218 ();
 sg13g2_decap_4 FILLER_76_2240 ();
 sg13g2_decap_4 FILLER_76_2248 ();
 sg13g2_fill_2 FILLER_76_2252 ();
 sg13g2_decap_4 FILLER_76_2317 ();
 sg13g2_fill_1 FILLER_76_2321 ();
 sg13g2_decap_8 FILLER_76_2338 ();
 sg13g2_fill_1 FILLER_76_2373 ();
 sg13g2_decap_8 FILLER_76_2399 ();
 sg13g2_decap_8 FILLER_76_2422 ();
 sg13g2_decap_4 FILLER_76_2429 ();
 sg13g2_fill_1 FILLER_76_2433 ();
 sg13g2_fill_2 FILLER_76_2450 ();
 sg13g2_fill_1 FILLER_76_2455 ();
 sg13g2_fill_1 FILLER_76_2474 ();
 sg13g2_fill_2 FILLER_76_2479 ();
 sg13g2_decap_8 FILLER_76_2489 ();
 sg13g2_decap_8 FILLER_76_2496 ();
 sg13g2_fill_1 FILLER_76_2503 ();
 sg13g2_fill_1 FILLER_76_2509 ();
 sg13g2_decap_4 FILLER_76_2518 ();
 sg13g2_fill_1 FILLER_76_2522 ();
 sg13g2_decap_8 FILLER_76_2542 ();
 sg13g2_decap_4 FILLER_76_2549 ();
 sg13g2_fill_1 FILLER_76_2553 ();
 sg13g2_fill_1 FILLER_76_2567 ();
 sg13g2_fill_1 FILLER_76_2573 ();
 sg13g2_fill_2 FILLER_76_2610 ();
 sg13g2_fill_2 FILLER_76_2625 ();
 sg13g2_decap_4 FILLER_76_2637 ();
 sg13g2_fill_1 FILLER_76_2641 ();
 sg13g2_fill_2 FILLER_76_2649 ();
 sg13g2_fill_1 FILLER_76_2660 ();
 sg13g2_decap_8 FILLER_76_2674 ();
 sg13g2_decap_4 FILLER_76_2681 ();
 sg13g2_fill_2 FILLER_76_2685 ();
 sg13g2_decap_8 FILLER_76_2691 ();
 sg13g2_decap_8 FILLER_76_2698 ();
 sg13g2_fill_2 FILLER_76_2705 ();
 sg13g2_fill_1 FILLER_76_2707 ();
 sg13g2_decap_4 FILLER_76_2750 ();
 sg13g2_decap_4 FILLER_76_2772 ();
 sg13g2_decap_4 FILLER_76_2835 ();
 sg13g2_fill_1 FILLER_76_2839 ();
 sg13g2_fill_1 FILLER_76_2868 ();
 sg13g2_fill_2 FILLER_76_2884 ();
 sg13g2_fill_1 FILLER_76_2886 ();
 sg13g2_decap_8 FILLER_76_2898 ();
 sg13g2_fill_2 FILLER_76_2905 ();
 sg13g2_fill_1 FILLER_76_2907 ();
 sg13g2_fill_2 FILLER_76_2943 ();
 sg13g2_fill_2 FILLER_76_2977 ();
 sg13g2_fill_2 FILLER_76_2984 ();
 sg13g2_fill_1 FILLER_76_2986 ();
 sg13g2_fill_2 FILLER_76_3000 ();
 sg13g2_decap_8 FILLER_76_3043 ();
 sg13g2_decap_8 FILLER_76_3059 ();
 sg13g2_fill_2 FILLER_76_3066 ();
 sg13g2_fill_2 FILLER_76_3084 ();
 sg13g2_decap_8 FILLER_76_3103 ();
 sg13g2_fill_2 FILLER_76_3110 ();
 sg13g2_fill_2 FILLER_76_3117 ();
 sg13g2_decap_8 FILLER_76_3132 ();
 sg13g2_fill_2 FILLER_76_3139 ();
 sg13g2_fill_1 FILLER_76_3160 ();
 sg13g2_decap_4 FILLER_76_3167 ();
 sg13g2_fill_2 FILLER_76_3185 ();
 sg13g2_fill_1 FILLER_76_3192 ();
 sg13g2_fill_2 FILLER_76_3197 ();
 sg13g2_fill_1 FILLER_76_3199 ();
 sg13g2_decap_8 FILLER_76_3218 ();
 sg13g2_decap_8 FILLER_76_3225 ();
 sg13g2_fill_2 FILLER_76_3232 ();
 sg13g2_fill_2 FILLER_76_3257 ();
 sg13g2_decap_4 FILLER_76_3331 ();
 sg13g2_decap_8 FILLER_76_3362 ();
 sg13g2_decap_8 FILLER_76_3369 ();
 sg13g2_decap_8 FILLER_76_3376 ();
 sg13g2_decap_8 FILLER_76_3383 ();
 sg13g2_decap_8 FILLER_76_3390 ();
 sg13g2_decap_8 FILLER_76_3397 ();
 sg13g2_decap_8 FILLER_76_3404 ();
 sg13g2_decap_8 FILLER_76_3411 ();
 sg13g2_decap_8 FILLER_76_3418 ();
 sg13g2_decap_8 FILLER_76_3425 ();
 sg13g2_decap_8 FILLER_76_3432 ();
 sg13g2_decap_8 FILLER_76_3439 ();
 sg13g2_decap_8 FILLER_76_3446 ();
 sg13g2_decap_8 FILLER_76_3453 ();
 sg13g2_decap_8 FILLER_76_3460 ();
 sg13g2_decap_8 FILLER_76_3467 ();
 sg13g2_decap_8 FILLER_76_3474 ();
 sg13g2_decap_8 FILLER_76_3481 ();
 sg13g2_decap_8 FILLER_76_3488 ();
 sg13g2_decap_8 FILLER_76_3495 ();
 sg13g2_decap_8 FILLER_76_3502 ();
 sg13g2_decap_8 FILLER_76_3509 ();
 sg13g2_decap_8 FILLER_76_3516 ();
 sg13g2_decap_8 FILLER_76_3523 ();
 sg13g2_decap_8 FILLER_76_3530 ();
 sg13g2_decap_8 FILLER_76_3537 ();
 sg13g2_decap_8 FILLER_76_3544 ();
 sg13g2_decap_8 FILLER_76_3551 ();
 sg13g2_decap_8 FILLER_76_3558 ();
 sg13g2_decap_8 FILLER_76_3565 ();
 sg13g2_decap_8 FILLER_76_3572 ();
 sg13g2_fill_1 FILLER_76_3579 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_4 FILLER_77_245 ();
 sg13g2_fill_1 FILLER_77_249 ();
 sg13g2_fill_1 FILLER_77_327 ();
 sg13g2_fill_1 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_77_410 ();
 sg13g2_decap_8 FILLER_77_417 ();
 sg13g2_decap_4 FILLER_77_424 ();
 sg13g2_fill_2 FILLER_77_441 ();
 sg13g2_fill_1 FILLER_77_443 ();
 sg13g2_fill_2 FILLER_77_500 ();
 sg13g2_decap_8 FILLER_77_506 ();
 sg13g2_fill_1 FILLER_77_513 ();
 sg13g2_decap_8 FILLER_77_578 ();
 sg13g2_fill_2 FILLER_77_585 ();
 sg13g2_fill_1 FILLER_77_587 ();
 sg13g2_fill_2 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_647 ();
 sg13g2_fill_2 FILLER_77_669 ();
 sg13g2_fill_1 FILLER_77_671 ();
 sg13g2_fill_2 FILLER_77_746 ();
 sg13g2_fill_1 FILLER_77_748 ();
 sg13g2_fill_2 FILLER_77_758 ();
 sg13g2_decap_4 FILLER_77_808 ();
 sg13g2_fill_2 FILLER_77_812 ();
 sg13g2_decap_4 FILLER_77_819 ();
 sg13g2_fill_2 FILLER_77_843 ();
 sg13g2_decap_8 FILLER_77_869 ();
 sg13g2_fill_2 FILLER_77_876 ();
 sg13g2_fill_1 FILLER_77_878 ();
 sg13g2_fill_2 FILLER_77_883 ();
 sg13g2_fill_1 FILLER_77_885 ();
 sg13g2_fill_2 FILLER_77_901 ();
 sg13g2_decap_8 FILLER_77_923 ();
 sg13g2_decap_8 FILLER_77_930 ();
 sg13g2_fill_1 FILLER_77_937 ();
 sg13g2_fill_2 FILLER_77_943 ();
 sg13g2_fill_1 FILLER_77_945 ();
 sg13g2_fill_1 FILLER_77_958 ();
 sg13g2_fill_1 FILLER_77_968 ();
 sg13g2_decap_4 FILLER_77_1000 ();
 sg13g2_fill_2 FILLER_77_1004 ();
 sg13g2_fill_2 FILLER_77_1038 ();
 sg13g2_fill_2 FILLER_77_1053 ();
 sg13g2_fill_1 FILLER_77_1055 ();
 sg13g2_fill_1 FILLER_77_1074 ();
 sg13g2_fill_2 FILLER_77_1078 ();
 sg13g2_fill_1 FILLER_77_1084 ();
 sg13g2_fill_2 FILLER_77_1094 ();
 sg13g2_decap_8 FILLER_77_1127 ();
 sg13g2_fill_2 FILLER_77_1134 ();
 sg13g2_decap_4 FILLER_77_1146 ();
 sg13g2_fill_2 FILLER_77_1174 ();
 sg13g2_decap_8 FILLER_77_1204 ();
 sg13g2_decap_4 FILLER_77_1211 ();
 sg13g2_fill_1 FILLER_77_1215 ();
 sg13g2_fill_1 FILLER_77_1244 ();
 sg13g2_fill_1 FILLER_77_1332 ();
 sg13g2_fill_1 FILLER_77_1353 ();
 sg13g2_decap_8 FILLER_77_1381 ();
 sg13g2_decap_4 FILLER_77_1388 ();
 sg13g2_fill_2 FILLER_77_1392 ();
 sg13g2_decap_4 FILLER_77_1414 ();
 sg13g2_decap_8 FILLER_77_1450 ();
 sg13g2_decap_4 FILLER_77_1457 ();
 sg13g2_fill_1 FILLER_77_1461 ();
 sg13g2_fill_2 FILLER_77_1489 ();
 sg13g2_fill_1 FILLER_77_1491 ();
 sg13g2_fill_1 FILLER_77_1510 ();
 sg13g2_decap_8 FILLER_77_1531 ();
 sg13g2_decap_8 FILLER_77_1538 ();
 sg13g2_fill_1 FILLER_77_1545 ();
 sg13g2_decap_8 FILLER_77_1598 ();
 sg13g2_fill_1 FILLER_77_1605 ();
 sg13g2_fill_1 FILLER_77_1643 ();
 sg13g2_fill_1 FILLER_77_1658 ();
 sg13g2_decap_4 FILLER_77_1663 ();
 sg13g2_fill_1 FILLER_77_1667 ();
 sg13g2_decap_4 FILLER_77_1676 ();
 sg13g2_decap_4 FILLER_77_1685 ();
 sg13g2_fill_1 FILLER_77_1689 ();
 sg13g2_fill_1 FILLER_77_1718 ();
 sg13g2_decap_8 FILLER_77_1736 ();
 sg13g2_fill_1 FILLER_77_1743 ();
 sg13g2_decap_4 FILLER_77_1773 ();
 sg13g2_decap_8 FILLER_77_1809 ();
 sg13g2_fill_2 FILLER_77_1816 ();
 sg13g2_fill_1 FILLER_77_1818 ();
 sg13g2_fill_1 FILLER_77_1840 ();
 sg13g2_fill_2 FILLER_77_1846 ();
 sg13g2_fill_1 FILLER_77_1848 ();
 sg13g2_fill_1 FILLER_77_1857 ();
 sg13g2_decap_8 FILLER_77_1867 ();
 sg13g2_fill_2 FILLER_77_1874 ();
 sg13g2_decap_8 FILLER_77_1885 ();
 sg13g2_decap_8 FILLER_77_1892 ();
 sg13g2_fill_1 FILLER_77_1931 ();
 sg13g2_decap_4 FILLER_77_1937 ();
 sg13g2_fill_2 FILLER_77_1941 ();
 sg13g2_fill_1 FILLER_77_1953 ();
 sg13g2_fill_2 FILLER_77_1979 ();
 sg13g2_decap_4 FILLER_77_2015 ();
 sg13g2_fill_2 FILLER_77_2035 ();
 sg13g2_decap_8 FILLER_77_2069 ();
 sg13g2_fill_1 FILLER_77_2076 ();
 sg13g2_decap_8 FILLER_77_2081 ();
 sg13g2_decap_8 FILLER_77_2088 ();
 sg13g2_decap_8 FILLER_77_2120 ();
 sg13g2_decap_4 FILLER_77_2127 ();
 sg13g2_decap_8 FILLER_77_2148 ();
 sg13g2_decap_8 FILLER_77_2155 ();
 sg13g2_decap_4 FILLER_77_2162 ();
 sg13g2_fill_1 FILLER_77_2170 ();
 sg13g2_decap_4 FILLER_77_2181 ();
 sg13g2_fill_1 FILLER_77_2185 ();
 sg13g2_fill_2 FILLER_77_2202 ();
 sg13g2_fill_1 FILLER_77_2204 ();
 sg13g2_fill_2 FILLER_77_2232 ();
 sg13g2_fill_1 FILLER_77_2234 ();
 sg13g2_fill_1 FILLER_77_2238 ();
 sg13g2_fill_2 FILLER_77_2267 ();
 sg13g2_fill_1 FILLER_77_2269 ();
 sg13g2_fill_1 FILLER_77_2283 ();
 sg13g2_fill_2 FILLER_77_2301 ();
 sg13g2_fill_2 FILLER_77_2313 ();
 sg13g2_decap_8 FILLER_77_2338 ();
 sg13g2_decap_8 FILLER_77_2345 ();
 sg13g2_fill_1 FILLER_77_2352 ();
 sg13g2_fill_1 FILLER_77_2358 ();
 sg13g2_fill_2 FILLER_77_2388 ();
 sg13g2_fill_1 FILLER_77_2390 ();
 sg13g2_decap_4 FILLER_77_2396 ();
 sg13g2_decap_4 FILLER_77_2420 ();
 sg13g2_fill_2 FILLER_77_2424 ();
 sg13g2_fill_2 FILLER_77_2481 ();
 sg13g2_fill_1 FILLER_77_2483 ();
 sg13g2_decap_8 FILLER_77_2493 ();
 sg13g2_fill_2 FILLER_77_2500 ();
 sg13g2_fill_1 FILLER_77_2520 ();
 sg13g2_fill_2 FILLER_77_2609 ();
 sg13g2_fill_1 FILLER_77_2611 ();
 sg13g2_decap_4 FILLER_77_2621 ();
 sg13g2_fill_1 FILLER_77_2625 ();
 sg13g2_fill_1 FILLER_77_2634 ();
 sg13g2_fill_2 FILLER_77_2647 ();
 sg13g2_decap_8 FILLER_77_2671 ();
 sg13g2_decap_4 FILLER_77_2678 ();
 sg13g2_decap_4 FILLER_77_2751 ();
 sg13g2_fill_1 FILLER_77_2755 ();
 sg13g2_decap_8 FILLER_77_2767 ();
 sg13g2_decap_8 FILLER_77_2774 ();
 sg13g2_fill_2 FILLER_77_2781 ();
 sg13g2_fill_1 FILLER_77_2783 ();
 sg13g2_decap_4 FILLER_77_2803 ();
 sg13g2_fill_2 FILLER_77_2807 ();
 sg13g2_fill_2 FILLER_77_2817 ();
 sg13g2_decap_8 FILLER_77_2828 ();
 sg13g2_decap_8 FILLER_77_2835 ();
 sg13g2_decap_8 FILLER_77_2842 ();
 sg13g2_fill_2 FILLER_77_2849 ();
 sg13g2_fill_1 FILLER_77_2851 ();
 sg13g2_decap_4 FILLER_77_2856 ();
 sg13g2_fill_1 FILLER_77_2860 ();
 sg13g2_fill_2 FILLER_77_2911 ();
 sg13g2_decap_8 FILLER_77_2917 ();
 sg13g2_decap_4 FILLER_77_2924 ();
 sg13g2_fill_2 FILLER_77_2928 ();
 sg13g2_fill_2 FILLER_77_2936 ();
 sg13g2_fill_1 FILLER_77_2943 ();
 sg13g2_decap_4 FILLER_77_2948 ();
 sg13g2_fill_1 FILLER_77_2952 ();
 sg13g2_fill_1 FILLER_77_2978 ();
 sg13g2_decap_8 FILLER_77_3000 ();
 sg13g2_fill_1 FILLER_77_3007 ();
 sg13g2_decap_4 FILLER_77_3012 ();
 sg13g2_decap_8 FILLER_77_3052 ();
 sg13g2_decap_4 FILLER_77_3059 ();
 sg13g2_fill_2 FILLER_77_3063 ();
 sg13g2_decap_4 FILLER_77_3081 ();
 sg13g2_decap_4 FILLER_77_3102 ();
 sg13g2_fill_1 FILLER_77_3118 ();
 sg13g2_decap_4 FILLER_77_3131 ();
 sg13g2_fill_1 FILLER_77_3135 ();
 sg13g2_decap_8 FILLER_77_3227 ();
 sg13g2_decap_4 FILLER_77_3234 ();
 sg13g2_decap_4 FILLER_77_3242 ();
 sg13g2_fill_1 FILLER_77_3246 ();
 sg13g2_decap_4 FILLER_77_3274 ();
 sg13g2_fill_2 FILLER_77_3278 ();
 sg13g2_decap_8 FILLER_77_3284 ();
 sg13g2_decap_8 FILLER_77_3291 ();
 sg13g2_decap_8 FILLER_77_3298 ();
 sg13g2_decap_8 FILLER_77_3305 ();
 sg13g2_decap_8 FILLER_77_3312 ();
 sg13g2_fill_1 FILLER_77_3319 ();
 sg13g2_decap_8 FILLER_77_3324 ();
 sg13g2_decap_8 FILLER_77_3331 ();
 sg13g2_fill_2 FILLER_77_3338 ();
 sg13g2_fill_1 FILLER_77_3340 ();
 sg13g2_decap_8 FILLER_77_3345 ();
 sg13g2_decap_8 FILLER_77_3352 ();
 sg13g2_decap_8 FILLER_77_3359 ();
 sg13g2_decap_8 FILLER_77_3366 ();
 sg13g2_decap_8 FILLER_77_3373 ();
 sg13g2_decap_8 FILLER_77_3380 ();
 sg13g2_decap_8 FILLER_77_3387 ();
 sg13g2_decap_8 FILLER_77_3394 ();
 sg13g2_decap_8 FILLER_77_3401 ();
 sg13g2_decap_8 FILLER_77_3408 ();
 sg13g2_decap_8 FILLER_77_3415 ();
 sg13g2_decap_8 FILLER_77_3422 ();
 sg13g2_decap_8 FILLER_77_3429 ();
 sg13g2_decap_8 FILLER_77_3436 ();
 sg13g2_decap_8 FILLER_77_3443 ();
 sg13g2_decap_8 FILLER_77_3450 ();
 sg13g2_decap_8 FILLER_77_3457 ();
 sg13g2_decap_8 FILLER_77_3464 ();
 sg13g2_decap_8 FILLER_77_3471 ();
 sg13g2_decap_8 FILLER_77_3478 ();
 sg13g2_decap_8 FILLER_77_3485 ();
 sg13g2_decap_8 FILLER_77_3492 ();
 sg13g2_decap_8 FILLER_77_3499 ();
 sg13g2_decap_8 FILLER_77_3506 ();
 sg13g2_decap_8 FILLER_77_3513 ();
 sg13g2_decap_8 FILLER_77_3520 ();
 sg13g2_decap_8 FILLER_77_3527 ();
 sg13g2_decap_8 FILLER_77_3534 ();
 sg13g2_decap_8 FILLER_77_3541 ();
 sg13g2_decap_8 FILLER_77_3548 ();
 sg13g2_decap_8 FILLER_77_3555 ();
 sg13g2_decap_8 FILLER_77_3562 ();
 sg13g2_decap_8 FILLER_77_3569 ();
 sg13g2_decap_4 FILLER_77_3576 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_4 FILLER_78_273 ();
 sg13g2_decap_4 FILLER_78_286 ();
 sg13g2_fill_1 FILLER_78_322 ();
 sg13g2_fill_2 FILLER_78_373 ();
 sg13g2_decap_4 FILLER_78_394 ();
 sg13g2_fill_1 FILLER_78_398 ();
 sg13g2_decap_8 FILLER_78_412 ();
 sg13g2_decap_8 FILLER_78_419 ();
 sg13g2_decap_4 FILLER_78_426 ();
 sg13g2_fill_2 FILLER_78_430 ();
 sg13g2_decap_8 FILLER_78_436 ();
 sg13g2_decap_4 FILLER_78_443 ();
 sg13g2_fill_2 FILLER_78_447 ();
 sg13g2_decap_8 FILLER_78_453 ();
 sg13g2_decap_8 FILLER_78_460 ();
 sg13g2_decap_8 FILLER_78_467 ();
 sg13g2_fill_2 FILLER_78_474 ();
 sg13g2_fill_1 FILLER_78_476 ();
 sg13g2_decap_8 FILLER_78_481 ();
 sg13g2_decap_4 FILLER_78_497 ();
 sg13g2_fill_1 FILLER_78_501 ();
 sg13g2_decap_8 FILLER_78_530 ();
 sg13g2_fill_2 FILLER_78_537 ();
 sg13g2_fill_1 FILLER_78_539 ();
 sg13g2_fill_2 FILLER_78_558 ();
 sg13g2_decap_4 FILLER_78_576 ();
 sg13g2_fill_2 FILLER_78_580 ();
 sg13g2_fill_2 FILLER_78_589 ();
 sg13g2_fill_2 FILLER_78_600 ();
 sg13g2_fill_2 FILLER_78_614 ();
 sg13g2_fill_2 FILLER_78_653 ();
 sg13g2_fill_1 FILLER_78_655 ();
 sg13g2_fill_2 FILLER_78_683 ();
 sg13g2_fill_1 FILLER_78_685 ();
 sg13g2_fill_2 FILLER_78_690 ();
 sg13g2_decap_8 FILLER_78_701 ();
 sg13g2_decap_8 FILLER_78_708 ();
 sg13g2_fill_2 FILLER_78_733 ();
 sg13g2_fill_1 FILLER_78_748 ();
 sg13g2_fill_2 FILLER_78_760 ();
 sg13g2_fill_2 FILLER_78_770 ();
 sg13g2_fill_2 FILLER_78_817 ();
 sg13g2_fill_1 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_879 ();
 sg13g2_fill_2 FILLER_78_886 ();
 sg13g2_fill_1 FILLER_78_888 ();
 sg13g2_fill_2 FILLER_78_956 ();
 sg13g2_decap_8 FILLER_78_966 ();
 sg13g2_decap_4 FILLER_78_973 ();
 sg13g2_decap_4 FILLER_78_1005 ();
 sg13g2_fill_2 FILLER_78_1009 ();
 sg13g2_decap_8 FILLER_78_1015 ();
 sg13g2_decap_4 FILLER_78_1022 ();
 sg13g2_fill_2 FILLER_78_1026 ();
 sg13g2_decap_4 FILLER_78_1037 ();
 sg13g2_fill_2 FILLER_78_1041 ();
 sg13g2_fill_2 FILLER_78_1086 ();
 sg13g2_decap_4 FILLER_78_1109 ();
 sg13g2_fill_2 FILLER_78_1113 ();
 sg13g2_decap_4 FILLER_78_1119 ();
 sg13g2_decap_8 FILLER_78_1162 ();
 sg13g2_fill_2 FILLER_78_1169 ();
 sg13g2_fill_1 FILLER_78_1174 ();
 sg13g2_decap_8 FILLER_78_1216 ();
 sg13g2_fill_2 FILLER_78_1223 ();
 sg13g2_fill_2 FILLER_78_1280 ();
 sg13g2_fill_2 FILLER_78_1310 ();
 sg13g2_fill_1 FILLER_78_1315 ();
 sg13g2_fill_1 FILLER_78_1333 ();
 sg13g2_decap_4 FILLER_78_1385 ();
 sg13g2_fill_2 FILLER_78_1400 ();
 sg13g2_decap_8 FILLER_78_1406 ();
 sg13g2_fill_2 FILLER_78_1413 ();
 sg13g2_fill_2 FILLER_78_1436 ();
 sg13g2_fill_1 FILLER_78_1465 ();
 sg13g2_decap_8 FILLER_78_1479 ();
 sg13g2_fill_2 FILLER_78_1486 ();
 sg13g2_fill_1 FILLER_78_1488 ();
 sg13g2_fill_1 FILLER_78_1558 ();
 sg13g2_fill_2 FILLER_78_1605 ();
 sg13g2_decap_4 FILLER_78_1620 ();
 sg13g2_fill_2 FILLER_78_1624 ();
 sg13g2_fill_2 FILLER_78_1682 ();
 sg13g2_fill_1 FILLER_78_1684 ();
 sg13g2_fill_1 FILLER_78_1713 ();
 sg13g2_decap_4 FILLER_78_1741 ();
 sg13g2_fill_1 FILLER_78_1745 ();
 sg13g2_decap_8 FILLER_78_1789 ();
 sg13g2_fill_2 FILLER_78_1796 ();
 sg13g2_fill_1 FILLER_78_1798 ();
 sg13g2_fill_1 FILLER_78_1865 ();
 sg13g2_decap_4 FILLER_78_1874 ();
 sg13g2_fill_2 FILLER_78_1878 ();
 sg13g2_fill_1 FILLER_78_1920 ();
 sg13g2_decap_4 FILLER_78_1933 ();
 sg13g2_fill_1 FILLER_78_1957 ();
 sg13g2_fill_1 FILLER_78_1976 ();
 sg13g2_decap_8 FILLER_78_1990 ();
 sg13g2_fill_2 FILLER_78_1997 ();
 sg13g2_fill_1 FILLER_78_2023 ();
 sg13g2_decap_8 FILLER_78_2034 ();
 sg13g2_fill_1 FILLER_78_2041 ();
 sg13g2_fill_1 FILLER_78_2070 ();
 sg13g2_fill_1 FILLER_78_2114 ();
 sg13g2_fill_1 FILLER_78_2123 ();
 sg13g2_fill_2 FILLER_78_2136 ();
 sg13g2_fill_2 FILLER_78_2142 ();
 sg13g2_fill_2 FILLER_78_2147 ();
 sg13g2_fill_1 FILLER_78_2149 ();
 sg13g2_decap_4 FILLER_78_2178 ();
 sg13g2_fill_1 FILLER_78_2182 ();
 sg13g2_fill_1 FILLER_78_2192 ();
 sg13g2_decap_8 FILLER_78_2215 ();
 sg13g2_fill_1 FILLER_78_2250 ();
 sg13g2_decap_4 FILLER_78_2260 ();
 sg13g2_fill_1 FILLER_78_2264 ();
 sg13g2_fill_2 FILLER_78_2293 ();
 sg13g2_fill_1 FILLER_78_2295 ();
 sg13g2_fill_2 FILLER_78_2338 ();
 sg13g2_fill_2 FILLER_78_2356 ();
 sg13g2_decap_4 FILLER_78_2361 ();
 sg13g2_fill_2 FILLER_78_2393 ();
 sg13g2_decap_8 FILLER_78_2413 ();
 sg13g2_decap_8 FILLER_78_2420 ();
 sg13g2_decap_4 FILLER_78_2427 ();
 sg13g2_fill_1 FILLER_78_2431 ();
 sg13g2_fill_1 FILLER_78_2454 ();
 sg13g2_fill_2 FILLER_78_2469 ();
 sg13g2_fill_2 FILLER_78_2504 ();
 sg13g2_fill_1 FILLER_78_2506 ();
 sg13g2_decap_8 FILLER_78_2516 ();
 sg13g2_fill_2 FILLER_78_2523 ();
 sg13g2_fill_1 FILLER_78_2525 ();
 sg13g2_decap_8 FILLER_78_2530 ();
 sg13g2_decap_4 FILLER_78_2537 ();
 sg13g2_fill_1 FILLER_78_2541 ();
 sg13g2_decap_8 FILLER_78_2546 ();
 sg13g2_decap_8 FILLER_78_2610 ();
 sg13g2_fill_2 FILLER_78_2617 ();
 sg13g2_fill_1 FILLER_78_2623 ();
 sg13g2_fill_1 FILLER_78_2643 ();
 sg13g2_decap_4 FILLER_78_2678 ();
 sg13g2_fill_2 FILLER_78_2682 ();
 sg13g2_fill_1 FILLER_78_2721 ();
 sg13g2_fill_1 FILLER_78_2731 ();
 sg13g2_decap_4 FILLER_78_2779 ();
 sg13g2_fill_1 FILLER_78_2783 ();
 sg13g2_decap_4 FILLER_78_2811 ();
 sg13g2_fill_2 FILLER_78_2815 ();
 sg13g2_fill_2 FILLER_78_2844 ();
 sg13g2_fill_1 FILLER_78_2846 ();
 sg13g2_fill_2 FILLER_78_2880 ();
 sg13g2_fill_1 FILLER_78_2882 ();
 sg13g2_decap_8 FILLER_78_2911 ();
 sg13g2_decap_4 FILLER_78_2918 ();
 sg13g2_decap_4 FILLER_78_2935 ();
 sg13g2_fill_2 FILLER_78_2939 ();
 sg13g2_fill_1 FILLER_78_2958 ();
 sg13g2_decap_4 FILLER_78_2994 ();
 sg13g2_fill_1 FILLER_78_2998 ();
 sg13g2_decap_8 FILLER_78_3027 ();
 sg13g2_decap_8 FILLER_78_3034 ();
 sg13g2_fill_1 FILLER_78_3041 ();
 sg13g2_decap_4 FILLER_78_3086 ();
 sg13g2_fill_2 FILLER_78_3096 ();
 sg13g2_decap_8 FILLER_78_3127 ();
 sg13g2_decap_8 FILLER_78_3134 ();
 sg13g2_decap_4 FILLER_78_3141 ();
 sg13g2_fill_1 FILLER_78_3145 ();
 sg13g2_fill_1 FILLER_78_3232 ();
 sg13g2_decap_8 FILLER_78_3289 ();
 sg13g2_decap_8 FILLER_78_3296 ();
 sg13g2_decap_8 FILLER_78_3303 ();
 sg13g2_decap_8 FILLER_78_3310 ();
 sg13g2_decap_8 FILLER_78_3317 ();
 sg13g2_decap_8 FILLER_78_3324 ();
 sg13g2_decap_8 FILLER_78_3331 ();
 sg13g2_decap_8 FILLER_78_3338 ();
 sg13g2_decap_8 FILLER_78_3345 ();
 sg13g2_decap_8 FILLER_78_3352 ();
 sg13g2_decap_8 FILLER_78_3359 ();
 sg13g2_decap_8 FILLER_78_3366 ();
 sg13g2_decap_8 FILLER_78_3373 ();
 sg13g2_decap_8 FILLER_78_3380 ();
 sg13g2_decap_8 FILLER_78_3387 ();
 sg13g2_decap_8 FILLER_78_3394 ();
 sg13g2_decap_8 FILLER_78_3401 ();
 sg13g2_decap_8 FILLER_78_3408 ();
 sg13g2_decap_8 FILLER_78_3415 ();
 sg13g2_decap_8 FILLER_78_3422 ();
 sg13g2_decap_8 FILLER_78_3429 ();
 sg13g2_decap_8 FILLER_78_3436 ();
 sg13g2_decap_8 FILLER_78_3443 ();
 sg13g2_decap_8 FILLER_78_3450 ();
 sg13g2_decap_8 FILLER_78_3457 ();
 sg13g2_decap_8 FILLER_78_3464 ();
 sg13g2_decap_8 FILLER_78_3471 ();
 sg13g2_decap_8 FILLER_78_3478 ();
 sg13g2_decap_8 FILLER_78_3485 ();
 sg13g2_decap_8 FILLER_78_3492 ();
 sg13g2_decap_8 FILLER_78_3499 ();
 sg13g2_decap_8 FILLER_78_3506 ();
 sg13g2_decap_8 FILLER_78_3513 ();
 sg13g2_decap_8 FILLER_78_3520 ();
 sg13g2_decap_8 FILLER_78_3527 ();
 sg13g2_decap_8 FILLER_78_3534 ();
 sg13g2_decap_8 FILLER_78_3541 ();
 sg13g2_decap_8 FILLER_78_3548 ();
 sg13g2_decap_8 FILLER_78_3555 ();
 sg13g2_decap_8 FILLER_78_3562 ();
 sg13g2_decap_8 FILLER_78_3569 ();
 sg13g2_decap_4 FILLER_78_3576 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_fill_2 FILLER_79_308 ();
 sg13g2_fill_2 FILLER_79_355 ();
 sg13g2_fill_2 FILLER_79_387 ();
 sg13g2_fill_1 FILLER_79_389 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_fill_2 FILLER_79_504 ();
 sg13g2_fill_1 FILLER_79_506 ();
 sg13g2_decap_8 FILLER_79_511 ();
 sg13g2_decap_8 FILLER_79_518 ();
 sg13g2_decap_8 FILLER_79_525 ();
 sg13g2_decap_8 FILLER_79_532 ();
 sg13g2_fill_2 FILLER_79_539 ();
 sg13g2_decap_8 FILLER_79_568 ();
 sg13g2_decap_4 FILLER_79_575 ();
 sg13g2_fill_1 FILLER_79_579 ();
 sg13g2_fill_2 FILLER_79_608 ();
 sg13g2_fill_1 FILLER_79_610 ();
 sg13g2_fill_1 FILLER_79_628 ();
 sg13g2_decap_8 FILLER_79_642 ();
 sg13g2_decap_8 FILLER_79_649 ();
 sg13g2_decap_4 FILLER_79_656 ();
 sg13g2_fill_1 FILLER_79_660 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_8 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_679 ();
 sg13g2_decap_8 FILLER_79_686 ();
 sg13g2_decap_8 FILLER_79_693 ();
 sg13g2_decap_8 FILLER_79_700 ();
 sg13g2_decap_4 FILLER_79_707 ();
 sg13g2_fill_1 FILLER_79_711 ();
 sg13g2_fill_1 FILLER_79_757 ();
 sg13g2_decap_4 FILLER_79_765 ();
 sg13g2_fill_2 FILLER_79_797 ();
 sg13g2_decap_4 FILLER_79_829 ();
 sg13g2_decap_8 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_79_868 ();
 sg13g2_decap_8 FILLER_79_875 ();
 sg13g2_decap_8 FILLER_79_882 ();
 sg13g2_decap_4 FILLER_79_889 ();
 sg13g2_fill_1 FILLER_79_893 ();
 sg13g2_decap_4 FILLER_79_898 ();
 sg13g2_fill_2 FILLER_79_902 ();
 sg13g2_decap_8 FILLER_79_907 ();
 sg13g2_decap_8 FILLER_79_914 ();
 sg13g2_decap_8 FILLER_79_921 ();
 sg13g2_decap_4 FILLER_79_956 ();
 sg13g2_fill_1 FILLER_79_960 ();
 sg13g2_decap_8 FILLER_79_970 ();
 sg13g2_decap_4 FILLER_79_977 ();
 sg13g2_fill_1 FILLER_79_981 ();
 sg13g2_decap_8 FILLER_79_1010 ();
 sg13g2_decap_8 FILLER_79_1017 ();
 sg13g2_decap_8 FILLER_79_1024 ();
 sg13g2_decap_8 FILLER_79_1031 ();
 sg13g2_decap_8 FILLER_79_1038 ();
 sg13g2_decap_8 FILLER_79_1045 ();
 sg13g2_decap_8 FILLER_79_1052 ();
 sg13g2_decap_8 FILLER_79_1059 ();
 sg13g2_decap_4 FILLER_79_1066 ();
 sg13g2_fill_2 FILLER_79_1106 ();
 sg13g2_fill_1 FILLER_79_1108 ();
 sg13g2_fill_2 FILLER_79_1146 ();
 sg13g2_fill_1 FILLER_79_1148 ();
 sg13g2_decap_8 FILLER_79_1199 ();
 sg13g2_decap_8 FILLER_79_1206 ();
 sg13g2_decap_8 FILLER_79_1213 ();
 sg13g2_decap_8 FILLER_79_1220 ();
 sg13g2_decap_4 FILLER_79_1227 ();
 sg13g2_decap_4 FILLER_79_1235 ();
 sg13g2_decap_8 FILLER_79_1248 ();
 sg13g2_decap_8 FILLER_79_1255 ();
 sg13g2_decap_8 FILLER_79_1262 ();
 sg13g2_fill_2 FILLER_79_1347 ();
 sg13g2_fill_1 FILLER_79_1349 ();
 sg13g2_fill_2 FILLER_79_1390 ();
 sg13g2_fill_1 FILLER_79_1392 ();
 sg13g2_decap_8 FILLER_79_1443 ();
 sg13g2_decap_8 FILLER_79_1450 ();
 sg13g2_decap_8 FILLER_79_1457 ();
 sg13g2_decap_8 FILLER_79_1464 ();
 sg13g2_decap_8 FILLER_79_1471 ();
 sg13g2_decap_8 FILLER_79_1478 ();
 sg13g2_decap_8 FILLER_79_1485 ();
 sg13g2_decap_4 FILLER_79_1492 ();
 sg13g2_fill_1 FILLER_79_1496 ();
 sg13g2_fill_1 FILLER_79_1525 ();
 sg13g2_decap_8 FILLER_79_1539 ();
 sg13g2_fill_2 FILLER_79_1546 ();
 sg13g2_fill_1 FILLER_79_1548 ();
 sg13g2_decap_4 FILLER_79_1553 ();
 sg13g2_fill_1 FILLER_79_1557 ();
 sg13g2_fill_1 FILLER_79_1562 ();
 sg13g2_fill_1 FILLER_79_1619 ();
 sg13g2_decap_4 FILLER_79_1651 ();
 sg13g2_fill_1 FILLER_79_1655 ();
 sg13g2_decap_8 FILLER_79_1693 ();
 sg13g2_fill_1 FILLER_79_1700 ();
 sg13g2_decap_4 FILLER_79_1770 ();
 sg13g2_decap_8 FILLER_79_1783 ();
 sg13g2_decap_8 FILLER_79_1790 ();
 sg13g2_decap_8 FILLER_79_1797 ();
 sg13g2_fill_1 FILLER_79_1804 ();
 sg13g2_decap_8 FILLER_79_1809 ();
 sg13g2_decap_8 FILLER_79_1816 ();
 sg13g2_decap_4 FILLER_79_1879 ();
 sg13g2_fill_2 FILLER_79_1883 ();
 sg13g2_decap_8 FILLER_79_1889 ();
 sg13g2_fill_2 FILLER_79_1905 ();
 sg13g2_fill_1 FILLER_79_1907 ();
 sg13g2_fill_2 FILLER_79_1914 ();
 sg13g2_decap_4 FILLER_79_1920 ();
 sg13g2_fill_2 FILLER_79_1924 ();
 sg13g2_fill_2 FILLER_79_1935 ();
 sg13g2_decap_4 FILLER_79_1991 ();
 sg13g2_fill_1 FILLER_79_1995 ();
 sg13g2_decap_8 FILLER_79_2037 ();
 sg13g2_fill_2 FILLER_79_2044 ();
 sg13g2_fill_1 FILLER_79_2046 ();
 sg13g2_fill_1 FILLER_79_2051 ();
 sg13g2_fill_2 FILLER_79_2061 ();
 sg13g2_fill_1 FILLER_79_2076 ();
 sg13g2_decap_8 FILLER_79_2081 ();
 sg13g2_decap_8 FILLER_79_2088 ();
 sg13g2_fill_2 FILLER_79_2095 ();
 sg13g2_fill_1 FILLER_79_2110 ();
 sg13g2_decap_8 FILLER_79_2114 ();
 sg13g2_decap_4 FILLER_79_2121 ();
 sg13g2_fill_2 FILLER_79_2125 ();
 sg13g2_decap_8 FILLER_79_2162 ();
 sg13g2_decap_8 FILLER_79_2169 ();
 sg13g2_decap_8 FILLER_79_2235 ();
 sg13g2_decap_8 FILLER_79_2242 ();
 sg13g2_decap_8 FILLER_79_2249 ();
 sg13g2_decap_8 FILLER_79_2256 ();
 sg13g2_decap_8 FILLER_79_2263 ();
 sg13g2_decap_8 FILLER_79_2270 ();
 sg13g2_fill_1 FILLER_79_2277 ();
 sg13g2_fill_1 FILLER_79_2306 ();
 sg13g2_fill_2 FILLER_79_2341 ();
 sg13g2_fill_1 FILLER_79_2343 ();
 sg13g2_decap_8 FILLER_79_2357 ();
 sg13g2_fill_1 FILLER_79_2364 ();
 sg13g2_decap_8 FILLER_79_2374 ();
 sg13g2_fill_1 FILLER_79_2381 ();
 sg13g2_decap_8 FILLER_79_2386 ();
 sg13g2_decap_8 FILLER_79_2421 ();
 sg13g2_decap_8 FILLER_79_2428 ();
 sg13g2_decap_4 FILLER_79_2435 ();
 sg13g2_fill_2 FILLER_79_2439 ();
 sg13g2_fill_2 FILLER_79_2469 ();
 sg13g2_decap_8 FILLER_79_2519 ();
 sg13g2_decap_8 FILLER_79_2526 ();
 sg13g2_decap_4 FILLER_79_2533 ();
 sg13g2_fill_1 FILLER_79_2574 ();
 sg13g2_fill_2 FILLER_79_2602 ();
 sg13g2_fill_1 FILLER_79_2617 ();
 sg13g2_fill_1 FILLER_79_2646 ();
 sg13g2_fill_1 FILLER_79_2688 ();
 sg13g2_decap_8 FILLER_79_2693 ();
 sg13g2_fill_2 FILLER_79_2748 ();
 sg13g2_decap_4 FILLER_79_2763 ();
 sg13g2_decap_8 FILLER_79_2776 ();
 sg13g2_decap_4 FILLER_79_2783 ();
 sg13g2_fill_1 FILLER_79_2787 ();
 sg13g2_fill_2 FILLER_79_2792 ();
 sg13g2_decap_8 FILLER_79_2826 ();
 sg13g2_decap_8 FILLER_79_2833 ();
 sg13g2_decap_8 FILLER_79_2840 ();
 sg13g2_decap_8 FILLER_79_2847 ();
 sg13g2_decap_8 FILLER_79_2854 ();
 sg13g2_decap_8 FILLER_79_2861 ();
 sg13g2_decap_8 FILLER_79_2868 ();
 sg13g2_decap_4 FILLER_79_2892 ();
 sg13g2_decap_8 FILLER_79_2900 ();
 sg13g2_fill_1 FILLER_79_2907 ();
 sg13g2_fill_2 FILLER_79_2917 ();
 sg13g2_fill_1 FILLER_79_2955 ();
 sg13g2_decap_8 FILLER_79_3030 ();
 sg13g2_decap_8 FILLER_79_3037 ();
 sg13g2_fill_2 FILLER_79_3044 ();
 sg13g2_fill_1 FILLER_79_3046 ();
 sg13g2_decap_8 FILLER_79_3051 ();
 sg13g2_decap_4 FILLER_79_3058 ();
 sg13g2_fill_1 FILLER_79_3062 ();
 sg13g2_fill_2 FILLER_79_3067 ();
 sg13g2_fill_2 FILLER_79_3091 ();
 sg13g2_decap_8 FILLER_79_3134 ();
 sg13g2_decap_8 FILLER_79_3141 ();
 sg13g2_fill_2 FILLER_79_3148 ();
 sg13g2_fill_1 FILLER_79_3150 ();
 sg13g2_decap_4 FILLER_79_3155 ();
 sg13g2_fill_2 FILLER_79_3227 ();
 sg13g2_decap_8 FILLER_79_3233 ();
 sg13g2_decap_8 FILLER_79_3240 ();
 sg13g2_decap_8 FILLER_79_3247 ();
 sg13g2_decap_4 FILLER_79_3254 ();
 sg13g2_fill_2 FILLER_79_3258 ();
 sg13g2_decap_8 FILLER_79_3264 ();
 sg13g2_fill_2 FILLER_79_3271 ();
 sg13g2_decap_8 FILLER_79_3282 ();
 sg13g2_decap_8 FILLER_79_3289 ();
 sg13g2_decap_8 FILLER_79_3296 ();
 sg13g2_decap_8 FILLER_79_3303 ();
 sg13g2_decap_8 FILLER_79_3310 ();
 sg13g2_decap_8 FILLER_79_3317 ();
 sg13g2_decap_8 FILLER_79_3324 ();
 sg13g2_decap_8 FILLER_79_3331 ();
 sg13g2_decap_8 FILLER_79_3338 ();
 sg13g2_decap_8 FILLER_79_3345 ();
 sg13g2_decap_8 FILLER_79_3352 ();
 sg13g2_decap_8 FILLER_79_3359 ();
 sg13g2_decap_8 FILLER_79_3366 ();
 sg13g2_decap_8 FILLER_79_3373 ();
 sg13g2_decap_8 FILLER_79_3380 ();
 sg13g2_decap_8 FILLER_79_3387 ();
 sg13g2_decap_8 FILLER_79_3394 ();
 sg13g2_decap_8 FILLER_79_3401 ();
 sg13g2_decap_8 FILLER_79_3408 ();
 sg13g2_decap_8 FILLER_79_3415 ();
 sg13g2_decap_8 FILLER_79_3422 ();
 sg13g2_decap_8 FILLER_79_3429 ();
 sg13g2_decap_8 FILLER_79_3436 ();
 sg13g2_decap_8 FILLER_79_3443 ();
 sg13g2_decap_8 FILLER_79_3450 ();
 sg13g2_decap_8 FILLER_79_3457 ();
 sg13g2_decap_8 FILLER_79_3464 ();
 sg13g2_decap_8 FILLER_79_3471 ();
 sg13g2_decap_8 FILLER_79_3478 ();
 sg13g2_decap_8 FILLER_79_3485 ();
 sg13g2_decap_8 FILLER_79_3492 ();
 sg13g2_decap_8 FILLER_79_3499 ();
 sg13g2_decap_8 FILLER_79_3506 ();
 sg13g2_decap_8 FILLER_79_3513 ();
 sg13g2_decap_8 FILLER_79_3520 ();
 sg13g2_decap_8 FILLER_79_3527 ();
 sg13g2_decap_8 FILLER_79_3534 ();
 sg13g2_decap_8 FILLER_79_3541 ();
 sg13g2_decap_8 FILLER_79_3548 ();
 sg13g2_decap_8 FILLER_79_3555 ();
 sg13g2_decap_8 FILLER_79_3562 ();
 sg13g2_decap_8 FILLER_79_3569 ();
 sg13g2_decap_4 FILLER_79_3576 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_8 FILLER_80_164 ();
 sg13g2_decap_8 FILLER_80_171 ();
 sg13g2_decap_8 FILLER_80_178 ();
 sg13g2_decap_8 FILLER_80_185 ();
 sg13g2_decap_8 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_213 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_227 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_decap_8 FILLER_80_241 ();
 sg13g2_decap_8 FILLER_80_248 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_269 ();
 sg13g2_decap_4 FILLER_80_276 ();
 sg13g2_decap_4 FILLER_80_284 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_fill_2 FILLER_80_299 ();
 sg13g2_fill_1 FILLER_80_358 ();
 sg13g2_fill_2 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_decap_8 FILLER_80_406 ();
 sg13g2_decap_8 FILLER_80_413 ();
 sg13g2_decap_8 FILLER_80_420 ();
 sg13g2_decap_8 FILLER_80_427 ();
 sg13g2_decap_8 FILLER_80_434 ();
 sg13g2_decap_8 FILLER_80_441 ();
 sg13g2_decap_8 FILLER_80_448 ();
 sg13g2_decap_8 FILLER_80_455 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_decap_8 FILLER_80_469 ();
 sg13g2_decap_8 FILLER_80_476 ();
 sg13g2_decap_8 FILLER_80_483 ();
 sg13g2_decap_8 FILLER_80_490 ();
 sg13g2_decap_8 FILLER_80_497 ();
 sg13g2_decap_8 FILLER_80_504 ();
 sg13g2_decap_8 FILLER_80_511 ();
 sg13g2_decap_8 FILLER_80_518 ();
 sg13g2_decap_4 FILLER_80_525 ();
 sg13g2_fill_2 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_decap_8 FILLER_80_570 ();
 sg13g2_fill_1 FILLER_80_577 ();
 sg13g2_decap_4 FILLER_80_610 ();
 sg13g2_decap_8 FILLER_80_642 ();
 sg13g2_decap_8 FILLER_80_649 ();
 sg13g2_decap_8 FILLER_80_656 ();
 sg13g2_decap_8 FILLER_80_663 ();
 sg13g2_decap_8 FILLER_80_670 ();
 sg13g2_decap_8 FILLER_80_677 ();
 sg13g2_decap_8 FILLER_80_684 ();
 sg13g2_decap_8 FILLER_80_691 ();
 sg13g2_decap_8 FILLER_80_698 ();
 sg13g2_decap_8 FILLER_80_705 ();
 sg13g2_decap_4 FILLER_80_712 ();
 sg13g2_fill_1 FILLER_80_716 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_4 FILLER_80_728 ();
 sg13g2_fill_2 FILLER_80_732 ();
 sg13g2_fill_2 FILLER_80_771 ();
 sg13g2_fill_1 FILLER_80_773 ();
 sg13g2_decap_8 FILLER_80_778 ();
 sg13g2_fill_1 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_4 FILLER_80_835 ();
 sg13g2_fill_2 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_decap_8 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_910 ();
 sg13g2_decap_8 FILLER_80_917 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_fill_2 FILLER_80_931 ();
 sg13g2_decap_4 FILLER_80_937 ();
 sg13g2_decap_8 FILLER_80_977 ();
 sg13g2_fill_2 FILLER_80_984 ();
 sg13g2_fill_1 FILLER_80_986 ();
 sg13g2_decap_8 FILLER_80_991 ();
 sg13g2_decap_8 FILLER_80_998 ();
 sg13g2_decap_8 FILLER_80_1005 ();
 sg13g2_decap_8 FILLER_80_1012 ();
 sg13g2_decap_8 FILLER_80_1019 ();
 sg13g2_decap_8 FILLER_80_1026 ();
 sg13g2_decap_8 FILLER_80_1033 ();
 sg13g2_decap_8 FILLER_80_1040 ();
 sg13g2_decap_8 FILLER_80_1047 ();
 sg13g2_decap_8 FILLER_80_1054 ();
 sg13g2_decap_8 FILLER_80_1061 ();
 sg13g2_decap_4 FILLER_80_1068 ();
 sg13g2_decap_8 FILLER_80_1088 ();
 sg13g2_decap_4 FILLER_80_1095 ();
 sg13g2_fill_1 FILLER_80_1099 ();
 sg13g2_decap_8 FILLER_80_1104 ();
 sg13g2_fill_2 FILLER_80_1111 ();
 sg13g2_fill_1 FILLER_80_1113 ();
 sg13g2_decap_8 FILLER_80_1118 ();
 sg13g2_fill_2 FILLER_80_1125 ();
 sg13g2_decap_4 FILLER_80_1158 ();
 sg13g2_fill_1 FILLER_80_1162 ();
 sg13g2_decap_8 FILLER_80_1167 ();
 sg13g2_decap_8 FILLER_80_1174 ();
 sg13g2_decap_8 FILLER_80_1181 ();
 sg13g2_decap_8 FILLER_80_1188 ();
 sg13g2_decap_8 FILLER_80_1195 ();
 sg13g2_decap_8 FILLER_80_1202 ();
 sg13g2_decap_8 FILLER_80_1209 ();
 sg13g2_decap_8 FILLER_80_1216 ();
 sg13g2_decap_8 FILLER_80_1223 ();
 sg13g2_decap_8 FILLER_80_1230 ();
 sg13g2_decap_8 FILLER_80_1237 ();
 sg13g2_decap_8 FILLER_80_1244 ();
 sg13g2_decap_8 FILLER_80_1251 ();
 sg13g2_decap_8 FILLER_80_1262 ();
 sg13g2_decap_4 FILLER_80_1269 ();
 sg13g2_fill_1 FILLER_80_1273 ();
 sg13g2_fill_2 FILLER_80_1278 ();
 sg13g2_fill_1 FILLER_80_1280 ();
 sg13g2_fill_1 FILLER_80_1290 ();
 sg13g2_decap_4 FILLER_80_1294 ();
 sg13g2_fill_1 FILLER_80_1330 ();
 sg13g2_fill_2 FILLER_80_1363 ();
 sg13g2_fill_1 FILLER_80_1365 ();
 sg13g2_decap_4 FILLER_80_1406 ();
 sg13g2_fill_1 FILLER_80_1410 ();
 sg13g2_decap_8 FILLER_80_1415 ();
 sg13g2_decap_8 FILLER_80_1422 ();
 sg13g2_decap_4 FILLER_80_1429 ();
 sg13g2_fill_1 FILLER_80_1433 ();
 sg13g2_decap_8 FILLER_80_1437 ();
 sg13g2_decap_8 FILLER_80_1444 ();
 sg13g2_decap_8 FILLER_80_1451 ();
 sg13g2_decap_8 FILLER_80_1458 ();
 sg13g2_decap_8 FILLER_80_1465 ();
 sg13g2_decap_8 FILLER_80_1472 ();
 sg13g2_decap_8 FILLER_80_1479 ();
 sg13g2_decap_8 FILLER_80_1486 ();
 sg13g2_decap_8 FILLER_80_1493 ();
 sg13g2_fill_2 FILLER_80_1500 ();
 sg13g2_decap_8 FILLER_80_1506 ();
 sg13g2_decap_8 FILLER_80_1513 ();
 sg13g2_decap_8 FILLER_80_1520 ();
 sg13g2_decap_8 FILLER_80_1527 ();
 sg13g2_decap_8 FILLER_80_1534 ();
 sg13g2_fill_2 FILLER_80_1541 ();
 sg13g2_fill_2 FILLER_80_1571 ();
 sg13g2_decap_4 FILLER_80_1577 ();
 sg13g2_fill_1 FILLER_80_1585 ();
 sg13g2_fill_2 FILLER_80_1595 ();
 sg13g2_decap_8 FILLER_80_1601 ();
 sg13g2_decap_8 FILLER_80_1608 ();
 sg13g2_decap_8 FILLER_80_1615 ();
 sg13g2_fill_2 FILLER_80_1622 ();
 sg13g2_fill_1 FILLER_80_1624 ();
 sg13g2_decap_8 FILLER_80_1629 ();
 sg13g2_decap_8 FILLER_80_1636 ();
 sg13g2_fill_2 FILLER_80_1643 ();
 sg13g2_fill_1 FILLER_80_1645 ();
 sg13g2_decap_8 FILLER_80_1650 ();
 sg13g2_decap_8 FILLER_80_1657 ();
 sg13g2_decap_4 FILLER_80_1664 ();
 sg13g2_fill_2 FILLER_80_1668 ();
 sg13g2_decap_8 FILLER_80_1674 ();
 sg13g2_decap_8 FILLER_80_1681 ();
 sg13g2_fill_2 FILLER_80_1688 ();
 sg13g2_decap_8 FILLER_80_1694 ();
 sg13g2_fill_2 FILLER_80_1701 ();
 sg13g2_decap_8 FILLER_80_1724 ();
 sg13g2_decap_4 FILLER_80_1731 ();
 sg13g2_decap_8 FILLER_80_1739 ();
 sg13g2_decap_8 FILLER_80_1746 ();
 sg13g2_decap_8 FILLER_80_1753 ();
 sg13g2_decap_8 FILLER_80_1760 ();
 sg13g2_decap_8 FILLER_80_1767 ();
 sg13g2_decap_8 FILLER_80_1774 ();
 sg13g2_decap_8 FILLER_80_1781 ();
 sg13g2_decap_8 FILLER_80_1788 ();
 sg13g2_decap_8 FILLER_80_1795 ();
 sg13g2_decap_8 FILLER_80_1802 ();
 sg13g2_decap_8 FILLER_80_1809 ();
 sg13g2_decap_8 FILLER_80_1816 ();
 sg13g2_decap_4 FILLER_80_1823 ();
 sg13g2_fill_1 FILLER_80_1827 ();
 sg13g2_decap_8 FILLER_80_1832 ();
 sg13g2_decap_8 FILLER_80_1839 ();
 sg13g2_decap_8 FILLER_80_1846 ();
 sg13g2_fill_1 FILLER_80_1853 ();
 sg13g2_fill_2 FILLER_80_1858 ();
 sg13g2_fill_1 FILLER_80_1860 ();
 sg13g2_decap_8 FILLER_80_1870 ();
 sg13g2_decap_8 FILLER_80_1877 ();
 sg13g2_decap_8 FILLER_80_1884 ();
 sg13g2_decap_8 FILLER_80_1891 ();
 sg13g2_decap_4 FILLER_80_1898 ();
 sg13g2_fill_2 FILLER_80_1902 ();
 sg13g2_fill_2 FILLER_80_1908 ();
 sg13g2_fill_1 FILLER_80_1910 ();
 sg13g2_fill_1 FILLER_80_1938 ();
 sg13g2_fill_2 FILLER_80_1967 ();
 sg13g2_decap_8 FILLER_80_1973 ();
 sg13g2_decap_8 FILLER_80_1989 ();
 sg13g2_decap_4 FILLER_80_1996 ();
 sg13g2_fill_2 FILLER_80_2000 ();
 sg13g2_decap_8 FILLER_80_2006 ();
 sg13g2_decap_8 FILLER_80_2013 ();
 sg13g2_fill_2 FILLER_80_2020 ();
 sg13g2_decap_8 FILLER_80_2081 ();
 sg13g2_decap_4 FILLER_80_2088 ();
 sg13g2_fill_1 FILLER_80_2092 ();
 sg13g2_fill_2 FILLER_80_2121 ();
 sg13g2_fill_1 FILLER_80_2123 ();
 sg13g2_decap_8 FILLER_80_2165 ();
 sg13g2_decap_8 FILLER_80_2172 ();
 sg13g2_decap_4 FILLER_80_2179 ();
 sg13g2_decap_8 FILLER_80_2187 ();
 sg13g2_decap_8 FILLER_80_2194 ();
 sg13g2_decap_8 FILLER_80_2201 ();
 sg13g2_decap_8 FILLER_80_2212 ();
 sg13g2_fill_2 FILLER_80_2219 ();
 sg13g2_fill_1 FILLER_80_2221 ();
 sg13g2_decap_8 FILLER_80_2231 ();
 sg13g2_decap_8 FILLER_80_2238 ();
 sg13g2_decap_8 FILLER_80_2245 ();
 sg13g2_decap_8 FILLER_80_2252 ();
 sg13g2_decap_8 FILLER_80_2259 ();
 sg13g2_decap_8 FILLER_80_2266 ();
 sg13g2_decap_8 FILLER_80_2273 ();
 sg13g2_decap_4 FILLER_80_2280 ();
 sg13g2_decap_8 FILLER_80_2288 ();
 sg13g2_decap_8 FILLER_80_2295 ();
 sg13g2_decap_8 FILLER_80_2302 ();
 sg13g2_fill_2 FILLER_80_2309 ();
 sg13g2_fill_1 FILLER_80_2311 ();
 sg13g2_decap_4 FILLER_80_2340 ();
 sg13g2_decap_4 FILLER_80_2372 ();
 sg13g2_fill_1 FILLER_80_2376 ();
 sg13g2_fill_1 FILLER_80_2405 ();
 sg13g2_decap_8 FILLER_80_2415 ();
 sg13g2_decap_8 FILLER_80_2422 ();
 sg13g2_decap_8 FILLER_80_2429 ();
 sg13g2_decap_8 FILLER_80_2436 ();
 sg13g2_fill_2 FILLER_80_2443 ();
 sg13g2_fill_1 FILLER_80_2445 ();
 sg13g2_decap_8 FILLER_80_2450 ();
 sg13g2_decap_8 FILLER_80_2457 ();
 sg13g2_fill_2 FILLER_80_2464 ();
 sg13g2_fill_1 FILLER_80_2466 ();
 sg13g2_decap_8 FILLER_80_2495 ();
 sg13g2_decap_8 FILLER_80_2502 ();
 sg13g2_decap_8 FILLER_80_2509 ();
 sg13g2_decap_8 FILLER_80_2516 ();
 sg13g2_decap_8 FILLER_80_2523 ();
 sg13g2_decap_8 FILLER_80_2530 ();
 sg13g2_decap_8 FILLER_80_2537 ();
 sg13g2_fill_2 FILLER_80_2544 ();
 sg13g2_decap_8 FILLER_80_2591 ();
 sg13g2_fill_2 FILLER_80_2598 ();
 sg13g2_fill_1 FILLER_80_2600 ();
 sg13g2_decap_4 FILLER_80_2629 ();
 sg13g2_fill_1 FILLER_80_2633 ();
 sg13g2_fill_2 FILLER_80_2662 ();
 sg13g2_fill_1 FILLER_80_2664 ();
 sg13g2_decap_8 FILLER_80_2669 ();
 sg13g2_decap_8 FILLER_80_2676 ();
 sg13g2_decap_8 FILLER_80_2683 ();
 sg13g2_decap_8 FILLER_80_2690 ();
 sg13g2_decap_4 FILLER_80_2697 ();
 sg13g2_decap_4 FILLER_80_2742 ();
 sg13g2_decap_4 FILLER_80_2778 ();
 sg13g2_fill_1 FILLER_80_2782 ();
 sg13g2_decap_8 FILLER_80_2820 ();
 sg13g2_decap_8 FILLER_80_2827 ();
 sg13g2_decap_8 FILLER_80_2834 ();
 sg13g2_decap_8 FILLER_80_2841 ();
 sg13g2_decap_8 FILLER_80_2848 ();
 sg13g2_decap_8 FILLER_80_2855 ();
 sg13g2_decap_8 FILLER_80_2862 ();
 sg13g2_decap_8 FILLER_80_2869 ();
 sg13g2_decap_8 FILLER_80_2876 ();
 sg13g2_decap_8 FILLER_80_2883 ();
 sg13g2_fill_1 FILLER_80_2890 ();
 sg13g2_decap_8 FILLER_80_2919 ();
 sg13g2_fill_2 FILLER_80_2926 ();
 sg13g2_fill_1 FILLER_80_2973 ();
 sg13g2_fill_2 FILLER_80_3002 ();
 sg13g2_decap_8 FILLER_80_3008 ();
 sg13g2_decap_8 FILLER_80_3015 ();
 sg13g2_decap_8 FILLER_80_3022 ();
 sg13g2_decap_8 FILLER_80_3029 ();
 sg13g2_decap_8 FILLER_80_3036 ();
 sg13g2_decap_8 FILLER_80_3043 ();
 sg13g2_decap_8 FILLER_80_3050 ();
 sg13g2_fill_1 FILLER_80_3057 ();
 sg13g2_fill_2 FILLER_80_3095 ();
 sg13g2_fill_1 FILLER_80_3097 ();
 sg13g2_decap_8 FILLER_80_3126 ();
 sg13g2_decap_8 FILLER_80_3133 ();
 sg13g2_decap_8 FILLER_80_3140 ();
 sg13g2_decap_8 FILLER_80_3147 ();
 sg13g2_decap_8 FILLER_80_3154 ();
 sg13g2_fill_2 FILLER_80_3161 ();
 sg13g2_fill_1 FILLER_80_3163 ();
 sg13g2_decap_8 FILLER_80_3168 ();
 sg13g2_decap_8 FILLER_80_3175 ();
 sg13g2_decap_8 FILLER_80_3182 ();
 sg13g2_decap_4 FILLER_80_3193 ();
 sg13g2_fill_1 FILLER_80_3197 ();
 sg13g2_decap_8 FILLER_80_3247 ();
 sg13g2_decap_8 FILLER_80_3254 ();
 sg13g2_decap_8 FILLER_80_3261 ();
 sg13g2_decap_8 FILLER_80_3268 ();
 sg13g2_decap_8 FILLER_80_3275 ();
 sg13g2_decap_8 FILLER_80_3282 ();
 sg13g2_decap_8 FILLER_80_3289 ();
 sg13g2_decap_8 FILLER_80_3296 ();
 sg13g2_decap_8 FILLER_80_3303 ();
 sg13g2_decap_8 FILLER_80_3310 ();
 sg13g2_decap_8 FILLER_80_3317 ();
 sg13g2_decap_8 FILLER_80_3324 ();
 sg13g2_decap_8 FILLER_80_3331 ();
 sg13g2_decap_8 FILLER_80_3338 ();
 sg13g2_decap_8 FILLER_80_3345 ();
 sg13g2_decap_8 FILLER_80_3352 ();
 sg13g2_decap_8 FILLER_80_3359 ();
 sg13g2_decap_8 FILLER_80_3366 ();
 sg13g2_decap_8 FILLER_80_3373 ();
 sg13g2_decap_8 FILLER_80_3380 ();
 sg13g2_decap_8 FILLER_80_3387 ();
 sg13g2_decap_8 FILLER_80_3394 ();
 sg13g2_decap_8 FILLER_80_3401 ();
 sg13g2_decap_8 FILLER_80_3408 ();
 sg13g2_decap_8 FILLER_80_3415 ();
 sg13g2_decap_8 FILLER_80_3422 ();
 sg13g2_decap_8 FILLER_80_3429 ();
 sg13g2_decap_8 FILLER_80_3436 ();
 sg13g2_decap_8 FILLER_80_3443 ();
 sg13g2_decap_8 FILLER_80_3450 ();
 sg13g2_decap_8 FILLER_80_3457 ();
 sg13g2_decap_8 FILLER_80_3464 ();
 sg13g2_decap_8 FILLER_80_3471 ();
 sg13g2_decap_8 FILLER_80_3478 ();
 sg13g2_decap_8 FILLER_80_3485 ();
 sg13g2_decap_8 FILLER_80_3492 ();
 sg13g2_decap_8 FILLER_80_3499 ();
 sg13g2_decap_8 FILLER_80_3506 ();
 sg13g2_decap_8 FILLER_80_3513 ();
 sg13g2_decap_8 FILLER_80_3520 ();
 sg13g2_decap_8 FILLER_80_3527 ();
 sg13g2_decap_8 FILLER_80_3534 ();
 sg13g2_decap_8 FILLER_80_3541 ();
 sg13g2_decap_8 FILLER_80_3548 ();
 sg13g2_decap_8 FILLER_80_3555 ();
 sg13g2_decap_8 FILLER_80_3562 ();
 sg13g2_decap_8 FILLER_80_3569 ();
 sg13g2_decap_4 FILLER_80_3576 ();
 assign uio_oe[0] = net1062;
 assign uio_oe[1] = net1063;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
endmodule
