module tt_um_jalcim (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire clknet_0_clk;
 wire \cam.found ;
 wire \cam.mem[0][0] ;
 wire \cam.mem[0][1] ;
 wire \cam.mem[0][2] ;
 wire \cam.mem[0][3] ;
 wire \cam.mem[0][4] ;
 wire \cam.mem[0][5] ;
 wire \cam.mem[0][6] ;
 wire \cam.mem[0][7] ;
 wire \cam.mem[10][0] ;
 wire \cam.mem[10][1] ;
 wire \cam.mem[10][2] ;
 wire \cam.mem[10][3] ;
 wire \cam.mem[10][4] ;
 wire \cam.mem[10][5] ;
 wire \cam.mem[10][6] ;
 wire \cam.mem[10][7] ;
 wire \cam.mem[11][0] ;
 wire \cam.mem[11][1] ;
 wire \cam.mem[11][2] ;
 wire \cam.mem[11][3] ;
 wire \cam.mem[11][4] ;
 wire \cam.mem[11][5] ;
 wire \cam.mem[11][6] ;
 wire \cam.mem[11][7] ;
 wire \cam.mem[12][0] ;
 wire \cam.mem[12][1] ;
 wire \cam.mem[12][2] ;
 wire \cam.mem[12][3] ;
 wire \cam.mem[12][4] ;
 wire \cam.mem[12][5] ;
 wire \cam.mem[12][6] ;
 wire \cam.mem[12][7] ;
 wire \cam.mem[13][0] ;
 wire \cam.mem[13][1] ;
 wire \cam.mem[13][2] ;
 wire \cam.mem[13][3] ;
 wire \cam.mem[13][4] ;
 wire \cam.mem[13][5] ;
 wire \cam.mem[13][6] ;
 wire \cam.mem[13][7] ;
 wire \cam.mem[14][0] ;
 wire \cam.mem[14][1] ;
 wire \cam.mem[14][2] ;
 wire \cam.mem[14][3] ;
 wire \cam.mem[14][4] ;
 wire \cam.mem[14][5] ;
 wire \cam.mem[14][6] ;
 wire \cam.mem[14][7] ;
 wire \cam.mem[15][0] ;
 wire \cam.mem[15][1] ;
 wire \cam.mem[15][2] ;
 wire \cam.mem[15][3] ;
 wire \cam.mem[15][4] ;
 wire \cam.mem[15][5] ;
 wire \cam.mem[15][6] ;
 wire \cam.mem[15][7] ;
 wire \cam.mem[1][0] ;
 wire \cam.mem[1][1] ;
 wire \cam.mem[1][2] ;
 wire \cam.mem[1][3] ;
 wire \cam.mem[1][4] ;
 wire \cam.mem[1][5] ;
 wire \cam.mem[1][6] ;
 wire \cam.mem[1][7] ;
 wire \cam.mem[2][0] ;
 wire \cam.mem[2][1] ;
 wire \cam.mem[2][2] ;
 wire \cam.mem[2][3] ;
 wire \cam.mem[2][4] ;
 wire \cam.mem[2][5] ;
 wire \cam.mem[2][6] ;
 wire \cam.mem[2][7] ;
 wire \cam.mem[3][0] ;
 wire \cam.mem[3][1] ;
 wire \cam.mem[3][2] ;
 wire \cam.mem[3][3] ;
 wire \cam.mem[3][4] ;
 wire \cam.mem[3][5] ;
 wire \cam.mem[3][6] ;
 wire \cam.mem[3][7] ;
 wire \cam.mem[4][0] ;
 wire \cam.mem[4][1] ;
 wire \cam.mem[4][2] ;
 wire \cam.mem[4][3] ;
 wire \cam.mem[4][4] ;
 wire \cam.mem[4][5] ;
 wire \cam.mem[4][6] ;
 wire \cam.mem[4][7] ;
 wire \cam.mem[5][0] ;
 wire \cam.mem[5][1] ;
 wire \cam.mem[5][2] ;
 wire \cam.mem[5][3] ;
 wire \cam.mem[5][4] ;
 wire \cam.mem[5][5] ;
 wire \cam.mem[5][6] ;
 wire \cam.mem[5][7] ;
 wire \cam.mem[6][0] ;
 wire \cam.mem[6][1] ;
 wire \cam.mem[6][2] ;
 wire \cam.mem[6][3] ;
 wire \cam.mem[6][4] ;
 wire \cam.mem[6][5] ;
 wire \cam.mem[6][6] ;
 wire \cam.mem[6][7] ;
 wire \cam.mem[7][0] ;
 wire \cam.mem[7][1] ;
 wire \cam.mem[7][2] ;
 wire \cam.mem[7][3] ;
 wire \cam.mem[7][4] ;
 wire \cam.mem[7][5] ;
 wire \cam.mem[7][6] ;
 wire \cam.mem[7][7] ;
 wire \cam.mem[8][0] ;
 wire \cam.mem[8][1] ;
 wire \cam.mem[8][2] ;
 wire \cam.mem[8][3] ;
 wire \cam.mem[8][4] ;
 wire \cam.mem[8][5] ;
 wire \cam.mem[8][6] ;
 wire \cam.mem[8][7] ;
 wire \cam.mem[9][0] ;
 wire \cam.mem[9][1] ;
 wire \cam.mem[9][2] ;
 wire \cam.mem[9][3] ;
 wire \cam.mem[9][4] ;
 wire \cam.mem[9][5] ;
 wire \cam.mem[9][6] ;
 wire \cam.mem[9][7] ;
 wire \fourhalt_latch.reg_n ;
 wire \fourhalt_latch.reg_p ;
 wire \onehalt_latch.reg_n ;
 wire \onehalt_latch.reg_p ;
 wire \treehalt_latch.reg_n ;
 wire \treehalt_latch.reg_p ;
 wire \twohalt_latch.reg_n ;
 wire \twohalt_latch.reg_p ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire \vga.counter[0] ;
 wire \vga.counter[1] ;
 wire \vga.counter[2] ;
 wire \vga.counter[3] ;
 wire \vga.counter[4] ;
 wire \vga.counter[5] ;
 wire \vga.counter[6] ;
 wire \vga.counter[7] ;
 wire \vga.hsync ;
 wire \vga.hvsync_gen.hpos[0] ;
 wire \vga.hvsync_gen.hpos[1] ;
 wire \vga.hvsync_gen.hpos[2] ;
 wire \vga.hvsync_gen.hpos[3] ;
 wire \vga.hvsync_gen.hpos[4] ;
 wire \vga.hvsync_gen.hpos[5] ;
 wire \vga.hvsync_gen.hpos[6] ;
 wire \vga.hvsync_gen.hpos[7] ;
 wire \vga.hvsync_gen.hpos[8] ;
 wire \vga.hvsync_gen.hpos[9] ;
 wire \vga.hvsync_gen.vpos[0] ;
 wire \vga.hvsync_gen.vpos[1] ;
 wire \vga.hvsync_gen.vpos[2] ;
 wire \vga.hvsync_gen.vpos[3] ;
 wire \vga.hvsync_gen.vpos[4] ;
 wire \vga.hvsync_gen.vpos[5] ;
 wire \vga.hvsync_gen.vpos[6] ;
 wire \vga.hvsync_gen.vpos[7] ;
 wire \vga.hvsync_gen.vpos[8] ;
 wire \vga.hvsync_gen.vpos[9] ;
 wire \vga.hvsync_gen.vsync ;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;

 sg13g2_inv_1 _0735_ (.Y(_0002_),
    .A(\vga.counter[0] ));
 sg13g2_inv_1 _0736_ (.Y(_0167_),
    .A(net188));
 sg13g2_inv_1 _0737_ (.Y(_0168_),
    .A(net190));
 sg13g2_inv_2 _0738_ (.Y(_0169_),
    .A(net172));
 sg13g2_inv_2 _0739_ (.Y(_0170_),
    .A(net168));
 sg13g2_inv_2 _0740_ (.Y(_0171_),
    .A(net154));
 sg13g2_inv_1 _0741_ (.Y(_0172_),
    .A(net151));
 sg13g2_inv_1 _0742_ (.Y(_0173_),
    .A(net275));
 sg13g2_inv_1 _0743_ (.Y(_0174_),
    .A(net285));
 sg13g2_inv_1 _0744_ (.Y(_0175_),
    .A(net274));
 sg13g2_inv_1 _0745_ (.Y(_0176_),
    .A(net251));
 sg13g2_inv_1 _0746_ (.Y(_0177_),
    .A(net292));
 sg13g2_inv_2 _0747_ (.Y(_0178_),
    .A(net246));
 sg13g2_inv_1 _0748_ (.Y(_0179_),
    .A(\vga.hvsync_gen.hpos[3] ));
 sg13g2_inv_1 _0749_ (.Y(_0180_),
    .A(\onehalt_latch.reg_p ));
 sg13g2_inv_1 _0750_ (.Y(_0181_),
    .A(\vga.counter[3] ));
 sg13g2_inv_1 _0751_ (.Y(_0182_),
    .A(net261));
 sg13g2_and3_1 _0752_ (.X(_0183_),
    .A(\vga.hvsync_gen.hpos[6] ),
    .B(\vga.hvsync_gen.hpos[5] ),
    .C(net407));
 sg13g2_nand2_1 _0753_ (.Y(_0184_),
    .A(\vga.hvsync_gen.hpos[7] ),
    .B(\vga.hvsync_gen.hpos[9] ));
 sg13g2_nor3_1 _0754_ (.A(\vga.hvsync_gen.hpos[6] ),
    .B(\vga.hvsync_gen.hpos[5] ),
    .C(net141),
    .Y(_0185_));
 sg13g2_nor4_1 _0755_ (.A(net249),
    .B(_0183_),
    .C(_0184_),
    .D(_0185_),
    .Y(_0000_));
 sg13g2_nand4_1 _0756_ (.B(\vga.hvsync_gen.vpos[6] ),
    .C(\vga.hvsync_gen.vpos[7] ),
    .A(\vga.hvsync_gen.vpos[5] ),
    .Y(_0186_),
    .D(\vga.hvsync_gen.vpos[8] ));
 sg13g2_nand2_1 _0757_ (.Y(_0187_),
    .A(\vga.hvsync_gen.vpos[3] ),
    .B(_0176_));
 sg13g2_nand2b_1 _0758_ (.Y(_0188_),
    .B(\vga.hvsync_gen.vpos[1] ),
    .A_N(\vga.hvsync_gen.vpos[2] ));
 sg13g2_nor4_1 _0759_ (.A(net246),
    .B(_0186_),
    .C(_0187_),
    .D(_0188_),
    .Y(_0001_));
 sg13g2_nor2_1 _0760_ (.A(\vga.hvsync_gen.hpos[5] ),
    .B(\vga.counter[5] ),
    .Y(_0189_));
 sg13g2_nand2_1 _0761_ (.Y(_0190_),
    .A(\vga.hvsync_gen.hpos[5] ),
    .B(\vga.counter[5] ));
 sg13g2_xor2_1 _0762_ (.B(\vga.counter[5] ),
    .A(\vga.hvsync_gen.hpos[5] ),
    .X(_0191_));
 sg13g2_nand2_1 _0763_ (.Y(_0192_),
    .A(net141),
    .B(\vga.counter[4] ));
 sg13g2_inv_1 _0764_ (.Y(_0193_),
    .A(_0192_));
 sg13g2_or2_1 _0765_ (.X(_0194_),
    .B(\vga.counter[4] ),
    .A(net141));
 sg13g2_a22oi_1 _0766_ (.Y(_0195_),
    .B1(\vga.hvsync_gen.hpos[1] ),
    .B2(\vga.counter[1] ),
    .A2(\vga.hvsync_gen.hpos[0] ),
    .A1(\vga.counter[0] ));
 sg13g2_nor2_1 _0767_ (.A(\vga.hvsync_gen.hpos[1] ),
    .B(\vga.counter[1] ),
    .Y(_0196_));
 sg13g2_nor2_1 _0768_ (.A(\vga.hvsync_gen.hpos[2] ),
    .B(\vga.counter[2] ),
    .Y(_0197_));
 sg13g2_or3_1 _0769_ (.A(_0195_),
    .B(_0196_),
    .C(_0197_),
    .X(_0198_));
 sg13g2_a22oi_1 _0770_ (.Y(_0199_),
    .B1(\vga.counter[2] ),
    .B2(\vga.hvsync_gen.hpos[2] ),
    .A2(\vga.counter[3] ),
    .A1(\vga.hvsync_gen.hpos[3] ));
 sg13g2_a22oi_1 _0771_ (.Y(_0200_),
    .B1(_0198_),
    .B2(_0199_),
    .A2(_0181_),
    .A1(_0179_));
 sg13g2_o21ai_1 _0772_ (.B1(_0194_),
    .Y(_0201_),
    .A1(_0193_),
    .A2(_0200_));
 sg13g2_nand2_1 _0773_ (.Y(_0202_),
    .A(\vga.hvsync_gen.hpos[9] ),
    .B(\vga.hvsync_gen.hpos[8] ));
 sg13g2_and4_1 _0774_ (.A(_0178_),
    .B(_0184_),
    .C(_0186_),
    .D(_0202_),
    .X(_0203_));
 sg13g2_nor2b_1 _0775_ (.A(net189),
    .B_N(_0203_),
    .Y(_0204_));
 sg13g2_xnor2_1 _0776_ (.Y(_0205_),
    .A(_0191_),
    .B(_0201_));
 sg13g2_and2_1 _0777_ (.A(net188),
    .B(net189),
    .X(_0206_));
 sg13g2_nand2_1 _0778_ (.Y(_0207_),
    .A(net6),
    .B(net145));
 sg13g2_and2_1 _0779_ (.A(net7),
    .B(_0207_),
    .X(_0208_));
 sg13g2_xor2_1 _0780_ (.B(\cam.mem[5][7] ),
    .A(net152),
    .X(_0209_));
 sg13g2_xor2_1 _0781_ (.B(\cam.mem[5][6] ),
    .A(net155),
    .X(_0210_));
 sg13g2_xor2_1 _0782_ (.B(\cam.mem[5][5] ),
    .A(net160),
    .X(_0211_));
 sg13g2_xor2_1 _0783_ (.B(\cam.mem[5][1] ),
    .A(net179),
    .X(_0212_));
 sg13g2_xor2_1 _0784_ (.B(\cam.mem[5][3] ),
    .A(net169),
    .X(_0213_));
 sg13g2_xor2_1 _0785_ (.B(\cam.mem[5][2] ),
    .A(net174),
    .X(_0214_));
 sg13g2_xor2_1 _0786_ (.B(\cam.mem[5][0] ),
    .A(net185),
    .X(_0215_));
 sg13g2_xor2_1 _0787_ (.B(\cam.mem[5][4] ),
    .A(net165),
    .X(_0216_));
 sg13g2_nor4_1 _0788_ (.A(_0209_),
    .B(_0210_),
    .C(_0213_),
    .D(_0215_),
    .Y(_0217_));
 sg13g2_nor4_2 _0789_ (.A(_0211_),
    .B(_0212_),
    .C(_0214_),
    .Y(_0218_),
    .D(_0216_));
 sg13g2_xor2_1 _0790_ (.B(net185),
    .A(\cam.mem[15][0] ),
    .X(_0219_));
 sg13g2_xor2_1 _0791_ (.B(\cam.mem[15][4] ),
    .A(net165),
    .X(_0220_));
 sg13g2_xor2_1 _0792_ (.B(\cam.mem[15][5] ),
    .A(net162),
    .X(_0221_));
 sg13g2_xor2_1 _0793_ (.B(net174),
    .A(\cam.mem[15][2] ),
    .X(_0222_));
 sg13g2_xor2_1 _0794_ (.B(\cam.mem[15][7] ),
    .A(net151),
    .X(_0223_));
 sg13g2_xor2_1 _0795_ (.B(\cam.mem[15][6] ),
    .A(net155),
    .X(_0224_));
 sg13g2_xor2_1 _0796_ (.B(net169),
    .A(\cam.mem[15][3] ),
    .X(_0225_));
 sg13g2_xor2_1 _0797_ (.B(net179),
    .A(\cam.mem[15][1] ),
    .X(_0226_));
 sg13g2_nor4_1 _0798_ (.A(_0221_),
    .B(_0223_),
    .C(_0224_),
    .D(_0225_),
    .Y(_0227_));
 sg13g2_nor4_2 _0799_ (.A(_0219_),
    .B(_0220_),
    .C(_0222_),
    .Y(_0228_),
    .D(_0226_));
 sg13g2_and2_1 _0800_ (.A(_0227_),
    .B(_0228_),
    .X(_0229_));
 sg13g2_a22oi_1 _0801_ (.Y(_0230_),
    .B1(_0227_),
    .B2(_0228_),
    .A2(_0218_),
    .A1(_0217_));
 sg13g2_xor2_1 _0802_ (.B(\cam.mem[13][3] ),
    .A(net168),
    .X(_0231_));
 sg13g2_xor2_1 _0803_ (.B(\cam.mem[13][7] ),
    .A(net149),
    .X(_0232_));
 sg13g2_xor2_1 _0804_ (.B(\cam.mem[13][1] ),
    .A(net176),
    .X(_0233_));
 sg13g2_xor2_1 _0805_ (.B(\cam.mem[13][6] ),
    .A(net154),
    .X(_0234_));
 sg13g2_xor2_1 _0806_ (.B(\cam.mem[13][2] ),
    .A(net172),
    .X(_0235_));
 sg13g2_xor2_1 _0807_ (.B(\cam.mem[13][4] ),
    .A(net163),
    .X(_0236_));
 sg13g2_xor2_1 _0808_ (.B(\cam.mem[13][5] ),
    .A(net158),
    .X(_0237_));
 sg13g2_xnor2_1 _0809_ (.Y(_0238_),
    .A(net183),
    .B(\cam.mem[13][0] ));
 sg13g2_nor4_1 _0810_ (.A(_0233_),
    .B(_0234_),
    .C(_0235_),
    .D(_0237_),
    .Y(_0239_));
 sg13g2_nor3_1 _0811_ (.A(_0231_),
    .B(_0232_),
    .C(_0236_),
    .Y(_0240_));
 sg13g2_nand3_1 _0812_ (.B(_0239_),
    .C(_0240_),
    .A(_0238_),
    .Y(_0241_));
 sg13g2_xor2_1 _0813_ (.B(\cam.mem[3][2] ),
    .A(net175),
    .X(_0242_));
 sg13g2_xor2_1 _0814_ (.B(\cam.mem[3][3] ),
    .A(net169),
    .X(_0243_));
 sg13g2_xor2_1 _0815_ (.B(\cam.mem[3][5] ),
    .A(net160),
    .X(_0244_));
 sg13g2_xor2_1 _0816_ (.B(\cam.mem[3][1] ),
    .A(net181),
    .X(_0245_));
 sg13g2_xor2_1 _0817_ (.B(\cam.mem[3][7] ),
    .A(net153),
    .X(_0246_));
 sg13g2_xor2_1 _0818_ (.B(\cam.mem[3][6] ),
    .A(net155),
    .X(_0247_));
 sg13g2_xnor2_1 _0819_ (.Y(_0248_),
    .A(net187),
    .B(\cam.mem[3][0] ));
 sg13g2_xor2_1 _0820_ (.B(\cam.mem[3][4] ),
    .A(net166),
    .X(_0249_));
 sg13g2_nor3_1 _0821_ (.A(_0242_),
    .B(_0246_),
    .C(_0247_),
    .Y(_0250_));
 sg13g2_nor4_1 _0822_ (.A(_0243_),
    .B(_0244_),
    .C(_0245_),
    .D(_0249_),
    .Y(_0251_));
 sg13g2_nand3_1 _0823_ (.B(_0250_),
    .C(_0251_),
    .A(_0248_),
    .Y(_0252_));
 sg13g2_nand3_1 _0824_ (.B(_0241_),
    .C(_0252_),
    .A(_0230_),
    .Y(_0253_));
 sg13g2_xor2_1 _0825_ (.B(\cam.mem[7][6] ),
    .A(net156),
    .X(_0254_));
 sg13g2_xor2_1 _0826_ (.B(\cam.mem[7][4] ),
    .A(net166),
    .X(_0255_));
 sg13g2_xnor2_1 _0827_ (.Y(_0256_),
    .A(net161),
    .B(\cam.mem[7][5] ));
 sg13g2_xor2_1 _0828_ (.B(\cam.mem[7][1] ),
    .A(net180),
    .X(_0257_));
 sg13g2_xor2_1 _0829_ (.B(\cam.mem[7][3] ),
    .A(net171),
    .X(_0258_));
 sg13g2_xor2_1 _0830_ (.B(\cam.mem[7][0] ),
    .A(net186),
    .X(_0259_));
 sg13g2_xor2_1 _0831_ (.B(\cam.mem[7][7] ),
    .A(net151),
    .X(_0260_));
 sg13g2_xor2_1 _0832_ (.B(\cam.mem[7][2] ),
    .A(net173),
    .X(_0261_));
 sg13g2_nor4_1 _0833_ (.A(_0254_),
    .B(_0255_),
    .C(_0258_),
    .D(_0260_),
    .Y(_0262_));
 sg13g2_nor3_1 _0834_ (.A(_0257_),
    .B(_0259_),
    .C(_0261_),
    .Y(_0263_));
 sg13g2_nand3_1 _0835_ (.B(_0262_),
    .C(_0263_),
    .A(_0256_),
    .Y(_0264_));
 sg13g2_xnor2_1 _0836_ (.Y(_0265_),
    .A(net175),
    .B(\cam.mem[1][2] ));
 sg13g2_xnor2_1 _0837_ (.Y(_0266_),
    .A(net184),
    .B(\cam.mem[1][0] ));
 sg13g2_xnor2_1 _0838_ (.Y(_0267_),
    .A(net150),
    .B(\cam.mem[1][7] ));
 sg13g2_xnor2_1 _0839_ (.Y(_0268_),
    .A(net159),
    .B(\cam.mem[1][5] ));
 sg13g2_xnor2_1 _0840_ (.Y(_0269_),
    .A(net164),
    .B(\cam.mem[1][4] ));
 sg13g2_xnor2_1 _0841_ (.Y(_0270_),
    .A(net171),
    .B(\cam.mem[1][3] ));
 sg13g2_xnor2_1 _0842_ (.Y(_0271_),
    .A(net157),
    .B(\cam.mem[1][6] ));
 sg13g2_xnor2_1 _0843_ (.Y(_0272_),
    .A(net178),
    .B(\cam.mem[1][1] ));
 sg13g2_nand4_1 _0844_ (.B(_0266_),
    .C(_0267_),
    .A(_0265_),
    .Y(_0273_),
    .D(_0271_));
 sg13g2_nand4_1 _0845_ (.B(_0269_),
    .C(_0270_),
    .A(_0268_),
    .Y(_0274_),
    .D(_0272_));
 sg13g2_o21ai_1 _0846_ (.B1(_0264_),
    .Y(_0275_),
    .A1(_0273_),
    .A2(_0274_));
 sg13g2_xor2_1 _0847_ (.B(\cam.mem[11][3] ),
    .A(net169),
    .X(_0276_));
 sg13g2_xor2_1 _0848_ (.B(\cam.mem[11][6] ),
    .A(net155),
    .X(_0277_));
 sg13g2_xnor2_1 _0849_ (.Y(_0278_),
    .A(net165),
    .B(\cam.mem[11][4] ));
 sg13g2_xor2_1 _0850_ (.B(\cam.mem[11][2] ),
    .A(net174),
    .X(_0279_));
 sg13g2_xor2_1 _0851_ (.B(\cam.mem[11][0] ),
    .A(net187),
    .X(_0280_));
 sg13g2_xor2_1 _0852_ (.B(\cam.mem[11][5] ),
    .A(net160),
    .X(_0281_));
 sg13g2_xor2_1 _0853_ (.B(\cam.mem[11][1] ),
    .A(net181),
    .X(_0282_));
 sg13g2_xor2_1 _0854_ (.B(\cam.mem[11][7] ),
    .A(net152),
    .X(_0283_));
 sg13g2_nor3_1 _0855_ (.A(_0276_),
    .B(_0280_),
    .C(_0282_),
    .Y(_0284_));
 sg13g2_nor4_1 _0856_ (.A(_0277_),
    .B(_0279_),
    .C(_0281_),
    .D(_0283_),
    .Y(_0285_));
 sg13g2_nand3_1 _0857_ (.B(_0284_),
    .C(_0285_),
    .A(_0278_),
    .Y(_0286_));
 sg13g2_xnor2_1 _0858_ (.Y(_0287_),
    .A(net179),
    .B(\cam.mem[9][1] ));
 sg13g2_xnor2_1 _0859_ (.Y(_0288_),
    .A(net185),
    .B(\cam.mem[9][0] ));
 sg13g2_xnor2_1 _0860_ (.Y(_0289_),
    .A(net152),
    .B(\cam.mem[9][7] ));
 sg13g2_xnor2_1 _0861_ (.Y(_0290_),
    .A(net160),
    .B(\cam.mem[9][5] ));
 sg13g2_xnor2_1 _0862_ (.Y(_0291_),
    .A(net169),
    .B(\cam.mem[9][3] ));
 sg13g2_xnor2_1 _0863_ (.Y(_0292_),
    .A(net165),
    .B(\cam.mem[9][4] ));
 sg13g2_xnor2_1 _0864_ (.Y(_0293_),
    .A(net155),
    .B(\cam.mem[9][6] ));
 sg13g2_xnor2_1 _0865_ (.Y(_0294_),
    .A(net174),
    .B(\cam.mem[9][2] ));
 sg13g2_nand4_1 _0866_ (.B(_0288_),
    .C(_0289_),
    .A(_0287_),
    .Y(_0295_),
    .D(_0293_));
 sg13g2_nand4_1 _0867_ (.B(_0291_),
    .C(_0292_),
    .A(_0290_),
    .Y(_0296_),
    .D(_0294_));
 sg13g2_o21ai_1 _0868_ (.B1(_0286_),
    .Y(_0297_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_or3_1 _0869_ (.A(_0253_),
    .B(_0275_),
    .C(_0297_),
    .X(_0298_));
 sg13g2_a22oi_1 _0870_ (.Y(_0299_),
    .B1(_0208_),
    .B2(_0298_),
    .A2(_0205_),
    .A1(_0204_));
 sg13g2_nor2_2 _0871_ (.A(net188),
    .B(net189),
    .Y(_0300_));
 sg13g2_or2_1 _0872_ (.X(_0301_),
    .B(net189),
    .A(net188));
 sg13g2_or2_1 _0873_ (.X(_0302_),
    .B(net186),
    .A(net2));
 sg13g2_nand2_1 _0874_ (.Y(_0303_),
    .A(net2),
    .B(net186));
 sg13g2_nand3_1 _0875_ (.B(_0302_),
    .C(_0303_),
    .A(_0300_),
    .Y(_0304_));
 sg13g2_or2_1 _0876_ (.X(_0305_),
    .B(_0304_),
    .A(_0172_));
 sg13g2_a21oi_1 _0877_ (.A1(_0172_),
    .A2(_0304_),
    .Y(_0306_),
    .B1(net189));
 sg13g2_and2_1 _0878_ (.A(net189),
    .B(\onehalt_latch.reg_n ),
    .X(_0307_));
 sg13g2_a221oi_1 _0879_ (.B2(_0180_),
    .C1(net188),
    .B1(_0307_),
    .A1(_0305_),
    .Y(_0308_),
    .A2(_0306_));
 sg13g2_a21oi_1 _0880_ (.A1(net188),
    .A2(_0299_),
    .Y(uo_out[0]),
    .B1(_0308_));
 sg13g2_nand3_1 _0881_ (.B(_0192_),
    .C(_0194_),
    .A(_0191_),
    .Y(_0309_));
 sg13g2_a221oi_1 _0882_ (.B2(_0199_),
    .C1(_0309_),
    .B1(_0198_),
    .A1(_0179_),
    .Y(_0310_),
    .A2(_0181_));
 sg13g2_o21ai_1 _0883_ (.B1(_0190_),
    .Y(_0311_),
    .A1(_0189_),
    .A2(_0192_));
 sg13g2_nand2_1 _0884_ (.Y(_0312_),
    .A(\vga.hvsync_gen.hpos[6] ),
    .B(\vga.counter[6] ));
 sg13g2_xor2_1 _0885_ (.B(\vga.counter[6] ),
    .A(\vga.hvsync_gen.hpos[6] ),
    .X(_0313_));
 sg13g2_o21ai_1 _0886_ (.B1(_0313_),
    .Y(_0314_),
    .A1(_0310_),
    .A2(_0311_));
 sg13g2_nor3_1 _0887_ (.A(_0310_),
    .B(_0311_),
    .C(_0313_),
    .Y(_0315_));
 sg13g2_nand3b_1 _0888_ (.B(_0204_),
    .C(_0314_),
    .Y(_0316_),
    .A_N(_0315_));
 sg13g2_xor2_1 _0889_ (.B(\cam.mem[6][3] ),
    .A(net170),
    .X(_0317_));
 sg13g2_xor2_1 _0890_ (.B(\cam.mem[6][6] ),
    .A(net156),
    .X(_0318_));
 sg13g2_xor2_1 _0891_ (.B(\cam.mem[6][5] ),
    .A(net161),
    .X(_0319_));
 sg13g2_xor2_1 _0892_ (.B(\cam.mem[6][7] ),
    .A(net151),
    .X(_0320_));
 sg13g2_xor2_1 _0893_ (.B(\cam.mem[6][0] ),
    .A(net186),
    .X(_0321_));
 sg13g2_xor2_1 _0894_ (.B(\cam.mem[6][2] ),
    .A(net173),
    .X(_0322_));
 sg13g2_xor2_1 _0895_ (.B(\cam.mem[6][4] ),
    .A(net166),
    .X(_0323_));
 sg13g2_xor2_1 _0896_ (.B(\cam.mem[6][1] ),
    .A(net180),
    .X(_0324_));
 sg13g2_nor4_1 _0897_ (.A(_0317_),
    .B(_0319_),
    .C(_0320_),
    .D(_0323_),
    .Y(_0325_));
 sg13g2_nor4_1 _0898_ (.A(_0318_),
    .B(_0321_),
    .C(_0322_),
    .D(_0324_),
    .Y(_0326_));
 sg13g2_a22oi_1 _0899_ (.Y(_0327_),
    .B1(_0325_),
    .B2(_0326_),
    .A2(_0228_),
    .A1(_0227_));
 sg13g2_xor2_1 _0900_ (.B(\cam.mem[2][3] ),
    .A(net170),
    .X(_0328_));
 sg13g2_xor2_1 _0901_ (.B(\cam.mem[2][0] ),
    .A(net186),
    .X(_0329_));
 sg13g2_xor2_1 _0902_ (.B(\cam.mem[2][6] ),
    .A(net156),
    .X(_0330_));
 sg13g2_xor2_1 _0903_ (.B(\cam.mem[2][7] ),
    .A(net151),
    .X(_0331_));
 sg13g2_xor2_1 _0904_ (.B(\cam.mem[2][2] ),
    .A(net173),
    .X(_0332_));
 sg13g2_xor2_1 _0905_ (.B(\cam.mem[2][4] ),
    .A(net166),
    .X(_0333_));
 sg13g2_xor2_1 _0906_ (.B(\cam.mem[2][5] ),
    .A(net161),
    .X(_0334_));
 sg13g2_xnor2_1 _0907_ (.Y(_0335_),
    .A(net180),
    .B(\cam.mem[2][1] ));
 sg13g2_nor4_1 _0908_ (.A(_0328_),
    .B(_0329_),
    .C(_0330_),
    .D(_0334_),
    .Y(_0336_));
 sg13g2_nor3_1 _0909_ (.A(_0331_),
    .B(_0332_),
    .C(_0333_),
    .Y(_0337_));
 sg13g2_nand3_1 _0910_ (.B(_0336_),
    .C(_0337_),
    .A(_0335_),
    .Y(_0338_));
 sg13g2_xor2_1 _0911_ (.B(\cam.mem[14][4] ),
    .A(net164),
    .X(_0339_));
 sg13g2_xor2_1 _0912_ (.B(\cam.mem[14][0] ),
    .A(net183),
    .X(_0340_));
 sg13g2_xor2_1 _0913_ (.B(\cam.mem[14][1] ),
    .A(net177),
    .X(_0341_));
 sg13g2_xor2_1 _0914_ (.B(\cam.mem[14][6] ),
    .A(net154),
    .X(_0342_));
 sg13g2_xor2_1 _0915_ (.B(\cam.mem[14][5] ),
    .A(net159),
    .X(_0343_));
 sg13g2_xor2_1 _0916_ (.B(\cam.mem[14][3] ),
    .A(net168),
    .X(_0344_));
 sg13g2_xnor2_1 _0917_ (.Y(_0345_),
    .A(net172),
    .B(\cam.mem[14][2] ));
 sg13g2_xor2_1 _0918_ (.B(\cam.mem[14][7] ),
    .A(net149),
    .X(_0346_));
 sg13g2_nor3_1 _0919_ (.A(_0339_),
    .B(_0341_),
    .C(_0343_),
    .Y(_0347_));
 sg13g2_nor4_1 _0920_ (.A(_0340_),
    .B(_0342_),
    .C(_0344_),
    .D(_0346_),
    .Y(_0348_));
 sg13g2_nand3_1 _0921_ (.B(_0347_),
    .C(_0348_),
    .A(_0345_),
    .Y(_0349_));
 sg13g2_xor2_1 _0922_ (.B(\cam.mem[10][4] ),
    .A(net165),
    .X(_0350_));
 sg13g2_xor2_1 _0923_ (.B(\cam.mem[10][1] ),
    .A(net179),
    .X(_0351_));
 sg13g2_xnor2_1 _0924_ (.Y(_0352_),
    .A(net169),
    .B(\cam.mem[10][3] ));
 sg13g2_xor2_1 _0925_ (.B(\cam.mem[10][5] ),
    .A(net160),
    .X(_0353_));
 sg13g2_xor2_1 _0926_ (.B(\cam.mem[10][2] ),
    .A(net174),
    .X(_0354_));
 sg13g2_xor2_1 _0927_ (.B(\cam.mem[10][0] ),
    .A(net185),
    .X(_0355_));
 sg13g2_xor2_1 _0928_ (.B(\cam.mem[10][6] ),
    .A(net155),
    .X(_0356_));
 sg13g2_xor2_1 _0929_ (.B(\cam.mem[10][7] ),
    .A(net152),
    .X(_0357_));
 sg13g2_nor3_1 _0930_ (.A(_0354_),
    .B(_0356_),
    .C(_0357_),
    .Y(_0358_));
 sg13g2_nor4_1 _0931_ (.A(_0350_),
    .B(_0351_),
    .C(_0353_),
    .D(_0355_),
    .Y(_0359_));
 sg13g2_nand3_1 _0932_ (.B(_0358_),
    .C(_0359_),
    .A(_0352_),
    .Y(_0360_));
 sg13g2_nand3_1 _0933_ (.B(_0327_),
    .C(_0349_),
    .A(_0264_),
    .Y(_0361_));
 sg13g2_and4_1 _0934_ (.A(_0252_),
    .B(_0286_),
    .C(_0338_),
    .D(_0360_),
    .X(_0362_));
 sg13g2_nand2b_1 _0935_ (.Y(_0363_),
    .B(_0362_),
    .A_N(_0361_));
 sg13g2_a21oi_1 _0936_ (.A1(_0208_),
    .A2(_0363_),
    .Y(_0364_),
    .B1(_0167_));
 sg13g2_nand2_1 _0937_ (.Y(_0365_),
    .A(net3),
    .B(net180));
 sg13g2_nor2_1 _0938_ (.A(net3),
    .B(net180),
    .Y(_0366_));
 sg13g2_nand3b_1 _0939_ (.B(_0300_),
    .C(_0365_),
    .Y(_0367_),
    .A_N(_0366_));
 sg13g2_o21ai_1 _0940_ (.B1(_0305_),
    .Y(_0368_),
    .A1(_0301_),
    .A2(_0303_));
 sg13g2_nor2b_1 _0941_ (.A(\onehalt_latch.reg_n ),
    .B_N(net7),
    .Y(_0369_));
 sg13g2_a21oi_1 _0942_ (.A1(\onehalt_latch.reg_p ),
    .A2(_0369_),
    .Y(_0370_),
    .B1(net188));
 sg13g2_xor2_1 _0943_ (.B(_0368_),
    .A(_0367_),
    .X(_0371_));
 sg13g2_a22oi_1 _0944_ (.Y(uo_out[1]),
    .B1(_0370_),
    .B2(_0371_),
    .A2(_0364_),
    .A1(_0316_));
 sg13g2_xnor2_1 _0945_ (.Y(_0372_),
    .A(\vga.hvsync_gen.hpos[7] ),
    .B(\vga.counter[7] ));
 sg13g2_a21o_1 _0946_ (.A2(_0314_),
    .A1(_0312_),
    .B1(_0372_),
    .X(_0373_));
 sg13g2_nand3_1 _0947_ (.B(_0314_),
    .C(_0372_),
    .A(_0312_),
    .Y(_0374_));
 sg13g2_nand3_1 _0948_ (.B(_0373_),
    .C(_0374_),
    .A(_0204_),
    .Y(_0375_));
 sg13g2_xor2_1 _0949_ (.B(\cam.mem[4][5] ),
    .A(net158),
    .X(_0376_));
 sg13g2_xor2_1 _0950_ (.B(\cam.mem[4][3] ),
    .A(net168),
    .X(_0377_));
 sg13g2_xor2_1 _0951_ (.B(\cam.mem[4][6] ),
    .A(net154),
    .X(_0378_));
 sg13g2_xor2_1 _0952_ (.B(\cam.mem[4][2] ),
    .A(net172),
    .X(_0379_));
 sg13g2_xor2_1 _0953_ (.B(\cam.mem[4][7] ),
    .A(net150),
    .X(_0380_));
 sg13g2_xor2_1 _0954_ (.B(\cam.mem[4][0] ),
    .A(net182),
    .X(_0381_));
 sg13g2_xor2_1 _0955_ (.B(\cam.mem[4][1] ),
    .A(net177),
    .X(_0382_));
 sg13g2_xor2_1 _0956_ (.B(\cam.mem[4][4] ),
    .A(net163),
    .X(_0383_));
 sg13g2_nor4_1 _0957_ (.A(_0378_),
    .B(_0379_),
    .C(_0380_),
    .D(_0381_),
    .Y(_0384_));
 sg13g2_nor4_1 _0958_ (.A(_0376_),
    .B(_0377_),
    .C(_0382_),
    .D(_0383_),
    .Y(_0385_));
 sg13g2_a22oi_1 _0959_ (.Y(_0386_),
    .B1(_0384_),
    .B2(_0385_),
    .A2(_0218_),
    .A1(_0217_));
 sg13g2_xor2_1 _0960_ (.B(\cam.mem[12][3] ),
    .A(net168),
    .X(_0387_));
 sg13g2_xnor2_1 _0961_ (.Y(_0388_),
    .A(net163),
    .B(\cam.mem[12][4] ));
 sg13g2_xor2_1 _0962_ (.B(\cam.mem[12][6] ),
    .A(net154),
    .X(_0389_));
 sg13g2_xor2_1 _0963_ (.B(\cam.mem[12][5] ),
    .A(net158),
    .X(_0390_));
 sg13g2_xor2_1 _0964_ (.B(\cam.mem[12][2] ),
    .A(net172),
    .X(_0391_));
 sg13g2_xor2_1 _0965_ (.B(\cam.mem[12][0] ),
    .A(net182),
    .X(_0392_));
 sg13g2_xor2_1 _0966_ (.B(\cam.mem[12][7] ),
    .A(net149),
    .X(_0393_));
 sg13g2_xor2_1 _0967_ (.B(\cam.mem[12][1] ),
    .A(net176),
    .X(_0394_));
 sg13g2_nor4_1 _0968_ (.A(_0387_),
    .B(_0391_),
    .C(_0392_),
    .D(_0393_),
    .Y(_0395_));
 sg13g2_nor3_1 _0969_ (.A(_0389_),
    .B(_0390_),
    .C(_0394_),
    .Y(_0396_));
 sg13g2_nand3_1 _0970_ (.B(_0395_),
    .C(_0396_),
    .A(_0388_),
    .Y(_0397_));
 sg13g2_nand3_1 _0971_ (.B(_0386_),
    .C(_0397_),
    .A(_0241_),
    .Y(_0398_));
 sg13g2_o21ai_1 _0972_ (.B1(_0208_),
    .Y(_0399_),
    .A1(_0361_),
    .A2(_0398_));
 sg13g2_and2_1 _0973_ (.A(net188),
    .B(_0399_),
    .X(_0400_));
 sg13g2_and2_1 _0974_ (.A(net4),
    .B(net173),
    .X(_0401_));
 sg13g2_nor2_1 _0975_ (.A(_0301_),
    .B(_0401_),
    .Y(_0402_));
 sg13g2_o21ai_1 _0976_ (.B1(_0402_),
    .Y(_0403_),
    .A1(net4),
    .A2(net173));
 sg13g2_inv_1 _0977_ (.Y(_0404_),
    .A(_0403_));
 sg13g2_nand2_1 _0978_ (.Y(_0405_),
    .A(_0303_),
    .B(_0365_));
 sg13g2_nand3b_1 _0979_ (.B(_0405_),
    .C(_0300_),
    .Y(_0406_),
    .A_N(_0366_));
 sg13g2_o21ai_1 _0980_ (.B1(_0406_),
    .Y(_0407_),
    .A1(_0305_),
    .A2(_0367_));
 sg13g2_xnor2_1 _0981_ (.Y(_0408_),
    .A(_0403_),
    .B(_0407_));
 sg13g2_nand3b_1 _0982_ (.B(\twohalt_latch.reg_n ),
    .C(net189),
    .Y(_0409_),
    .A_N(\twohalt_latch.reg_p ));
 sg13g2_nor2b_1 _0983_ (.A(_0408_),
    .B_N(_0409_),
    .Y(_0410_));
 sg13g2_a22oi_1 _0984_ (.Y(uo_out[2]),
    .B1(_0410_),
    .B2(_0167_),
    .A2(_0400_),
    .A1(_0375_));
 sg13g2_or2_1 _0985_ (.X(_0411_),
    .B(net170),
    .A(net5));
 sg13g2_nand2_1 _0986_ (.Y(_0412_),
    .A(net5),
    .B(net170));
 sg13g2_nand3_1 _0987_ (.B(_0411_),
    .C(_0412_),
    .A(_0300_),
    .Y(_0413_));
 sg13g2_a22oi_1 _0988_ (.Y(_0414_),
    .B1(_0404_),
    .B2(_0407_),
    .A2(_0401_),
    .A1(_0300_));
 sg13g2_xnor2_1 _0989_ (.Y(_0415_),
    .A(_0413_),
    .B(_0414_));
 sg13g2_xnor2_1 _0990_ (.Y(_0416_),
    .A(net154),
    .B(\cam.mem[8][6] ));
 sg13g2_xnor2_1 _0991_ (.Y(_0417_),
    .A(net168),
    .B(\cam.mem[8][3] ));
 sg13g2_xnor2_1 _0992_ (.Y(_0418_),
    .A(net158),
    .B(\cam.mem[8][5] ));
 sg13g2_xnor2_1 _0993_ (.Y(_0419_),
    .A(net176),
    .B(\cam.mem[8][1] ));
 sg13g2_xnor2_1 _0994_ (.Y(_0420_),
    .A(net172),
    .B(\cam.mem[8][2] ));
 sg13g2_xnor2_1 _0995_ (.Y(_0421_),
    .A(net182),
    .B(\cam.mem[8][0] ));
 sg13g2_xor2_1 _0996_ (.B(\cam.mem[8][4] ),
    .A(net163),
    .X(_0422_));
 sg13g2_xnor2_1 _0997_ (.Y(_0423_),
    .A(net149),
    .B(\cam.mem[8][7] ));
 sg13g2_nand4_1 _0998_ (.B(_0418_),
    .C(_0420_),
    .A(_0416_),
    .Y(_0424_),
    .D(_0421_));
 sg13g2_nand3_1 _0999_ (.B(_0419_),
    .C(_0423_),
    .A(_0417_),
    .Y(_0425_));
 sg13g2_nor3_1 _1000_ (.A(_0422_),
    .B(_0424_),
    .C(_0425_),
    .Y(_0426_));
 sg13g2_nand4_1 _1001_ (.B(_0349_),
    .C(_0360_),
    .A(_0241_),
    .Y(_0427_),
    .D(_0397_));
 sg13g2_or3_1 _1002_ (.A(_0297_),
    .B(_0426_),
    .C(_0427_),
    .X(_0428_));
 sg13g2_nor2b_1 _1003_ (.A(net6),
    .B_N(net145),
    .Y(_0429_));
 sg13g2_o21ai_1 _1004_ (.B1(_0429_),
    .Y(_0430_),
    .A1(_0229_),
    .A2(_0428_));
 sg13g2_nor2_2 _1005_ (.A(_0167_),
    .B(net189),
    .Y(_0431_));
 sg13g2_nor2b_1 _1006_ (.A(net8),
    .B_N(net7),
    .Y(_0432_));
 sg13g2_nor2b_1 _1007_ (.A(\twohalt_latch.reg_n ),
    .B_N(\twohalt_latch.reg_p ),
    .Y(_0433_));
 sg13g2_a22oi_1 _1008_ (.Y(_0434_),
    .B1(net143),
    .B2(_0433_),
    .A2(_0431_),
    .A1(net142));
 sg13g2_nand3_1 _1009_ (.B(_0430_),
    .C(_0434_),
    .A(_0415_),
    .Y(uo_out[3]));
 sg13g2_o21ai_1 _1010_ (.B1(_0412_),
    .Y(_0435_),
    .A1(_0413_),
    .A2(_0414_));
 sg13g2_nand3b_1 _1011_ (.B(net143),
    .C(\treehalt_latch.reg_n ),
    .Y(_0436_),
    .A_N(\treehalt_latch.reg_p ));
 sg13g2_nand3_1 _1012_ (.B(_0203_),
    .C(_0431_),
    .A(\vga.hvsync_gen.vpos[2] ),
    .Y(_0437_));
 sg13g2_nand2_1 _1013_ (.Y(_0438_),
    .A(_0436_),
    .B(_0437_));
 sg13g2_a21o_2 _1014_ (.A2(_0435_),
    .A1(_0300_),
    .B1(_0438_),
    .X(uo_out[4]));
 sg13g2_nor2b_1 _1015_ (.A(\treehalt_latch.reg_n ),
    .B_N(\treehalt_latch.reg_p ),
    .Y(_0439_));
 sg13g2_a22oi_1 _1016_ (.Y(_0440_),
    .B1(net144),
    .B2(_0439_),
    .A2(_0206_),
    .A1(\cam.found ));
 sg13g2_nand2_1 _1017_ (.Y(uo_out[5]),
    .A(_0437_),
    .B(_0440_));
 sg13g2_nand2_1 _1018_ (.Y(_0441_),
    .A(\fourhalt_latch.reg_n ),
    .B(net143));
 sg13g2_nand3_1 _1019_ (.B(_0203_),
    .C(_0431_),
    .A(\vga.hvsync_gen.vpos[5] ),
    .Y(_0442_));
 sg13g2_o21ai_1 _1020_ (.B1(_0442_),
    .Y(uo_out[6]),
    .A1(\fourhalt_latch.reg_p ),
    .A2(_0441_));
 sg13g2_nor2b_1 _1021_ (.A(\fourhalt_latch.reg_n ),
    .B_N(\fourhalt_latch.reg_p ),
    .Y(_0443_));
 sg13g2_a22oi_1 _1022_ (.Y(_0444_),
    .B1(net143),
    .B2(_0443_),
    .A2(_0431_),
    .A1(\vga.hsync ));
 sg13g2_inv_1 _1023_ (.Y(uo_out[7]),
    .A(_0444_));
 sg13g2_xor2_1 _1024_ (.B(\vga.counter[1] ),
    .A(\vga.counter[0] ),
    .X(_0003_));
 sg13g2_nand3_1 _1025_ (.B(\vga.counter[2] ),
    .C(\vga.counter[1] ),
    .A(\vga.counter[0] ),
    .Y(_0445_));
 sg13g2_a21o_1 _1026_ (.A2(\vga.counter[1] ),
    .A1(\vga.counter[0] ),
    .B1(\vga.counter[2] ),
    .X(_0446_));
 sg13g2_and2_1 _1027_ (.A(_0445_),
    .B(_0446_),
    .X(_0004_));
 sg13g2_nor2_2 _1028_ (.A(_0181_),
    .B(_0445_),
    .Y(_0447_));
 sg13g2_xnor2_1 _1029_ (.Y(_0005_),
    .A(\vga.counter[3] ),
    .B(_0445_));
 sg13g2_xor2_1 _1030_ (.B(_0447_),
    .A(\vga.counter[4] ),
    .X(_0006_));
 sg13g2_nand3_1 _1031_ (.B(\vga.counter[4] ),
    .C(_0447_),
    .A(\vga.counter[5] ),
    .Y(_0448_));
 sg13g2_a21o_1 _1032_ (.A2(_0447_),
    .A1(\vga.counter[4] ),
    .B1(\vga.counter[5] ),
    .X(_0449_));
 sg13g2_and2_1 _1033_ (.A(_0448_),
    .B(_0449_),
    .X(_0007_));
 sg13g2_nand4_1 _1034_ (.B(\vga.counter[4] ),
    .C(\vga.counter[6] ),
    .A(\vga.counter[5] ),
    .Y(_0450_),
    .D(_0447_));
 sg13g2_xnor2_1 _1035_ (.Y(_0008_),
    .A(\vga.counter[6] ),
    .B(_0448_));
 sg13g2_xnor2_1 _1036_ (.Y(_0009_),
    .A(\vga.counter[7] ),
    .B(_0450_));
 sg13g2_and2_1 _1037_ (.A(net171),
    .B(net143),
    .X(_0010_));
 sg13g2_and2_1 _1038_ (.A(net248),
    .B(net389),
    .X(_0451_));
 sg13g2_and3_2 _1039_ (.X(_0452_),
    .A(net297),
    .B(net262),
    .C(_0451_));
 sg13g2_nor4_1 _1040_ (.A(\vga.hvsync_gen.hpos[7] ),
    .B(\vga.hvsync_gen.hpos[6] ),
    .C(\vga.hvsync_gen.hpos[5] ),
    .D(_0202_),
    .Y(_0453_));
 sg13g2_nand3_1 _1041_ (.B(_0452_),
    .C(_0453_),
    .A(net141),
    .Y(_0454_));
 sg13g2_nor4_1 _1042_ (.A(\vga.hvsync_gen.vpos[6] ),
    .B(\vga.hvsync_gen.vpos[7] ),
    .C(\vga.hvsync_gen.vpos[8] ),
    .D(_0178_),
    .Y(_0455_));
 sg13g2_nand2b_1 _1043_ (.Y(_0456_),
    .B(\vga.hvsync_gen.vpos[2] ),
    .A_N(\vga.hvsync_gen.vpos[5] ));
 sg13g2_nor4_1 _1044_ (.A(\vga.hvsync_gen.vpos[0] ),
    .B(\vga.hvsync_gen.vpos[1] ),
    .C(_0187_),
    .D(_0456_),
    .Y(_0457_));
 sg13g2_a21o_1 _1045_ (.A2(_0457_),
    .A1(_0455_),
    .B1(_0168_),
    .X(_0458_));
 sg13g2_nor2_1 _1046_ (.A(_0454_),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_or2_1 _1047_ (.X(_0460_),
    .B(_0458_),
    .A(_0454_));
 sg13g2_nor2_1 _1048_ (.A(net296),
    .B(_0459_),
    .Y(_0461_));
 sg13g2_and2_1 _1049_ (.A(net190),
    .B(_0454_),
    .X(_0462_));
 sg13g2_nand2_2 _1050_ (.Y(_0463_),
    .A(net190),
    .B(_0454_));
 sg13g2_a21oi_1 _1051_ (.A1(net296),
    .A2(_0463_),
    .Y(_0011_),
    .B1(_0461_));
 sg13g2_nand2_1 _1052_ (.Y(_0464_),
    .A(net380),
    .B(net136));
 sg13g2_xnor2_1 _1053_ (.Y(_0465_),
    .A(net296),
    .B(net380));
 sg13g2_o21ai_1 _1054_ (.B1(_0464_),
    .Y(_0012_),
    .A1(_0460_),
    .A2(_0465_));
 sg13g2_nand2_1 _1055_ (.Y(_0466_),
    .A(net374),
    .B(net136));
 sg13g2_a21oi_1 _1056_ (.A1(net296),
    .A2(\vga.hvsync_gen.vpos[1] ),
    .Y(_0467_),
    .B1(net374));
 sg13g2_nand3_1 _1057_ (.B(\vga.hvsync_gen.vpos[1] ),
    .C(net374),
    .A(net296),
    .Y(_0468_));
 sg13g2_nand2b_1 _1058_ (.Y(_0469_),
    .B(_0468_),
    .A_N(_0467_));
 sg13g2_o21ai_1 _1059_ (.B1(_0466_),
    .Y(_0013_),
    .A1(_0460_),
    .A2(_0469_));
 sg13g2_nand2_1 _1060_ (.Y(_0470_),
    .A(net280),
    .B(net136));
 sg13g2_nand4_1 _1061_ (.B(net380),
    .C(net374),
    .A(net296),
    .Y(_0471_),
    .D(net280));
 sg13g2_xor2_1 _1062_ (.B(_0468_),
    .A(net280),
    .X(_0472_));
 sg13g2_o21ai_1 _1063_ (.B1(_0470_),
    .Y(_0014_),
    .A1(_0460_),
    .A2(_0472_));
 sg13g2_nand2_1 _1064_ (.Y(_0473_),
    .A(net251),
    .B(net136));
 sg13g2_nor2_1 _1065_ (.A(_0176_),
    .B(_0471_),
    .Y(_0474_));
 sg13g2_xnor2_1 _1066_ (.Y(_0475_),
    .A(_0176_),
    .B(_0471_));
 sg13g2_o21ai_1 _1067_ (.B1(_0473_),
    .Y(_0015_),
    .A1(_0460_),
    .A2(_0475_));
 sg13g2_nand2_1 _1068_ (.Y(_0476_),
    .A(net294),
    .B(net136));
 sg13g2_xnor2_1 _1069_ (.Y(_0477_),
    .A(net294),
    .B(_0474_));
 sg13g2_o21ai_1 _1070_ (.B1(_0476_),
    .Y(_0016_),
    .A1(_0460_),
    .A2(_0477_));
 sg13g2_nand2_1 _1071_ (.Y(_0478_),
    .A(net287),
    .B(net136));
 sg13g2_nand3_1 _1072_ (.B(net287),
    .C(_0474_),
    .A(net294),
    .Y(_0479_));
 sg13g2_a21o_1 _1073_ (.A2(_0474_),
    .A1(\vga.hvsync_gen.vpos[5] ),
    .B1(net287),
    .X(_0480_));
 sg13g2_nand2_1 _1074_ (.Y(_0481_),
    .A(_0479_),
    .B(_0480_));
 sg13g2_o21ai_1 _1075_ (.B1(_0478_),
    .Y(_0017_),
    .A1(_0460_),
    .A2(_0481_));
 sg13g2_nand2_1 _1076_ (.Y(_0482_),
    .A(net292),
    .B(net136));
 sg13g2_nor2_1 _1077_ (.A(_0177_),
    .B(_0479_),
    .Y(_0483_));
 sg13g2_xor2_1 _1078_ (.B(_0479_),
    .A(net292),
    .X(_0484_));
 sg13g2_o21ai_1 _1079_ (.B1(_0482_),
    .Y(_0018_),
    .A1(_0460_),
    .A2(_0484_));
 sg13g2_nand2_1 _1080_ (.Y(_0485_),
    .A(net282),
    .B(_0483_));
 sg13g2_a21oi_1 _1081_ (.A1(_0459_),
    .A2(_0485_),
    .Y(_0486_),
    .B1(_0462_));
 sg13g2_a21oi_1 _1082_ (.A1(_0459_),
    .A2(_0483_),
    .Y(_0487_),
    .B1(net282));
 sg13g2_nor2_1 _1083_ (.A(_0486_),
    .B(net283),
    .Y(_0019_));
 sg13g2_nand4_1 _1084_ (.B(_0178_),
    .C(_0459_),
    .A(net282),
    .Y(_0488_),
    .D(_0483_));
 sg13g2_o21ai_1 _1085_ (.B1(_0488_),
    .Y(_0020_),
    .A1(_0178_),
    .A2(_0486_));
 sg13g2_nand2_1 _1086_ (.Y(_0489_),
    .A(net5),
    .B(net145));
 sg13g2_nor2_2 _1087_ (.A(net4),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_nand4_1 _1088_ (.B(net1),
    .C(net192),
    .A(net6),
    .Y(_0491_),
    .D(net145));
 sg13g2_inv_1 _1089_ (.Y(_0492_),
    .A(_0491_));
 sg13g2_nand2_2 _1090_ (.Y(_0493_),
    .A(net3),
    .B(_0492_));
 sg13g2_nor2_2 _1091_ (.A(net2),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_nand2_2 _1092_ (.Y(_0495_),
    .A(_0490_),
    .B(_0494_));
 sg13g2_mux2_1 _1093_ (.A0(net185),
    .A1(net337),
    .S(_0495_),
    .X(_0021_));
 sg13g2_mux2_1 _1094_ (.A0(net179),
    .A1(net307),
    .S(_0495_),
    .X(_0022_));
 sg13g2_mux2_1 _1095_ (.A0(net174),
    .A1(net382),
    .S(_0495_),
    .X(_0023_));
 sg13g2_mux2_1 _1096_ (.A0(net169),
    .A1(net329),
    .S(_0495_),
    .X(_0024_));
 sg13g2_mux2_1 _1097_ (.A0(net166),
    .A1(net312),
    .S(_0495_),
    .X(_0025_));
 sg13g2_mux2_1 _1098_ (.A0(net161),
    .A1(net391),
    .S(_0495_),
    .X(_0026_));
 sg13g2_mux2_1 _1099_ (.A0(net155),
    .A1(net342),
    .S(_0495_),
    .X(_0027_));
 sg13g2_mux2_1 _1100_ (.A0(net152),
    .A1(net377),
    .S(_0495_),
    .X(_0028_));
 sg13g2_nand2_1 _1101_ (.Y(_0496_),
    .A(net4),
    .B(net145));
 sg13g2_nand3_1 _1102_ (.B(net5),
    .C(net145),
    .A(net4),
    .Y(_0497_));
 sg13g2_nand2_2 _1103_ (.Y(_0498_),
    .A(net2),
    .B(net145));
 sg13g2_inv_1 _1104_ (.Y(_0499_),
    .A(_0498_));
 sg13g2_nor3_2 _1105_ (.A(net3),
    .B(_0491_),
    .C(_0499_),
    .Y(_0500_));
 sg13g2_nor2b_2 _1106_ (.A(_0497_),
    .B_N(_0500_),
    .Y(_0501_));
 sg13g2_mux2_1 _1107_ (.A0(net305),
    .A1(net182),
    .S(net135),
    .X(_0029_));
 sg13g2_mux2_1 _1108_ (.A0(net385),
    .A1(net176),
    .S(net135),
    .X(_0030_));
 sg13g2_nor2_1 _1109_ (.A(net286),
    .B(net135),
    .Y(_0502_));
 sg13g2_a21oi_1 _1110_ (.A1(net148),
    .A2(net135),
    .Y(_0031_),
    .B1(_0502_));
 sg13g2_nor2_1 _1111_ (.A(net276),
    .B(net135),
    .Y(_0503_));
 sg13g2_a21oi_1 _1112_ (.A1(net147),
    .A2(_0501_),
    .Y(_0032_),
    .B1(_0503_));
 sg13g2_mux2_1 _1113_ (.A0(net343),
    .A1(net163),
    .S(net135),
    .X(_0033_));
 sg13g2_mux2_1 _1114_ (.A0(net360),
    .A1(net158),
    .S(net135),
    .X(_0034_));
 sg13g2_nor2_1 _1115_ (.A(net291),
    .B(_0501_),
    .Y(_0504_));
 sg13g2_a21oi_1 _1116_ (.A1(net146),
    .A2(_0501_),
    .Y(_0035_),
    .B1(_0504_));
 sg13g2_mux2_1 _1117_ (.A0(net353),
    .A1(net149),
    .S(net135),
    .X(_0036_));
 sg13g2_nor3_2 _1118_ (.A(net3),
    .B(_0491_),
    .C(_0498_),
    .Y(_0505_));
 sg13g2_nand2_2 _1119_ (.Y(_0506_),
    .A(_0490_),
    .B(_0505_));
 sg13g2_mux2_1 _1120_ (.A0(net185),
    .A1(net315),
    .S(_0506_),
    .X(_0037_));
 sg13g2_mux2_1 _1121_ (.A0(net179),
    .A1(net384),
    .S(net140),
    .X(_0038_));
 sg13g2_nand2_1 _1122_ (.Y(_0507_),
    .A(net254),
    .B(net140));
 sg13g2_o21ai_1 _1123_ (.B1(_0507_),
    .Y(_0039_),
    .A1(net148),
    .A2(net140));
 sg13g2_nand2_1 _1124_ (.Y(_0508_),
    .A(net266),
    .B(net140));
 sg13g2_o21ai_1 _1125_ (.B1(_0508_),
    .Y(_0040_),
    .A1(net147),
    .A2(net140));
 sg13g2_mux2_1 _1126_ (.A0(net165),
    .A1(net313),
    .S(net140),
    .X(_0041_));
 sg13g2_mux2_1 _1127_ (.A0(net160),
    .A1(net334),
    .S(_0506_),
    .X(_0042_));
 sg13g2_nand2_1 _1128_ (.Y(_0509_),
    .A(net270),
    .B(net140));
 sg13g2_o21ai_1 _1129_ (.B1(_0509_),
    .Y(_0043_),
    .A1(net146),
    .A2(net140));
 sg13g2_mux2_1 _1130_ (.A0(net152),
    .A1(net388),
    .S(_0506_),
    .X(_0044_));
 sg13g2_nand2_2 _1131_ (.Y(_0510_),
    .A(_0490_),
    .B(_0500_));
 sg13g2_mux2_1 _1132_ (.A0(net182),
    .A1(net393),
    .S(net134),
    .X(_0045_));
 sg13g2_mux2_1 _1133_ (.A0(net176),
    .A1(net326),
    .S(net134),
    .X(_0046_));
 sg13g2_nand2_1 _1134_ (.Y(_0511_),
    .A(net255),
    .B(net134));
 sg13g2_o21ai_1 _1135_ (.B1(_0511_),
    .Y(_0047_),
    .A1(net148),
    .A2(net134));
 sg13g2_nand2_1 _1136_ (.Y(_0512_),
    .A(net269),
    .B(net134));
 sg13g2_o21ai_1 _1137_ (.B1(_0512_),
    .Y(_0048_),
    .A1(net147),
    .A2(_0510_));
 sg13g2_mux2_1 _1138_ (.A0(net163),
    .A1(net328),
    .S(net134),
    .X(_0049_));
 sg13g2_mux2_1 _1139_ (.A0(net158),
    .A1(net308),
    .S(net134),
    .X(_0050_));
 sg13g2_nand2_1 _1140_ (.Y(_0513_),
    .A(net267),
    .B(_0510_));
 sg13g2_o21ai_1 _1141_ (.B1(_0513_),
    .Y(_0051_),
    .A1(net146),
    .A2(_0510_));
 sg13g2_mux2_1 _1142_ (.A0(net149),
    .A1(net349),
    .S(net134),
    .X(_0052_));
 sg13g2_nor2_2 _1143_ (.A(net5),
    .B(_0496_),
    .Y(_0514_));
 sg13g2_nor2_2 _1144_ (.A(_0493_),
    .B(_0498_),
    .Y(_0515_));
 sg13g2_nand2_2 _1145_ (.Y(_0516_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_mux2_1 _1146_ (.A0(net186),
    .A1(net323),
    .S(_0516_),
    .X(_0053_));
 sg13g2_mux2_1 _1147_ (.A0(net180),
    .A1(net361),
    .S(_0516_),
    .X(_0054_));
 sg13g2_mux2_1 _1148_ (.A0(net173),
    .A1(net376),
    .S(_0516_),
    .X(_0055_));
 sg13g2_mux2_1 _1149_ (.A0(net171),
    .A1(net338),
    .S(_0516_),
    .X(_0056_));
 sg13g2_mux2_1 _1150_ (.A0(net166),
    .A1(net395),
    .S(_0516_),
    .X(_0057_));
 sg13g2_mux2_1 _1151_ (.A0(net161),
    .A1(net316),
    .S(_0516_),
    .X(_0058_));
 sg13g2_mux2_1 _1152_ (.A0(net156),
    .A1(net392),
    .S(_0516_),
    .X(_0059_));
 sg13g2_mux2_1 _1153_ (.A0(net151),
    .A1(net369),
    .S(_0516_),
    .X(_0060_));
 sg13g2_nand2_2 _1154_ (.Y(_0517_),
    .A(_0494_),
    .B(_0514_));
 sg13g2_mux2_1 _1155_ (.A0(net186),
    .A1(net368),
    .S(_0517_),
    .X(_0061_));
 sg13g2_mux2_1 _1156_ (.A0(net180),
    .A1(net394),
    .S(_0517_),
    .X(_0062_));
 sg13g2_mux2_1 _1157_ (.A0(net173),
    .A1(net317),
    .S(_0517_),
    .X(_0063_));
 sg13g2_mux2_1 _1158_ (.A0(net170),
    .A1(net331),
    .S(_0517_),
    .X(_0064_));
 sg13g2_mux2_1 _1159_ (.A0(net167),
    .A1(net345),
    .S(_0517_),
    .X(_0065_));
 sg13g2_mux2_1 _1160_ (.A0(net162),
    .A1(net355),
    .S(_0517_),
    .X(_0066_));
 sg13g2_mux2_1 _1161_ (.A0(net156),
    .A1(net390),
    .S(_0517_),
    .X(_0067_));
 sg13g2_mux2_1 _1162_ (.A0(net151),
    .A1(net299),
    .S(_0517_),
    .X(_0068_));
 sg13g2_nand2b_2 _1163_ (.Y(_0518_),
    .B(_0505_),
    .A_N(_0497_));
 sg13g2_mux2_1 _1164_ (.A0(net183),
    .A1(net346),
    .S(net139),
    .X(_0069_));
 sg13g2_mux2_1 _1165_ (.A0(net176),
    .A1(net319),
    .S(net139),
    .X(_0070_));
 sg13g2_nand2_1 _1166_ (.Y(_0519_),
    .A(net257),
    .B(_0518_));
 sg13g2_o21ai_1 _1167_ (.B1(_0519_),
    .Y(_0071_),
    .A1(net148),
    .A2(net139));
 sg13g2_nand2_1 _1168_ (.Y(_0520_),
    .A(net256),
    .B(_0518_));
 sg13g2_o21ai_1 _1169_ (.B1(_0520_),
    .Y(_0072_),
    .A1(net147),
    .A2(net139));
 sg13g2_mux2_1 _1170_ (.A0(net163),
    .A1(net383),
    .S(net139),
    .X(_0073_));
 sg13g2_mux2_1 _1171_ (.A0(net158),
    .A1(net352),
    .S(net139),
    .X(_0074_));
 sg13g2_nand2_1 _1172_ (.Y(_0521_),
    .A(net253),
    .B(_0518_));
 sg13g2_o21ai_1 _1173_ (.B1(_0521_),
    .Y(_0075_),
    .A1(net146),
    .A2(net139));
 sg13g2_mux2_1 _1174_ (.A0(net149),
    .A1(net356),
    .S(net139),
    .X(_0076_));
 sg13g2_nand2_2 _1175_ (.Y(_0522_),
    .A(_0505_),
    .B(_0514_));
 sg13g2_mux2_1 _1176_ (.A0(net185),
    .A1(net340),
    .S(net138),
    .X(_0077_));
 sg13g2_mux2_1 _1177_ (.A0(net179),
    .A1(net398),
    .S(net138),
    .X(_0078_));
 sg13g2_nand2_1 _1178_ (.Y(_0523_),
    .A(net271),
    .B(net138));
 sg13g2_o21ai_1 _1179_ (.B1(_0523_),
    .Y(_0079_),
    .A1(_0169_),
    .A2(net138));
 sg13g2_nand2_1 _1180_ (.Y(_0524_),
    .A(net260),
    .B(_0522_));
 sg13g2_o21ai_1 _1181_ (.B1(_0524_),
    .Y(_0080_),
    .A1(_0170_),
    .A2(net138));
 sg13g2_mux2_1 _1182_ (.A0(net165),
    .A1(net379),
    .S(net138),
    .X(_0081_));
 sg13g2_mux2_1 _1183_ (.A0(net160),
    .A1(net350),
    .S(net138),
    .X(_0082_));
 sg13g2_nand2_1 _1184_ (.Y(_0525_),
    .A(net265),
    .B(_0522_));
 sg13g2_o21ai_1 _1185_ (.B1(_0525_),
    .Y(_0083_),
    .A1(net146),
    .A2(_0522_));
 sg13g2_mux2_1 _1186_ (.A0(net152),
    .A1(net378),
    .S(net138),
    .X(_0084_));
 sg13g2_nand2_2 _1187_ (.Y(_0526_),
    .A(_0500_),
    .B(_0514_));
 sg13g2_mux2_1 _1188_ (.A0(net182),
    .A1(net324),
    .S(net133),
    .X(_0085_));
 sg13g2_mux2_1 _1189_ (.A0(net177),
    .A1(net381),
    .S(net133),
    .X(_0086_));
 sg13g2_nand2_1 _1190_ (.Y(_0527_),
    .A(net268),
    .B(_0526_));
 sg13g2_o21ai_1 _1191_ (.B1(_0527_),
    .Y(_0087_),
    .A1(_0169_),
    .A2(net133));
 sg13g2_nand2_1 _1192_ (.Y(_0528_),
    .A(net264),
    .B(net133));
 sg13g2_o21ai_1 _1193_ (.B1(_0528_),
    .Y(_0088_),
    .A1(_0170_),
    .A2(net133));
 sg13g2_mux2_1 _1194_ (.A0(net163),
    .A1(net364),
    .S(net133),
    .X(_0089_));
 sg13g2_mux2_1 _1195_ (.A0(net158),
    .A1(net333),
    .S(net133),
    .X(_0090_));
 sg13g2_nand2_1 _1196_ (.Y(_0529_),
    .A(net259),
    .B(_0526_));
 sg13g2_o21ai_1 _1197_ (.B1(_0529_),
    .Y(_0091_),
    .A1(_0171_),
    .A2(_0526_));
 sg13g2_mux2_1 _1198_ (.A0(net150),
    .A1(net310),
    .S(net133),
    .X(_0092_));
 sg13g2_nand2_2 _1199_ (.Y(_0530_),
    .A(_0490_),
    .B(_0515_));
 sg13g2_mux2_1 _1200_ (.A0(net187),
    .A1(net300),
    .S(_0530_),
    .X(_0093_));
 sg13g2_mux2_1 _1201_ (.A0(net181),
    .A1(net318),
    .S(_0530_),
    .X(_0094_));
 sg13g2_mux2_1 _1202_ (.A0(net174),
    .A1(net335),
    .S(_0530_),
    .X(_0095_));
 sg13g2_mux2_1 _1203_ (.A0(net170),
    .A1(net303),
    .S(_0530_),
    .X(_0096_));
 sg13g2_mux2_1 _1204_ (.A0(net166),
    .A1(net400),
    .S(_0530_),
    .X(_0097_));
 sg13g2_mux2_1 _1205_ (.A0(net161),
    .A1(net309),
    .S(_0530_),
    .X(_0098_));
 sg13g2_mux2_1 _1206_ (.A0(net155),
    .A1(net362),
    .S(_0530_),
    .X(_0099_));
 sg13g2_mux2_1 _1207_ (.A0(net152),
    .A1(net396),
    .S(_0530_),
    .X(_0100_));
 sg13g2_o21ai_1 _1208_ (.B1(net145),
    .Y(_0531_),
    .A1(net4),
    .A2(net5));
 sg13g2_and2_1 _1209_ (.A(_0515_),
    .B(_0531_),
    .X(_0532_));
 sg13g2_mux2_1 _1210_ (.A0(net301),
    .A1(net187),
    .S(_0532_),
    .X(_0101_));
 sg13g2_mux2_1 _1211_ (.A0(net311),
    .A1(net181),
    .S(_0532_),
    .X(_0102_));
 sg13g2_mux2_1 _1212_ (.A0(net302),
    .A1(net175),
    .S(_0532_),
    .X(_0103_));
 sg13g2_mux2_1 _1213_ (.A0(net367),
    .A1(net169),
    .S(_0532_),
    .X(_0104_));
 sg13g2_mux2_1 _1214_ (.A0(net371),
    .A1(net167),
    .S(_0532_),
    .X(_0105_));
 sg13g2_mux2_1 _1215_ (.A0(net358),
    .A1(net160),
    .S(_0532_),
    .X(_0106_));
 sg13g2_mux2_1 _1216_ (.A0(net372),
    .A1(net156),
    .S(_0532_),
    .X(_0107_));
 sg13g2_mux2_1 _1217_ (.A0(net306),
    .A1(net153),
    .S(_0532_),
    .X(_0108_));
 sg13g2_and2_1 _1218_ (.A(_0494_),
    .B(_0531_),
    .X(_0533_));
 sg13g2_mux2_1 _1219_ (.A0(net304),
    .A1(net187),
    .S(_0533_),
    .X(_0109_));
 sg13g2_mux2_1 _1220_ (.A0(net336),
    .A1(net180),
    .S(_0533_),
    .X(_0110_));
 sg13g2_mux2_1 _1221_ (.A0(net387),
    .A1(net173),
    .S(_0533_),
    .X(_0111_));
 sg13g2_mux2_1 _1222_ (.A0(net354),
    .A1(net170),
    .S(_0533_),
    .X(_0112_));
 sg13g2_mux2_1 _1223_ (.A0(net397),
    .A1(net167),
    .S(_0533_),
    .X(_0113_));
 sg13g2_mux2_1 _1224_ (.A0(net322),
    .A1(net161),
    .S(_0533_),
    .X(_0114_));
 sg13g2_mux2_1 _1225_ (.A0(net320),
    .A1(net156),
    .S(_0533_),
    .X(_0115_));
 sg13g2_mux2_1 _1226_ (.A0(net348),
    .A1(net153),
    .S(_0533_),
    .X(_0116_));
 sg13g2_nor3_2 _1227_ (.A(net2),
    .B(_0493_),
    .C(_0497_),
    .Y(_0534_));
 sg13g2_mux2_1 _1228_ (.A0(net359),
    .A1(net183),
    .S(net132),
    .X(_0117_));
 sg13g2_mux2_1 _1229_ (.A0(net339),
    .A1(net177),
    .S(_0534_),
    .X(_0118_));
 sg13g2_nor2_1 _1230_ (.A(net277),
    .B(net132),
    .Y(_0535_));
 sg13g2_a21oi_1 _1231_ (.A1(net148),
    .A2(_0534_),
    .Y(_0119_),
    .B1(_0535_));
 sg13g2_nor2_1 _1232_ (.A(net279),
    .B(net132),
    .Y(_0536_));
 sg13g2_a21oi_1 _1233_ (.A1(net147),
    .A2(net132),
    .Y(_0120_),
    .B1(_0536_));
 sg13g2_mux2_1 _1234_ (.A0(net330),
    .A1(net164),
    .S(net132),
    .X(_0121_));
 sg13g2_mux2_1 _1235_ (.A0(net351),
    .A1(net159),
    .S(_0534_),
    .X(_0122_));
 sg13g2_nor2_1 _1236_ (.A(net289),
    .B(net132),
    .Y(_0537_));
 sg13g2_a21oi_1 _1237_ (.A1(net146),
    .A2(net132),
    .Y(_0123_),
    .B1(_0537_));
 sg13g2_mux2_1 _1238_ (.A0(net365),
    .A1(net149),
    .S(net132),
    .X(_0124_));
 sg13g2_nand2_2 _1239_ (.Y(_0538_),
    .A(_0505_),
    .B(_0531_));
 sg13g2_mux2_1 _1240_ (.A0(net184),
    .A1(net325),
    .S(_0538_),
    .X(_0125_));
 sg13g2_mux2_1 _1241_ (.A0(net178),
    .A1(net373),
    .S(net137),
    .X(_0126_));
 sg13g2_nand2_1 _1242_ (.Y(_0539_),
    .A(net272),
    .B(net137));
 sg13g2_o21ai_1 _1243_ (.B1(_0539_),
    .Y(_0127_),
    .A1(net148),
    .A2(net137));
 sg13g2_nand2_1 _1244_ (.Y(_0540_),
    .A(net258),
    .B(net137));
 sg13g2_o21ai_1 _1245_ (.B1(_0540_),
    .Y(_0128_),
    .A1(net147),
    .A2(net137));
 sg13g2_mux2_1 _1246_ (.A0(net164),
    .A1(net363),
    .S(_0538_),
    .X(_0129_));
 sg13g2_mux2_1 _1247_ (.A0(net159),
    .A1(net341),
    .S(_0538_),
    .X(_0130_));
 sg13g2_nand2_1 _1248_ (.Y(_0541_),
    .A(net273),
    .B(net137));
 sg13g2_o21ai_1 _1249_ (.B1(_0541_),
    .Y(_0131_),
    .A1(net146),
    .A2(net137));
 sg13g2_mux2_1 _1250_ (.A0(net150),
    .A1(net321),
    .S(net137),
    .X(_0132_));
 sg13g2_nand2_2 _1251_ (.Y(_0542_),
    .A(_0500_),
    .B(_0531_));
 sg13g2_mux2_1 _1252_ (.A0(net182),
    .A1(net327),
    .S(net131),
    .X(_0133_));
 sg13g2_mux2_1 _1253_ (.A0(net176),
    .A1(net332),
    .S(net131),
    .X(_0134_));
 sg13g2_nor2_1 _1254_ (.A(net172),
    .B(net131),
    .Y(_0543_));
 sg13g2_a21oi_1 _1255_ (.A1(_0173_),
    .A2(net131),
    .Y(_0135_),
    .B1(_0543_));
 sg13g2_nor2_1 _1256_ (.A(net168),
    .B(net131),
    .Y(_0544_));
 sg13g2_a21oi_1 _1257_ (.A1(_0174_),
    .A2(net131),
    .Y(_0136_),
    .B1(_0544_));
 sg13g2_mux2_1 _1258_ (.A0(net164),
    .A1(net386),
    .S(net131),
    .X(_0137_));
 sg13g2_mux2_1 _1259_ (.A0(net159),
    .A1(net347),
    .S(net131),
    .X(_0138_));
 sg13g2_nor2_1 _1260_ (.A(net154),
    .B(_0542_),
    .Y(_0545_));
 sg13g2_a21oi_1 _1261_ (.A1(_0175_),
    .A2(_0542_),
    .Y(_0139_),
    .B1(_0545_));
 sg13g2_mux2_1 _1262_ (.A0(net150),
    .A1(net344),
    .S(_0542_),
    .X(_0140_));
 sg13g2_nand2_1 _1263_ (.Y(_0546_),
    .A(net1),
    .B(_0207_));
 sg13g2_xor2_1 _1264_ (.B(\cam.mem[0][7] ),
    .A(net150),
    .X(_0547_));
 sg13g2_xnor2_1 _1265_ (.Y(_0548_),
    .A(net164),
    .B(\cam.mem[0][4] ));
 sg13g2_xor2_1 _1266_ (.B(\cam.mem[0][5] ),
    .A(net159),
    .X(_0549_));
 sg13g2_xor2_1 _1267_ (.B(\cam.mem[0][0] ),
    .A(net182),
    .X(_0550_));
 sg13g2_a221oi_1 _1268_ (.B2(net154),
    .C1(_0550_),
    .B1(_0175_),
    .A1(net148),
    .Y(_0551_),
    .A2(\cam.mem[0][2] ));
 sg13g2_a22oi_1 _1269_ (.Y(_0552_),
    .B1(\cam.mem[0][6] ),
    .B2(net146),
    .A2(_0174_),
    .A1(net168));
 sg13g2_xor2_1 _1270_ (.B(\cam.mem[0][1] ),
    .A(net176),
    .X(_0553_));
 sg13g2_a221oi_1 _1271_ (.B2(net147),
    .C1(_0553_),
    .B1(\cam.mem[0][3] ),
    .A1(net172),
    .Y(_0554_),
    .A2(_0173_));
 sg13g2_nand4_1 _1272_ (.B(_0551_),
    .C(_0552_),
    .A(_0548_),
    .Y(_0555_),
    .D(_0554_));
 sg13g2_nor3_1 _1273_ (.A(_0547_),
    .B(_0549_),
    .C(_0555_),
    .Y(_0556_));
 sg13g2_or3_1 _1274_ (.A(_0275_),
    .B(_0546_),
    .C(_0556_),
    .X(_0557_));
 sg13g2_nand4_1 _1275_ (.B(_0327_),
    .C(_0338_),
    .A(_0252_),
    .Y(_0558_),
    .D(_0386_));
 sg13g2_nor3_1 _1276_ (.A(_0428_),
    .B(_0557_),
    .C(_0558_),
    .Y(_0559_));
 sg13g2_a21oi_1 _1277_ (.A1(_0182_),
    .A2(_0546_),
    .Y(_0141_),
    .B1(_0559_));
 sg13g2_nor2_1 _1278_ (.A(net248),
    .B(_0463_),
    .Y(_0142_));
 sg13g2_nor2_1 _1279_ (.A(net248),
    .B(net389),
    .Y(_0560_));
 sg13g2_nor3_1 _1280_ (.A(_0451_),
    .B(_0463_),
    .C(_0560_),
    .Y(_0143_));
 sg13g2_o21ai_1 _1281_ (.B1(net136),
    .Y(_0561_),
    .A1(net262),
    .A2(_0451_));
 sg13g2_a21oi_1 _1282_ (.A1(net262),
    .A2(_0451_),
    .Y(_0144_),
    .B1(_0561_));
 sg13g2_a21oi_1 _1283_ (.A1(net262),
    .A2(_0451_),
    .Y(_0562_),
    .B1(net297));
 sg13g2_nor3_1 _1284_ (.A(_0168_),
    .B(_0452_),
    .C(net298),
    .Y(_0145_));
 sg13g2_o21ai_1 _1285_ (.B1(net190),
    .Y(_0563_),
    .A1(net141),
    .A2(_0452_));
 sg13g2_a21oi_1 _1286_ (.A1(net141),
    .A2(_0452_),
    .Y(_0146_),
    .B1(_0563_));
 sg13g2_and3_1 _1287_ (.X(_0564_),
    .A(net401),
    .B(net141),
    .C(_0452_));
 sg13g2_a21oi_1 _1288_ (.A1(net141),
    .A2(_0452_),
    .Y(_0565_),
    .B1(net401));
 sg13g2_nor3_1 _1289_ (.A(_0463_),
    .B(_0564_),
    .C(net402),
    .Y(_0147_));
 sg13g2_and2_1 _1290_ (.A(_0183_),
    .B(_0452_),
    .X(_0566_));
 sg13g2_nor2_1 _1291_ (.A(net405),
    .B(_0564_),
    .Y(_0567_));
 sg13g2_nor3_1 _1292_ (.A(_0463_),
    .B(_0566_),
    .C(net406),
    .Y(_0148_));
 sg13g2_xnor2_1 _1293_ (.Y(_0568_),
    .A(net295),
    .B(_0566_));
 sg13g2_nor2_1 _1294_ (.A(_0463_),
    .B(_0568_),
    .Y(_0149_));
 sg13g2_a21oi_1 _1295_ (.A1(net295),
    .A2(_0566_),
    .Y(_0569_),
    .B1(net249));
 sg13g2_and3_1 _1296_ (.X(_0570_),
    .A(net295),
    .B(net249),
    .C(_0566_));
 sg13g2_nor3_1 _1297_ (.A(_0463_),
    .B(_0569_),
    .C(_0570_),
    .Y(_0150_));
 sg13g2_a21oi_1 _1298_ (.A1(net404),
    .A2(_0570_),
    .Y(_0571_),
    .B1(_0463_));
 sg13g2_o21ai_1 _1299_ (.B1(_0571_),
    .Y(_0572_),
    .A1(net404),
    .A2(_0570_));
 sg13g2_inv_1 _1300_ (.Y(_0151_),
    .A(_0572_));
 sg13g2_and2_1 _1301_ (.A(net2),
    .B(net144),
    .X(_0152_));
 sg13g2_and2_1 _1302_ (.A(net186),
    .B(net144),
    .X(_0153_));
 sg13g2_and2_1 _1303_ (.A(net3),
    .B(net144),
    .X(_0154_));
 sg13g2_and2_1 _1304_ (.A(net178),
    .B(net143),
    .X(_0155_));
 sg13g2_and2_1 _1305_ (.A(net4),
    .B(net144),
    .X(_0156_));
 sg13g2_and2_1 _1306_ (.A(net175),
    .B(net143),
    .X(_0157_));
 sg13g2_and2_1 _1307_ (.A(net5),
    .B(net143),
    .X(_0158_));
 sg13g2_nor3_2 _1308_ (.A(_0493_),
    .B(_0497_),
    .C(_0498_),
    .Y(_0573_));
 sg13g2_mux2_1 _1309_ (.A0(net370),
    .A1(net185),
    .S(_0573_),
    .X(_0159_));
 sg13g2_mux2_1 _1310_ (.A0(net399),
    .A1(net179),
    .S(_0573_),
    .X(_0160_));
 sg13g2_nor2_1 _1311_ (.A(net290),
    .B(net130),
    .Y(_0574_));
 sg13g2_a21oi_1 _1312_ (.A1(net148),
    .A2(net130),
    .Y(_0161_),
    .B1(_0574_));
 sg13g2_nor2_1 _1313_ (.A(net278),
    .B(net130),
    .Y(_0575_));
 sg13g2_a21oi_1 _1314_ (.A1(net147),
    .A2(net130),
    .Y(_0162_),
    .B1(_0575_));
 sg13g2_mux2_1 _1315_ (.A0(net366),
    .A1(net165),
    .S(net130),
    .X(_0163_));
 sg13g2_mux2_1 _1316_ (.A0(net357),
    .A1(net162),
    .S(_0573_),
    .X(_0164_));
 sg13g2_nor2_1 _1317_ (.A(net284),
    .B(net130),
    .Y(_0576_));
 sg13g2_a21oi_1 _1318_ (.A1(_0171_),
    .A2(net130),
    .Y(_0165_),
    .B1(_0576_));
 sg13g2_mux2_1 _1319_ (.A0(net314),
    .A1(net151),
    .S(net130),
    .X(_0166_));
 sg13g2_dfrbpq_1 _1320_ (.RESET_B(net35),
    .D(_0010_),
    .Q(\fourhalt_latch.reg_n ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1321_ (.RESET_B(net26),
    .D(net247),
    .Q(\vga.hvsync_gen.vsync ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1322_ (.RESET_B(net50),
    .D(_0011_),
    .Q(\vga.hvsync_gen.vpos[0] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1323_ (.RESET_B(net48),
    .D(_0012_),
    .Q(\vga.hvsync_gen.vpos[1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _1324_ (.RESET_B(net46),
    .D(net375),
    .Q(\vga.hvsync_gen.vpos[2] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _1325_ (.RESET_B(net44),
    .D(net281),
    .Q(\vga.hvsync_gen.vpos[3] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1326_ (.RESET_B(net42),
    .D(net252),
    .Q(\vga.hvsync_gen.vpos[4] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1327_ (.RESET_B(net40),
    .D(_0016_),
    .Q(\vga.hvsync_gen.vpos[5] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _1328_ (.RESET_B(net38),
    .D(net288),
    .Q(\vga.hvsync_gen.vpos[6] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1329_ (.RESET_B(net33),
    .D(net293),
    .Q(\vga.hvsync_gen.vpos[7] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1330_ (.RESET_B(net31),
    .D(_0019_),
    .Q(\vga.hvsync_gen.vpos[8] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1331_ (.RESET_B(net36),
    .D(_0020_),
    .Q(\vga.hvsync_gen.vpos[9] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1332_ (.RESET_B(net37),
    .D(net250),
    .Q(\vga.hsync ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1333_ (.RESET_B(net190),
    .D(_0002_),
    .Q(\vga.counter[0] ),
    .CLK(net142));
 sg13g2_dfrbpq_2 _1334_ (.RESET_B(net190),
    .D(_0003_),
    .Q(\vga.counter[1] ),
    .CLK(net142));
 sg13g2_dfrbpq_1 _1335_ (.RESET_B(net190),
    .D(_0004_),
    .Q(\vga.counter[2] ),
    .CLK(net142));
 sg13g2_dfrbpq_1 _1336_ (.RESET_B(net190),
    .D(_0005_),
    .Q(\vga.counter[3] ),
    .CLK(net142));
 sg13g2_dfrbpq_2 _1337_ (.RESET_B(net191),
    .D(_0006_),
    .Q(\vga.counter[4] ),
    .CLK(net142));
 sg13g2_dfrbpq_2 _1338_ (.RESET_B(net191),
    .D(_0007_),
    .Q(\vga.counter[5] ),
    .CLK(net142));
 sg13g2_dfrbpq_2 _1339_ (.RESET_B(net191),
    .D(_0008_),
    .Q(\vga.counter[6] ),
    .CLK(net142));
 sg13g2_dfrbpq_1 _1340_ (.RESET_B(net191),
    .D(_0009_),
    .Q(\vga.counter[7] ),
    .CLK(\vga.hvsync_gen.vsync ));
 sg13g2_dfrbpq_1 _1341_ (.RESET_B(net29),
    .D(_0021_),
    .Q(\cam.mem[10][0] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1342_ (.RESET_B(net28),
    .D(_0022_),
    .Q(\cam.mem[10][1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1343_ (.RESET_B(net27),
    .D(_0023_),
    .Q(\cam.mem[10][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1344_ (.RESET_B(net25),
    .D(_0024_),
    .Q(\cam.mem[10][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1345_ (.RESET_B(net245),
    .D(_0025_),
    .Q(\cam.mem[10][4] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1346_ (.RESET_B(net244),
    .D(_0026_),
    .Q(\cam.mem[10][5] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1347_ (.RESET_B(net243),
    .D(_0027_),
    .Q(\cam.mem[10][6] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1348_ (.RESET_B(net242),
    .D(_0028_),
    .Q(\cam.mem[10][7] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1349_ (.RESET_B(net241),
    .D(_0029_),
    .Q(\cam.mem[12][0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1350_ (.RESET_B(net240),
    .D(_0030_),
    .Q(\cam.mem[12][1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1351_ (.RESET_B(net239),
    .D(_0031_),
    .Q(\cam.mem[12][2] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1352_ (.RESET_B(net238),
    .D(_0032_),
    .Q(\cam.mem[12][3] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1353_ (.RESET_B(net237),
    .D(_0033_),
    .Q(\cam.mem[12][4] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1354_ (.RESET_B(net236),
    .D(_0034_),
    .Q(\cam.mem[12][5] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1355_ (.RESET_B(net235),
    .D(_0035_),
    .Q(\cam.mem[12][6] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1356_ (.RESET_B(net234),
    .D(_0036_),
    .Q(\cam.mem[12][7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1357_ (.RESET_B(net233),
    .D(_0037_),
    .Q(\cam.mem[9][0] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1358_ (.RESET_B(net232),
    .D(_0038_),
    .Q(\cam.mem[9][1] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1359_ (.RESET_B(net231),
    .D(_0039_),
    .Q(\cam.mem[9][2] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1360_ (.RESET_B(net230),
    .D(_0040_),
    .Q(\cam.mem[9][3] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1361_ (.RESET_B(net229),
    .D(_0041_),
    .Q(\cam.mem[9][4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1362_ (.RESET_B(net228),
    .D(_0042_),
    .Q(\cam.mem[9][5] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1363_ (.RESET_B(net227),
    .D(_0043_),
    .Q(\cam.mem[9][6] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1364_ (.RESET_B(net226),
    .D(_0044_),
    .Q(\cam.mem[9][7] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1365_ (.RESET_B(net225),
    .D(_0045_),
    .Q(\cam.mem[8][0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1366_ (.RESET_B(net224),
    .D(_0046_),
    .Q(\cam.mem[8][1] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1367_ (.RESET_B(net223),
    .D(_0047_),
    .Q(\cam.mem[8][2] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1368_ (.RESET_B(net222),
    .D(_0048_),
    .Q(\cam.mem[8][3] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1369_ (.RESET_B(net221),
    .D(_0049_),
    .Q(\cam.mem[8][4] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1370_ (.RESET_B(net220),
    .D(_0050_),
    .Q(\cam.mem[8][5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1371_ (.RESET_B(net219),
    .D(_0051_),
    .Q(\cam.mem[8][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1372_ (.RESET_B(net218),
    .D(_0052_),
    .Q(\cam.mem[8][7] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1373_ (.RESET_B(net217),
    .D(_0053_),
    .Q(\cam.mem[7][0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1374_ (.RESET_B(net216),
    .D(_0054_),
    .Q(\cam.mem[7][1] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1375_ (.RESET_B(net215),
    .D(_0055_),
    .Q(\cam.mem[7][2] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1376_ (.RESET_B(net214),
    .D(_0056_),
    .Q(\cam.mem[7][3] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1377_ (.RESET_B(net213),
    .D(_0057_),
    .Q(\cam.mem[7][4] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1378_ (.RESET_B(net212),
    .D(_0058_),
    .Q(\cam.mem[7][5] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1379_ (.RESET_B(net211),
    .D(_0059_),
    .Q(\cam.mem[7][6] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1380_ (.RESET_B(net210),
    .D(_0060_),
    .Q(\cam.mem[7][7] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1381_ (.RESET_B(net209),
    .D(_0061_),
    .Q(\cam.mem[6][0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1382_ (.RESET_B(net208),
    .D(_0062_),
    .Q(\cam.mem[6][1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1383_ (.RESET_B(net207),
    .D(_0063_),
    .Q(\cam.mem[6][2] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1384_ (.RESET_B(net206),
    .D(_0064_),
    .Q(\cam.mem[6][3] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1385_ (.RESET_B(net205),
    .D(_0065_),
    .Q(\cam.mem[6][4] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1386_ (.RESET_B(net204),
    .D(_0066_),
    .Q(\cam.mem[6][5] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net203),
    .D(_0067_),
    .Q(\cam.mem[6][6] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1388_ (.RESET_B(net202),
    .D(_0068_),
    .Q(\cam.mem[6][7] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1389_ (.RESET_B(net201),
    .D(_0069_),
    .Q(\cam.mem[13][0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1390_ (.RESET_B(net200),
    .D(_0070_),
    .Q(\cam.mem[13][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net199),
    .D(_0071_),
    .Q(\cam.mem[13][2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1392_ (.RESET_B(net198),
    .D(_0072_),
    .Q(\cam.mem[13][3] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1393_ (.RESET_B(net197),
    .D(_0073_),
    .Q(\cam.mem[13][4] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1394_ (.RESET_B(net196),
    .D(_0074_),
    .Q(\cam.mem[13][5] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1395_ (.RESET_B(net195),
    .D(_0075_),
    .Q(\cam.mem[13][6] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1396_ (.RESET_B(net194),
    .D(_0076_),
    .Q(\cam.mem[13][7] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1397_ (.RESET_B(net193),
    .D(_0077_),
    .Q(\cam.mem[5][0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1398_ (.RESET_B(net129),
    .D(_0078_),
    .Q(\cam.mem[5][1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1399_ (.RESET_B(net128),
    .D(_0079_),
    .Q(\cam.mem[5][2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1400_ (.RESET_B(net127),
    .D(_0080_),
    .Q(\cam.mem[5][3] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1401_ (.RESET_B(net126),
    .D(_0081_),
    .Q(\cam.mem[5][4] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1402_ (.RESET_B(net125),
    .D(_0082_),
    .Q(\cam.mem[5][5] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1403_ (.RESET_B(net124),
    .D(_0083_),
    .Q(\cam.mem[5][6] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1404_ (.RESET_B(net123),
    .D(_0084_),
    .Q(\cam.mem[5][7] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1405_ (.RESET_B(net122),
    .D(_0085_),
    .Q(\cam.mem[4][0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1406_ (.RESET_B(net121),
    .D(_0086_),
    .Q(\cam.mem[4][1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1407_ (.RESET_B(net120),
    .D(_0087_),
    .Q(\cam.mem[4][2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1408_ (.RESET_B(net119),
    .D(_0088_),
    .Q(\cam.mem[4][3] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1409_ (.RESET_B(net118),
    .D(_0089_),
    .Q(\cam.mem[4][4] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1410_ (.RESET_B(net117),
    .D(_0090_),
    .Q(\cam.mem[4][5] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1411_ (.RESET_B(net116),
    .D(_0091_),
    .Q(\cam.mem[4][6] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1412_ (.RESET_B(net115),
    .D(_0092_),
    .Q(\cam.mem[4][7] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1413_ (.RESET_B(net114),
    .D(_0093_),
    .Q(\cam.mem[11][0] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1414_ (.RESET_B(net113),
    .D(_0094_),
    .Q(\cam.mem[11][1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1415_ (.RESET_B(net112),
    .D(_0095_),
    .Q(\cam.mem[11][2] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1416_ (.RESET_B(net111),
    .D(_0096_),
    .Q(\cam.mem[11][3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net110),
    .D(_0097_),
    .Q(\cam.mem[11][4] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1418_ (.RESET_B(net109),
    .D(_0098_),
    .Q(\cam.mem[11][5] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1419_ (.RESET_B(net108),
    .D(_0099_),
    .Q(\cam.mem[11][6] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net107),
    .D(_0100_),
    .Q(\cam.mem[11][7] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1421_ (.RESET_B(net106),
    .D(_0101_),
    .Q(\cam.mem[3][0] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net105),
    .D(_0102_),
    .Q(\cam.mem[3][1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1423_ (.RESET_B(net104),
    .D(_0103_),
    .Q(\cam.mem[3][2] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net103),
    .D(_0104_),
    .Q(\cam.mem[3][3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1425_ (.RESET_B(net102),
    .D(_0105_),
    .Q(\cam.mem[3][4] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1426_ (.RESET_B(net101),
    .D(_0106_),
    .Q(\cam.mem[3][5] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net100),
    .D(_0107_),
    .Q(\cam.mem[3][6] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net99),
    .D(_0108_),
    .Q(\cam.mem[3][7] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net98),
    .D(_0109_),
    .Q(\cam.mem[2][0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1430_ (.RESET_B(net97),
    .D(_0110_),
    .Q(\cam.mem[2][1] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1431_ (.RESET_B(net96),
    .D(_0111_),
    .Q(\cam.mem[2][2] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1432_ (.RESET_B(net95),
    .D(_0112_),
    .Q(\cam.mem[2][3] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1433_ (.RESET_B(net94),
    .D(_0113_),
    .Q(\cam.mem[2][4] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1434_ (.RESET_B(net93),
    .D(_0114_),
    .Q(\cam.mem[2][5] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1435_ (.RESET_B(net92),
    .D(_0115_),
    .Q(\cam.mem[2][6] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1436_ (.RESET_B(net91),
    .D(_0116_),
    .Q(\cam.mem[2][7] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1437_ (.RESET_B(net90),
    .D(_0117_),
    .Q(\cam.mem[14][0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1438_ (.RESET_B(net89),
    .D(_0118_),
    .Q(\cam.mem[14][1] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1439_ (.RESET_B(net88),
    .D(_0119_),
    .Q(\cam.mem[14][2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1440_ (.RESET_B(net87),
    .D(_0120_),
    .Q(\cam.mem[14][3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1441_ (.RESET_B(net86),
    .D(_0121_),
    .Q(\cam.mem[14][4] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1442_ (.RESET_B(net85),
    .D(_0122_),
    .Q(\cam.mem[14][5] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1443_ (.RESET_B(net84),
    .D(_0123_),
    .Q(\cam.mem[14][6] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1444_ (.RESET_B(net83),
    .D(_0124_),
    .Q(\cam.mem[14][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net82),
    .D(_0125_),
    .Q(\cam.mem[1][0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net81),
    .D(_0126_),
    .Q(\cam.mem[1][1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net80),
    .D(_0127_),
    .Q(\cam.mem[1][2] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1448_ (.RESET_B(net79),
    .D(_0128_),
    .Q(\cam.mem[1][3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1449_ (.RESET_B(net78),
    .D(_0129_),
    .Q(\cam.mem[1][4] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net77),
    .D(_0130_),
    .Q(\cam.mem[1][5] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1451_ (.RESET_B(net76),
    .D(_0131_),
    .Q(\cam.mem[1][6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1452_ (.RESET_B(net75),
    .D(_0132_),
    .Q(\cam.mem[1][7] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1453_ (.RESET_B(net74),
    .D(_0133_),
    .Q(\cam.mem[0][0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net73),
    .D(_0134_),
    .Q(\cam.mem[0][1] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net72),
    .D(_0135_),
    .Q(\cam.mem[0][2] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1456_ (.RESET_B(net71),
    .D(_0136_),
    .Q(\cam.mem[0][3] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net70),
    .D(_0137_),
    .Q(\cam.mem[0][4] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net69),
    .D(_0138_),
    .Q(\cam.mem[0][5] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1459_ (.RESET_B(net68),
    .D(_0139_),
    .Q(\cam.mem[0][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1460_ (.RESET_B(net67),
    .D(_0140_),
    .Q(\cam.mem[0][7] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1461_ (.RESET_B(net192),
    .D(_0141_),
    .Q(\cam.found ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1462_ (.RESET_B(net66),
    .D(_0142_),
    .Q(\vga.hvsync_gen.hpos[0] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1463_ (.RESET_B(net65),
    .D(_0143_),
    .Q(\vga.hvsync_gen.hpos[1] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1464_ (.RESET_B(net64),
    .D(net263),
    .Q(\vga.hvsync_gen.hpos[2] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1465_ (.RESET_B(net63),
    .D(_0145_),
    .Q(\vga.hvsync_gen.hpos[3] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1466_ (.RESET_B(net62),
    .D(_0146_),
    .Q(\vga.hvsync_gen.hpos[4] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1467_ (.RESET_B(net61),
    .D(net403),
    .Q(\vga.hvsync_gen.hpos[5] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1468_ (.RESET_B(net60),
    .D(_0148_),
    .Q(\vga.hvsync_gen.hpos[6] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1469_ (.RESET_B(net59),
    .D(_0149_),
    .Q(\vga.hvsync_gen.hpos[7] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1470_ (.RESET_B(net58),
    .D(_0150_),
    .Q(\vga.hvsync_gen.hpos[8] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1471_ (.RESET_B(net57),
    .D(_0151_),
    .Q(\vga.hvsync_gen.hpos[9] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1472_ (.RESET_B(net56),
    .D(_0152_),
    .Q(\onehalt_latch.reg_p ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1473_ (.RESET_B(net55),
    .D(_0153_),
    .Q(\onehalt_latch.reg_n ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1474_ (.RESET_B(net54),
    .D(_0154_),
    .Q(\twohalt_latch.reg_p ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1475_ (.RESET_B(net53),
    .D(_0155_),
    .Q(\twohalt_latch.reg_n ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1476_ (.RESET_B(net52),
    .D(_0156_),
    .Q(\treehalt_latch.reg_p ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1477_ (.RESET_B(net51),
    .D(_0157_),
    .Q(\treehalt_latch.reg_n ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1478_ (.RESET_B(net49),
    .D(_0158_),
    .Q(\fourhalt_latch.reg_p ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1479_ (.RESET_B(net47),
    .D(_0159_),
    .Q(\cam.mem[15][0] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1480_ (.RESET_B(net45),
    .D(_0160_),
    .Q(\cam.mem[15][1] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1481_ (.RESET_B(net43),
    .D(_0161_),
    .Q(\cam.mem[15][2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net41),
    .D(_0162_),
    .Q(\cam.mem[15][3] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1483_ (.RESET_B(net39),
    .D(_0163_),
    .Q(\cam.mem[15][4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1484_ (.RESET_B(net34),
    .D(_0164_),
    .Q(\cam.mem[15][5] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1485_ (.RESET_B(net32),
    .D(_0165_),
    .Q(\cam.mem[15][6] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1486_ (.RESET_B(net30),
    .D(_0166_),
    .Q(\cam.mem[15][7] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_tiehi _1321__26 (.L_HI(net26));
 sg13g2_tiehi _1343__27 (.L_HI(net27));
 sg13g2_tiehi _1342__28 (.L_HI(net28));
 sg13g2_tiehi _1341__29 (.L_HI(net29));
 sg13g2_tiehi _1486__30 (.L_HI(net30));
 sg13g2_tiehi _1330__31 (.L_HI(net31));
 sg13g2_tiehi _1485__32 (.L_HI(net32));
 sg13g2_tiehi _1329__33 (.L_HI(net33));
 sg13g2_tiehi _1484__34 (.L_HI(net34));
 sg13g2_tiehi _1320__35 (.L_HI(net35));
 sg13g2_tiehi _1331__36 (.L_HI(net36));
 sg13g2_tiehi _1332__37 (.L_HI(net37));
 sg13g2_tiehi _1328__38 (.L_HI(net38));
 sg13g2_tiehi _1483__39 (.L_HI(net39));
 sg13g2_tiehi _1327__40 (.L_HI(net40));
 sg13g2_tiehi _1482__41 (.L_HI(net41));
 sg13g2_tiehi _1326__42 (.L_HI(net42));
 sg13g2_tiehi _1481__43 (.L_HI(net43));
 sg13g2_tiehi _1325__44 (.L_HI(net44));
 sg13g2_tiehi _1480__45 (.L_HI(net45));
 sg13g2_tiehi _1324__46 (.L_HI(net46));
 sg13g2_tiehi _1479__47 (.L_HI(net47));
 sg13g2_tiehi _1323__48 (.L_HI(net48));
 sg13g2_tiehi _1478__49 (.L_HI(net49));
 sg13g2_tiehi _1322__50 (.L_HI(net50));
 sg13g2_tiehi _1477__51 (.L_HI(net51));
 sg13g2_tiehi _1476__52 (.L_HI(net52));
 sg13g2_tiehi _1475__53 (.L_HI(net53));
 sg13g2_tiehi _1474__54 (.L_HI(net54));
 sg13g2_tiehi _1473__55 (.L_HI(net55));
 sg13g2_tiehi _1472__56 (.L_HI(net56));
 sg13g2_tiehi _1471__57 (.L_HI(net57));
 sg13g2_tiehi _1470__58 (.L_HI(net58));
 sg13g2_tiehi _1469__59 (.L_HI(net59));
 sg13g2_tiehi _1468__60 (.L_HI(net60));
 sg13g2_tiehi _1467__61 (.L_HI(net61));
 sg13g2_tiehi _1466__62 (.L_HI(net62));
 sg13g2_tiehi _1465__63 (.L_HI(net63));
 sg13g2_tiehi _1464__64 (.L_HI(net64));
 sg13g2_tiehi _1463__65 (.L_HI(net65));
 sg13g2_tiehi _1462__66 (.L_HI(net66));
 sg13g2_tiehi _1460__67 (.L_HI(net67));
 sg13g2_tiehi _1459__68 (.L_HI(net68));
 sg13g2_tiehi _1458__69 (.L_HI(net69));
 sg13g2_tiehi _1457__70 (.L_HI(net70));
 sg13g2_tiehi _1456__71 (.L_HI(net71));
 sg13g2_tiehi _1455__72 (.L_HI(net72));
 sg13g2_tiehi _1454__73 (.L_HI(net73));
 sg13g2_tiehi _1453__74 (.L_HI(net74));
 sg13g2_tiehi _1452__75 (.L_HI(net75));
 sg13g2_tiehi _1451__76 (.L_HI(net76));
 sg13g2_tiehi _1450__77 (.L_HI(net77));
 sg13g2_tiehi _1449__78 (.L_HI(net78));
 sg13g2_tiehi _1448__79 (.L_HI(net79));
 sg13g2_tiehi _1447__80 (.L_HI(net80));
 sg13g2_tiehi _1446__81 (.L_HI(net81));
 sg13g2_tiehi _1445__82 (.L_HI(net82));
 sg13g2_tiehi _1444__83 (.L_HI(net83));
 sg13g2_tiehi _1443__84 (.L_HI(net84));
 sg13g2_tiehi _1442__85 (.L_HI(net85));
 sg13g2_tiehi _1441__86 (.L_HI(net86));
 sg13g2_tiehi _1440__87 (.L_HI(net87));
 sg13g2_tiehi _1439__88 (.L_HI(net88));
 sg13g2_tiehi _1438__89 (.L_HI(net89));
 sg13g2_tiehi _1437__90 (.L_HI(net90));
 sg13g2_tiehi _1436__91 (.L_HI(net91));
 sg13g2_tiehi _1435__92 (.L_HI(net92));
 sg13g2_tiehi _1434__93 (.L_HI(net93));
 sg13g2_tiehi _1433__94 (.L_HI(net94));
 sg13g2_tiehi _1432__95 (.L_HI(net95));
 sg13g2_tiehi _1431__96 (.L_HI(net96));
 sg13g2_tiehi _1430__97 (.L_HI(net97));
 sg13g2_tiehi _1429__98 (.L_HI(net98));
 sg13g2_tiehi _1428__99 (.L_HI(net99));
 sg13g2_tiehi _1427__100 (.L_HI(net100));
 sg13g2_tiehi _1426__101 (.L_HI(net101));
 sg13g2_tiehi _1425__102 (.L_HI(net102));
 sg13g2_tiehi _1424__103 (.L_HI(net103));
 sg13g2_tiehi _1423__104 (.L_HI(net104));
 sg13g2_tiehi _1422__105 (.L_HI(net105));
 sg13g2_tiehi _1421__106 (.L_HI(net106));
 sg13g2_tiehi _1420__107 (.L_HI(net107));
 sg13g2_tiehi _1419__108 (.L_HI(net108));
 sg13g2_tiehi _1418__109 (.L_HI(net109));
 sg13g2_tiehi _1417__110 (.L_HI(net110));
 sg13g2_tiehi _1416__111 (.L_HI(net111));
 sg13g2_tiehi _1415__112 (.L_HI(net112));
 sg13g2_tiehi _1414__113 (.L_HI(net113));
 sg13g2_tiehi _1413__114 (.L_HI(net114));
 sg13g2_tiehi _1412__115 (.L_HI(net115));
 sg13g2_tiehi _1411__116 (.L_HI(net116));
 sg13g2_tiehi _1410__117 (.L_HI(net117));
 sg13g2_tiehi _1409__118 (.L_HI(net118));
 sg13g2_tiehi _1408__119 (.L_HI(net119));
 sg13g2_tiehi _1407__120 (.L_HI(net120));
 sg13g2_tiehi _1406__121 (.L_HI(net121));
 sg13g2_tiehi _1405__122 (.L_HI(net122));
 sg13g2_tiehi _1404__123 (.L_HI(net123));
 sg13g2_tiehi _1403__124 (.L_HI(net124));
 sg13g2_tiehi _1402__125 (.L_HI(net125));
 sg13g2_tiehi _1401__126 (.L_HI(net126));
 sg13g2_tiehi _1400__127 (.L_HI(net127));
 sg13g2_tiehi _1399__128 (.L_HI(net128));
 sg13g2_tiehi _1398__129 (.L_HI(net129));
 sg13g2_tiehi _1397__130 (.L_HI(net193));
 sg13g2_tiehi _1396__131 (.L_HI(net194));
 sg13g2_tiehi _1395__132 (.L_HI(net195));
 sg13g2_tiehi _1394__133 (.L_HI(net196));
 sg13g2_tiehi _1393__134 (.L_HI(net197));
 sg13g2_tiehi _1392__135 (.L_HI(net198));
 sg13g2_tiehi _1391__136 (.L_HI(net199));
 sg13g2_tiehi _1390__137 (.L_HI(net200));
 sg13g2_tiehi _1389__138 (.L_HI(net201));
 sg13g2_tiehi _1388__139 (.L_HI(net202));
 sg13g2_tiehi _1387__140 (.L_HI(net203));
 sg13g2_tiehi _1386__141 (.L_HI(net204));
 sg13g2_tiehi _1385__142 (.L_HI(net205));
 sg13g2_tiehi _1384__143 (.L_HI(net206));
 sg13g2_tiehi _1383__144 (.L_HI(net207));
 sg13g2_tiehi _1382__145 (.L_HI(net208));
 sg13g2_tiehi _1381__146 (.L_HI(net209));
 sg13g2_tiehi _1380__147 (.L_HI(net210));
 sg13g2_tiehi _1379__148 (.L_HI(net211));
 sg13g2_tiehi _1378__149 (.L_HI(net212));
 sg13g2_tiehi _1377__150 (.L_HI(net213));
 sg13g2_tiehi _1376__151 (.L_HI(net214));
 sg13g2_tiehi _1375__152 (.L_HI(net215));
 sg13g2_tiehi _1374__153 (.L_HI(net216));
 sg13g2_tiehi _1373__154 (.L_HI(net217));
 sg13g2_tiehi _1372__155 (.L_HI(net218));
 sg13g2_tiehi _1371__156 (.L_HI(net219));
 sg13g2_tiehi _1370__157 (.L_HI(net220));
 sg13g2_tiehi _1369__158 (.L_HI(net221));
 sg13g2_tiehi _1368__159 (.L_HI(net222));
 sg13g2_tiehi _1367__160 (.L_HI(net223));
 sg13g2_tiehi _1366__161 (.L_HI(net224));
 sg13g2_tiehi _1365__162 (.L_HI(net225));
 sg13g2_tiehi _1364__163 (.L_HI(net226));
 sg13g2_tiehi _1363__164 (.L_HI(net227));
 sg13g2_tiehi _1362__165 (.L_HI(net228));
 sg13g2_tiehi _1361__166 (.L_HI(net229));
 sg13g2_tiehi _1360__167 (.L_HI(net230));
 sg13g2_tiehi _1359__168 (.L_HI(net231));
 sg13g2_tiehi _1358__169 (.L_HI(net232));
 sg13g2_tiehi _1357__170 (.L_HI(net233));
 sg13g2_tiehi _1356__171 (.L_HI(net234));
 sg13g2_tiehi _1355__172 (.L_HI(net235));
 sg13g2_tiehi _1354__173 (.L_HI(net236));
 sg13g2_tiehi _1353__174 (.L_HI(net237));
 sg13g2_tiehi _1352__175 (.L_HI(net238));
 sg13g2_tiehi _1351__176 (.L_HI(net239));
 sg13g2_tiehi _1350__177 (.L_HI(net240));
 sg13g2_tiehi _1349__178 (.L_HI(net241));
 sg13g2_tiehi _1348__179 (.L_HI(net242));
 sg13g2_tiehi _1347__180 (.L_HI(net243));
 sg13g2_tiehi _1346__181 (.L_HI(net244));
 sg13g2_tiehi _1345__182 (.L_HI(net245));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_jalcim_10 (.L_LO(net10));
 sg13g2_tielo tt_um_jalcim_11 (.L_LO(net11));
 sg13g2_tielo tt_um_jalcim_12 (.L_LO(net12));
 sg13g2_tielo tt_um_jalcim_13 (.L_LO(net13));
 sg13g2_tielo tt_um_jalcim_14 (.L_LO(net14));
 sg13g2_tielo tt_um_jalcim_15 (.L_LO(net15));
 sg13g2_tielo tt_um_jalcim_16 (.L_LO(net16));
 sg13g2_tielo tt_um_jalcim_17 (.L_LO(net17));
 sg13g2_tielo tt_um_jalcim_18 (.L_LO(net18));
 sg13g2_tielo tt_um_jalcim_19 (.L_LO(net19));
 sg13g2_tielo tt_um_jalcim_20 (.L_LO(net20));
 sg13g2_tielo tt_um_jalcim_21 (.L_LO(net21));
 sg13g2_tielo tt_um_jalcim_22 (.L_LO(net22));
 sg13g2_tielo tt_um_jalcim_23 (.L_LO(net23));
 sg13g2_tielo tt_um_jalcim_24 (.L_LO(net24));
 sg13g2_tiehi _1344__25 (.L_HI(net25));
 sg13g2_buf_8 fanout130 (.A(_0573_),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(_0542_),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(_0534_),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(_0526_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(_0510_),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(_0501_),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(_0462_),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(_0538_),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(_0522_),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(_0518_),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(_0506_),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(net407),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(\vga.hvsync_gen.vsync ),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(_0432_),
    .X(net143));
 sg13g2_buf_1 fanout144 (.A(_0432_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0206_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(_0171_),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(_0170_),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(_0169_),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(uio_in[7]),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net153),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(uio_in[7]),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(uio_in[7]),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(net157),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net157),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(uio_in[6]),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(net159),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(net162),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(uio_in[5]),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(net167),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(uio_in[4]),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net171),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(uio_in[3]),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net175),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(uio_in[2]),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(net178),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(uio_in[1]),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(net181),
    .X(net179));
 sg13g2_buf_8 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(uio_in[1]),
    .X(net181));
 sg13g2_buf_8 fanout182 (.A(net184),
    .X(net182));
 sg13g2_buf_1 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(uio_in[0]),
    .X(net184));
 sg13g2_buf_8 fanout185 (.A(net187),
    .X(net185));
 sg13g2_buf_8 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_8 fanout187 (.A(uio_in[0]),
    .X(net187));
 sg13g2_buf_8 fanout188 (.A(net8),
    .X(net188));
 sg13g2_buf_8 fanout189 (.A(net7),
    .X(net189));
 sg13g2_buf_8 fanout190 (.A(net192),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_8 fanout192 (.A(rst_n),
    .X(net192));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_jalcim_9 (.L_LO(net9));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vga.hvsync_gen.vpos[9] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0001_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold3 (.A(\vga.hvsync_gen.hpos[0] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold4 (.A(\vga.hvsync_gen.hpos[8] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0000_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold6 (.A(\vga.hvsync_gen.vpos[4] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0015_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cam.mem[13][6] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cam.mem[9][2] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cam.mem[8][2] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cam.mem[13][3] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cam.mem[13][2] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold13 (.A(\cam.mem[1][3] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cam.mem[4][6] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold15 (.A(\cam.mem[5][3] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cam.found ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold17 (.A(\vga.hvsync_gen.hpos[2] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0144_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold19 (.A(\cam.mem[4][3] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold20 (.A(\cam.mem[5][6] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cam.mem[9][3] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold22 (.A(\cam.mem[8][6] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cam.mem[4][2] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cam.mem[8][3] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold25 (.A(\cam.mem[9][6] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cam.mem[5][2] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cam.mem[1][2] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold28 (.A(\cam.mem[1][6] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cam.mem[0][6] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cam.mem[0][2] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cam.mem[12][3] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cam.mem[14][2] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold33 (.A(\cam.mem[15][3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cam.mem[14][3] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold35 (.A(\vga.hvsync_gen.vpos[3] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0014_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold37 (.A(\vga.hvsync_gen.vpos[8] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0487_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cam.mem[15][6] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cam.mem[0][3] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cam.mem[12][2] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold42 (.A(\vga.hvsync_gen.vpos[6] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0017_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cam.mem[14][6] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold45 (.A(\cam.mem[15][2] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cam.mem[12][6] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold47 (.A(\vga.hvsync_gen.vpos[7] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0018_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold49 (.A(\vga.hvsync_gen.vpos[5] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold50 (.A(\vga.hvsync_gen.hpos[7] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold51 (.A(\vga.hvsync_gen.vpos[0] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold52 (.A(\vga.hvsync_gen.hpos[3] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0562_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cam.mem[6][7] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cam.mem[11][0] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cam.mem[3][0] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cam.mem[3][2] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cam.mem[11][3] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cam.mem[2][0] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cam.mem[12][0] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cam.mem[3][7] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cam.mem[10][1] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cam.mem[8][5] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold64 (.A(\cam.mem[11][5] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cam.mem[4][7] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold66 (.A(\cam.mem[3][1] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cam.mem[10][4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cam.mem[9][4] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cam.mem[15][7] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cam.mem[9][0] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cam.mem[7][5] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cam.mem[6][2] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cam.mem[11][1] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cam.mem[13][1] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cam.mem[2][6] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold76 (.A(\cam.mem[1][7] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold77 (.A(\cam.mem[2][5] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cam.mem[7][0] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cam.mem[4][0] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cam.mem[1][0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cam.mem[8][1] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cam.mem[0][0] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cam.mem[8][4] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cam.mem[10][3] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cam.mem[14][4] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cam.mem[6][3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cam.mem[0][1] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cam.mem[4][5] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cam.mem[9][5] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cam.mem[11][2] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cam.mem[2][1] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cam.mem[10][0] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cam.mem[7][3] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cam.mem[14][1] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cam.mem[5][0] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cam.mem[1][5] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cam.mem[10][6] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cam.mem[12][4] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cam.mem[0][7] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cam.mem[6][4] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cam.mem[13][0] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cam.mem[0][5] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cam.mem[2][7] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cam.mem[8][7] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cam.mem[5][5] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cam.mem[14][5] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cam.mem[13][5] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cam.mem[12][7] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cam.mem[2][3] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cam.mem[6][5] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cam.mem[13][7] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cam.mem[15][5] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cam.mem[3][5] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cam.mem[14][0] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cam.mem[12][5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cam.mem[7][1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cam.mem[11][6] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cam.mem[1][4] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cam.mem[4][4] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cam.mem[14][7] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold121 (.A(\cam.mem[15][4] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cam.mem[3][3] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cam.mem[6][0] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cam.mem[7][7] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cam.mem[15][0] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cam.mem[3][4] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cam.mem[3][6] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cam.mem[1][1] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold129 (.A(\vga.hvsync_gen.vpos[2] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0013_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cam.mem[7][2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cam.mem[10][7] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cam.mem[5][7] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cam.mem[5][4] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold135 (.A(\vga.hvsync_gen.vpos[1] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold136 (.A(\cam.mem[4][1] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cam.mem[10][2] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cam.mem[13][4] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cam.mem[9][1] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cam.mem[12][1] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cam.mem[0][4] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cam.mem[2][2] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cam.mem[9][7] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold144 (.A(\vga.hvsync_gen.hpos[1] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cam.mem[6][6] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cam.mem[10][5] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cam.mem[7][6] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cam.mem[8][0] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cam.mem[6][1] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cam.mem[7][4] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cam.mem[11][7] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cam.mem[2][4] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cam.mem[5][1] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cam.mem[15][1] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cam.mem[11][4] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold156 (.A(\vga.hvsync_gen.hpos[5] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0565_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0147_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold159 (.A(\vga.hvsync_gen.hpos[9] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold160 (.A(\vga.hvsync_gen.hpos[6] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0567_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold162 (.A(\vga.hvsync_gen.hpos[4] ),
    .X(net407));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_4 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_169 ();
 sg13g2_decap_8 FILLER_0_176 ();
 sg13g2_decap_8 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_197 ();
 sg13g2_decap_8 FILLER_0_204 ();
 sg13g2_decap_8 FILLER_0_211 ();
 sg13g2_decap_8 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_fill_1 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_255 ();
 sg13g2_decap_4 FILLER_0_262 ();
 sg13g2_fill_1 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_fill_1 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_fill_2 FILLER_1_112 ();
 sg13g2_fill_1 FILLER_1_114 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_fill_1 FILLER_1_154 ();
 sg13g2_fill_1 FILLER_1_159 ();
 sg13g2_decap_8 FILLER_1_199 ();
 sg13g2_decap_8 FILLER_1_206 ();
 sg13g2_decap_8 FILLER_1_213 ();
 sg13g2_fill_2 FILLER_1_220 ();
 sg13g2_fill_1 FILLER_1_222 ();
 sg13g2_decap_4 FILLER_1_227 ();
 sg13g2_decap_8 FILLER_1_293 ();
 sg13g2_decap_8 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_4 FILLER_2_105 ();
 sg13g2_fill_1 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_4 FILLER_2_144 ();
 sg13g2_fill_1 FILLER_2_148 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_fill_2 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_4 FILLER_3_98 ();
 sg13g2_fill_1 FILLER_3_102 ();
 sg13g2_fill_2 FILLER_3_107 ();
 sg13g2_fill_1 FILLER_3_109 ();
 sg13g2_fill_2 FILLER_3_148 ();
 sg13g2_fill_2 FILLER_3_180 ();
 sg13g2_fill_1 FILLER_3_205 ();
 sg13g2_fill_2 FILLER_3_243 ();
 sg13g2_decap_4 FILLER_3_278 ();
 sg13g2_fill_1 FILLER_3_282 ();
 sg13g2_fill_2 FILLER_3_293 ();
 sg13g2_decap_8 FILLER_3_345 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_fill_2 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_4 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_22 ();
 sg13g2_decap_8 FILLER_4_43 ();
 sg13g2_fill_1 FILLER_4_50 ();
 sg13g2_fill_2 FILLER_4_88 ();
 sg13g2_fill_1 FILLER_4_90 ();
 sg13g2_fill_1 FILLER_4_148 ();
 sg13g2_decap_4 FILLER_4_179 ();
 sg13g2_fill_1 FILLER_4_183 ();
 sg13g2_decap_8 FILLER_4_205 ();
 sg13g2_decap_4 FILLER_4_212 ();
 sg13g2_fill_2 FILLER_4_216 ();
 sg13g2_fill_2 FILLER_4_236 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_fill_2 FILLER_4_279 ();
 sg13g2_decap_4 FILLER_4_306 ();
 sg13g2_fill_2 FILLER_4_310 ();
 sg13g2_decap_4 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_11 ();
 sg13g2_fill_1 FILLER_5_54 ();
 sg13g2_fill_2 FILLER_5_59 ();
 sg13g2_decap_4 FILLER_5_75 ();
 sg13g2_fill_2 FILLER_5_88 ();
 sg13g2_fill_1 FILLER_5_90 ();
 sg13g2_fill_1 FILLER_5_131 ();
 sg13g2_fill_2 FILLER_5_164 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_213 ();
 sg13g2_fill_1 FILLER_5_220 ();
 sg13g2_fill_2 FILLER_5_247 ();
 sg13g2_fill_1 FILLER_5_249 ();
 sg13g2_decap_4 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_263 ();
 sg13g2_fill_1 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_fill_2 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_4 FILLER_5_368 ();
 sg13g2_fill_1 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_11 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_fill_1 FILLER_6_57 ();
 sg13g2_fill_1 FILLER_6_96 ();
 sg13g2_fill_2 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_137 ();
 sg13g2_fill_1 FILLER_6_139 ();
 sg13g2_decap_8 FILLER_6_157 ();
 sg13g2_decap_8 FILLER_6_164 ();
 sg13g2_fill_2 FILLER_6_175 ();
 sg13g2_decap_4 FILLER_6_185 ();
 sg13g2_fill_2 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_4 FILLER_6_207 ();
 sg13g2_fill_2 FILLER_6_211 ();
 sg13g2_fill_2 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_229 ();
 sg13g2_decap_8 FILLER_6_275 ();
 sg13g2_decap_8 FILLER_6_282 ();
 sg13g2_decap_4 FILLER_6_289 ();
 sg13g2_fill_2 FILLER_6_293 ();
 sg13g2_decap_4 FILLER_6_303 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_34 ();
 sg13g2_decap_8 FILLER_7_64 ();
 sg13g2_fill_1 FILLER_7_71 ();
 sg13g2_decap_4 FILLER_7_81 ();
 sg13g2_fill_2 FILLER_7_85 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_128 ();
 sg13g2_fill_2 FILLER_7_150 ();
 sg13g2_fill_1 FILLER_7_152 ();
 sg13g2_decap_8 FILLER_7_157 ();
 sg13g2_decap_8 FILLER_7_164 ();
 sg13g2_fill_2 FILLER_7_171 ();
 sg13g2_fill_2 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_fill_2 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_fill_1 FILLER_7_348 ();
 sg13g2_fill_2 FILLER_7_357 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_85 ();
 sg13g2_decap_4 FILLER_8_92 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_224 ();
 sg13g2_fill_2 FILLER_8_340 ();
 sg13g2_fill_2 FILLER_8_357 ();
 sg13g2_fill_2 FILLER_8_381 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_fill_2 FILLER_9_81 ();
 sg13g2_fill_1 FILLER_9_83 ();
 sg13g2_decap_4 FILLER_9_169 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_220 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_decap_4 FILLER_9_234 ();
 sg13g2_fill_1 FILLER_9_238 ();
 sg13g2_fill_1 FILLER_9_247 ();
 sg13g2_fill_2 FILLER_9_275 ();
 sg13g2_fill_2 FILLER_9_286 ();
 sg13g2_decap_4 FILLER_9_296 ();
 sg13g2_fill_2 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_decap_4 FILLER_9_333 ();
 sg13g2_fill_2 FILLER_9_337 ();
 sg13g2_fill_2 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_4 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_18 ();
 sg13g2_fill_1 FILLER_10_23 ();
 sg13g2_fill_2 FILLER_10_55 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_fill_1 FILLER_10_115 ();
 sg13g2_fill_1 FILLER_10_125 ();
 sg13g2_fill_1 FILLER_10_150 ();
 sg13g2_decap_4 FILLER_10_168 ();
 sg13g2_fill_2 FILLER_10_172 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_232 ();
 sg13g2_decap_4 FILLER_10_239 ();
 sg13g2_fill_1 FILLER_10_243 ();
 sg13g2_decap_4 FILLER_10_271 ();
 sg13g2_decap_8 FILLER_10_288 ();
 sg13g2_fill_2 FILLER_10_295 ();
 sg13g2_fill_1 FILLER_10_297 ();
 sg13g2_decap_4 FILLER_10_308 ();
 sg13g2_fill_2 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_fill_2 FILLER_11_48 ();
 sg13g2_decap_8 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_fill_2 FILLER_11_95 ();
 sg13g2_fill_1 FILLER_11_97 ();
 sg13g2_decap_8 FILLER_11_125 ();
 sg13g2_decap_8 FILLER_11_132 ();
 sg13g2_decap_8 FILLER_11_139 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_decap_4 FILLER_11_166 ();
 sg13g2_fill_2 FILLER_11_210 ();
 sg13g2_decap_4 FILLER_11_221 ();
 sg13g2_fill_1 FILLER_11_225 ();
 sg13g2_fill_1 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_fill_1 FILLER_11_293 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_decap_4 FILLER_11_358 ();
 sg13g2_fill_2 FILLER_11_362 ();
 sg13g2_fill_2 FILLER_11_374 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_58 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_fill_2 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_decap_4 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_180 ();
 sg13g2_fill_1 FILLER_12_218 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_decap_4 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_293 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_decap_4 FILLER_12_345 ();
 sg13g2_fill_2 FILLER_12_357 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_9 ();
 sg13g2_fill_2 FILLER_13_50 ();
 sg13g2_fill_1 FILLER_13_101 ();
 sg13g2_decap_4 FILLER_13_181 ();
 sg13g2_decap_4 FILLER_13_219 ();
 sg13g2_fill_2 FILLER_13_302 ();
 sg13g2_fill_1 FILLER_13_304 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_4 FILLER_13_358 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_61 ();
 sg13g2_fill_2 FILLER_14_84 ();
 sg13g2_decap_4 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_fill_2 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_159 ();
 sg13g2_decap_4 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_174 ();
 sg13g2_decap_8 FILLER_14_181 ();
 sg13g2_decap_8 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_215 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_fill_1 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_4 FILLER_14_301 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_2 FILLER_14_333 ();
 sg13g2_fill_1 FILLER_14_335 ();
 sg13g2_fill_2 FILLER_14_344 ();
 sg13g2_fill_1 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_374 ();
 sg13g2_fill_1 FILLER_14_376 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_fill_2 FILLER_15_41 ();
 sg13g2_fill_1 FILLER_15_43 ();
 sg13g2_fill_2 FILLER_15_68 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_103 ();
 sg13g2_decap_8 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_117 ();
 sg13g2_decap_4 FILLER_15_122 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_fill_2 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_262 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_336 ();
 sg13g2_decap_4 FILLER_15_346 ();
 sg13g2_fill_2 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_fill_2 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_299 ();
 sg13g2_decap_4 FILLER_16_345 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_fill_2 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_43 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_4 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_74 ();
 sg13g2_decap_8 FILLER_17_92 ();
 sg13g2_decap_8 FILLER_17_99 ();
 sg13g2_decap_8 FILLER_17_106 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_fill_1 FILLER_17_214 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_2 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_4 FILLER_17_320 ();
 sg13g2_fill_2 FILLER_17_351 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_79 ();
 sg13g2_decap_8 FILLER_18_89 ();
 sg13g2_decap_4 FILLER_18_106 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_2 FILLER_18_138 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_decap_8 FILLER_18_195 ();
 sg13g2_decap_8 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_4 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_236 ();
 sg13g2_decap_8 FILLER_18_243 ();
 sg13g2_decap_8 FILLER_18_250 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_fill_1 FILLER_18_274 ();
 sg13g2_fill_2 FILLER_18_288 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_4 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_315 ();
 sg13g2_fill_1 FILLER_18_343 ();
 sg13g2_decap_4 FILLER_18_361 ();
 sg13g2_fill_2 FILLER_18_365 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_118 ();
 sg13g2_decap_4 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_142 ();
 sg13g2_decap_4 FILLER_19_149 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_fill_2 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_220 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_244 ();
 sg13g2_decap_4 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_fill_2 FILLER_19_292 ();
 sg13g2_fill_1 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_4 FILLER_19_308 ();
 sg13g2_fill_1 FILLER_19_312 ();
 sg13g2_decap_4 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_decap_4 FILLER_19_362 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_22 ();
 sg13g2_fill_1 FILLER_20_33 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_4 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_decap_4 FILLER_20_118 ();
 sg13g2_fill_2 FILLER_20_127 ();
 sg13g2_fill_2 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_fill_2 FILLER_20_145 ();
 sg13g2_decap_4 FILLER_20_174 ();
 sg13g2_decap_4 FILLER_20_203 ();
 sg13g2_decap_4 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_fill_2 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_decap_8 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_314 ();
 sg13g2_fill_2 FILLER_20_318 ();
 sg13g2_decap_4 FILLER_20_330 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_48 ();
 sg13g2_fill_1 FILLER_21_50 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_75 ();
 sg13g2_decap_8 FILLER_21_82 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_decap_8 FILLER_21_101 ();
 sg13g2_decap_4 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_fill_2 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_142 ();
 sg13g2_decap_4 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_184 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_decap_4 FILLER_21_254 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_266 ();
 sg13g2_decap_4 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_311 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_30 ();
 sg13g2_fill_1 FILLER_22_37 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_fill_1 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_2 FILLER_22_179 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_decap_4 FILLER_22_196 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_4 FILLER_22_259 ();
 sg13g2_decap_4 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_51 ();
 sg13g2_fill_2 FILLER_23_60 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_decap_4 FILLER_23_90 ();
 sg13g2_fill_1 FILLER_23_94 ();
 sg13g2_fill_2 FILLER_23_131 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_decap_4 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_decap_4 FILLER_23_251 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_decap_4 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_fill_1 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_30 ();
 sg13g2_decap_8 FILLER_24_48 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_92 ();
 sg13g2_fill_1 FILLER_24_121 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_170 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_fill_1 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_23 ();
 sg13g2_fill_1 FILLER_25_29 ();
 sg13g2_fill_2 FILLER_25_37 ();
 sg13g2_decap_8 FILLER_25_43 ();
 sg13g2_decap_4 FILLER_25_50 ();
 sg13g2_fill_2 FILLER_25_54 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_67 ();
 sg13g2_decap_8 FILLER_25_72 ();
 sg13g2_decap_8 FILLER_25_79 ();
 sg13g2_decap_8 FILLER_25_86 ();
 sg13g2_fill_2 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_fill_2 FILLER_25_104 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_162 ();
 sg13g2_decap_4 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_173 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_decap_4 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_263 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_4 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_4 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_decap_4 FILLER_25_373 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_fill_2 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_4 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_4 FILLER_26_168 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_fill_2 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_decap_4 FILLER_26_240 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_4 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_373 ();
 sg13g2_fill_1 FILLER_26_375 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_89 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_fill_2 FILLER_27_110 ();
 sg13g2_decap_8 FILLER_27_125 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_decap_4 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_234 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_decap_4 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_fill_2 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_1 FILLER_28_36 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_58 ();
 sg13g2_fill_2 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_fill_2 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_4 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_fill_2 FILLER_28_372 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_fill_2 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_26 ();
 sg13g2_fill_2 FILLER_29_55 ();
 sg13g2_fill_1 FILLER_29_57 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_115 ();
 sg13g2_fill_1 FILLER_29_117 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_165 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_decap_4 FILLER_29_314 ();
 sg13g2_fill_2 FILLER_29_318 ();
 sg13g2_decap_4 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_357 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_79 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_decap_4 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_decap_4 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_decap_8 FILLER_30_180 ();
 sg13g2_decap_8 FILLER_30_187 ();
 sg13g2_decap_4 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_241 ();
 sg13g2_decap_4 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_65 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_125 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_decap_4 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_decap_4 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_fill_2 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_45 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_1 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_decap_8 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_155 ();
 sg13g2_decap_8 FILLER_32_162 ();
 sg13g2_decap_8 FILLER_32_169 ();
 sg13g2_decap_4 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_decap_8 FILLER_32_232 ();
 sg13g2_fill_2 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_264 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_decap_4 FILLER_32_331 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_118 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_181 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_decap_8 FILLER_33_241 ();
 sg13g2_decap_4 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_256 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_decap_8 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_315 ();
 sg13g2_decap_4 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_decap_4 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_1 FILLER_34_36 ();
 sg13g2_decap_8 FILLER_34_142 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_255 ();
 sg13g2_decap_8 FILLER_34_262 ();
 sg13g2_fill_1 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_decap_4 FILLER_34_296 ();
 sg13g2_fill_2 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_96 ();
 sg13g2_fill_1 FILLER_35_107 ();
 sg13g2_decap_4 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_decap_4 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_35_239 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_312 ();
 sg13g2_decap_4 FILLER_35_323 ();
 sg13g2_fill_1 FILLER_35_327 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_362 ();
 sg13g2_decap_4 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_383 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_69 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_113 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_fill_1 FILLER_36_146 ();
 sg13g2_decap_4 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_195 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_decap_8 FILLER_36_247 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_fill_2 FILLER_37_74 ();
 sg13g2_fill_1 FILLER_37_76 ();
 sg13g2_fill_1 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_191 ();
 sg13g2_decap_4 FILLER_37_198 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_fill_1 FILLER_37_254 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_decap_4 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_25 ();
 sg13g2_fill_1 FILLER_38_30 ();
 sg13g2_fill_2 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_46 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_134 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_4 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_decap_8 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_251 ();
 sg13g2_decap_8 FILLER_38_258 ();
 sg13g2_decap_4 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_325 ();
 sg13g2_fill_2 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
